module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_inv ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _15030_ (.A(\cpu.dec.r_op[5] ),
    .X(_08295_));
 sg13g2_buf_1 _15031_ (.A(_08295_),
    .X(_08296_));
 sg13g2_buf_8 _15032_ (.A(\cpu.addr[13] ),
    .X(_08297_));
 sg13g2_buf_8 _15033_ (.A(net1156),
    .X(_08298_));
 sg13g2_buf_8 _15034_ (.A(\cpu.addr[12] ),
    .X(_08299_));
 sg13g2_buf_8 _15035_ (.A(_08299_),
    .X(_08300_));
 sg13g2_buf_2 _15036_ (.A(\cpu.addr[14] ),
    .X(_08301_));
 sg13g2_buf_8 _15037_ (.A(_08301_),
    .X(_08302_));
 sg13g2_buf_8 _15038_ (.A(net1095),
    .X(_08303_));
 sg13g2_mux4_1 _15039_ (.S0(net1096),
    .A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net937),
    .X(_08304_));
 sg13g2_mux4_1 _15040_ (.S0(net1096),
    .A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(net937),
    .X(_08305_));
 sg13g2_mux4_1 _15041_ (.S0(net1096),
    .A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(net937),
    .X(_08306_));
 sg13g2_mux4_1 _15042_ (.S0(net1096),
    .A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(_08303_),
    .X(_08307_));
 sg13g2_buf_2 _15043_ (.A(_00193_),
    .X(_08308_));
 sg13g2_inv_2 _15044_ (.Y(_08309_),
    .A(_08308_));
 sg13g2_buf_8 _15045_ (.A(\cpu.ex.ifetch ),
    .X(_08310_));
 sg13g2_buf_2 _15046_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08311_));
 sg13g2_nand2b_1 _15047_ (.Y(_08312_),
    .B(_08311_),
    .A_N(_08310_));
 sg13g2_nand2_1 _15048_ (.Y(_08313_),
    .A(_08309_),
    .B(_08312_));
 sg13g2_buf_8 _15049_ (.A(_08313_),
    .X(_08314_));
 sg13g2_buf_8 _15050_ (.A(\cpu.addr[15] ),
    .X(_08315_));
 sg13g2_buf_8 _15051_ (.A(_08315_),
    .X(_08316_));
 sg13g2_mux4_1 _15052_ (.S0(net824),
    .A0(_08304_),
    .A1(_08305_),
    .A2(_08306_),
    .A3(_08307_),
    .S1(net1094),
    .X(_08317_));
 sg13g2_nand2_1 _15053_ (.Y(_08318_),
    .A(_08298_),
    .B(_08317_));
 sg13g2_nor2_1 _15054_ (.A(_08299_),
    .B(net1094),
    .Y(_08319_));
 sg13g2_nand2b_1 _15055_ (.Y(_08320_),
    .B(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A_N(net1095));
 sg13g2_nand2_1 _15056_ (.Y(_08321_),
    .A(_08303_),
    .B(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_nand3_1 _15057_ (.B(_08320_),
    .C(_08321_),
    .A(_08319_),
    .Y(_08322_));
 sg13g2_nand2_1 _15058_ (.Y(_08323_),
    .A(_08299_),
    .B(_08315_));
 sg13g2_mux2_1 _15059_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S(_08301_),
    .X(_08324_));
 sg13g2_nor2_1 _15060_ (.A(_08323_),
    .B(_08324_),
    .Y(_08325_));
 sg13g2_nand2b_1 _15061_ (.Y(_08326_),
    .B(_08299_),
    .A_N(_08315_));
 sg13g2_buf_1 _15062_ (.A(_08326_),
    .X(_08327_));
 sg13g2_mux2_1 _15063_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S(_08301_),
    .X(_08328_));
 sg13g2_nor2_1 _15064_ (.A(_08327_),
    .B(_08328_),
    .Y(_08329_));
 sg13g2_nand2b_1 _15065_ (.Y(_08330_),
    .B(net1094),
    .A_N(_08299_));
 sg13g2_mux2_1 _15066_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .S(net1095),
    .X(_08331_));
 sg13g2_nor2_1 _15067_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sg13g2_inv_1 _15068_ (.Y(_08333_),
    .A(\cpu.addr[13] ));
 sg13g2_buf_1 _15069_ (.A(_08333_),
    .X(_08334_));
 sg13g2_nand3_1 _15070_ (.B(_08309_),
    .C(_08312_),
    .A(net1093),
    .Y(_08335_));
 sg13g2_nor4_1 _15071_ (.A(_08325_),
    .B(_08329_),
    .C(_08332_),
    .D(_08335_),
    .Y(_08336_));
 sg13g2_nand2b_1 _15072_ (.Y(_08337_),
    .B(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A_N(net937));
 sg13g2_nand2_1 _15073_ (.Y(_08338_),
    .A(net937),
    .B(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_nand3_1 _15074_ (.B(_08337_),
    .C(_08338_),
    .A(_08319_),
    .Y(_08339_));
 sg13g2_mux2_1 _15075_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S(net1095),
    .X(_08340_));
 sg13g2_nor2_1 _15076_ (.A(_08323_),
    .B(_08340_),
    .Y(_08341_));
 sg13g2_mux2_1 _15077_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S(_08302_),
    .X(_08342_));
 sg13g2_nor2_1 _15078_ (.A(_08327_),
    .B(_08342_),
    .Y(_08343_));
 sg13g2_mux2_1 _15079_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .S(_08302_),
    .X(_08344_));
 sg13g2_nor2_1 _15080_ (.A(_08330_),
    .B(_08344_),
    .Y(_08345_));
 sg13g2_nor2b_1 _15081_ (.A(_08310_),
    .B_N(_08311_),
    .Y(_08346_));
 sg13g2_o21ai_1 _15082_ (.B1(net1093),
    .Y(_08347_),
    .A1(_08308_),
    .A2(_08346_));
 sg13g2_nor4_1 _15083_ (.A(_08341_),
    .B(_08343_),
    .C(_08345_),
    .D(_08347_),
    .Y(_08348_));
 sg13g2_buf_8 _15084_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08349_));
 sg13g2_buf_2 _15085_ (.A(\cpu.ex.io_access ),
    .X(_08350_));
 sg13g2_buf_2 _15086_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08351_));
 sg13g2_buf_8 _15087_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08352_));
 sg13g2_nor2_1 _15088_ (.A(_08351_),
    .B(net1154),
    .Y(_08353_));
 sg13g2_buf_2 _15089_ (.A(_08353_),
    .X(_08354_));
 sg13g2_nor2_2 _15090_ (.A(_08350_),
    .B(_08354_),
    .Y(_08355_));
 sg13g2_nand2_1 _15091_ (.Y(_08356_),
    .A(net1155),
    .B(_08355_));
 sg13g2_a221oi_1 _15092_ (.B2(_08348_),
    .C1(_08356_),
    .B1(_08339_),
    .A1(_08322_),
    .Y(_08357_),
    .A2(_08336_));
 sg13g2_buf_1 _15093_ (.A(_08357_),
    .X(_08358_));
 sg13g2_nand2_1 _15094_ (.Y(_08359_),
    .A(_08318_),
    .B(_08358_));
 sg13g2_inv_1 _15095_ (.Y(_08360_),
    .A(_08359_));
 sg13g2_buf_1 _15096_ (.A(\cpu.ex.r_read_stall ),
    .X(_08361_));
 sg13g2_buf_1 _15097_ (.A(_08361_),
    .X(_08362_));
 sg13g2_nor2b_1 _15098_ (.A(net1092),
    .B_N(_00189_),
    .Y(_08363_));
 sg13g2_buf_2 _15099_ (.A(\cpu.dec.supmode ),
    .X(_08364_));
 sg13g2_nand3_1 _15100_ (.B(net1155),
    .C(_08310_),
    .A(_08364_),
    .Y(_08365_));
 sg13g2_buf_2 _15101_ (.A(\cpu.ex.pc[13] ),
    .X(_08366_));
 sg13g2_buf_8 _15102_ (.A(_08366_),
    .X(_08367_));
 sg13g2_buf_1 _15103_ (.A(\cpu.ex.pc[14] ),
    .X(_08368_));
 sg13g2_buf_8 _15104_ (.A(_08368_),
    .X(_08369_));
 sg13g2_mux4_1 _15105_ (.S0(net1091),
    .A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S1(net1090),
    .X(_08370_));
 sg13g2_mux4_1 _15106_ (.S0(_08366_),
    .A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S1(net1090),
    .X(_08371_));
 sg13g2_buf_8 _15107_ (.A(\cpu.ex.pc[12] ),
    .X(_08372_));
 sg13g2_inv_2 _15108_ (.Y(_08373_),
    .A(_08372_));
 sg13g2_mux2_1 _15109_ (.A0(_08370_),
    .A1(_08371_),
    .S(_08373_),
    .X(_08374_));
 sg13g2_buf_2 _15110_ (.A(\cpu.ex.pc[15] ),
    .X(_08375_));
 sg13g2_inv_1 _15111_ (.Y(_08376_),
    .A(_08375_));
 sg13g2_buf_1 _15112_ (.A(_08376_),
    .X(_08377_));
 sg13g2_o21ai_1 _15113_ (.B1(net936),
    .Y(_08378_),
    .A1(_08365_),
    .A2(_08374_));
 sg13g2_mux4_1 _15114_ (.S0(_08366_),
    .A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S1(net1090),
    .X(_08379_));
 sg13g2_nor2_1 _15115_ (.A(net1153),
    .B(_08379_),
    .Y(_08380_));
 sg13g2_nand2b_1 _15116_ (.Y(_08381_),
    .B(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A_N(_08368_));
 sg13g2_nand2_1 _15117_ (.Y(_08382_),
    .A(net1090),
    .B(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_and4_1 _15118_ (.A(net1153),
    .B(net1091),
    .C(_08381_),
    .D(_08382_),
    .X(_08383_));
 sg13g2_mux2_1 _15119_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(net1090),
    .X(_08384_));
 sg13g2_nor3_1 _15120_ (.A(_08373_),
    .B(net1091),
    .C(_08384_),
    .Y(_08385_));
 sg13g2_nor4_1 _15121_ (.A(_08377_),
    .B(_08380_),
    .C(_08383_),
    .D(_08385_),
    .Y(_08386_));
 sg13g2_nand2_1 _15122_ (.Y(_08387_),
    .A(net1155),
    .B(_08310_));
 sg13g2_mux4_1 _15123_ (.S0(net1153),
    .A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S1(net1090),
    .X(_08388_));
 sg13g2_mux4_1 _15124_ (.S0(net1153),
    .A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S1(_08368_),
    .X(_08389_));
 sg13g2_mux2_1 _15125_ (.A0(_08388_),
    .A1(_08389_),
    .S(net1091),
    .X(_08390_));
 sg13g2_or3_1 _15126_ (.A(_08364_),
    .B(_08387_),
    .C(_08390_),
    .X(_08391_));
 sg13g2_o21ai_1 _15127_ (.B1(_08391_),
    .Y(_08392_),
    .A1(_08365_),
    .A2(_08386_));
 sg13g2_mux4_1 _15128_ (.S0(_08367_),
    .A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S1(_08369_),
    .X(_08393_));
 sg13g2_mux4_1 _15129_ (.S0(_08367_),
    .A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S1(_08369_),
    .X(_08394_));
 sg13g2_mux2_1 _15130_ (.A0(_08393_),
    .A1(_08394_),
    .S(_08373_),
    .X(_08395_));
 sg13g2_nor4_1 _15131_ (.A(_08375_),
    .B(_08364_),
    .C(_08387_),
    .D(_08395_),
    .Y(_08396_));
 sg13g2_a21oi_1 _15132_ (.A1(_08378_),
    .A2(_08392_),
    .Y(_08397_),
    .B1(_08396_));
 sg13g2_buf_1 _15133_ (.A(_08397_),
    .X(_08398_));
 sg13g2_inv_1 _15134_ (.Y(_08399_),
    .A(_00197_));
 sg13g2_buf_1 _15135_ (.A(_00198_),
    .X(_08400_));
 sg13g2_inv_1 _15136_ (.Y(_08401_),
    .A(net1152));
 sg13g2_buf_1 _15137_ (.A(\cpu.cond[0] ),
    .X(_08402_));
 sg13g2_buf_8 _15138_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08403_));
 sg13g2_or2_1 _15139_ (.X(_08404_),
    .B(net1152),
    .A(net1151));
 sg13g2_nand2_1 _15140_ (.Y(_08405_),
    .A(net1151),
    .B(_08361_));
 sg13g2_nand3_1 _15141_ (.B(_08404_),
    .C(_08405_),
    .A(_08402_),
    .Y(_08406_));
 sg13g2_o21ai_1 _15142_ (.B1(_08406_),
    .Y(_08407_),
    .A1(_08401_),
    .A2(_08361_));
 sg13g2_buf_2 _15143_ (.A(_08407_),
    .X(_08408_));
 sg13g2_inv_1 _15144_ (.Y(_08409_),
    .A(_08355_));
 sg13g2_o21ai_1 _15145_ (.B1(_08409_),
    .Y(_08410_),
    .A1(_08399_),
    .A2(_08408_));
 sg13g2_buf_8 _15146_ (.A(net937),
    .X(_08411_));
 sg13g2_nand2_1 _15147_ (.Y(_08412_),
    .A(net1093),
    .B(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_nand2_1 _15148_ (.Y(_08413_),
    .A(net1156),
    .B(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_nand3_1 _15149_ (.B(_08412_),
    .C(_08413_),
    .A(_08319_),
    .Y(_08414_));
 sg13g2_mux2_1 _15150_ (.A0(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S(net1156),
    .X(_08415_));
 sg13g2_nor2_1 _15151_ (.A(_08323_),
    .B(_08415_),
    .Y(_08416_));
 sg13g2_mux2_1 _15152_ (.A0(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S(_08297_),
    .X(_08417_));
 sg13g2_nor2_1 _15153_ (.A(_08327_),
    .B(_08417_),
    .Y(_08418_));
 sg13g2_mux2_1 _15154_ (.A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[14] ),
    .S(net1156),
    .X(_08419_));
 sg13g2_nor2_1 _15155_ (.A(_08330_),
    .B(_08419_),
    .Y(_08420_));
 sg13g2_nor3_1 _15156_ (.A(_08416_),
    .B(_08418_),
    .C(_08420_),
    .Y(_08421_));
 sg13g2_nand4_1 _15157_ (.B(net824),
    .C(_08414_),
    .A(net823),
    .Y(_08422_),
    .D(_08421_));
 sg13g2_mux4_1 _15158_ (.S0(_08299_),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net937),
    .X(_08423_));
 sg13g2_or2_1 _15159_ (.X(_08424_),
    .B(_08423_),
    .A(net1156));
 sg13g2_inv_2 _15160_ (.Y(_08425_),
    .A(_08316_));
 sg13g2_mux2_1 _15161_ (.A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[30] ),
    .S(net1095),
    .X(_08426_));
 sg13g2_nor3_1 _15162_ (.A(net1096),
    .B(net1093),
    .C(_08426_),
    .Y(_08427_));
 sg13g2_inv_2 _15163_ (.Y(_08428_),
    .A(net1096));
 sg13g2_mux2_1 _15164_ (.A0(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S(net1095),
    .X(_08429_));
 sg13g2_nor3_1 _15165_ (.A(_08428_),
    .B(net1093),
    .C(_08429_),
    .Y(_08430_));
 sg13g2_nor4_1 _15166_ (.A(_08425_),
    .B(net824),
    .C(_08427_),
    .D(_08430_),
    .Y(_08431_));
 sg13g2_mux4_1 _15167_ (.S0(_08299_),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(net937),
    .X(_08432_));
 sg13g2_or2_1 _15168_ (.X(_08433_),
    .B(_08432_),
    .A(net1156));
 sg13g2_mux2_1 _15169_ (.A0(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S(net1095),
    .X(_08434_));
 sg13g2_nor3_1 _15170_ (.A(_08428_),
    .B(_08334_),
    .C(_08434_),
    .Y(_08435_));
 sg13g2_mux2_1 _15171_ (.A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[22] ),
    .S(net1095),
    .X(_08436_));
 sg13g2_nor3_1 _15172_ (.A(net1096),
    .B(_08334_),
    .C(_08436_),
    .Y(_08437_));
 sg13g2_nor4_1 _15173_ (.A(net1094),
    .B(net824),
    .C(_08435_),
    .D(_08437_),
    .Y(_08438_));
 sg13g2_a22oi_1 _15174_ (.Y(_08439_),
    .B1(_08433_),
    .B2(_08438_),
    .A2(_08431_),
    .A1(_08424_));
 sg13g2_mux4_1 _15175_ (.S0(net1096),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(net1156),
    .X(_08440_));
 sg13g2_nand2b_1 _15176_ (.Y(_08441_),
    .B(net1094),
    .A_N(_08440_));
 sg13g2_nor2_1 _15177_ (.A(_08308_),
    .B(_08346_),
    .Y(_08442_));
 sg13g2_buf_8 _15178_ (.A(_08442_),
    .X(_08443_));
 sg13g2_mux2_1 _15179_ (.A0(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S(net1156),
    .X(_08444_));
 sg13g2_nor2_1 _15180_ (.A(_08327_),
    .B(_08444_),
    .Y(_08445_));
 sg13g2_mux2_1 _15181_ (.A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ),
    .S(_08297_),
    .X(_08446_));
 sg13g2_nor2b_1 _15182_ (.A(_08446_),
    .B_N(_08319_),
    .Y(_08447_));
 sg13g2_nor4_1 _15183_ (.A(net823),
    .B(net822),
    .C(_08445_),
    .D(_08447_),
    .Y(_08448_));
 sg13g2_inv_2 _15184_ (.Y(_08449_),
    .A(_08349_));
 sg13g2_a21oi_1 _15185_ (.A1(_08441_),
    .A2(_08448_),
    .Y(_08450_),
    .B1(_08449_));
 sg13g2_nand4_1 _15186_ (.B(_08422_),
    .C(_08439_),
    .A(_08410_),
    .Y(_08451_),
    .D(_08450_));
 sg13g2_buf_8 _15187_ (.A(_08451_),
    .X(_08452_));
 sg13g2_a22oi_1 _15188_ (.Y(_08453_),
    .B1(net490),
    .B2(_08452_),
    .A2(_08363_),
    .A1(_08354_));
 sg13g2_buf_2 _15189_ (.A(_08453_),
    .X(_08454_));
 sg13g2_nor2_1 _15190_ (.A(_08360_),
    .B(_08454_),
    .Y(_08455_));
 sg13g2_buf_1 _15191_ (.A(_08455_),
    .X(_08456_));
 sg13g2_inv_2 _15192_ (.Y(_08457_),
    .A(net275));
 sg13g2_nor2_1 _15193_ (.A(_00189_),
    .B(_08457_),
    .Y(_08458_));
 sg13g2_buf_2 _15194_ (.A(_00192_),
    .X(_08459_));
 sg13g2_buf_1 _15195_ (.A(_08459_),
    .X(_08460_));
 sg13g2_buf_2 _15196_ (.A(net1153),
    .X(_08461_));
 sg13g2_buf_2 _15197_ (.A(net1088),
    .X(_08462_));
 sg13g2_buf_2 _15198_ (.A(net935),
    .X(_08463_));
 sg13g2_buf_1 _15199_ (.A(net1091),
    .X(_08464_));
 sg13g2_buf_2 _15200_ (.A(_08464_),
    .X(_08465_));
 sg13g2_buf_1 _15201_ (.A(net820),
    .X(_08466_));
 sg13g2_mux4_1 _15202_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net714),
    .X(_08467_));
 sg13g2_mux4_1 _15203_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net714),
    .X(_08468_));
 sg13g2_buf_2 _15204_ (.A(net935),
    .X(_08469_));
 sg13g2_buf_2 _15205_ (.A(net820),
    .X(_08470_));
 sg13g2_mux4_1 _15206_ (.S0(_08469_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net713),
    .X(_08471_));
 sg13g2_mux4_1 _15207_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(_08470_),
    .X(_08472_));
 sg13g2_buf_2 _15208_ (.A(net936),
    .X(_08473_));
 sg13g2_buf_2 _15209_ (.A(net818),
    .X(_08474_));
 sg13g2_buf_1 _15210_ (.A(net1090),
    .X(_08475_));
 sg13g2_buf_1 _15211_ (.A(net933),
    .X(_08476_));
 sg13g2_mux4_1 _15212_ (.S0(net712),
    .A0(_08467_),
    .A1(_08468_),
    .A2(_08471_),
    .A3(_08472_),
    .S1(net817),
    .X(_08477_));
 sg13g2_mux4_1 _15213_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net713),
    .X(_08478_));
 sg13g2_mux4_1 _15214_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net714),
    .X(_08479_));
 sg13g2_mux4_1 _15215_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net713),
    .X(_08480_));
 sg13g2_mux4_1 _15216_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(net713),
    .X(_08481_));
 sg13g2_mux4_1 _15217_ (.S0(net712),
    .A0(_08478_),
    .A1(_08479_),
    .A2(_08480_),
    .A3(_08481_),
    .S1(net817),
    .X(_08482_));
 sg13g2_buf_1 _15218_ (.A(_08364_),
    .X(_08483_));
 sg13g2_buf_1 _15219_ (.A(net1087),
    .X(_08484_));
 sg13g2_mux2_1 _15220_ (.A0(_08477_),
    .A1(_08482_),
    .S(net932),
    .X(_08485_));
 sg13g2_nand2b_1 _15221_ (.Y(_08486_),
    .B(_08485_),
    .A_N(net1089));
 sg13g2_buf_1 _15222_ (.A(_08486_),
    .X(_08487_));
 sg13g2_buf_2 _15223_ (.A(_00190_),
    .X(_08488_));
 sg13g2_buf_1 _15224_ (.A(_08488_),
    .X(_08489_));
 sg13g2_buf_2 _15225_ (.A(\cpu.ex.pc[2] ),
    .X(_08490_));
 sg13g2_buf_1 _15226_ (.A(\cpu.ex.pc[4] ),
    .X(_08491_));
 sg13g2_buf_8 _15227_ (.A(\cpu.ex.pc[3] ),
    .X(_08492_));
 sg13g2_nor2b_1 _15228_ (.A(net1150),
    .B_N(net1149),
    .Y(_08493_));
 sg13g2_nand2b_1 _15229_ (.Y(_08494_),
    .B(net1150),
    .A_N(net1149));
 sg13g2_o21ai_1 _15230_ (.B1(_08494_),
    .Y(_08495_),
    .A1(_08490_),
    .A2(_08493_));
 sg13g2_nand2_1 _15231_ (.Y(_08496_),
    .A(net1086),
    .B(_08495_));
 sg13g2_buf_2 _15232_ (.A(_08496_),
    .X(_08497_));
 sg13g2_buf_1 _15233_ (.A(_08497_),
    .X(_08498_));
 sg13g2_buf_1 _15234_ (.A(net637),
    .X(_08499_));
 sg13g2_buf_1 _15235_ (.A(_08499_),
    .X(_08500_));
 sg13g2_inv_2 _15236_ (.Y(_08501_),
    .A(_08490_));
 sg13g2_and2_1 _15237_ (.A(_08501_),
    .B(_08493_),
    .X(_08502_));
 sg13g2_buf_2 _15238_ (.A(_08502_),
    .X(_08503_));
 sg13g2_buf_1 _15239_ (.A(_08503_),
    .X(_08504_));
 sg13g2_buf_1 _15240_ (.A(_08504_),
    .X(_08505_));
 sg13g2_buf_1 _15241_ (.A(net636),
    .X(_08506_));
 sg13g2_nor3_1 _15242_ (.A(_08490_),
    .B(net1149),
    .C(_08488_),
    .Y(_08507_));
 sg13g2_buf_1 _15243_ (.A(_08507_),
    .X(_08508_));
 sg13g2_buf_1 _15244_ (.A(net931),
    .X(_08509_));
 sg13g2_buf_1 _15245_ (.A(net816),
    .X(_08510_));
 sg13g2_buf_1 _15246_ (.A(net710),
    .X(_08511_));
 sg13g2_a22oi_1 _15247_ (.Y(_08512_),
    .B1(net635),
    .B2(\cpu.icache.r_tag[4][21] ),
    .A2(net550),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_nor3_1 _15248_ (.A(_08501_),
    .B(net1149),
    .C(net1150),
    .Y(_08513_));
 sg13g2_buf_2 _15249_ (.A(_08513_),
    .X(_08514_));
 sg13g2_buf_1 _15250_ (.A(_08514_),
    .X(_08515_));
 sg13g2_buf_1 _15251_ (.A(net709),
    .X(_08516_));
 sg13g2_and2_1 _15252_ (.A(_08490_),
    .B(_08492_),
    .X(_08517_));
 sg13g2_buf_2 _15253_ (.A(_08517_),
    .X(_08518_));
 sg13g2_and2_1 _15254_ (.A(_08488_),
    .B(_08518_),
    .X(_08519_));
 sg13g2_buf_1 _15255_ (.A(_08519_),
    .X(_08520_));
 sg13g2_buf_2 _15256_ (.A(net708),
    .X(_08521_));
 sg13g2_buf_1 _15257_ (.A(net633),
    .X(_08522_));
 sg13g2_a22oi_1 _15258_ (.Y(_08523_),
    .B1(net549),
    .B2(\cpu.icache.r_tag[3][21] ),
    .A2(net634),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_buf_1 _15259_ (.A(_08489_),
    .X(_08524_));
 sg13g2_buf_1 _15260_ (.A(net930),
    .X(_08525_));
 sg13g2_buf_2 _15261_ (.A(_08490_),
    .X(_08526_));
 sg13g2_nor2b_1 _15262_ (.A(_08526_),
    .B_N(net1149),
    .Y(_08527_));
 sg13g2_buf_1 _15263_ (.A(_08527_),
    .X(_08528_));
 sg13g2_buf_2 _15264_ (.A(net1149),
    .X(_08529_));
 sg13g2_buf_2 _15265_ (.A(net1084),
    .X(_08530_));
 sg13g2_buf_1 _15266_ (.A(net929),
    .X(_08531_));
 sg13g2_mux2_1 _15267_ (.A0(\cpu.icache.r_tag[5][21] ),
    .A1(\cpu.icache.r_tag[7][21] ),
    .S(net813),
    .X(_08532_));
 sg13g2_buf_1 _15268_ (.A(net1085),
    .X(_08533_));
 sg13g2_buf_1 _15269_ (.A(_08533_),
    .X(_08534_));
 sg13g2_a22oi_1 _15270_ (.Y(_08535_),
    .B1(_08532_),
    .B2(net812),
    .A2(net814),
    .A1(\cpu.icache.r_tag[6][21] ));
 sg13g2_or2_1 _15271_ (.X(_08536_),
    .B(_08535_),
    .A(net815));
 sg13g2_nand4_1 _15272_ (.B(_08512_),
    .C(_08523_),
    .A(net489),
    .Y(_08537_),
    .D(_08536_));
 sg13g2_o21ai_1 _15273_ (.B1(_08537_),
    .Y(_08538_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net489));
 sg13g2_xor2_1 _15274_ (.B(_08538_),
    .A(net396),
    .X(_08539_));
 sg13g2_buf_1 _15275_ (.A(net1155),
    .X(_08540_));
 sg13g2_buf_2 _15276_ (.A(net1153),
    .X(_08541_));
 sg13g2_buf_1 _15277_ (.A(net1091),
    .X(_08542_));
 sg13g2_mux4_1 _15278_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net927),
    .X(_08543_));
 sg13g2_mux4_1 _15279_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net927),
    .X(_08544_));
 sg13g2_mux4_1 _15280_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(net934),
    .X(_08545_));
 sg13g2_mux4_1 _15281_ (.S0(_08541_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(_08542_),
    .X(_08546_));
 sg13g2_mux4_1 _15282_ (.S0(net936),
    .A0(_08543_),
    .A1(_08544_),
    .A2(_08545_),
    .A3(_08546_),
    .S1(net933),
    .X(_08547_));
 sg13g2_mux4_1 _15283_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net927),
    .X(_08548_));
 sg13g2_mux4_1 _15284_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net927),
    .X(_08549_));
 sg13g2_mux4_1 _15285_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net934),
    .X(_08550_));
 sg13g2_mux4_1 _15286_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net934),
    .X(_08551_));
 sg13g2_mux4_1 _15287_ (.S0(net936),
    .A0(_08548_),
    .A1(_08549_),
    .A2(_08550_),
    .A3(_08551_),
    .S1(net933),
    .X(_08552_));
 sg13g2_mux2_1 _15288_ (.A0(_08547_),
    .A1(_08552_),
    .S(net1087),
    .X(_08553_));
 sg13g2_nor2_1 _15289_ (.A(_08373_),
    .B(net1083),
    .Y(_08554_));
 sg13g2_a21oi_1 _15290_ (.A1(net1083),
    .A2(_08553_),
    .Y(_08555_),
    .B1(_08554_));
 sg13g2_buf_2 _15291_ (.A(_08555_),
    .X(_08556_));
 sg13g2_buf_1 _15292_ (.A(_08497_),
    .X(_08557_));
 sg13g2_nor2_1 _15293_ (.A(net1149),
    .B(_08488_),
    .Y(_08558_));
 sg13g2_and2_1 _15294_ (.A(net1085),
    .B(_08558_),
    .X(_08559_));
 sg13g2_buf_1 _15295_ (.A(_08559_),
    .X(_08560_));
 sg13g2_buf_1 _15296_ (.A(_08514_),
    .X(_08561_));
 sg13g2_a22oi_1 _15297_ (.Y(_08562_),
    .B1(net707),
    .B2(\cpu.icache.r_tag[1][12] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][12] ));
 sg13g2_a22oi_1 _15298_ (.Y(_08563_),
    .B1(net708),
    .B2(\cpu.icache.r_tag[3][12] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_mux2_1 _15299_ (.A0(\cpu.icache.r_tag[4][12] ),
    .A1(\cpu.icache.r_tag[6][12] ),
    .S(net1084),
    .X(_08564_));
 sg13g2_buf_2 _15300_ (.A(_08501_),
    .X(_08565_));
 sg13g2_a22oi_1 _15301_ (.Y(_08566_),
    .B1(_08564_),
    .B2(net926),
    .A2(_08518_),
    .A1(\cpu.icache.r_tag[7][12] ));
 sg13g2_or2_1 _15302_ (.X(_08567_),
    .B(_08566_),
    .A(net930));
 sg13g2_nand4_1 _15303_ (.B(_08562_),
    .C(_08563_),
    .A(net632),
    .Y(_08568_),
    .D(_08567_));
 sg13g2_o21ai_1 _15304_ (.B1(_08568_),
    .Y(_08569_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net551));
 sg13g2_xnor2_1 _15305_ (.Y(_08570_),
    .A(net488),
    .B(_08569_));
 sg13g2_mux4_1 _15306_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net934),
    .X(_08571_));
 sg13g2_mux4_1 _15307_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net934),
    .X(_08572_));
 sg13g2_mux4_1 _15308_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net934),
    .X(_08573_));
 sg13g2_mux4_1 _15309_ (.S0(_08461_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(_08464_),
    .X(_08574_));
 sg13g2_mux4_1 _15310_ (.S0(net936),
    .A0(_08571_),
    .A1(_08572_),
    .A2(_08573_),
    .A3(_08574_),
    .S1(net933),
    .X(_08575_));
 sg13g2_nand2_1 _15311_ (.Y(_08576_),
    .A(net1087),
    .B(_08575_));
 sg13g2_mux4_1 _15312_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net934),
    .X(_08577_));
 sg13g2_mux4_1 _15313_ (.S0(_08461_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net934),
    .X(_08578_));
 sg13g2_buf_2 _15314_ (.A(net1153),
    .X(_08579_));
 sg13g2_buf_2 _15315_ (.A(net1091),
    .X(_08580_));
 sg13g2_mux4_1 _15316_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(net925),
    .X(_08581_));
 sg13g2_mux4_1 _15317_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net925),
    .X(_08582_));
 sg13g2_mux4_1 _15318_ (.S0(net936),
    .A0(_08577_),
    .A1(_08578_),
    .A2(_08581_),
    .A3(_08582_),
    .S1(net933),
    .X(_08583_));
 sg13g2_nand2b_1 _15319_ (.Y(_08584_),
    .B(_08583_),
    .A_N(net1087));
 sg13g2_nand3_1 _15320_ (.B(_08576_),
    .C(_08584_),
    .A(net1083),
    .Y(_08585_));
 sg13g2_o21ai_1 _15321_ (.B1(_08585_),
    .Y(_08586_),
    .A1(net714),
    .A2(net1083));
 sg13g2_buf_2 _15322_ (.A(_08586_),
    .X(_08587_));
 sg13g2_buf_1 _15323_ (.A(_08497_),
    .X(_08588_));
 sg13g2_a22oi_1 _15324_ (.Y(_08589_),
    .B1(net707),
    .B2(\cpu.icache.r_tag[1][13] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][13] ));
 sg13g2_nor2_2 _15325_ (.A(_08490_),
    .B(_08488_),
    .Y(_08590_));
 sg13g2_and2_1 _15326_ (.A(net1084),
    .B(_08590_),
    .X(_08591_));
 sg13g2_buf_1 _15327_ (.A(_08591_),
    .X(_08592_));
 sg13g2_buf_1 _15328_ (.A(_08592_),
    .X(_08593_));
 sg13g2_a22oi_1 _15329_ (.Y(_08594_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][13] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][13] ));
 sg13g2_buf_1 _15330_ (.A(_08489_),
    .X(_08595_));
 sg13g2_mux2_1 _15331_ (.A0(\cpu.icache.r_tag[7][13] ),
    .A1(\cpu.icache.r_tag[3][13] ),
    .S(net924),
    .X(_08596_));
 sg13g2_buf_2 _15332_ (.A(_08518_),
    .X(_08597_));
 sg13g2_a22oi_1 _15333_ (.Y(_08598_),
    .B1(_08596_),
    .B2(net810),
    .A2(net816),
    .A1(\cpu.icache.r_tag[4][13] ));
 sg13g2_nand4_1 _15334_ (.B(_08589_),
    .C(_08594_),
    .A(net632),
    .Y(_08599_),
    .D(_08598_));
 sg13g2_o21ai_1 _15335_ (.B1(_08599_),
    .Y(_08600_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net631));
 sg13g2_xnor2_1 _15336_ (.Y(_08601_),
    .A(net437),
    .B(_08600_));
 sg13g2_nand2_1 _15337_ (.Y(_08602_),
    .A(_08570_),
    .B(_08601_));
 sg13g2_mux4_1 _15338_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net925),
    .X(_08603_));
 sg13g2_mux4_1 _15339_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net925),
    .X(_08604_));
 sg13g2_mux4_1 _15340_ (.S0(_08579_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(_08580_),
    .X(_08605_));
 sg13g2_mux4_1 _15341_ (.S0(_08579_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(_08580_),
    .X(_08606_));
 sg13g2_mux4_1 _15342_ (.S0(net936),
    .A0(_08603_),
    .A1(_08604_),
    .A2(_08605_),
    .A3(_08606_),
    .S1(_08475_),
    .X(_08607_));
 sg13g2_mux4_1 _15343_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net925),
    .X(_08608_));
 sg13g2_mux4_1 _15344_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net925),
    .X(_08609_));
 sg13g2_mux4_1 _15345_ (.S0(net1153),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1091),
    .X(_08610_));
 sg13g2_mux4_1 _15346_ (.S0(net1081),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net925),
    .X(_08611_));
 sg13g2_mux4_1 _15347_ (.S0(net936),
    .A0(_08608_),
    .A1(_08609_),
    .A2(_08610_),
    .A3(_08611_),
    .S1(net1090),
    .X(_08612_));
 sg13g2_mux2_1 _15348_ (.A0(_08607_),
    .A1(_08612_),
    .S(net1087),
    .X(_08613_));
 sg13g2_nand2b_1 _15349_ (.Y(_08614_),
    .B(_08613_),
    .A_N(net1089));
 sg13g2_buf_1 _15350_ (.A(_08614_),
    .X(_08615_));
 sg13g2_buf_1 _15351_ (.A(net631),
    .X(_08616_));
 sg13g2_buf_2 _15352_ (.A(_08530_),
    .X(_08617_));
 sg13g2_mux4_1 _15353_ (.S0(net928),
    .A0(\cpu.icache.r_tag[4][23] ),
    .A1(\cpu.icache.r_tag[5][23] ),
    .A2(\cpu.icache.r_tag[6][23] ),
    .A3(\cpu.icache.r_tag[7][23] ),
    .S1(net809),
    .X(_08618_));
 sg13g2_inv_1 _15354_ (.Y(_08619_),
    .A(net1086));
 sg13g2_buf_1 _15355_ (.A(_08503_),
    .X(_08620_));
 sg13g2_a22oi_1 _15356_ (.Y(_08621_),
    .B1(net708),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(net705),
    .A1(\cpu.icache.r_tag[2][23] ));
 sg13g2_inv_1 _15357_ (.Y(_08622_),
    .A(_08621_));
 sg13g2_a221oi_1 _15358_ (.B2(_08619_),
    .C1(_08622_),
    .B1(_08618_),
    .A1(\cpu.icache.r_tag[1][23] ),
    .Y(_08623_),
    .A2(net709));
 sg13g2_nor2_1 _15359_ (.A(\cpu.icache.r_tag[0][23] ),
    .B(net551),
    .Y(_08624_));
 sg13g2_a21oi_1 _15360_ (.A1(net548),
    .A2(_08623_),
    .Y(_08625_),
    .B1(_08624_));
 sg13g2_xnor2_1 _15361_ (.Y(_08626_),
    .A(net487),
    .B(_08625_));
 sg13g2_buf_2 _15362_ (.A(net935),
    .X(_08627_));
 sg13g2_buf_2 _15363_ (.A(net925),
    .X(_08628_));
 sg13g2_buf_2 _15364_ (.A(net807),
    .X(_08629_));
 sg13g2_mux4_1 _15365_ (.S0(_08627_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(_08629_),
    .X(_08630_));
 sg13g2_mux4_1 _15366_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net704),
    .X(_08631_));
 sg13g2_buf_1 _15367_ (.A(net1081),
    .X(_08632_));
 sg13g2_buf_2 _15368_ (.A(net923),
    .X(_08633_));
 sg13g2_buf_2 _15369_ (.A(net807),
    .X(_08634_));
 sg13g2_mux4_1 _15370_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net703),
    .X(_08635_));
 sg13g2_mux4_1 _15371_ (.S0(_08633_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(_08634_),
    .X(_08636_));
 sg13g2_buf_1 _15372_ (.A(net933),
    .X(_08637_));
 sg13g2_mux4_1 _15373_ (.S0(_08473_),
    .A0(_08630_),
    .A1(_08631_),
    .A2(_08635_),
    .A3(_08636_),
    .S1(net805),
    .X(_08638_));
 sg13g2_mux4_1 _15374_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net703),
    .X(_08639_));
 sg13g2_mux4_1 _15375_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net703),
    .X(_08640_));
 sg13g2_buf_2 _15376_ (.A(net923),
    .X(_08641_));
 sg13g2_buf_2 _15377_ (.A(net807),
    .X(_08642_));
 sg13g2_mux4_1 _15378_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net702),
    .X(_08643_));
 sg13g2_mux4_1 _15379_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net702),
    .X(_08644_));
 sg13g2_mux4_1 _15380_ (.S0(net818),
    .A0(_08639_),
    .A1(_08640_),
    .A2(_08643_),
    .A3(_08644_),
    .S1(net805),
    .X(_08645_));
 sg13g2_mux2_1 _15381_ (.A0(_08638_),
    .A1(_08645_),
    .S(net932),
    .X(_08646_));
 sg13g2_nand2b_1 _15382_ (.Y(_08647_),
    .B(_08646_),
    .A_N(net1089));
 sg13g2_buf_1 _15383_ (.A(_08647_),
    .X(_08648_));
 sg13g2_buf_1 _15384_ (.A(net811),
    .X(_08649_));
 sg13g2_a22oi_1 _15385_ (.Y(_08650_),
    .B1(net636),
    .B2(\cpu.icache.r_tag[2][18] ),
    .A2(net701),
    .A1(\cpu.icache.r_tag[5][18] ));
 sg13g2_a22oi_1 _15386_ (.Y(_08651_),
    .B1(net816),
    .B2(\cpu.icache.r_tag[4][18] ),
    .A2(net709),
    .A1(\cpu.icache.r_tag[1][18] ));
 sg13g2_mux2_1 _15387_ (.A0(\cpu.icache.r_tag[7][18] ),
    .A1(\cpu.icache.r_tag[3][18] ),
    .S(net924),
    .X(_08652_));
 sg13g2_a22oi_1 _15388_ (.Y(_08653_),
    .B1(_08652_),
    .B2(net928),
    .A2(_08590_),
    .A1(\cpu.icache.r_tag[6][18] ));
 sg13g2_nand2b_1 _15389_ (.Y(_08654_),
    .B(net809),
    .A_N(_08653_));
 sg13g2_nand3_1 _15390_ (.B(_08651_),
    .C(_08654_),
    .A(_08650_),
    .Y(_08655_));
 sg13g2_mux2_1 _15391_ (.A0(\cpu.icache.r_tag[0][18] ),
    .A1(_08655_),
    .S(net551),
    .X(_08656_));
 sg13g2_xnor2_1 _15392_ (.Y(_08657_),
    .A(_08648_),
    .B(_08656_));
 sg13g2_mux4_1 _15393_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(net807),
    .X(_08658_));
 sg13g2_mux4_1 _15394_ (.S0(_08632_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(_08628_),
    .X(_08659_));
 sg13g2_mux4_1 _15395_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(net807),
    .X(_08660_));
 sg13g2_mux4_1 _15396_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net807),
    .X(_08661_));
 sg13g2_mux4_1 _15397_ (.S0(net818),
    .A0(_08658_),
    .A1(_08659_),
    .A2(_08660_),
    .A3(_08661_),
    .S1(_08475_),
    .X(_08662_));
 sg13g2_mux4_1 _15398_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(_08628_),
    .X(_08663_));
 sg13g2_mux4_1 _15399_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net807),
    .X(_08664_));
 sg13g2_mux4_1 _15400_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net927),
    .X(_08665_));
 sg13g2_mux4_1 _15401_ (.S0(net923),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net807),
    .X(_08666_));
 sg13g2_mux4_1 _15402_ (.S0(net818),
    .A0(_08663_),
    .A1(_08664_),
    .A2(_08665_),
    .A3(_08666_),
    .S1(net933),
    .X(_08667_));
 sg13g2_mux2_1 _15403_ (.A0(_08662_),
    .A1(_08667_),
    .S(_08483_),
    .X(_08668_));
 sg13g2_nand2b_1 _15404_ (.Y(_08669_),
    .B(_08668_),
    .A_N(net1089));
 sg13g2_buf_1 _15405_ (.A(_08669_),
    .X(_08670_));
 sg13g2_mux4_1 _15406_ (.S0(net1085),
    .A0(\cpu.icache.r_tag[4][22] ),
    .A1(\cpu.icache.r_tag[5][22] ),
    .A2(\cpu.icache.r_tag[6][22] ),
    .A3(\cpu.icache.r_tag[7][22] ),
    .S1(net813),
    .X(_08671_));
 sg13g2_nand2_1 _15407_ (.Y(_08672_),
    .A(_08619_),
    .B(_08671_));
 sg13g2_a22oi_1 _15408_ (.Y(_08673_),
    .B1(net633),
    .B2(\cpu.icache.r_tag[3][22] ),
    .A2(net705),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_nand2_1 _15409_ (.Y(_08674_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net707));
 sg13g2_nand4_1 _15410_ (.B(_08672_),
    .C(_08673_),
    .A(net632),
    .Y(_08675_),
    .D(_08674_));
 sg13g2_o21ai_1 _15411_ (.B1(_08675_),
    .Y(_08676_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(net551));
 sg13g2_xnor2_1 _15412_ (.Y(_08677_),
    .A(net436),
    .B(_08676_));
 sg13g2_mux4_1 _15413_ (.S0(_08541_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(_08542_),
    .X(_08678_));
 sg13g2_mux4_1 _15414_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net927),
    .X(_08679_));
 sg13g2_mux4_1 _15415_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net927),
    .X(_08680_));
 sg13g2_mux4_1 _15416_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net927),
    .X(_08681_));
 sg13g2_mux4_1 _15417_ (.S0(_08375_),
    .A0(_08678_),
    .A1(_08679_),
    .A2(_08680_),
    .A3(_08681_),
    .S1(_08483_),
    .X(_08682_));
 sg13g2_nand2b_1 _15418_ (.Y(_08683_),
    .B(net1083),
    .A_N(_08682_));
 sg13g2_mux4_1 _15419_ (.S0(net935),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net820),
    .X(_08684_));
 sg13g2_mux4_1 _15420_ (.S0(net935),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net820),
    .X(_08685_));
 sg13g2_mux4_1 _15421_ (.S0(net935),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net820),
    .X(_08686_));
 sg13g2_mux4_1 _15422_ (.S0(_08462_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(_08465_),
    .X(_08687_));
 sg13g2_mux4_1 _15423_ (.S0(_08375_),
    .A0(_08684_),
    .A1(_08685_),
    .A2(_08686_),
    .A3(_08687_),
    .S1(net1087),
    .X(_08688_));
 sg13g2_nor2_1 _15424_ (.A(net817),
    .B(_08449_),
    .Y(_08689_));
 sg13g2_a22oi_1 _15425_ (.Y(_08690_),
    .B1(_08688_),
    .B2(_08689_),
    .A2(_08683_),
    .A1(net817));
 sg13g2_buf_2 _15426_ (.A(_08690_),
    .X(_08691_));
 sg13g2_mux4_1 _15427_ (.S0(net1085),
    .A0(\cpu.icache.r_tag[4][14] ),
    .A1(\cpu.icache.r_tag[5][14] ),
    .A2(\cpu.icache.r_tag[6][14] ),
    .A3(\cpu.icache.r_tag[7][14] ),
    .S1(net813),
    .X(_08692_));
 sg13g2_nand2_1 _15428_ (.Y(_08693_),
    .A(_08619_),
    .B(_08692_));
 sg13g2_a22oi_1 _15429_ (.Y(_08694_),
    .B1(net633),
    .B2(\cpu.icache.r_tag[3][14] ),
    .A2(net705),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_nand2_1 _15430_ (.Y(_08695_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(net707));
 sg13g2_nand4_1 _15431_ (.B(_08693_),
    .C(_08694_),
    .A(net632),
    .Y(_08696_),
    .D(_08695_));
 sg13g2_o21ai_1 _15432_ (.B1(_08696_),
    .Y(_08697_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net551));
 sg13g2_xnor2_1 _15433_ (.Y(_08698_),
    .A(net486),
    .B(_08697_));
 sg13g2_nand2_1 _15434_ (.Y(_08699_),
    .A(_08677_),
    .B(_08698_));
 sg13g2_or4_1 _15435_ (.A(_08602_),
    .B(_08626_),
    .C(_08657_),
    .D(_08699_),
    .X(_08700_));
 sg13g2_mux4_1 _15436_ (.S0(_08469_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(_08470_),
    .X(_08701_));
 sg13g2_mux4_1 _15437_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net713),
    .X(_08702_));
 sg13g2_buf_2 _15438_ (.A(net935),
    .X(_08703_));
 sg13g2_buf_2 _15439_ (.A(net820),
    .X(_08704_));
 sg13g2_mux4_1 _15440_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net700),
    .X(_08705_));
 sg13g2_mux4_1 _15441_ (.S0(_08703_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net700),
    .X(_08706_));
 sg13g2_mux4_1 _15442_ (.S0(net712),
    .A0(_08701_),
    .A1(_08702_),
    .A2(_08705_),
    .A3(_08706_),
    .S1(net817),
    .X(_08707_));
 sg13g2_mux4_1 _15443_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net700),
    .X(_08708_));
 sg13g2_mux4_1 _15444_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net700),
    .X(_08709_));
 sg13g2_mux4_1 _15445_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net704),
    .X(_08710_));
 sg13g2_mux4_1 _15446_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net704),
    .X(_08711_));
 sg13g2_mux4_1 _15447_ (.S0(net712),
    .A0(_08708_),
    .A1(_08709_),
    .A2(_08710_),
    .A3(_08711_),
    .S1(net805),
    .X(_08712_));
 sg13g2_mux2_1 _15448_ (.A0(_08707_),
    .A1(_08712_),
    .S(net932),
    .X(_08713_));
 sg13g2_nand2b_1 _15449_ (.Y(_08714_),
    .B(_08713_),
    .A_N(net1089));
 sg13g2_buf_2 _15450_ (.A(_08714_),
    .X(_08715_));
 sg13g2_buf_1 _15451_ (.A(net709),
    .X(_08716_));
 sg13g2_a22oi_1 _15452_ (.Y(_08717_),
    .B1(net710),
    .B2(\cpu.icache.r_tag[4][19] ),
    .A2(net630),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_a22oi_1 _15453_ (.Y(_08718_),
    .B1(net549),
    .B2(\cpu.icache.r_tag[3][19] ),
    .A2(net636),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_buf_1 _15454_ (.A(net930),
    .X(_08719_));
 sg13g2_mux2_1 _15455_ (.A0(\cpu.icache.r_tag[5][19] ),
    .A1(\cpu.icache.r_tag[7][19] ),
    .S(net929),
    .X(_08720_));
 sg13g2_a22oi_1 _15456_ (.Y(_08721_),
    .B1(net814),
    .B2(\cpu.icache.r_tag[6][19] ),
    .A2(_08720_),
    .A1(net928));
 sg13g2_or2_1 _15457_ (.X(_08722_),
    .B(_08721_),
    .A(net802));
 sg13g2_nand3_1 _15458_ (.B(_08718_),
    .C(_08722_),
    .A(_08717_),
    .Y(_08723_));
 sg13g2_mux2_1 _15459_ (.A0(\cpu.icache.r_tag[0][19] ),
    .A1(_08723_),
    .S(net548),
    .X(_08724_));
 sg13g2_xor2_1 _15460_ (.B(_08724_),
    .A(_08715_),
    .X(_08725_));
 sg13g2_mux4_1 _15461_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(_08704_),
    .X(_08726_));
 sg13g2_mux4_1 _15462_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net713),
    .X(_08727_));
 sg13g2_mux4_1 _15463_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net704),
    .X(_08728_));
 sg13g2_mux4_1 _15464_ (.S0(_08703_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(_08704_),
    .X(_08729_));
 sg13g2_mux4_1 _15465_ (.S0(net712),
    .A0(_08726_),
    .A1(_08727_),
    .A2(_08728_),
    .A3(_08729_),
    .S1(net817),
    .X(_08730_));
 sg13g2_mux4_1 _15466_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net700),
    .X(_08731_));
 sg13g2_mux4_1 _15467_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net700),
    .X(_08732_));
 sg13g2_mux4_1 _15468_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net704),
    .X(_08733_));
 sg13g2_mux4_1 _15469_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net704),
    .X(_08734_));
 sg13g2_mux4_1 _15470_ (.S0(net818),
    .A0(_08731_),
    .A1(_08732_),
    .A2(_08733_),
    .A3(_08734_),
    .S1(net805),
    .X(_08735_));
 sg13g2_mux2_1 _15471_ (.A0(_08730_),
    .A1(_08735_),
    .S(net932),
    .X(_08736_));
 sg13g2_nand2b_1 _15472_ (.Y(_08737_),
    .B(_08736_),
    .A_N(net1089));
 sg13g2_buf_2 _15473_ (.A(_08737_),
    .X(_08738_));
 sg13g2_buf_1 _15474_ (.A(net705),
    .X(_08739_));
 sg13g2_a22oi_1 _15475_ (.Y(_08740_),
    .B1(net629),
    .B2(\cpu.icache.r_tag[2][17] ),
    .A2(net630),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_a22oi_1 _15476_ (.Y(_08741_),
    .B1(net710),
    .B2(\cpu.icache.r_tag[4][17] ),
    .A2(net549),
    .A1(\cpu.icache.r_tag[3][17] ));
 sg13g2_mux2_1 _15477_ (.A0(\cpu.icache.r_tag[5][17] ),
    .A1(\cpu.icache.r_tag[7][17] ),
    .S(net929),
    .X(_08742_));
 sg13g2_buf_1 _15478_ (.A(_08533_),
    .X(_08743_));
 sg13g2_a22oi_1 _15479_ (.Y(_08744_),
    .B1(_08742_),
    .B2(net801),
    .A2(net814),
    .A1(\cpu.icache.r_tag[6][17] ));
 sg13g2_or2_1 _15480_ (.X(_08745_),
    .B(_08744_),
    .A(net802));
 sg13g2_nand4_1 _15481_ (.B(_08740_),
    .C(_08741_),
    .A(net548),
    .Y(_08746_),
    .D(_08745_));
 sg13g2_o21ai_1 _15482_ (.B1(_08746_),
    .Y(_08747_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(net489));
 sg13g2_xnor2_1 _15483_ (.Y(_08748_),
    .A(net394),
    .B(_08747_));
 sg13g2_nand2_1 _15484_ (.Y(_08749_),
    .A(_08725_),
    .B(_08748_));
 sg13g2_mux4_1 _15485_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net704),
    .X(_08750_));
 sg13g2_mux4_1 _15486_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net704),
    .X(_08751_));
 sg13g2_mux4_1 _15487_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net703),
    .X(_08752_));
 sg13g2_mux4_1 _15488_ (.S0(_08633_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(_08634_),
    .X(_08753_));
 sg13g2_mux4_1 _15489_ (.S0(net818),
    .A0(_08750_),
    .A1(_08751_),
    .A2(_08752_),
    .A3(_08753_),
    .S1(net805),
    .X(_08754_));
 sg13g2_mux4_1 _15490_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net703),
    .X(_08755_));
 sg13g2_mux4_1 _15491_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net703),
    .X(_08756_));
 sg13g2_mux4_1 _15492_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net702),
    .X(_08757_));
 sg13g2_mux4_1 _15493_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net702),
    .X(_08758_));
 sg13g2_mux4_1 _15494_ (.S0(net818),
    .A0(_08755_),
    .A1(_08756_),
    .A2(_08757_),
    .A3(_08758_),
    .S1(net805),
    .X(_08759_));
 sg13g2_mux2_1 _15495_ (.A0(_08754_),
    .A1(_08759_),
    .S(net932),
    .X(_08760_));
 sg13g2_nand2b_1 _15496_ (.Y(_08761_),
    .B(_08760_),
    .A_N(net1089));
 sg13g2_buf_2 _15497_ (.A(_08761_),
    .X(_08762_));
 sg13g2_mux2_1 _15498_ (.A0(\cpu.icache.r_tag[7][16] ),
    .A1(\cpu.icache.r_tag[3][16] ),
    .S(net930),
    .X(_08763_));
 sg13g2_a22oi_1 _15499_ (.Y(_08764_),
    .B1(_08763_),
    .B2(net810),
    .A2(net710),
    .A1(\cpu.icache.r_tag[4][16] ));
 sg13g2_a22oi_1 _15500_ (.Y(_08765_),
    .B1(net629),
    .B2(\cpu.icache.r_tag[2][16] ),
    .A2(net630),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_buf_2 _15501_ (.A(_08592_),
    .X(_08766_));
 sg13g2_a22oi_1 _15502_ (.Y(_08767_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(net701),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_nand4_1 _15503_ (.B(_08764_),
    .C(_08765_),
    .A(net548),
    .Y(_08768_),
    .D(_08767_));
 sg13g2_o21ai_1 _15504_ (.B1(_08768_),
    .Y(_08769_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net489));
 sg13g2_xnor2_1 _15505_ (.Y(_08770_),
    .A(_08762_),
    .B(_08769_));
 sg13g2_mux4_1 _15506_ (.S0(net808),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net703),
    .X(_08771_));
 sg13g2_mux4_1 _15507_ (.S0(_08627_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(_08629_),
    .X(_08772_));
 sg13g2_mux4_1 _15508_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net702),
    .X(_08773_));
 sg13g2_mux4_1 _15509_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net703),
    .X(_08774_));
 sg13g2_mux4_1 _15510_ (.S0(net933),
    .A0(_08771_),
    .A1(_08772_),
    .A2(_08773_),
    .A3(_08774_),
    .S1(net1087),
    .X(_08775_));
 sg13g2_a21oi_1 _15511_ (.A1(net1083),
    .A2(_08775_),
    .Y(_08776_),
    .B1(_08375_));
 sg13g2_mux4_1 _15512_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(net713),
    .X(_08777_));
 sg13g2_mux4_1 _15513_ (.S0(net819),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net713),
    .X(_08778_));
 sg13g2_mux4_1 _15514_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net700),
    .X(_08779_));
 sg13g2_mux4_1 _15515_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net700),
    .X(_08780_));
 sg13g2_mux4_1 _15516_ (.S0(net805),
    .A0(_08777_),
    .A1(_08778_),
    .A2(_08779_),
    .A3(_08780_),
    .S1(net1087),
    .X(_08781_));
 sg13g2_nor3_1 _15517_ (.A(net712),
    .B(_08449_),
    .C(_08781_),
    .Y(_08782_));
 sg13g2_or2_1 _15518_ (.X(_08783_),
    .B(_08782_),
    .A(_08776_));
 sg13g2_buf_2 _15519_ (.A(_08783_),
    .X(_08784_));
 sg13g2_a22oi_1 _15520_ (.Y(_08785_),
    .B1(net629),
    .B2(\cpu.icache.r_tag[2][15] ),
    .A2(net709),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_a22oi_1 _15521_ (.Y(_08786_),
    .B1(net710),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(net633),
    .A1(\cpu.icache.r_tag[3][15] ));
 sg13g2_mux2_1 _15522_ (.A0(\cpu.icache.r_tag[5][15] ),
    .A1(\cpu.icache.r_tag[7][15] ),
    .S(net929),
    .X(_08787_));
 sg13g2_a22oi_1 _15523_ (.Y(_08788_),
    .B1(_08787_),
    .B2(net928),
    .A2(net814),
    .A1(\cpu.icache.r_tag[6][15] ));
 sg13g2_or2_1 _15524_ (.X(_08789_),
    .B(_08788_),
    .A(net802));
 sg13g2_nand4_1 _15525_ (.B(_08785_),
    .C(_08786_),
    .A(net551),
    .Y(_08790_),
    .D(_08789_));
 sg13g2_o21ai_1 _15526_ (.B1(_08790_),
    .Y(_08791_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net489));
 sg13g2_xnor2_1 _15527_ (.Y(_08792_),
    .A(net392),
    .B(_08791_));
 sg13g2_mux4_1 _15528_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net702),
    .X(_08793_));
 sg13g2_mux4_1 _15529_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(_08642_),
    .X(_08794_));
 sg13g2_mux4_1 _15530_ (.S0(_08641_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(_08465_),
    .X(_08795_));
 sg13g2_mux4_1 _15531_ (.S0(_08641_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(_08642_),
    .X(_08796_));
 sg13g2_mux4_1 _15532_ (.S0(_08473_),
    .A0(_08793_),
    .A1(_08794_),
    .A2(_08795_),
    .A3(_08796_),
    .S1(_08637_),
    .X(_08797_));
 sg13g2_mux4_1 _15533_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net702),
    .X(_08798_));
 sg13g2_mux4_1 _15534_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(net702),
    .X(_08799_));
 sg13g2_mux4_1 _15535_ (.S0(net935),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net820),
    .X(_08800_));
 sg13g2_mux4_1 _15536_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(net820),
    .X(_08801_));
 sg13g2_mux4_1 _15537_ (.S0(net818),
    .A0(_08798_),
    .A1(_08799_),
    .A2(_08800_),
    .A3(_08801_),
    .S1(net805),
    .X(_08802_));
 sg13g2_mux2_1 _15538_ (.A0(_08797_),
    .A1(_08802_),
    .S(net932),
    .X(_08803_));
 sg13g2_nand2b_1 _15539_ (.Y(_08804_),
    .B(_08803_),
    .A_N(net1089));
 sg13g2_buf_1 _15540_ (.A(_08804_),
    .X(_08805_));
 sg13g2_a22oi_1 _15541_ (.Y(_08806_),
    .B1(net636),
    .B2(\cpu.icache.r_tag[2][20] ),
    .A2(net701),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_a22oi_1 _15542_ (.Y(_08807_),
    .B1(net710),
    .B2(\cpu.icache.r_tag[4][20] ),
    .A2(net709),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_mux2_1 _15543_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(net924),
    .X(_08808_));
 sg13g2_a22oi_1 _15544_ (.Y(_08809_),
    .B1(_08808_),
    .B2(net928),
    .A2(_08590_),
    .A1(\cpu.icache.r_tag[6][20] ));
 sg13g2_buf_1 _15545_ (.A(net809),
    .X(_08810_));
 sg13g2_nand2b_1 _15546_ (.Y(_08811_),
    .B(net698),
    .A_N(_08809_));
 sg13g2_nand3_1 _15547_ (.B(_08807_),
    .C(_08811_),
    .A(_08806_),
    .Y(_08812_));
 sg13g2_mux2_1 _15548_ (.A0(\cpu.icache.r_tag[0][20] ),
    .A1(_08812_),
    .S(net548),
    .X(_08813_));
 sg13g2_xor2_1 _15549_ (.B(_08813_),
    .A(_08805_),
    .X(_08814_));
 sg13g2_buf_2 _15550_ (.A(\cpu.ex.pc[5] ),
    .X(_08815_));
 sg13g2_mux2_1 _15551_ (.A0(\cpu.icache.r_tag[7][5] ),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net924),
    .X(_08816_));
 sg13g2_a22oi_1 _15552_ (.Y(_08817_),
    .B1(_08816_),
    .B2(net810),
    .A2(net931),
    .A1(\cpu.icache.r_tag[4][5] ));
 sg13g2_a22oi_1 _15553_ (.Y(_08818_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][5] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_buf_1 _15554_ (.A(_08514_),
    .X(_08819_));
 sg13g2_a22oi_1 _15555_ (.Y(_08820_),
    .B1(net697),
    .B2(\cpu.icache.r_tag[1][5] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][5] ));
 sg13g2_nand4_1 _15556_ (.B(_08817_),
    .C(_08818_),
    .A(net637),
    .Y(_08821_),
    .D(_08820_));
 sg13g2_o21ai_1 _15557_ (.B1(_08821_),
    .Y(_08822_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net631));
 sg13g2_xor2_1 _15558_ (.B(_08822_),
    .A(_08815_),
    .X(_08823_));
 sg13g2_buf_2 _15559_ (.A(\cpu.ex.pc[9] ),
    .X(_08824_));
 sg13g2_inv_1 _15560_ (.Y(_08825_),
    .A(_08824_));
 sg13g2_nand2_1 _15561_ (.Y(_08826_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(net697));
 sg13g2_a22oi_1 _15562_ (.Y(_08827_),
    .B1(net931),
    .B2(\cpu.icache.r_tag[4][9] ),
    .A2(net706),
    .A1(\cpu.icache.r_tag[6][9] ));
 sg13g2_and2_1 _15563_ (.A(_08619_),
    .B(_08518_),
    .X(_08828_));
 sg13g2_buf_2 _15564_ (.A(_08828_),
    .X(_08829_));
 sg13g2_and2_1 _15565_ (.A(net1084),
    .B(net1086),
    .X(_08830_));
 sg13g2_a22oi_1 _15566_ (.Y(_08831_),
    .B1(_08830_),
    .B2(\cpu.icache.r_tag[3][9] ),
    .A2(_08558_),
    .A1(\cpu.icache.r_tag[5][9] ));
 sg13g2_nor2_1 _15567_ (.A(net926),
    .B(_08831_),
    .Y(_08832_));
 sg13g2_a221oi_1 _15568_ (.B2(\cpu.icache.r_tag[7][9] ),
    .C1(_08832_),
    .B1(_08829_),
    .A1(\cpu.icache.r_tag[2][9] ),
    .Y(_08833_),
    .A2(_08503_));
 sg13g2_nand4_1 _15569_ (.B(_08826_),
    .C(_08827_),
    .A(net637),
    .Y(_08834_),
    .D(_08833_));
 sg13g2_o21ai_1 _15570_ (.B1(_08834_),
    .Y(_08835_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net631));
 sg13g2_xnor2_1 _15571_ (.Y(_08836_),
    .A(net1080),
    .B(_08835_));
 sg13g2_mux4_1 _15572_ (.S0(net801),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net698),
    .X(_08837_));
 sg13g2_mux4_1 _15573_ (.S0(net801),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net698),
    .X(_08838_));
 sg13g2_inv_1 _15574_ (.Y(_08839_),
    .A(_08491_));
 sg13g2_mux2_1 _15575_ (.A0(_08837_),
    .A1(_08838_),
    .S(_08839_),
    .X(_08840_));
 sg13g2_buf_1 _15576_ (.A(\cpu.ex.pc[10] ),
    .X(_08841_));
 sg13g2_a22oi_1 _15577_ (.Y(_08842_),
    .B1(net711),
    .B2(\cpu.icache.r_tag[2][10] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_a22oi_1 _15578_ (.Y(_08843_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][10] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][10] ));
 sg13g2_mux2_1 _15579_ (.A0(\cpu.icache.r_tag[7][10] ),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net1086),
    .X(_08844_));
 sg13g2_a22oi_1 _15580_ (.Y(_08845_),
    .B1(_08844_),
    .B2(_08518_),
    .A2(net931),
    .A1(\cpu.icache.r_tag[4][10] ));
 sg13g2_nand4_1 _15581_ (.B(_08842_),
    .C(_08843_),
    .A(net637),
    .Y(_08846_),
    .D(_08845_));
 sg13g2_o21ai_1 _15582_ (.B1(_08846_),
    .Y(_08847_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net632));
 sg13g2_xor2_1 _15583_ (.B(_08847_),
    .A(_08841_),
    .X(_08848_));
 sg13g2_nand4_1 _15584_ (.B(_08836_),
    .C(_08840_),
    .A(_08823_),
    .Y(_08849_),
    .D(_08848_));
 sg13g2_buf_1 _15585_ (.A(\cpu.ex.pc[8] ),
    .X(_08850_));
 sg13g2_inv_1 _15586_ (.Y(_08851_),
    .A(_08850_));
 sg13g2_buf_1 _15587_ (.A(_08851_),
    .X(_08852_));
 sg13g2_a22oi_1 _15588_ (.Y(_08853_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][8] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_a22oi_1 _15589_ (.Y(_08854_),
    .B1(net708),
    .B2(\cpu.icache.r_tag[3][8] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_nor2_1 _15590_ (.A(net1085),
    .B(net1084),
    .Y(_08855_));
 sg13g2_buf_2 _15591_ (.A(_08855_),
    .X(_08856_));
 sg13g2_mux2_1 _15592_ (.A0(\cpu.icache.r_tag[5][8] ),
    .A1(\cpu.icache.r_tag[7][8] ),
    .S(net1084),
    .X(_08857_));
 sg13g2_a22oi_1 _15593_ (.Y(_08858_),
    .B1(_08857_),
    .B2(net1085),
    .A2(_08856_),
    .A1(\cpu.icache.r_tag[4][8] ));
 sg13g2_or2_1 _15594_ (.X(_08859_),
    .B(_08858_),
    .A(net930));
 sg13g2_nand4_1 _15595_ (.B(_08853_),
    .C(_08854_),
    .A(net637),
    .Y(_08860_),
    .D(_08859_));
 sg13g2_o21ai_1 _15596_ (.B1(_08860_),
    .Y(_08861_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net631));
 sg13g2_xnor2_1 _15597_ (.Y(_08862_),
    .A(net922),
    .B(_08861_));
 sg13g2_buf_1 _15598_ (.A(\cpu.ex.pc[6] ),
    .X(_08863_));
 sg13g2_a22oi_1 _15599_ (.Y(_08864_),
    .B1(net697),
    .B2(\cpu.icache.r_tag[1][6] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_a22oi_1 _15600_ (.Y(_08865_),
    .B1(net708),
    .B2(\cpu.icache.r_tag[3][6] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][6] ));
 sg13g2_mux2_1 _15601_ (.A0(\cpu.icache.r_tag[4][6] ),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net1084),
    .X(_08866_));
 sg13g2_a22oi_1 _15602_ (.Y(_08867_),
    .B1(_08866_),
    .B2(_08501_),
    .A2(_08518_),
    .A1(\cpu.icache.r_tag[7][6] ));
 sg13g2_or2_1 _15603_ (.X(_08868_),
    .B(_08867_),
    .A(net930));
 sg13g2_nand4_1 _15604_ (.B(_08864_),
    .C(_08865_),
    .A(net637),
    .Y(_08869_),
    .D(_08868_));
 sg13g2_o21ai_1 _15605_ (.B1(_08869_),
    .Y(_08870_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net631));
 sg13g2_xor2_1 _15606_ (.B(_08870_),
    .A(_08863_),
    .X(_08871_));
 sg13g2_inv_1 _15607_ (.Y(_08872_),
    .A(\cpu.ex.pc[7] ));
 sg13g2_a22oi_1 _15608_ (.Y(_08873_),
    .B1(net931),
    .B2(\cpu.icache.r_tag[4][7] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_a22oi_1 _15609_ (.Y(_08874_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][7] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_buf_1 _15610_ (.A(_08558_),
    .X(_08875_));
 sg13g2_mux2_1 _15611_ (.A0(\cpu.icache.r_tag[7][7] ),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net1086),
    .X(_08876_));
 sg13g2_a22oi_1 _15612_ (.Y(_08877_),
    .B1(_08876_),
    .B2(net929),
    .A2(net921),
    .A1(\cpu.icache.r_tag[5][7] ));
 sg13g2_nand2b_1 _15613_ (.Y(_08878_),
    .B(net928),
    .A_N(_08877_));
 sg13g2_nand4_1 _15614_ (.B(_08873_),
    .C(_08874_),
    .A(net637),
    .Y(_08879_),
    .D(_08878_));
 sg13g2_o21ai_1 _15615_ (.B1(_08879_),
    .Y(_08880_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net631));
 sg13g2_xnor2_1 _15616_ (.Y(_08881_),
    .A(_08872_),
    .B(_08880_));
 sg13g2_inv_1 _15617_ (.Y(_08882_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15618_ (.A(_08882_),
    .X(_08883_));
 sg13g2_a22oi_1 _15619_ (.Y(_08884_),
    .B1(net697),
    .B2(\cpu.icache.r_tag[1][11] ),
    .A2(net811),
    .A1(\cpu.icache.r_tag[5][11] ));
 sg13g2_a22oi_1 _15620_ (.Y(_08885_),
    .B1(net706),
    .B2(\cpu.icache.r_tag[6][11] ),
    .A2(net711),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_mux2_1 _15621_ (.A0(\cpu.icache.r_tag[7][11] ),
    .A1(\cpu.icache.r_tag[3][11] ),
    .S(net924),
    .X(_08886_));
 sg13g2_a22oi_1 _15622_ (.Y(_08887_),
    .B1(_08886_),
    .B2(net810),
    .A2(net931),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_nand4_1 _15623_ (.B(_08884_),
    .C(_08885_),
    .A(net637),
    .Y(_08888_),
    .D(_08887_));
 sg13g2_o21ai_1 _15624_ (.B1(_08888_),
    .Y(_08889_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net632));
 sg13g2_xnor2_1 _15625_ (.Y(_08890_),
    .A(net1079),
    .B(_08889_));
 sg13g2_nand4_1 _15626_ (.B(_08871_),
    .C(_08881_),
    .A(_08862_),
    .Y(_08891_),
    .D(_08890_));
 sg13g2_nor2_1 _15627_ (.A(_08849_),
    .B(_08891_),
    .Y(_08892_));
 sg13g2_nand4_1 _15628_ (.B(_08792_),
    .C(_08814_),
    .A(_08770_),
    .Y(_08893_),
    .D(_08892_));
 sg13g2_nor4_2 _15629_ (.A(_08539_),
    .B(_08700_),
    .C(_08749_),
    .Y(_08894_),
    .D(_08893_));
 sg13g2_nand2_1 _15630_ (.Y(_08895_),
    .A(_08458_),
    .B(_08894_));
 sg13g2_buf_1 _15631_ (.A(_08895_),
    .X(_08896_));
 sg13g2_buf_1 _15632_ (.A(net174),
    .X(_08897_));
 sg13g2_buf_1 _15633_ (.A(\cpu.ex.pc[1] ),
    .X(_08898_));
 sg13g2_buf_1 _15634_ (.A(_08898_),
    .X(_08899_));
 sg13g2_nor2_1 _15635_ (.A(_00206_),
    .B(net632),
    .Y(_08900_));
 sg13g2_mux2_1 _15636_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(net930),
    .X(_08901_));
 sg13g2_a22oi_1 _15637_ (.Y(_08902_),
    .B1(_08901_),
    .B2(net809),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][17] ));
 sg13g2_nor2_1 _15638_ (.A(net926),
    .B(_08902_),
    .Y(_08903_));
 sg13g2_a22oi_1 _15639_ (.Y(_08904_),
    .B1(net636),
    .B2(\cpu.icache.r_data[2][17] ),
    .A2(net707),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_a22oi_1 _15640_ (.Y(_08905_),
    .B1(net816),
    .B2(\cpu.icache.r_data[4][17] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[6][17] ));
 sg13g2_nand2_1 _15641_ (.Y(_08906_),
    .A(_08904_),
    .B(_08905_));
 sg13g2_nor3_1 _15642_ (.A(_08900_),
    .B(_08903_),
    .C(_08906_),
    .Y(_08907_));
 sg13g2_and2_1 _15643_ (.A(net1086),
    .B(_08495_),
    .X(_08908_));
 sg13g2_buf_1 _15644_ (.A(_08908_),
    .X(_08909_));
 sg13g2_nand2_1 _15645_ (.Y(_08910_),
    .A(_00205_),
    .B(_08909_));
 sg13g2_mux2_1 _15646_ (.A0(\cpu.icache.r_data[4][1] ),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(net929),
    .X(_08911_));
 sg13g2_a22oi_1 _15647_ (.Y(_08912_),
    .B1(_08590_),
    .B2(_08911_),
    .A2(net633),
    .A1(\cpu.icache.r_data[3][1] ));
 sg13g2_a22oi_1 _15648_ (.Y(_08913_),
    .B1(net707),
    .B2(\cpu.icache.r_data[1][1] ),
    .A2(net701),
    .A1(\cpu.icache.r_data[5][1] ));
 sg13g2_a22oi_1 _15649_ (.Y(_08914_),
    .B1(_08829_),
    .B2(\cpu.icache.r_data[7][1] ),
    .A2(net705),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_nand4_1 _15650_ (.B(_08912_),
    .C(_08913_),
    .A(net632),
    .Y(_08915_),
    .D(_08914_));
 sg13g2_a21oi_1 _15651_ (.A1(_08910_),
    .A2(_08915_),
    .Y(_08916_),
    .B1(net1078));
 sg13g2_a21oi_1 _15652_ (.A1(net1078),
    .A2(_08907_),
    .Y(_08917_),
    .B1(_08916_));
 sg13g2_buf_1 _15653_ (.A(_08917_),
    .X(_08918_));
 sg13g2_buf_1 _15654_ (.A(net1078),
    .X(_08919_));
 sg13g2_buf_1 _15655_ (.A(net920),
    .X(_08920_));
 sg13g2_nor2_1 _15656_ (.A(_00204_),
    .B(net489),
    .Y(_08921_));
 sg13g2_mux2_1 _15657_ (.A0(\cpu.icache.r_data[5][16] ),
    .A1(\cpu.icache.r_data[7][16] ),
    .S(net809),
    .X(_08922_));
 sg13g2_a22oi_1 _15658_ (.Y(_08923_),
    .B1(_08922_),
    .B2(net812),
    .A2(_08856_),
    .A1(\cpu.icache.r_data[4][16] ));
 sg13g2_nor2_1 _15659_ (.A(net815),
    .B(_08923_),
    .Y(_08924_));
 sg13g2_buf_1 _15660_ (.A(net699),
    .X(_08925_));
 sg13g2_a22oi_1 _15661_ (.Y(_08926_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net550),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_a22oi_1 _15662_ (.Y(_08927_),
    .B1(net549),
    .B2(\cpu.icache.r_data[3][16] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][16] ));
 sg13g2_nand2_1 _15663_ (.Y(_08928_),
    .A(_08926_),
    .B(_08927_));
 sg13g2_nor3_1 _15664_ (.A(_08921_),
    .B(_08924_),
    .C(_08928_),
    .Y(_08929_));
 sg13g2_buf_1 _15665_ (.A(_08909_),
    .X(_08930_));
 sg13g2_buf_1 _15666_ (.A(net627),
    .X(_08931_));
 sg13g2_nand2_1 _15667_ (.Y(_08932_),
    .A(_00203_),
    .B(net547));
 sg13g2_a22oi_1 _15668_ (.Y(_08933_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][0] ),
    .A2(net550),
    .A1(\cpu.icache.r_data[2][0] ));
 sg13g2_a22oi_1 _15669_ (.Y(_08934_),
    .B1(net549),
    .B2(\cpu.icache.r_data[3][0] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_mux2_1 _15670_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(\cpu.icache.r_data[7][0] ),
    .S(net813),
    .X(_08935_));
 sg13g2_a22oi_1 _15671_ (.Y(_08936_),
    .B1(_08935_),
    .B2(net801),
    .A2(net814),
    .A1(\cpu.icache.r_data[6][0] ));
 sg13g2_or2_1 _15672_ (.X(_08937_),
    .B(_08936_),
    .A(net815));
 sg13g2_nand4_1 _15673_ (.B(_08933_),
    .C(_08934_),
    .A(net489),
    .Y(_08938_),
    .D(_08937_));
 sg13g2_a21oi_1 _15674_ (.A1(_08932_),
    .A2(_08938_),
    .Y(_08939_),
    .B1(_08919_));
 sg13g2_a21o_1 _15675_ (.A2(_08929_),
    .A1(net800),
    .B1(_08939_),
    .X(_08940_));
 sg13g2_buf_1 _15676_ (.A(_08940_),
    .X(_08941_));
 sg13g2_nor2_1 _15677_ (.A(net347),
    .B(_08941_),
    .Y(_08942_));
 sg13g2_buf_2 _15678_ (.A(_08942_),
    .X(_08943_));
 sg13g2_nor2_1 _15679_ (.A(_00202_),
    .B(net548),
    .Y(_08944_));
 sg13g2_mux2_1 _15680_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(net802),
    .X(_08945_));
 sg13g2_a22oi_1 _15681_ (.Y(_08946_),
    .B1(_08945_),
    .B2(net698),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][31] ));
 sg13g2_nor2_1 _15682_ (.A(net926),
    .B(_08946_),
    .Y(_08947_));
 sg13g2_a22oi_1 _15683_ (.Y(_08948_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][31] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_a22oi_1 _15684_ (.Y(_08949_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][31] ),
    .A2(net629),
    .A1(\cpu.icache.r_data[2][31] ));
 sg13g2_nand2_1 _15685_ (.Y(_08950_),
    .A(_08948_),
    .B(_08949_));
 sg13g2_nor3_1 _15686_ (.A(_08944_),
    .B(_08947_),
    .C(_08950_),
    .Y(_08951_));
 sg13g2_nand2_1 _15687_ (.Y(_08952_),
    .A(_00201_),
    .B(net547));
 sg13g2_and2_1 _15688_ (.A(\cpu.icache.r_data[5][15] ),
    .B(net701),
    .X(_08953_));
 sg13g2_a221oi_1 _15689_ (.B2(\cpu.icache.r_data[3][15] ),
    .C1(_08953_),
    .B1(net549),
    .A1(\cpu.icache.r_data[1][15] ),
    .Y(_08954_),
    .A2(net630));
 sg13g2_a22oi_1 _15690_ (.Y(_08955_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][15] ),
    .A2(_08739_),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_buf_1 _15691_ (.A(_08829_),
    .X(_08956_));
 sg13g2_a22oi_1 _15692_ (.Y(_08957_),
    .B1(net626),
    .B2(\cpu.icache.r_data[7][15] ),
    .A2(net628),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_nand4_1 _15693_ (.B(_08954_),
    .C(_08955_),
    .A(_08616_),
    .Y(_08958_),
    .D(_08957_));
 sg13g2_a21oi_1 _15694_ (.A1(_08952_),
    .A2(_08958_),
    .Y(_08959_),
    .B1(net920));
 sg13g2_a21o_1 _15695_ (.A2(_08951_),
    .A1(net800),
    .B1(_08959_),
    .X(_08960_));
 sg13g2_buf_1 _15696_ (.A(_08960_),
    .X(_08961_));
 sg13g2_a22oi_1 _15697_ (.Y(_08962_),
    .B1(_08925_),
    .B2(\cpu.icache.r_data[6][30] ),
    .A2(net629),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_mux2_1 _15698_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net802),
    .X(_08963_));
 sg13g2_a22oi_1 _15699_ (.Y(_08964_),
    .B1(net810),
    .B2(_08963_),
    .A2(_08716_),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_a22oi_1 _15700_ (.Y(_08965_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][30] ),
    .A2(net701),
    .A1(\cpu.icache.r_data[5][30] ));
 sg13g2_nand2_1 _15701_ (.Y(_08966_),
    .A(\cpu.icache.r_data[0][30] ),
    .B(_08930_));
 sg13g2_nand4_1 _15702_ (.B(_08964_),
    .C(_08965_),
    .A(_08962_),
    .Y(_08967_),
    .D(_08966_));
 sg13g2_a22oi_1 _15703_ (.Y(_08968_),
    .B1(net709),
    .B2(\cpu.icache.r_data[1][14] ),
    .A2(net701),
    .A1(\cpu.icache.r_data[5][14] ));
 sg13g2_a22oi_1 _15704_ (.Y(_08969_),
    .B1(net633),
    .B2(\cpu.icache.r_data[3][14] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][14] ));
 sg13g2_mux2_1 _15705_ (.A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(net929),
    .X(_08970_));
 sg13g2_a22oi_1 _15706_ (.Y(_08971_),
    .B1(_08970_),
    .B2(net926),
    .A2(_08518_),
    .A1(\cpu.icache.r_data[7][14] ));
 sg13g2_or2_1 _15707_ (.X(_08972_),
    .B(_08971_),
    .A(net930));
 sg13g2_nand4_1 _15708_ (.B(_08968_),
    .C(_08969_),
    .A(_08588_),
    .Y(_08973_),
    .D(_08972_));
 sg13g2_o21ai_1 _15709_ (.B1(_08973_),
    .Y(_08974_),
    .A1(\cpu.icache.r_data[0][14] ),
    .A2(net551));
 sg13g2_nor2_1 _15710_ (.A(net920),
    .B(_08974_),
    .Y(_08975_));
 sg13g2_a21oi_1 _15711_ (.A1(net920),
    .A2(_08967_),
    .Y(_08976_),
    .B1(_08975_));
 sg13g2_buf_1 _15712_ (.A(_08976_),
    .X(_08977_));
 sg13g2_mux2_1 _15713_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(net924),
    .X(_08978_));
 sg13g2_a22oi_1 _15714_ (.Y(_08979_),
    .B1(_08978_),
    .B2(net809),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][29] ));
 sg13g2_nand2b_1 _15715_ (.Y(_08980_),
    .B(net801),
    .A_N(_08979_));
 sg13g2_a22oi_1 _15716_ (.Y(_08981_),
    .B1(_08505_),
    .B2(\cpu.icache.r_data[2][29] ),
    .A2(_08515_),
    .A1(\cpu.icache.r_data[1][29] ));
 sg13g2_a22oi_1 _15717_ (.Y(_08982_),
    .B1(net816),
    .B2(\cpu.icache.r_data[4][29] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[6][29] ));
 sg13g2_nand3_1 _15718_ (.B(_08981_),
    .C(_08982_),
    .A(_08980_),
    .Y(_08983_));
 sg13g2_a21oi_1 _15719_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net627),
    .Y(_08984_),
    .B1(_08983_));
 sg13g2_nand2b_1 _15720_ (.Y(_08985_),
    .B(net627),
    .A_N(\cpu.icache.r_data[0][13] ));
 sg13g2_and2_1 _15721_ (.A(\cpu.icache.r_data[5][13] ),
    .B(net811),
    .X(_08986_));
 sg13g2_a221oi_1 _15722_ (.B2(\cpu.icache.r_data[3][13] ),
    .C1(_08986_),
    .B1(net633),
    .A1(\cpu.icache.r_data[1][13] ),
    .Y(_08987_),
    .A2(net707));
 sg13g2_a22oi_1 _15723_ (.Y(_08988_),
    .B1(net816),
    .B2(\cpu.icache.r_data[4][13] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_a22oi_1 _15724_ (.Y(_08989_),
    .B1(_08829_),
    .B2(\cpu.icache.r_data[7][13] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[6][13] ));
 sg13g2_nand4_1 _15725_ (.B(_08987_),
    .C(_08988_),
    .A(_08588_),
    .Y(_08990_),
    .D(_08989_));
 sg13g2_a21oi_1 _15726_ (.A1(_08985_),
    .A2(_08990_),
    .Y(_08991_),
    .B1(net1078));
 sg13g2_a21o_1 _15727_ (.A2(_08984_),
    .A1(net920),
    .B1(_08991_),
    .X(_08992_));
 sg13g2_buf_1 _15728_ (.A(_08992_),
    .X(_08993_));
 sg13g2_nand2_1 _15729_ (.Y(_08994_),
    .A(_08977_),
    .B(net346));
 sg13g2_nor2_1 _15730_ (.A(_08961_),
    .B(_08994_),
    .Y(_08995_));
 sg13g2_buf_2 _15731_ (.A(_08995_),
    .X(_08996_));
 sg13g2_buf_1 _15732_ (.A(_08996_),
    .X(_08997_));
 sg13g2_nand2_1 _15733_ (.Y(_08998_),
    .A(_08943_),
    .B(net173));
 sg13g2_a22oi_1 _15734_ (.Y(_08999_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][27] ),
    .A2(net550),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_mux2_1 _15735_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net815),
    .X(_09000_));
 sg13g2_a22oi_1 _15736_ (.Y(_09001_),
    .B1(net810),
    .B2(_09000_),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][27] ));
 sg13g2_buf_2 _15737_ (.A(net701),
    .X(_09002_));
 sg13g2_a22oi_1 _15738_ (.Y(_09003_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][27] ),
    .A2(net625),
    .A1(\cpu.icache.r_data[5][27] ));
 sg13g2_nand2b_1 _15739_ (.Y(_09004_),
    .B(net547),
    .A_N(_00210_));
 sg13g2_nand4_1 _15740_ (.B(_09001_),
    .C(_09003_),
    .A(_08999_),
    .Y(_09005_),
    .D(_09004_));
 sg13g2_inv_1 _15741_ (.Y(_09006_),
    .A(_08898_));
 sg13g2_nand2_1 _15742_ (.Y(_09007_),
    .A(_00209_),
    .B(net547));
 sg13g2_mux2_1 _15743_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(\cpu.icache.r_data[3][11] ),
    .S(net802),
    .X(_09008_));
 sg13g2_a22oi_1 _15744_ (.Y(_09009_),
    .B1(_09008_),
    .B2(_08597_),
    .A2(_08510_),
    .A1(\cpu.icache.r_data[4][11] ));
 sg13g2_a22oi_1 _15745_ (.Y(_09010_),
    .B1(net629),
    .B2(\cpu.icache.r_data[2][11] ),
    .A2(net630),
    .A1(\cpu.icache.r_data[1][11] ));
 sg13g2_a22oi_1 _15746_ (.Y(_09011_),
    .B1(_08925_),
    .B2(\cpu.icache.r_data[6][11] ),
    .A2(_08649_),
    .A1(\cpu.icache.r_data[5][11] ));
 sg13g2_nand4_1 _15747_ (.B(_09009_),
    .C(_09010_),
    .A(_08616_),
    .Y(_09012_),
    .D(_09011_));
 sg13g2_and3_1 _15748_ (.X(_09013_),
    .A(net1077),
    .B(_09007_),
    .C(_09012_));
 sg13g2_a21o_1 _15749_ (.A2(_09005_),
    .A1(net800),
    .B1(_09013_),
    .X(_09014_));
 sg13g2_buf_1 _15750_ (.A(_09014_),
    .X(_09015_));
 sg13g2_nor2_1 _15751_ (.A(_00208_),
    .B(net489),
    .Y(_09016_));
 sg13g2_mux2_1 _15752_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(\cpu.icache.r_data[7][26] ),
    .S(net809),
    .X(_09017_));
 sg13g2_a22oi_1 _15753_ (.Y(_09018_),
    .B1(_09017_),
    .B2(net812),
    .A2(_08856_),
    .A1(\cpu.icache.r_data[4][26] ));
 sg13g2_nor2_1 _15754_ (.A(net815),
    .B(_09018_),
    .Y(_09019_));
 sg13g2_a22oi_1 _15755_ (.Y(_09020_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][26] ),
    .A2(net550),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_buf_1 _15756_ (.A(net633),
    .X(_09021_));
 sg13g2_a22oi_1 _15757_ (.Y(_09022_),
    .B1(net546),
    .B2(\cpu.icache.r_data[3][26] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_nand2_1 _15758_ (.Y(_09023_),
    .A(_09020_),
    .B(_09022_));
 sg13g2_nor3_1 _15759_ (.A(_09016_),
    .B(_09019_),
    .C(_09023_),
    .Y(_09024_));
 sg13g2_nand2_1 _15760_ (.Y(_09025_),
    .A(_00207_),
    .B(_08931_));
 sg13g2_a22oi_1 _15761_ (.Y(_09026_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][10] ),
    .A2(net550),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_a22oi_1 _15762_ (.Y(_09027_),
    .B1(net549),
    .B2(\cpu.icache.r_data[3][10] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[1][10] ));
 sg13g2_mux2_1 _15763_ (.A0(\cpu.icache.r_data[5][10] ),
    .A1(\cpu.icache.r_data[7][10] ),
    .S(net813),
    .X(_09028_));
 sg13g2_a22oi_1 _15764_ (.Y(_09029_),
    .B1(_09028_),
    .B2(net801),
    .A2(net814),
    .A1(\cpu.icache.r_data[6][10] ));
 sg13g2_or2_1 _15765_ (.X(_09030_),
    .B(_09029_),
    .A(net815));
 sg13g2_nand4_1 _15766_ (.B(_09026_),
    .C(_09027_),
    .A(_08500_),
    .Y(_09031_),
    .D(_09030_));
 sg13g2_a21oi_1 _15767_ (.A1(_09025_),
    .A2(_09031_),
    .Y(_09032_),
    .B1(_08920_));
 sg13g2_a21oi_1 _15768_ (.A1(net800),
    .A2(_09024_),
    .Y(_09033_),
    .B1(_09032_));
 sg13g2_buf_1 _15769_ (.A(_09033_),
    .X(_09034_));
 sg13g2_inv_1 _15770_ (.Y(_09035_),
    .A(_09034_));
 sg13g2_nor4_1 _15771_ (.A(net174),
    .B(_08998_),
    .C(net345),
    .D(_09035_),
    .Y(_09036_));
 sg13g2_a21o_1 _15772_ (.A2(net143),
    .A1(net1097),
    .B1(_09036_),
    .X(_00016_));
 sg13g2_buf_1 _15773_ (.A(\cpu.dec.r_op[4] ),
    .X(_09037_));
 sg13g2_buf_1 _15774_ (.A(net1148),
    .X(_09038_));
 sg13g2_inv_1 _15775_ (.Y(_09039_),
    .A(net1076));
 sg13g2_nand4_1 _15776_ (.B(_08862_),
    .C(_08871_),
    .A(_08823_),
    .Y(_09040_),
    .D(_08881_));
 sg13g2_nand4_1 _15777_ (.B(_08890_),
    .C(_08840_),
    .A(_08836_),
    .Y(_09041_),
    .D(_08848_));
 sg13g2_nor2_1 _15778_ (.A(_09040_),
    .B(_09041_),
    .Y(_09042_));
 sg13g2_nand4_1 _15779_ (.B(_08725_),
    .C(_08698_),
    .A(_08677_),
    .Y(_09043_),
    .D(_09042_));
 sg13g2_nand2_1 _15780_ (.Y(_09044_),
    .A(_08770_),
    .B(_08792_));
 sg13g2_nor3_1 _15781_ (.A(_08626_),
    .B(_08539_),
    .C(_09044_),
    .Y(_09045_));
 sg13g2_buf_1 _15782_ (.A(_08648_),
    .X(_09046_));
 sg13g2_xor2_1 _15783_ (.B(_08656_),
    .A(net344),
    .X(_09047_));
 sg13g2_nand4_1 _15784_ (.B(_08814_),
    .C(_09047_),
    .A(_09045_),
    .Y(_09048_),
    .D(_08748_));
 sg13g2_nor3_1 _15785_ (.A(_08602_),
    .B(_09043_),
    .C(_09048_),
    .Y(_09049_));
 sg13g2_and2_1 _15786_ (.A(_08458_),
    .B(_09049_),
    .X(_09050_));
 sg13g2_buf_1 _15787_ (.A(_09050_),
    .X(_09051_));
 sg13g2_buf_1 _15788_ (.A(_09051_),
    .X(_09052_));
 sg13g2_a22oi_1 _15789_ (.Y(_09053_),
    .B1(net931),
    .B2(\cpu.icache.r_data[4][12] ),
    .A2(_08503_),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15790_ (.Y(_09054_),
    .B1(net708),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_data[1][12] ));
 sg13g2_mux2_1 _15791_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(\cpu.icache.r_data[7][12] ),
    .S(net1149),
    .X(_09055_));
 sg13g2_a22oi_1 _15792_ (.Y(_09056_),
    .B1(_09055_),
    .B2(net1085),
    .A2(_08527_),
    .A1(\cpu.icache.r_data[6][12] ));
 sg13g2_or2_1 _15793_ (.X(_09057_),
    .B(_09056_),
    .A(net1086));
 sg13g2_and4_1 _15794_ (.A(_08497_),
    .B(_09053_),
    .C(_09054_),
    .D(_09057_),
    .X(_09058_));
 sg13g2_a21oi_1 _15795_ (.A1(_00215_),
    .A2(_08909_),
    .Y(_09059_),
    .B1(_09058_));
 sg13g2_nor2_1 _15796_ (.A(_00216_),
    .B(_08497_),
    .Y(_09060_));
 sg13g2_mux2_1 _15797_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(\cpu.icache.r_data[7][28] ),
    .S(net1084),
    .X(_09061_));
 sg13g2_a22oi_1 _15798_ (.Y(_09062_),
    .B1(_09061_),
    .B2(_08526_),
    .A2(_08856_),
    .A1(\cpu.icache.r_data[4][28] ));
 sg13g2_nor2_1 _15799_ (.A(net924),
    .B(_09062_),
    .Y(_09063_));
 sg13g2_a22oi_1 _15800_ (.Y(_09064_),
    .B1(_08592_),
    .B2(\cpu.icache.r_data[6][28] ),
    .A2(_08503_),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_a22oi_1 _15801_ (.Y(_09065_),
    .B1(net708),
    .B2(\cpu.icache.r_data[3][28] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_data[1][28] ));
 sg13g2_nand2_1 _15802_ (.Y(_09066_),
    .A(_09064_),
    .B(_09065_));
 sg13g2_or4_1 _15803_ (.A(net1077),
    .B(_09060_),
    .C(_09063_),
    .D(_09066_),
    .X(_09067_));
 sg13g2_o21ai_1 _15804_ (.B1(_09067_),
    .Y(_09068_),
    .A1(_08898_),
    .A2(_09059_));
 sg13g2_buf_1 _15805_ (.A(_09068_),
    .X(_09069_));
 sg13g2_inv_1 _15806_ (.Y(_09070_),
    .A(net390));
 sg13g2_buf_1 _15807_ (.A(_09070_),
    .X(_09071_));
 sg13g2_nor2_1 _15808_ (.A(_00214_),
    .B(_08497_),
    .Y(_09072_));
 sg13g2_mux2_1 _15809_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(net1086),
    .X(_09073_));
 sg13g2_a22oi_1 _15810_ (.Y(_09074_),
    .B1(_09073_),
    .B2(net813),
    .A2(_08875_),
    .A1(\cpu.icache.r_data[5][22] ));
 sg13g2_nor2_1 _15811_ (.A(net926),
    .B(_09074_),
    .Y(_09075_));
 sg13g2_a22oi_1 _15812_ (.Y(_09076_),
    .B1(net706),
    .B2(\cpu.icache.r_data[6][22] ),
    .A2(net697),
    .A1(\cpu.icache.r_data[1][22] ));
 sg13g2_a22oi_1 _15813_ (.Y(_09077_),
    .B1(net931),
    .B2(\cpu.icache.r_data[4][22] ),
    .A2(_08504_),
    .A1(\cpu.icache.r_data[2][22] ));
 sg13g2_nand2_1 _15814_ (.Y(_09078_),
    .A(_09076_),
    .B(_09077_));
 sg13g2_nor3_1 _15815_ (.A(_09072_),
    .B(_09075_),
    .C(_09078_),
    .Y(_09079_));
 sg13g2_nand2_1 _15816_ (.Y(_09080_),
    .A(_00213_),
    .B(_08909_));
 sg13g2_a22oi_1 _15817_ (.Y(_09081_),
    .B1(_08508_),
    .B2(\cpu.icache.r_data[4][6] ),
    .A2(_08503_),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_a22oi_1 _15818_ (.Y(_09082_),
    .B1(net708),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_mux2_1 _15819_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(\cpu.icache.r_data[7][6] ),
    .S(_08529_),
    .X(_09083_));
 sg13g2_a22oi_1 _15820_ (.Y(_09084_),
    .B1(_09083_),
    .B2(net1085),
    .A2(net814),
    .A1(\cpu.icache.r_data[6][6] ));
 sg13g2_or2_1 _15821_ (.X(_09085_),
    .B(_09084_),
    .A(_08524_));
 sg13g2_nand4_1 _15822_ (.B(_09081_),
    .C(_09082_),
    .A(_08498_),
    .Y(_09086_),
    .D(_09085_));
 sg13g2_a21oi_1 _15823_ (.A1(_09080_),
    .A2(_09086_),
    .Y(_09087_),
    .B1(net1078));
 sg13g2_a21oi_1 _15824_ (.A1(net1078),
    .A2(_09079_),
    .Y(_09088_),
    .B1(_09087_));
 sg13g2_buf_2 _15825_ (.A(_09088_),
    .X(_09089_));
 sg13g2_nor2_1 _15826_ (.A(_00212_),
    .B(_08498_),
    .Y(_09090_));
 sg13g2_mux2_1 _15827_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(net924),
    .X(_09091_));
 sg13g2_a22oi_1 _15828_ (.Y(_09092_),
    .B1(_09091_),
    .B2(_08617_),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][21] ));
 sg13g2_nor2_1 _15829_ (.A(net926),
    .B(_09092_),
    .Y(_09093_));
 sg13g2_a22oi_1 _15830_ (.Y(_09094_),
    .B1(net699),
    .B2(\cpu.icache.r_data[6][21] ),
    .A2(_08819_),
    .A1(\cpu.icache.r_data[1][21] ));
 sg13g2_a22oi_1 _15831_ (.Y(_09095_),
    .B1(net816),
    .B2(\cpu.icache.r_data[4][21] ),
    .A2(net705),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_nand2_1 _15832_ (.Y(_09096_),
    .A(_09094_),
    .B(_09095_));
 sg13g2_nor3_1 _15833_ (.A(_09090_),
    .B(_09093_),
    .C(_09096_),
    .Y(_09097_));
 sg13g2_nand2_1 _15834_ (.Y(_09098_),
    .A(_00211_),
    .B(_08909_));
 sg13g2_a22oi_1 _15835_ (.Y(_09099_),
    .B1(net705),
    .B2(\cpu.icache.r_data[2][5] ),
    .A2(_08819_),
    .A1(\cpu.icache.r_data[1][5] ));
 sg13g2_nand2_1 _15836_ (.Y(_09100_),
    .A(\cpu.icache.r_data[6][5] ),
    .B(_08593_));
 sg13g2_a22oi_1 _15837_ (.Y(_09101_),
    .B1(_08830_),
    .B2(\cpu.icache.r_data[3][5] ),
    .A2(_08558_),
    .A1(\cpu.icache.r_data[5][5] ));
 sg13g2_nor2_1 _15838_ (.A(net926),
    .B(_09101_),
    .Y(_09102_));
 sg13g2_a221oi_1 _15839_ (.B2(\cpu.icache.r_data[7][5] ),
    .C1(_09102_),
    .B1(_08829_),
    .A1(\cpu.icache.r_data[4][5] ),
    .Y(_09103_),
    .A2(_08508_));
 sg13g2_nand4_1 _15840_ (.B(_09099_),
    .C(_09100_),
    .A(_08557_),
    .Y(_09104_),
    .D(_09103_));
 sg13g2_a21oi_1 _15841_ (.A1(_09098_),
    .A2(_09104_),
    .Y(_09105_),
    .B1(net1078));
 sg13g2_a21oi_1 _15842_ (.A1(net1078),
    .A2(_09097_),
    .Y(_09106_),
    .B1(_09105_));
 sg13g2_buf_1 _15843_ (.A(_09106_),
    .X(_09107_));
 sg13g2_nor2_1 _15844_ (.A(_09089_),
    .B(_09107_),
    .Y(_09108_));
 sg13g2_buf_1 _15845_ (.A(_09108_),
    .X(_09109_));
 sg13g2_inv_1 _15846_ (.Y(_09110_),
    .A(net347));
 sg13g2_buf_1 _15847_ (.A(_09110_),
    .X(_09111_));
 sg13g2_nor2_1 _15848_ (.A(net231),
    .B(_08941_),
    .Y(_09112_));
 sg13g2_buf_1 _15849_ (.A(_09112_),
    .X(_09113_));
 sg13g2_nand2_1 _15850_ (.Y(_09114_),
    .A(_08996_),
    .B(net194));
 sg13g2_nand2_1 _15851_ (.Y(_09115_),
    .A(net345),
    .B(_09034_));
 sg13g2_buf_1 _15852_ (.A(_09115_),
    .X(_09116_));
 sg13g2_nor2_1 _15853_ (.A(_09114_),
    .B(_09116_),
    .Y(_09117_));
 sg13g2_buf_2 _15854_ (.A(_09117_),
    .X(_09118_));
 sg13g2_nand4_1 _15855_ (.B(net274),
    .C(_09109_),
    .A(net142),
    .Y(_09119_),
    .D(_09118_));
 sg13g2_o21ai_1 _15856_ (.B1(_09119_),
    .Y(_00015_),
    .A1(_09039_),
    .A2(net108));
 sg13g2_buf_1 _15857_ (.A(net174),
    .X(_09120_));
 sg13g2_buf_1 _15858_ (.A(_09120_),
    .X(_09121_));
 sg13g2_buf_1 _15859_ (.A(net800),
    .X(_09122_));
 sg13g2_a21o_1 _15860_ (.A2(_09097_),
    .A1(net696),
    .B1(_09105_),
    .X(_09123_));
 sg13g2_buf_1 _15861_ (.A(_09123_),
    .X(_09124_));
 sg13g2_buf_1 _15862_ (.A(net390),
    .X(_09125_));
 sg13g2_nand2_1 _15863_ (.Y(_09126_),
    .A(_09125_),
    .B(_09089_));
 sg13g2_buf_1 _15864_ (.A(_09034_),
    .X(_09127_));
 sg13g2_o21ai_1 _15865_ (.B1(net230),
    .Y(_09128_),
    .A1(net389),
    .A2(_09126_));
 sg13g2_nand4_1 _15866_ (.B(net173),
    .C(net345),
    .A(_08943_),
    .Y(_09129_),
    .D(_09128_));
 sg13g2_buf_1 _15867_ (.A(\cpu.dec.r_op[2] ),
    .X(_09130_));
 sg13g2_buf_1 _15868_ (.A(net1147),
    .X(_09131_));
 sg13g2_buf_1 _15869_ (.A(net174),
    .X(_09132_));
 sg13g2_nand2_1 _15870_ (.Y(_09133_),
    .A(net1075),
    .B(net140));
 sg13g2_o21ai_1 _15871_ (.B1(_09133_),
    .Y(_00013_),
    .A1(net107),
    .A2(_09129_));
 sg13g2_nor3_1 _15872_ (.A(net274),
    .B(_09089_),
    .C(net389),
    .Y(_09134_));
 sg13g2_nor2_1 _15873_ (.A(_08998_),
    .B(_09116_),
    .Y(_09135_));
 sg13g2_inv_1 _15874_ (.Y(_09136_),
    .A(_09118_));
 sg13g2_inv_2 _15875_ (.Y(_09137_),
    .A(_09089_));
 sg13g2_nand3_1 _15876_ (.B(_09137_),
    .C(_09107_),
    .A(net274),
    .Y(_09138_));
 sg13g2_buf_1 _15877_ (.A(_09138_),
    .X(_09139_));
 sg13g2_nor2_1 _15878_ (.A(_00222_),
    .B(net548),
    .Y(_09140_));
 sg13g2_mux2_1 _15879_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(net802),
    .X(_09141_));
 sg13g2_a22oi_1 _15880_ (.Y(_09142_),
    .B1(_09141_),
    .B2(_08810_),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][20] ));
 sg13g2_nor2_1 _15881_ (.A(_08565_),
    .B(_09142_),
    .Y(_09143_));
 sg13g2_a22oi_1 _15882_ (.Y(_09144_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][20] ),
    .A2(net630),
    .A1(\cpu.icache.r_data[1][20] ));
 sg13g2_a22oi_1 _15883_ (.Y(_09145_),
    .B1(net710),
    .B2(\cpu.icache.r_data[4][20] ),
    .A2(_08739_),
    .A1(\cpu.icache.r_data[2][20] ));
 sg13g2_nand2_1 _15884_ (.Y(_09146_),
    .A(_09144_),
    .B(_09145_));
 sg13g2_nor3_1 _15885_ (.A(_09140_),
    .B(_09143_),
    .C(_09146_),
    .Y(_09147_));
 sg13g2_nand2_1 _15886_ (.Y(_09148_),
    .A(_00221_),
    .B(net547));
 sg13g2_a22oi_1 _15887_ (.Y(_09149_),
    .B1(net628),
    .B2(\cpu.icache.r_data[6][4] ),
    .A2(net629),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_a22oi_1 _15888_ (.Y(_09150_),
    .B1(net710),
    .B2(\cpu.icache.r_data[4][4] ),
    .A2(net630),
    .A1(\cpu.icache.r_data[1][4] ));
 sg13g2_mux2_1 _15889_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_08524_),
    .X(_09151_));
 sg13g2_a22oi_1 _15890_ (.Y(_09152_),
    .B1(_09151_),
    .B2(net809),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][4] ));
 sg13g2_nand2b_1 _15891_ (.Y(_09153_),
    .B(net812),
    .A_N(_09152_));
 sg13g2_nand4_1 _15892_ (.B(_09149_),
    .C(_09150_),
    .A(net548),
    .Y(_09154_),
    .D(_09153_));
 sg13g2_a21oi_1 _15893_ (.A1(_09148_),
    .A2(_09154_),
    .Y(_09155_),
    .B1(net920));
 sg13g2_a21oi_1 _15894_ (.A1(net696),
    .A2(_09147_),
    .Y(_09156_),
    .B1(_09155_));
 sg13g2_buf_1 _15895_ (.A(_09156_),
    .X(_09157_));
 sg13g2_buf_1 _15896_ (.A(_09157_),
    .X(_09158_));
 sg13g2_nor2_1 _15897_ (.A(_00220_),
    .B(_08557_),
    .Y(_09159_));
 sg13g2_mux2_1 _15898_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(\cpu.icache.r_data[7][19] ),
    .S(_08530_),
    .X(_09160_));
 sg13g2_a22oi_1 _15899_ (.Y(_09161_),
    .B1(_09160_),
    .B2(_08743_),
    .A2(_08856_),
    .A1(\cpu.icache.r_data[4][19] ));
 sg13g2_nor2_1 _15900_ (.A(_08719_),
    .B(_09161_),
    .Y(_09162_));
 sg13g2_a22oi_1 _15901_ (.Y(_09163_),
    .B1(net699),
    .B2(\cpu.icache.r_data[6][19] ),
    .A2(net705),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_a22oi_1 _15902_ (.Y(_09164_),
    .B1(_08521_),
    .B2(\cpu.icache.r_data[3][19] ),
    .A2(net707),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_nand2_1 _15903_ (.Y(_09165_),
    .A(_09163_),
    .B(_09164_));
 sg13g2_nor3_1 _15904_ (.A(_09159_),
    .B(_09162_),
    .C(_09165_),
    .Y(_09166_));
 sg13g2_nand2_1 _15905_ (.Y(_09167_),
    .A(_00219_),
    .B(net627));
 sg13g2_mux2_1 _15906_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_08595_),
    .X(_09168_));
 sg13g2_a22oi_1 _15907_ (.Y(_09169_),
    .B1(_09168_),
    .B2(_08597_),
    .A2(net816),
    .A1(\cpu.icache.r_data[4][3] ));
 sg13g2_a22oi_1 _15908_ (.Y(_09170_),
    .B1(_08620_),
    .B2(\cpu.icache.r_data[2][3] ),
    .A2(_08561_),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_a22oi_1 _15909_ (.Y(_09171_),
    .B1(_08766_),
    .B2(\cpu.icache.r_data[6][3] ),
    .A2(_08649_),
    .A1(\cpu.icache.r_data[5][3] ));
 sg13g2_nand4_1 _15910_ (.B(_09169_),
    .C(_09170_),
    .A(net631),
    .Y(_09172_),
    .D(_09171_));
 sg13g2_a21oi_1 _15911_ (.A1(_09167_),
    .A2(_09172_),
    .Y(_09173_),
    .B1(_08899_));
 sg13g2_a21oi_1 _15912_ (.A1(net920),
    .A2(_09166_),
    .Y(_09174_),
    .B1(_09173_));
 sg13g2_buf_1 _15913_ (.A(_09174_),
    .X(_09175_));
 sg13g2_nand2b_1 _15914_ (.Y(_09176_),
    .B(net627),
    .A_N(_00218_));
 sg13g2_mux2_1 _15915_ (.A0(\cpu.icache.r_data[5][18] ),
    .A1(\cpu.icache.r_data[7][18] ),
    .S(_08531_),
    .X(_09177_));
 sg13g2_a22oi_1 _15916_ (.Y(_09178_),
    .B1(_09177_),
    .B2(_08743_),
    .A2(_08856_),
    .A1(\cpu.icache.r_data[4][18] ));
 sg13g2_or2_1 _15917_ (.X(_09179_),
    .B(_09178_),
    .A(_08525_));
 sg13g2_a22oi_1 _15918_ (.Y(_09180_),
    .B1(_08522_),
    .B2(\cpu.icache.r_data[3][18] ),
    .A2(net629),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_a22oi_1 _15919_ (.Y(_09181_),
    .B1(_08766_),
    .B2(\cpu.icache.r_data[6][18] ),
    .A2(_08716_),
    .A1(\cpu.icache.r_data[1][18] ));
 sg13g2_nand4_1 _15920_ (.B(_09179_),
    .C(_09180_),
    .A(_09176_),
    .Y(_09182_),
    .D(_09181_));
 sg13g2_nand2_1 _15921_ (.Y(_09183_),
    .A(\cpu.icache.r_data[1][2] ),
    .B(_08561_));
 sg13g2_a22oi_1 _15922_ (.Y(_09184_),
    .B1(_08520_),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(_08560_),
    .A1(\cpu.icache.r_data[5][2] ));
 sg13g2_a22oi_1 _15923_ (.Y(_09185_),
    .B1(_08509_),
    .B2(\cpu.icache.r_data[4][2] ),
    .A2(_08620_),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_a22oi_1 _15924_ (.Y(_09186_),
    .B1(_08829_),
    .B2(\cpu.icache.r_data[7][2] ),
    .A2(_08593_),
    .A1(\cpu.icache.r_data[6][2] ));
 sg13g2_nand4_1 _15925_ (.B(_09184_),
    .C(_09185_),
    .A(_09183_),
    .Y(_09187_),
    .D(_09186_));
 sg13g2_nor2_1 _15926_ (.A(_08930_),
    .B(_09187_),
    .Y(_09188_));
 sg13g2_a21oi_1 _15927_ (.A1(_00217_),
    .A2(_08931_),
    .Y(_09189_),
    .B1(_09188_));
 sg13g2_mux2_1 _15928_ (.A0(_09182_),
    .A1(_09189_),
    .S(net1077),
    .X(_09190_));
 sg13g2_buf_2 _15929_ (.A(_09190_),
    .X(_09191_));
 sg13g2_nand2_1 _15930_ (.Y(_09192_),
    .A(net342),
    .B(_09191_));
 sg13g2_nor4_1 _15931_ (.A(_09136_),
    .B(_09139_),
    .C(net273),
    .D(_09192_),
    .Y(_09193_));
 sg13g2_a21oi_1 _15932_ (.A1(_09134_),
    .A2(_09135_),
    .Y(_09194_),
    .B1(_09193_));
 sg13g2_buf_2 _15933_ (.A(\cpu.dec.r_op[3] ),
    .X(_09195_));
 sg13g2_buf_1 _15934_ (.A(_09195_),
    .X(_09196_));
 sg13g2_nand2_1 _15935_ (.Y(_09197_),
    .A(net1074),
    .B(net140));
 sg13g2_o21ai_1 _15936_ (.B1(_09197_),
    .Y(_00014_),
    .A1(net107),
    .A2(_09194_));
 sg13g2_nor2_1 _15937_ (.A(net342),
    .B(_09191_),
    .Y(_09198_));
 sg13g2_nor2b_1 _15938_ (.A(_09139_),
    .B_N(_09198_),
    .Y(_09199_));
 sg13g2_and2_1 _15939_ (.A(net273),
    .B(_09199_),
    .X(_09200_));
 sg13g2_a22oi_1 _15940_ (.Y(_09201_),
    .B1(_09200_),
    .B2(_09118_),
    .A2(_09135_),
    .A1(_09109_));
 sg13g2_buf_2 _15941_ (.A(\cpu.dec.r_op[6] ),
    .X(_09202_));
 sg13g2_buf_1 _15942_ (.A(_09202_),
    .X(_09203_));
 sg13g2_nand2_1 _15943_ (.Y(_09204_),
    .A(net1073),
    .B(net140));
 sg13g2_o21ai_1 _15944_ (.B1(_09204_),
    .Y(_00017_),
    .A1(net107),
    .A2(_09201_));
 sg13g2_buf_1 _15945_ (.A(\cpu.spi.r_count[7] ),
    .X(_09205_));
 sg13g2_buf_1 _15946_ (.A(\cpu.spi.r_count[3] ),
    .X(_09206_));
 sg13g2_buf_1 _15947_ (.A(\cpu.spi.r_count[0] ),
    .X(_09207_));
 sg13g2_buf_1 _15948_ (.A(\cpu.spi.r_count[1] ),
    .X(_09208_));
 sg13g2_nor2_1 _15949_ (.A(_09207_),
    .B(_09208_),
    .Y(_09209_));
 sg13g2_nand2b_1 _15950_ (.Y(_09210_),
    .B(_09209_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _15951_ (.A(_09206_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09210_),
    .Y(_09211_));
 sg13g2_nor2b_1 _15952_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09211_),
    .Y(_09212_));
 sg13g2_nor2b_1 _15953_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09212_),
    .Y(_09213_));
 sg13g2_buf_1 _15954_ (.A(_09213_),
    .X(_09214_));
 sg13g2_nand2b_1 _15955_ (.Y(_09215_),
    .B(_09214_),
    .A_N(_09205_));
 sg13g2_buf_1 _15956_ (.A(_09215_),
    .X(_09216_));
 sg13g2_buf_1 _15957_ (.A(_09216_),
    .X(_09217_));
 sg13g2_buf_1 _15958_ (.A(\cpu.addr[3] ),
    .X(_09218_));
 sg13g2_buf_8 _15959_ (.A(net1146),
    .X(_09219_));
 sg13g2_buf_1 _15960_ (.A(_09219_),
    .X(_09220_));
 sg13g2_buf_1 _15961_ (.A(net919),
    .X(_09221_));
 sg13g2_buf_1 _15962_ (.A(_09221_),
    .X(_09222_));
 sg13g2_buf_1 _15963_ (.A(net695),
    .X(_09223_));
 sg13g2_buf_1 _15964_ (.A(\cpu.addr[6] ),
    .X(_09224_));
 sg13g2_buf_1 _15965_ (.A(_09224_),
    .X(_09225_));
 sg13g2_buf_1 _15966_ (.A(\cpu.addr[8] ),
    .X(_09226_));
 sg13g2_buf_1 _15967_ (.A(_09226_),
    .X(_09227_));
 sg13g2_buf_1 _15968_ (.A(\cpu.addr[7] ),
    .X(_09228_));
 sg13g2_buf_1 _15969_ (.A(_09228_),
    .X(_09229_));
 sg13g2_nor2b_1 _15970_ (.A(net1070),
    .B_N(net1069),
    .Y(_09230_));
 sg13g2_buf_1 _15971_ (.A(_09230_),
    .X(_09231_));
 sg13g2_nand2_2 _15972_ (.Y(_09232_),
    .A(net1071),
    .B(_09231_));
 sg13g2_buf_2 _15973_ (.A(\cpu.addr[2] ),
    .X(_09233_));
 sg13g2_buf_1 _15974_ (.A(_09233_),
    .X(_09234_));
 sg13g2_buf_1 _15975_ (.A(net1068),
    .X(_09235_));
 sg13g2_buf_2 _15976_ (.A(net918),
    .X(_09236_));
 sg13g2_buf_1 _15977_ (.A(net798),
    .X(_09237_));
 sg13g2_buf_2 _15978_ (.A(\cpu.addr[1] ),
    .X(_09238_));
 sg13g2_buf_1 _15979_ (.A(_09238_),
    .X(_09239_));
 sg13g2_nor2_2 _15980_ (.A(net694),
    .B(net1067),
    .Y(_09240_));
 sg13g2_buf_1 _15981_ (.A(\cpu.dec.r_trap ),
    .X(_09241_));
 sg13g2_buf_1 _15982_ (.A(\cpu.ex.r_ie ),
    .X(_09242_));
 sg13g2_inv_2 _15983_ (.Y(_09243_),
    .A(_09242_));
 sg13g2_buf_1 _15984_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09244_));
 sg13g2_buf_2 _15985_ (.A(ui_in[3]),
    .X(_09245_));
 sg13g2_buf_2 _15986_ (.A(ui_in[6]),
    .X(_09246_));
 sg13g2_a22oi_1 _15987_ (.Y(_09247_),
    .B1(\cpu.gpio.r_enable_in[6] ),
    .B2(_09246_),
    .A2(_09245_),
    .A1(\cpu.gpio.r_enable_in[3] ));
 sg13g2_buf_8 _15988_ (.A(ui_in[5]),
    .X(_09248_));
 sg13g2_buf_1 _15989_ (.A(uio_in[6]),
    .X(_09249_));
 sg13g2_a22oi_1 _15990_ (.Y(_09250_),
    .B1(\cpu.gpio.r_enable_io[6] ),
    .B2(_09249_),
    .A2(_09248_),
    .A1(\cpu.gpio.r_enable_in[5] ));
 sg13g2_buf_1 _15991_ (.A(\cpu.gpio.r_enable_in[7] ),
    .X(_09251_));
 sg13g2_buf_8 _15992_ (.A(ui_in[7]),
    .X(_09252_));
 sg13g2_buf_1 _15993_ (.A(uio_in[4]),
    .X(_09253_));
 sg13g2_a22oi_1 _15994_ (.Y(_09254_),
    .B1(\cpu.gpio.r_enable_io[4] ),
    .B2(_09253_),
    .A2(_09252_),
    .A1(_09251_));
 sg13g2_buf_8 _15995_ (.A(ui_in[0]),
    .X(_09255_));
 sg13g2_buf_1 _15996_ (.A(\cpu.gpio.r_enable_io[7] ),
    .X(_09256_));
 sg13g2_buf_2 _15997_ (.A(uio_in[7]),
    .X(_09257_));
 sg13g2_a22oi_1 _15998_ (.Y(_09258_),
    .B1(_09256_),
    .B2(_09257_),
    .A2(_09255_),
    .A1(\cpu.gpio.r_enable_in[0] ));
 sg13g2_nand4_1 _15999_ (.B(_09250_),
    .C(_09254_),
    .A(_09247_),
    .Y(_09259_),
    .D(_09258_));
 sg13g2_buf_2 _16000_ (.A(ui_in[2]),
    .X(_09260_));
 sg13g2_buf_1 _16001_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_09261_));
 sg13g2_buf_1 _16002_ (.A(ui_in[4]),
    .X(_09262_));
 sg13g2_a22oi_1 _16003_ (.Y(_09263_),
    .B1(_09261_),
    .B2(_09262_),
    .A2(_09260_),
    .A1(\cpu.gpio.r_enable_in[2] ));
 sg13g2_buf_2 _16004_ (.A(ui_in[1]),
    .X(_09264_));
 sg13g2_buf_1 _16005_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09265_));
 sg13g2_buf_1 _16006_ (.A(uio_in[5]),
    .X(_09266_));
 sg13g2_a22oi_1 _16007_ (.Y(_09267_),
    .B1(_09265_),
    .B2(_09266_),
    .A2(_09264_),
    .A1(\cpu.gpio.r_enable_in[1] ));
 sg13g2_nand2_1 _16008_ (.Y(_09268_),
    .A(_09263_),
    .B(_09267_));
 sg13g2_or2_1 _16009_ (.X(_09269_),
    .B(_09268_),
    .A(_09259_));
 sg13g2_buf_1 _16010_ (.A(\cpu.intr.r_timer ),
    .X(_09270_));
 sg13g2_buf_1 _16011_ (.A(\cpu.intr.r_enable[2] ),
    .X(_09271_));
 sg13g2_buf_1 _16012_ (.A(\cpu.intr.r_swi ),
    .X(_09272_));
 sg13g2_a22oi_1 _16013_ (.Y(_09273_),
    .B1(\cpu.intr.r_enable[3] ),
    .B2(_09272_),
    .A2(_09271_),
    .A1(_09270_));
 sg13g2_buf_1 _16014_ (.A(\cpu.intr.r_clock ),
    .X(_09274_));
 sg13g2_buf_1 _16015_ (.A(\cpu.intr.spi_intr ),
    .X(_09275_));
 sg13g2_buf_1 _16016_ (.A(\cpu.intr.r_enable[5] ),
    .X(_09276_));
 sg13g2_a22oi_1 _16017_ (.Y(_09277_),
    .B1(_09275_),
    .B2(_09276_),
    .A2(\cpu.intr.r_enable[1] ),
    .A1(_09274_));
 sg13g2_buf_2 _16018_ (.A(\cpu.uart.r_x_int ),
    .X(_09278_));
 sg13g2_buf_1 _16019_ (.A(\cpu.uart.r_r_int ),
    .X(_09279_));
 sg13g2_buf_1 _16020_ (.A(\cpu.intr.r_enable[0] ),
    .X(_09280_));
 sg13g2_o21ai_1 _16021_ (.B1(_09280_),
    .Y(_09281_),
    .A1(_09278_),
    .A2(_09279_));
 sg13g2_nand3_1 _16022_ (.B(_09277_),
    .C(_09281_),
    .A(_09273_),
    .Y(_09282_));
 sg13g2_a21oi_1 _16023_ (.A1(_09244_),
    .A2(_09269_),
    .Y(_09283_),
    .B1(_09282_));
 sg13g2_nor2_2 _16024_ (.A(_09243_),
    .B(_09283_),
    .Y(_09284_));
 sg13g2_and2_1 _16025_ (.A(_08364_),
    .B(_09284_),
    .X(_09285_));
 sg13g2_nor4_2 _16026_ (.A(_09241_),
    .B(_08360_),
    .C(_08454_),
    .Y(_09286_),
    .D(_09285_));
 sg13g2_nand3_1 _16027_ (.B(_09240_),
    .C(_09286_),
    .A(_08399_),
    .Y(_09287_));
 sg13g2_nor4_2 _16028_ (.A(net624),
    .B(_08408_),
    .C(_09232_),
    .Y(_09288_),
    .D(_09287_));
 sg13g2_buf_1 _16029_ (.A(\cpu.spi.r_state[1] ),
    .X(_09289_));
 sg13g2_inv_1 _16030_ (.Y(_09290_),
    .A(net1145));
 sg13g2_nand3b_1 _16031_ (.B(_09286_),
    .C(_08350_),
    .Y(_09291_),
    .A_N(_08354_));
 sg13g2_buf_2 _16032_ (.A(_09291_),
    .X(_09292_));
 sg13g2_or2_1 _16033_ (.X(_09293_),
    .B(_09292_),
    .A(_09232_));
 sg13g2_buf_2 _16034_ (.A(_09293_),
    .X(_09294_));
 sg13g2_nor2_1 _16035_ (.A(net695),
    .B(_09294_),
    .Y(_09295_));
 sg13g2_buf_2 _16036_ (.A(_09295_),
    .X(_09296_));
 sg13g2_nor2_1 _16037_ (.A(_09290_),
    .B(_09296_),
    .Y(_09297_));
 sg13g2_buf_1 _16038_ (.A(\cpu.spi.r_state[3] ),
    .X(_09298_));
 sg13g2_a21oi_1 _16039_ (.A1(_09288_),
    .A2(_09297_),
    .Y(_09299_),
    .B1(_09298_));
 sg13g2_buf_1 _16040_ (.A(\cpu.spi.r_state[0] ),
    .X(_09300_));
 sg13g2_nand2_1 _16041_ (.Y(_09301_),
    .A(_09240_),
    .B(_09296_));
 sg13g2_nand2b_1 _16042_ (.Y(_09302_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _16043_ (.A(_09302_),
    .X(_09303_));
 sg13g2_buf_1 _16044_ (.A(_09303_),
    .X(_09304_));
 sg13g2_a21oi_1 _16045_ (.A1(net1144),
    .A2(_09301_),
    .Y(_09305_),
    .B1(net917));
 sg13g2_o21ai_1 _16046_ (.B1(_09305_),
    .Y(_00029_),
    .A1(net388),
    .A2(_09299_));
 sg13g2_nor2b_1 _16047_ (.A(r_reset),
    .B_N(net1),
    .Y(_09306_));
 sg13g2_buf_1 _16048_ (.A(_09306_),
    .X(_09307_));
 sg13g2_buf_1 _16049_ (.A(net1066),
    .X(_09308_));
 sg13g2_buf_1 _16050_ (.A(net916),
    .X(_09309_));
 sg13g2_buf_1 _16051_ (.A(_09309_),
    .X(_09310_));
 sg13g2_buf_1 _16052_ (.A(net1145),
    .X(_09311_));
 sg13g2_inv_1 _16053_ (.Y(_09312_),
    .A(_09218_));
 sg13g2_buf_1 _16054_ (.A(_09312_),
    .X(_09313_));
 sg13g2_buf_1 _16055_ (.A(net915),
    .X(_09314_));
 sg13g2_nand2b_1 _16056_ (.Y(_09315_),
    .B(net796),
    .A_N(_09294_));
 sg13g2_nand2_1 _16057_ (.Y(_09316_),
    .A(_09311_),
    .B(_09315_));
 sg13g2_buf_1 _16058_ (.A(\cpu.spi.r_state[6] ),
    .X(_09317_));
 sg13g2_buf_1 _16059_ (.A(_09317_),
    .X(_09318_));
 sg13g2_nor2b_1 _16060_ (.A(_09205_),
    .B_N(_09214_),
    .Y(_09319_));
 sg13g2_buf_2 _16061_ (.A(_09319_),
    .X(_09320_));
 sg13g2_buf_1 _16062_ (.A(_09320_),
    .X(_09321_));
 sg13g2_buf_1 _16063_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09322_));
 sg13g2_buf_1 _16064_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09323_));
 sg13g2_nor3_1 _16065_ (.A(_09322_),
    .B(_09323_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09324_));
 sg13g2_buf_1 _16066_ (.A(\cpu.spi.r_timeout_count[7] ),
    .X(_09325_));
 sg13g2_buf_1 _16067_ (.A(\cpu.spi.r_timeout_count[0] ),
    .X(_09326_));
 sg13g2_buf_1 _16068_ (.A(\cpu.spi.r_timeout_count[1] ),
    .X(_09327_));
 sg13g2_or3_1 _16069_ (.A(_09326_),
    .B(_09327_),
    .C(\cpu.spi.r_timeout_count[2] ),
    .X(_09328_));
 sg13g2_buf_1 _16070_ (.A(_09328_),
    .X(_09329_));
 sg13g2_or2_1 _16071_ (.X(_09330_),
    .B(_09329_),
    .A(\cpu.spi.r_timeout_count[3] ));
 sg13g2_buf_1 _16072_ (.A(_09330_),
    .X(_09331_));
 sg13g2_or2_1 _16073_ (.X(_09332_),
    .B(_09331_),
    .A(\cpu.spi.r_timeout_count[4] ));
 sg13g2_buf_1 _16074_ (.A(_09332_),
    .X(_09333_));
 sg13g2_or2_1 _16075_ (.X(_09334_),
    .B(_09333_),
    .A(\cpu.spi.r_timeout_count[5] ));
 sg13g2_buf_1 _16076_ (.A(_09334_),
    .X(_09335_));
 sg13g2_or2_1 _16077_ (.X(_09336_),
    .B(_09335_),
    .A(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _16078_ (.A(_09336_),
    .X(_09337_));
 sg13g2_o21ai_1 _16079_ (.B1(\cpu.spi.r_searching ),
    .Y(_09338_),
    .A1(_09325_),
    .A2(_09337_));
 sg13g2_nand2_1 _16080_ (.Y(_09339_),
    .A(_09324_),
    .B(_09338_));
 sg13g2_buf_1 _16081_ (.A(\cpu.spi.r_in[3] ),
    .X(_09340_));
 sg13g2_buf_1 _16082_ (.A(\cpu.spi.r_in[6] ),
    .X(_09341_));
 sg13g2_buf_1 _16083_ (.A(\cpu.spi.r_in[1] ),
    .X(_09342_));
 sg13g2_buf_1 _16084_ (.A(\cpu.spi.r_in[0] ),
    .X(_09343_));
 sg13g2_nand2_1 _16085_ (.Y(_09344_),
    .A(_09342_),
    .B(_09343_));
 sg13g2_nand3_1 _16086_ (.B(_09341_),
    .C(_09344_),
    .A(_09340_),
    .Y(_09345_));
 sg13g2_buf_1 _16087_ (.A(\cpu.spi.r_in[2] ),
    .X(_09346_));
 sg13g2_buf_1 _16088_ (.A(\cpu.spi.r_in[5] ),
    .X(_09347_));
 sg13g2_buf_1 _16089_ (.A(\cpu.spi.r_in[4] ),
    .X(_09348_));
 sg13g2_nand4_1 _16090_ (.B(_09347_),
    .C(_09348_),
    .A(_09346_),
    .Y(_09349_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _16091_ (.A(_09345_),
    .B(_09349_),
    .Y(_09350_));
 sg13g2_o21ai_1 _16092_ (.B1(\cpu.spi.r_searching ),
    .Y(_09351_),
    .A1(_00224_),
    .A2(_09350_));
 sg13g2_nand2_1 _16093_ (.Y(_09352_),
    .A(_09339_),
    .B(_09351_));
 sg13g2_nand3_1 _16094_ (.B(_09321_),
    .C(_09352_),
    .A(net1064),
    .Y(_09353_));
 sg13g2_o21ai_1 _16095_ (.B1(_09353_),
    .Y(_09354_),
    .A1(_09288_),
    .A2(_09316_));
 sg13g2_and2_1 _16096_ (.A(net693),
    .B(_09354_),
    .X(_00030_));
 sg13g2_nand4_1 _16097_ (.B(net387),
    .C(_09339_),
    .A(net1064),
    .Y(_09355_),
    .D(_09351_));
 sg13g2_buf_1 _16098_ (.A(\cpu.spi.r_state[2] ),
    .X(_09356_));
 sg13g2_buf_1 _16099_ (.A(\cpu.spi.r_state[4] ),
    .X(_09357_));
 sg13g2_buf_1 _16100_ (.A(_09296_),
    .X(_09358_));
 sg13g2_buf_1 _16101_ (.A(_09358_),
    .X(_09359_));
 sg13g2_a21oi_1 _16102_ (.A1(_09311_),
    .A2(net87),
    .Y(_09360_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_nand3b_1 _16103_ (.B(net387),
    .C(_09360_),
    .Y(_09361_),
    .A_N(_09357_));
 sg13g2_o21ai_1 _16104_ (.B1(_09361_),
    .Y(_09362_),
    .A1(net1143),
    .A2(net387));
 sg13g2_buf_1 _16105_ (.A(net917),
    .X(_09363_));
 sg13g2_buf_1 _16106_ (.A(net795),
    .X(_09364_));
 sg13g2_a21oi_1 _16107_ (.A1(_09355_),
    .A2(_09362_),
    .Y(_00031_),
    .B1(net692));
 sg13g2_buf_1 _16108_ (.A(net795),
    .X(_09365_));
 sg13g2_nor3_1 _16109_ (.A(net691),
    .B(net387),
    .C(_09299_),
    .Y(_00032_));
 sg13g2_nand3_1 _16110_ (.B(_09240_),
    .C(net87),
    .A(net1144),
    .Y(_09366_));
 sg13g2_nand2_1 _16111_ (.Y(_09367_),
    .A(_09357_),
    .B(_09217_));
 sg13g2_buf_2 _16112_ (.A(net795),
    .X(_09368_));
 sg13g2_buf_1 _16113_ (.A(_09368_),
    .X(_09369_));
 sg13g2_a21oi_1 _16114_ (.A1(_09366_),
    .A2(_09367_),
    .Y(_00033_),
    .B1(net623));
 sg13g2_nor3_1 _16115_ (.A(net691),
    .B(net387),
    .C(_09360_),
    .Y(_00034_));
 sg13g2_nand2_1 _16116_ (.Y(_09370_),
    .A(net1064),
    .B(net388));
 sg13g2_nand2_1 _16117_ (.Y(_09371_),
    .A(net1143),
    .B(net387));
 sg13g2_a21oi_1 _16118_ (.A1(_09370_),
    .A2(_09371_),
    .Y(_00035_),
    .B1(net623));
 sg13g2_buf_1 _16119_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09372_));
 sg13g2_buf_1 _16120_ (.A(\cpu.dec.mult ),
    .X(_09373_));
 sg13g2_inv_1 _16121_ (.Y(_09374_),
    .A(_09373_));
 sg13g2_nand3b_1 _16122_ (.B(\cpu.dec.iready ),
    .C(_00199_),
    .Y(_09375_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_2 _16123_ (.A(_09375_),
    .X(_09376_));
 sg13g2_nor3_1 _16124_ (.A(_09374_),
    .B(_09303_),
    .C(_09376_),
    .Y(_09377_));
 sg13g2_inv_1 _16125_ (.Y(_09378_),
    .A(\cpu.dec.div ));
 sg13g2_nor3_1 _16126_ (.A(_09378_),
    .B(_09303_),
    .C(_09376_),
    .Y(_09379_));
 sg13g2_buf_2 _16127_ (.A(_09379_),
    .X(_09380_));
 sg13g2_nor2_1 _16128_ (.A(_09377_),
    .B(_09380_),
    .Y(_09381_));
 sg13g2_buf_1 _16129_ (.A(_09381_),
    .X(_09382_));
 sg13g2_and2_1 _16130_ (.A(net1142),
    .B(net622),
    .X(_09383_));
 sg13g2_buf_2 _16131_ (.A(_09383_),
    .X(_09384_));
 sg13g2_inv_2 _16132_ (.Y(\cpu.ex.c_mult_off[0] ),
    .A(_09384_));
 sg13g2_buf_2 _16133_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09385_));
 sg13g2_buf_2 _16134_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09386_));
 sg13g2_or3_1 _16135_ (.A(_09385_),
    .B(_09386_),
    .C(\cpu.ex.c_mult_off[0] ),
    .X(_09387_));
 sg13g2_buf_2 _16136_ (.A(_09387_),
    .X(_09388_));
 sg13g2_nor2_2 _16137_ (.A(\cpu.ex.r_mult_off[3] ),
    .B(_09388_),
    .Y(_09389_));
 sg13g2_buf_1 _16138_ (.A(_09380_),
    .X(_09390_));
 sg13g2_o21ai_1 _16139_ (.B1(_09306_),
    .Y(_09391_),
    .A1(\cpu.ex.r_div_running ),
    .A2(net690));
 sg13g2_a21oi_1 _16140_ (.A1(\cpu.ex.r_div_running ),
    .A2(_09389_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09391_));
 sg13g2_buf_1 _16141_ (.A(\cpu.ex.r_mult_running ),
    .X(_09392_));
 sg13g2_buf_1 _16142_ (.A(_09377_),
    .X(_09393_));
 sg13g2_buf_1 _16143_ (.A(_09393_),
    .X(_09394_));
 sg13g2_o21ai_1 _16144_ (.B1(net1066),
    .Y(_09395_),
    .A1(\cpu.ex.r_mult_running ),
    .A2(net689));
 sg13g2_a21oi_1 _16145_ (.A1(net1141),
    .A2(_09389_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09395_));
 sg13g2_inv_1 _16146_ (.Y(_09396_),
    .A(\cpu.qspi.r_state[17] ));
 sg13g2_inv_2 _16147_ (.Y(_09397_),
    .A(_08310_));
 sg13g2_buf_2 _16148_ (.A(\cpu.dcache.flush_write ),
    .X(_09398_));
 sg13g2_inv_1 _16149_ (.Y(_09399_),
    .A(_09398_));
 sg13g2_buf_8 _16150_ (.A(_08300_),
    .X(_09400_));
 sg13g2_buf_8 _16151_ (.A(net914),
    .X(_09401_));
 sg13g2_buf_8 _16152_ (.A(_08298_),
    .X(_09402_));
 sg13g2_buf_2 _16153_ (.A(net913),
    .X(_09403_));
 sg13g2_mux4_1 _16154_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net792),
    .X(_09404_));
 sg13g2_mux4_1 _16155_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net792),
    .X(_09405_));
 sg13g2_buf_8 _16156_ (.A(_08300_),
    .X(_09406_));
 sg13g2_buf_8 _16157_ (.A(_09406_),
    .X(_09407_));
 sg13g2_buf_2 _16158_ (.A(net913),
    .X(_09408_));
 sg13g2_mux4_1 _16159_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net790),
    .X(_09409_));
 sg13g2_buf_8 _16160_ (.A(_09406_),
    .X(_09410_));
 sg13g2_mux4_1 _16161_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net790),
    .X(_09411_));
 sg13g2_buf_2 _16162_ (.A(_08425_),
    .X(_09412_));
 sg13g2_buf_1 _16163_ (.A(net823),
    .X(_09413_));
 sg13g2_mux4_1 _16164_ (.S0(net788),
    .A0(_09404_),
    .A1(_09405_),
    .A2(_09409_),
    .A3(_09411_),
    .S1(net688),
    .X(_09414_));
 sg13g2_nand2_1 _16165_ (.Y(_09415_),
    .A(net822),
    .B(_09414_));
 sg13g2_buf_1 _16166_ (.A(net824),
    .X(_09416_));
 sg13g2_mux4_1 _16167_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(net790),
    .X(_09417_));
 sg13g2_mux4_1 _16168_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(_09403_),
    .X(_09418_));
 sg13g2_buf_2 _16169_ (.A(net913),
    .X(_09419_));
 sg13g2_mux4_1 _16170_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(_09419_),
    .X(_09420_));
 sg13g2_mux4_1 _16171_ (.S0(_09407_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net787),
    .X(_09421_));
 sg13g2_buf_2 _16172_ (.A(net823),
    .X(_09422_));
 sg13g2_mux4_1 _16173_ (.S0(net788),
    .A0(_09417_),
    .A1(_09418_),
    .A2(_09420_),
    .A3(_09421_),
    .S1(net686),
    .X(_09423_));
 sg13g2_nand2_1 _16174_ (.Y(_09424_),
    .A(net687),
    .B(_09423_));
 sg13g2_a21oi_1 _16175_ (.A1(_09415_),
    .A2(_09424_),
    .Y(_09425_),
    .B1(_08459_));
 sg13g2_buf_2 _16176_ (.A(_09425_),
    .X(_09426_));
 sg13g2_buf_2 _16177_ (.A(\cpu.addr[4] ),
    .X(_09427_));
 sg13g2_and3_1 _16178_ (.X(_09428_),
    .A(_09233_),
    .B(_09427_),
    .C(net1146));
 sg13g2_buf_1 _16179_ (.A(_09428_),
    .X(_09429_));
 sg13g2_buf_1 _16180_ (.A(_09429_),
    .X(_09430_));
 sg13g2_buf_1 _16181_ (.A(_00229_),
    .X(_09431_));
 sg13g2_nand2_1 _16182_ (.Y(_09432_),
    .A(_09233_),
    .B(_09431_));
 sg13g2_buf_2 _16183_ (.A(_09432_),
    .X(_09433_));
 sg13g2_nor2_1 _16184_ (.A(_09427_),
    .B(net1146),
    .Y(_09434_));
 sg13g2_buf_1 _16185_ (.A(_09434_),
    .X(_09435_));
 sg13g2_and2_1 _16186_ (.A(_09433_),
    .B(net912),
    .X(_09436_));
 sg13g2_buf_2 _16187_ (.A(_09436_),
    .X(_09437_));
 sg13g2_buf_1 _16188_ (.A(_09437_),
    .X(_09438_));
 sg13g2_inv_1 _16189_ (.Y(_09439_),
    .A(_00253_));
 sg13g2_a22oi_1 _16190_ (.Y(_09440_),
    .B1(net621),
    .B2(_09439_),
    .A2(net786),
    .A1(\cpu.dcache.r_tag[7][23] ));
 sg13g2_nor2_1 _16191_ (.A(net915),
    .B(_09433_),
    .Y(_09441_));
 sg13g2_buf_1 _16192_ (.A(_09441_),
    .X(_09442_));
 sg13g2_nor2b_1 _16193_ (.A(_09233_),
    .B_N(_09218_),
    .Y(_09443_));
 sg13g2_buf_1 _16194_ (.A(_09443_),
    .X(_09444_));
 sg13g2_and2_1 _16195_ (.A(net1140),
    .B(_09444_),
    .X(_09445_));
 sg13g2_buf_1 _16196_ (.A(_09445_),
    .X(_09446_));
 sg13g2_buf_1 _16197_ (.A(net684),
    .X(_09447_));
 sg13g2_a22oi_1 _16198_ (.Y(_09448_),
    .B1(net620),
    .B2(\cpu.dcache.r_tag[2][23] ),
    .A2(net685),
    .A1(\cpu.dcache.r_tag[3][23] ));
 sg13g2_buf_1 _16199_ (.A(net1146),
    .X(_09449_));
 sg13g2_nor2b_1 _16200_ (.A(_09233_),
    .B_N(_09427_),
    .Y(_09450_));
 sg13g2_buf_2 _16201_ (.A(_09450_),
    .X(_09451_));
 sg13g2_and2_1 _16202_ (.A(_09449_),
    .B(_09451_),
    .X(_09452_));
 sg13g2_buf_2 _16203_ (.A(_09452_),
    .X(_09453_));
 sg13g2_buf_1 _16204_ (.A(_09453_),
    .X(_09454_));
 sg13g2_nor2_1 _16205_ (.A(net1063),
    .B(_09433_),
    .Y(_09455_));
 sg13g2_buf_2 _16206_ (.A(_09455_),
    .X(_09456_));
 sg13g2_buf_1 _16207_ (.A(_09456_),
    .X(_09457_));
 sg13g2_nand2_1 _16208_ (.Y(_09458_),
    .A(net918),
    .B(\cpu.dcache.r_tag[5][23] ));
 sg13g2_inv_2 _16209_ (.Y(_09459_),
    .A(_09234_));
 sg13g2_buf_1 _16210_ (.A(_09459_),
    .X(_09460_));
 sg13g2_nand2_1 _16211_ (.Y(_09461_),
    .A(net785),
    .B(\cpu.dcache.r_tag[4][23] ));
 sg13g2_nand2b_1 _16212_ (.Y(_09462_),
    .B(_09427_),
    .A_N(net1146));
 sg13g2_buf_2 _16213_ (.A(_09462_),
    .X(_09463_));
 sg13g2_a21oi_1 _16214_ (.A1(_09458_),
    .A2(_09461_),
    .Y(_09464_),
    .B1(_09463_));
 sg13g2_a221oi_1 _16215_ (.B2(\cpu.dcache.r_tag[1][23] ),
    .C1(_09464_),
    .B1(net618),
    .A1(\cpu.dcache.r_tag[6][23] ),
    .Y(_09465_),
    .A2(net619));
 sg13g2_nand3_1 _16216_ (.B(_09448_),
    .C(_09465_),
    .A(_09440_),
    .Y(_09466_));
 sg13g2_xnor2_1 _16217_ (.Y(_09467_),
    .A(_09426_),
    .B(_09466_));
 sg13g2_mux4_1 _16218_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net787),
    .X(_09468_));
 sg13g2_mux4_1 _16219_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net787),
    .X(_09469_));
 sg13g2_buf_8 _16220_ (.A(_09406_),
    .X(_09470_));
 sg13g2_buf_2 _16221_ (.A(_08298_),
    .X(_09471_));
 sg13g2_mux4_1 _16222_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net911),
    .X(_09472_));
 sg13g2_buf_8 _16223_ (.A(_09406_),
    .X(_09473_));
 sg13g2_mux4_1 _16224_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net911),
    .X(_09474_));
 sg13g2_mux4_1 _16225_ (.S0(net788),
    .A0(_09468_),
    .A1(_09469_),
    .A2(_09472_),
    .A3(_09474_),
    .S1(net686),
    .X(_09475_));
 sg13g2_nand2_1 _16226_ (.Y(_09476_),
    .A(net822),
    .B(_09475_));
 sg13g2_mux4_1 _16227_ (.S0(_09473_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(net787),
    .X(_09477_));
 sg13g2_mux4_1 _16228_ (.S0(_09407_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(_09419_),
    .X(_09478_));
 sg13g2_buf_2 _16229_ (.A(_08298_),
    .X(_09479_));
 sg13g2_mux4_1 _16230_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(_09479_),
    .X(_09480_));
 sg13g2_mux4_1 _16231_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net910),
    .X(_09481_));
 sg13g2_mux4_1 _16232_ (.S0(_09412_),
    .A0(_09477_),
    .A1(_09478_),
    .A2(_09480_),
    .A3(_09481_),
    .S1(_09422_),
    .X(_09482_));
 sg13g2_nand2_1 _16233_ (.Y(_09483_),
    .A(net687),
    .B(_09482_));
 sg13g2_a21oi_2 _16234_ (.B1(_08459_),
    .Y(_09484_),
    .A2(_09483_),
    .A1(_09476_));
 sg13g2_buf_8 _16235_ (.A(_09484_),
    .X(_09485_));
 sg13g2_a22oi_1 _16236_ (.Y(_09486_),
    .B1(net684),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(net786),
    .A1(\cpu.dcache.r_tag[7][19] ));
 sg13g2_inv_1 _16237_ (.Y(_09487_),
    .A(_00252_));
 sg13g2_nor2_1 _16238_ (.A(_09459_),
    .B(_09463_),
    .Y(_09488_));
 sg13g2_buf_1 _16239_ (.A(_09488_),
    .X(_09489_));
 sg13g2_a22oi_1 _16240_ (.Y(_09490_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][19] ),
    .A2(_09437_),
    .A1(_09487_));
 sg13g2_and2_1 _16241_ (.A(net915),
    .B(_09451_),
    .X(_09491_));
 sg13g2_buf_2 _16242_ (.A(_09491_),
    .X(_09492_));
 sg13g2_buf_1 _16243_ (.A(_09492_),
    .X(_09493_));
 sg13g2_a22oi_1 _16244_ (.Y(_09494_),
    .B1(net617),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(net618),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_a22oi_1 _16245_ (.Y(_09495_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[3][19] ),
    .A2(net619),
    .A1(\cpu.dcache.r_tag[6][19] ));
 sg13g2_nand4_1 _16246_ (.B(_09490_),
    .C(_09494_),
    .A(_09486_),
    .Y(_09496_),
    .D(_09495_));
 sg13g2_xnor2_1 _16247_ (.Y(_09497_),
    .A(net435),
    .B(_09496_));
 sg13g2_mux4_1 _16248_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net911),
    .X(_09498_));
 sg13g2_mux4_1 _16249_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(_09471_),
    .X(_09499_));
 sg13g2_mux4_1 _16250_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net910),
    .X(_09500_));
 sg13g2_mux4_1 _16251_ (.S0(_09470_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net910),
    .X(_09501_));
 sg13g2_mux4_1 _16252_ (.S0(_09412_),
    .A0(_09498_),
    .A1(_09499_),
    .A2(_09500_),
    .A3(_09501_),
    .S1(net686),
    .X(_09502_));
 sg13g2_nand2_1 _16253_ (.Y(_09503_),
    .A(net822),
    .B(_09502_));
 sg13g2_mux4_1 _16254_ (.S0(_09470_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09471_),
    .X(_09504_));
 sg13g2_mux4_1 _16255_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net911),
    .X(_09505_));
 sg13g2_buf_8 _16256_ (.A(_09406_),
    .X(_09506_));
 sg13g2_mux4_1 _16257_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(_09479_),
    .X(_09507_));
 sg13g2_mux4_1 _16258_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net910),
    .X(_09508_));
 sg13g2_buf_2 _16259_ (.A(_08425_),
    .X(_09509_));
 sg13g2_mux4_1 _16260_ (.S0(_09509_),
    .A0(_09504_),
    .A1(_09505_),
    .A2(_09507_),
    .A3(_09508_),
    .S1(_09422_),
    .X(_09510_));
 sg13g2_nand2_1 _16261_ (.Y(_09511_),
    .A(net687),
    .B(_09510_));
 sg13g2_a21oi_2 _16262_ (.B1(_08459_),
    .Y(_09512_),
    .A2(_09511_),
    .A1(_09503_));
 sg13g2_buf_1 _16263_ (.A(_09512_),
    .X(_09513_));
 sg13g2_nand2_1 _16264_ (.Y(_09514_),
    .A(_09433_),
    .B(net912));
 sg13g2_buf_2 _16265_ (.A(_09514_),
    .X(_09515_));
 sg13g2_buf_1 _16266_ (.A(_09515_),
    .X(_09516_));
 sg13g2_a22oi_1 _16267_ (.Y(_09517_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[3][17] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][17] ));
 sg13g2_a22oi_1 _16268_ (.Y(_09518_),
    .B1(net684),
    .B2(\cpu.dcache.r_tag[2][17] ),
    .A2(_09456_),
    .A1(\cpu.dcache.r_tag[1][17] ));
 sg13g2_mux2_1 _16269_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(\cpu.dcache.r_tag[7][17] ),
    .S(net1063),
    .X(_09519_));
 sg13g2_nor2_1 _16270_ (.A(_09233_),
    .B(net1146),
    .Y(_09520_));
 sg13g2_buf_2 _16271_ (.A(_09520_),
    .X(_09521_));
 sg13g2_a22oi_1 _16272_ (.Y(_09522_),
    .B1(_09521_),
    .B2(\cpu.dcache.r_tag[4][17] ),
    .A2(_09519_),
    .A1(net1068));
 sg13g2_buf_1 _16273_ (.A(_09427_),
    .X(_09523_));
 sg13g2_buf_1 _16274_ (.A(_09523_),
    .X(_09524_));
 sg13g2_nand2b_1 _16275_ (.Y(_09525_),
    .B(net909),
    .A_N(_09522_));
 sg13g2_and4_1 _16276_ (.A(net616),
    .B(_09517_),
    .C(_09518_),
    .D(_09525_),
    .X(_09526_));
 sg13g2_a21oi_1 _16277_ (.A1(_00250_),
    .A2(net621),
    .Y(_09527_),
    .B1(_09526_));
 sg13g2_xnor2_1 _16278_ (.Y(_09528_),
    .A(net434),
    .B(_09527_));
 sg13g2_mux4_1 _16279_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net911),
    .X(_09529_));
 sg13g2_mux4_1 _16280_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net911),
    .X(_09530_));
 sg13g2_mux4_1 _16281_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net910),
    .X(_09531_));
 sg13g2_mux4_1 _16282_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net910),
    .X(_09532_));
 sg13g2_mux4_1 _16283_ (.S0(net781),
    .A0(_09529_),
    .A1(_09530_),
    .A2(_09531_),
    .A3(_09532_),
    .S1(net686),
    .X(_09533_));
 sg13g2_nand2_1 _16284_ (.Y(_09534_),
    .A(net822),
    .B(_09533_));
 sg13g2_mux4_1 _16285_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net911),
    .X(_09535_));
 sg13g2_mux4_1 _16286_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net911),
    .X(_09536_));
 sg13g2_buf_2 _16287_ (.A(_08298_),
    .X(_09537_));
 sg13g2_mux4_1 _16288_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net908),
    .X(_09538_));
 sg13g2_mux4_1 _16289_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net908),
    .X(_09539_));
 sg13g2_mux4_1 _16290_ (.S0(net781),
    .A0(_09535_),
    .A1(_09536_),
    .A2(_09538_),
    .A3(_09539_),
    .S1(net686),
    .X(_09540_));
 sg13g2_nand2_1 _16291_ (.Y(_09541_),
    .A(_09416_),
    .B(_09540_));
 sg13g2_a21oi_1 _16292_ (.A1(_09534_),
    .A2(_09541_),
    .Y(_09542_),
    .B1(_08459_));
 sg13g2_buf_1 _16293_ (.A(_09542_),
    .X(_09543_));
 sg13g2_a22oi_1 _16294_ (.Y(_09544_),
    .B1(net621),
    .B2(\cpu.dcache.r_tag[0][20] ),
    .A2(net786),
    .A1(\cpu.dcache.r_tag[7][20] ));
 sg13g2_a22oi_1 _16295_ (.Y(_09545_),
    .B1(net617),
    .B2(\cpu.dcache.r_tag[4][20] ),
    .A2(net618),
    .A1(\cpu.dcache.r_tag[1][20] ));
 sg13g2_a22oi_1 _16296_ (.Y(_09546_),
    .B1(_09489_),
    .B2(\cpu.dcache.r_tag[5][20] ),
    .A2(net619),
    .A1(\cpu.dcache.r_tag[6][20] ));
 sg13g2_buf_1 _16297_ (.A(net685),
    .X(_09547_));
 sg13g2_a22oi_1 _16298_ (.Y(_09548_),
    .B1(net620),
    .B2(\cpu.dcache.r_tag[2][20] ),
    .A2(net615),
    .A1(\cpu.dcache.r_tag[3][20] ));
 sg13g2_nand4_1 _16299_ (.B(_09545_),
    .C(_09546_),
    .A(_09544_),
    .Y(_09549_),
    .D(_09548_));
 sg13g2_xnor2_1 _16300_ (.Y(_09550_),
    .A(net433),
    .B(_09549_));
 sg13g2_nand4_1 _16301_ (.B(_09497_),
    .C(_09528_),
    .A(_09467_),
    .Y(_09551_),
    .D(_09550_));
 sg13g2_inv_1 _16302_ (.Y(_09552_),
    .A(_00248_));
 sg13g2_a22oi_1 _16303_ (.Y(_09553_),
    .B1(net617),
    .B2(\cpu.dcache.r_tag[4][15] ),
    .A2(_09438_),
    .A1(_09552_));
 sg13g2_a22oi_1 _16304_ (.Y(_09554_),
    .B1(net620),
    .B2(\cpu.dcache.r_tag[2][15] ),
    .A2(net618),
    .A1(\cpu.dcache.r_tag[1][15] ));
 sg13g2_a22oi_1 _16305_ (.Y(_09555_),
    .B1(net619),
    .B2(\cpu.dcache.r_tag[6][15] ),
    .A2(_09430_),
    .A1(\cpu.dcache.r_tag[7][15] ));
 sg13g2_a22oi_1 _16306_ (.Y(_09556_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][15] ),
    .A2(_09442_),
    .A1(\cpu.dcache.r_tag[3][15] ));
 sg13g2_nand4_1 _16307_ (.B(_09554_),
    .C(_09555_),
    .A(_09553_),
    .Y(_09557_),
    .D(_09556_));
 sg13g2_buf_1 _16308_ (.A(net1094),
    .X(_09558_));
 sg13g2_mux4_1 _16309_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net792),
    .X(_09559_));
 sg13g2_mux4_1 _16310_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net792),
    .X(_09560_));
 sg13g2_mux4_1 _16311_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net790),
    .X(_09561_));
 sg13g2_mux4_1 _16312_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(net790),
    .X(_09562_));
 sg13g2_mux4_1 _16313_ (.S0(net824),
    .A0(_09559_),
    .A1(_09560_),
    .A2(_09561_),
    .A3(_09562_),
    .S1(net686),
    .X(_09563_));
 sg13g2_nand2_1 _16314_ (.Y(_09564_),
    .A(net1155),
    .B(_09563_));
 sg13g2_buf_8 _16315_ (.A(net914),
    .X(_09565_));
 sg13g2_buf_2 _16316_ (.A(net913),
    .X(_09566_));
 sg13g2_mux4_1 _16317_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net779),
    .X(_09567_));
 sg13g2_mux4_1 _16318_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(net779),
    .X(_09568_));
 sg13g2_mux4_1 _16319_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net792),
    .X(_09569_));
 sg13g2_mux4_1 _16320_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net792),
    .X(_09570_));
 sg13g2_mux4_1 _16321_ (.S0(net824),
    .A0(_09567_),
    .A1(_09568_),
    .A2(_09569_),
    .A3(_09570_),
    .S1(net688),
    .X(_09571_));
 sg13g2_o21ai_1 _16322_ (.B1(net1094),
    .Y(_09572_),
    .A1(_08449_),
    .A2(_09571_));
 sg13g2_o21ai_1 _16323_ (.B1(_09572_),
    .Y(_09573_),
    .A1(net907),
    .A2(_09564_));
 sg13g2_buf_1 _16324_ (.A(_09573_),
    .X(_09574_));
 sg13g2_xnor2_1 _16325_ (.Y(_09575_),
    .A(_09557_),
    .B(_09574_));
 sg13g2_mux4_1 _16326_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net779),
    .X(_09576_));
 sg13g2_mux4_1 _16327_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net779),
    .X(_09577_));
 sg13g2_mux4_1 _16328_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net790),
    .X(_09578_));
 sg13g2_mux4_1 _16329_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net792),
    .X(_09579_));
 sg13g2_mux4_1 _16330_ (.S0(net788),
    .A0(_09576_),
    .A1(_09577_),
    .A2(_09578_),
    .A3(_09579_),
    .S1(net688),
    .X(_09580_));
 sg13g2_nand2_1 _16331_ (.Y(_09581_),
    .A(net822),
    .B(_09580_));
 sg13g2_mux4_1 _16332_ (.S0(_09401_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(_09403_),
    .X(_09582_));
 sg13g2_mux4_1 _16333_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(_09566_),
    .X(_09583_));
 sg13g2_mux4_1 _16334_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net790),
    .X(_09584_));
 sg13g2_mux4_1 _16335_ (.S0(_09410_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(_09408_),
    .X(_09585_));
 sg13g2_mux4_1 _16336_ (.S0(net788),
    .A0(_09582_),
    .A1(_09583_),
    .A2(_09584_),
    .A3(_09585_),
    .S1(net688),
    .X(_09586_));
 sg13g2_nand2_1 _16337_ (.Y(_09587_),
    .A(net687),
    .B(_09586_));
 sg13g2_a21oi_2 _16338_ (.B1(_08460_),
    .Y(_09588_),
    .A2(_09587_),
    .A1(_09581_));
 sg13g2_buf_1 _16339_ (.A(_09588_),
    .X(_09589_));
 sg13g2_nand2_1 _16340_ (.Y(_09590_),
    .A(\cpu.dcache.r_tag[4][22] ),
    .B(net617));
 sg13g2_a22oi_1 _16341_ (.Y(_09591_),
    .B1(net684),
    .B2(\cpu.dcache.r_tag[2][22] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][22] ));
 sg13g2_a22oi_1 _16342_ (.Y(_09592_),
    .B1(net618),
    .B2(\cpu.dcache.r_tag[1][22] ),
    .A2(_09429_),
    .A1(\cpu.dcache.r_tag[7][22] ));
 sg13g2_a22oi_1 _16343_ (.Y(_09593_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][22] ),
    .A2(net685),
    .A1(\cpu.dcache.r_tag[3][22] ));
 sg13g2_nand4_1 _16344_ (.B(_09591_),
    .C(_09592_),
    .A(_09590_),
    .Y(_09594_),
    .D(_09593_));
 sg13g2_mux2_1 _16345_ (.A0(\cpu.dcache.r_tag[0][22] ),
    .A1(_09594_),
    .S(net616),
    .X(_09595_));
 sg13g2_xnor2_1 _16346_ (.Y(_09596_),
    .A(net431),
    .B(_09595_));
 sg13g2_mux4_1 _16347_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net787),
    .X(_09597_));
 sg13g2_mux4_1 _16348_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net787),
    .X(_09598_));
 sg13g2_mux4_1 _16349_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net910),
    .X(_09599_));
 sg13g2_mux4_1 _16350_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net910),
    .X(_09600_));
 sg13g2_mux4_1 _16351_ (.S0(net824),
    .A0(_09597_),
    .A1(_09598_),
    .A2(_09599_),
    .A3(_09600_),
    .S1(_08316_),
    .X(_09601_));
 sg13g2_nand2_1 _16352_ (.Y(_09602_),
    .A(net1155),
    .B(_09601_));
 sg13g2_mux4_1 _16353_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net790),
    .X(_09603_));
 sg13g2_mux4_1 _16354_ (.S0(_09410_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(_09408_),
    .X(_09604_));
 sg13g2_mux4_1 _16355_ (.S0(net783),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net787),
    .X(_09605_));
 sg13g2_mux4_1 _16356_ (.S0(_09473_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(net787),
    .X(_09606_));
 sg13g2_mux4_1 _16357_ (.S0(_08314_),
    .A0(_09603_),
    .A1(_09604_),
    .A2(_09605_),
    .A3(_09606_),
    .S1(net1094),
    .X(_09607_));
 sg13g2_o21ai_1 _16358_ (.B1(net688),
    .Y(_09608_),
    .A1(_08449_),
    .A2(_09607_));
 sg13g2_o21ai_1 _16359_ (.B1(_09608_),
    .Y(_09609_),
    .A1(_09413_),
    .A2(_09602_));
 sg13g2_buf_1 _16360_ (.A(_09609_),
    .X(_09610_));
 sg13g2_a22oi_1 _16361_ (.Y(_09611_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][14] ),
    .A2(_09456_),
    .A1(\cpu.dcache.r_tag[1][14] ));
 sg13g2_and2_1 _16362_ (.A(\cpu.dcache.r_tag[7][14] ),
    .B(_09429_),
    .X(_09612_));
 sg13g2_a221oi_1 _16363_ (.B2(\cpu.dcache.r_tag[4][14] ),
    .C1(_09612_),
    .B1(_09492_),
    .A1(\cpu.dcache.r_tag[2][14] ),
    .Y(_09613_),
    .A2(net684));
 sg13g2_a22oi_1 _16364_ (.Y(_09614_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[3][14] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][14] ));
 sg13g2_and4_1 _16365_ (.A(_09516_),
    .B(_09611_),
    .C(_09613_),
    .D(_09614_),
    .X(_09615_));
 sg13g2_a21oi_1 _16366_ (.A1(_00247_),
    .A2(net621),
    .Y(_09616_),
    .B1(_09615_));
 sg13g2_xnor2_1 _16367_ (.Y(_09617_),
    .A(_09610_),
    .B(_09616_));
 sg13g2_nand3_1 _16368_ (.B(_09596_),
    .C(_09617_),
    .A(_09575_),
    .Y(_09618_));
 sg13g2_a22oi_1 _16369_ (.Y(_09619_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][13] ),
    .A2(_09454_),
    .A1(\cpu.dcache.r_tag[6][13] ));
 sg13g2_inv_1 _16370_ (.Y(_09620_),
    .A(_00246_));
 sg13g2_a22oi_1 _16371_ (.Y(_09621_),
    .B1(_09447_),
    .B2(\cpu.dcache.r_tag[2][13] ),
    .A2(net621),
    .A1(_09620_));
 sg13g2_a22oi_1 _16372_ (.Y(_09622_),
    .B1(_09457_),
    .B2(\cpu.dcache.r_tag[1][13] ),
    .A2(net786),
    .A1(\cpu.dcache.r_tag[7][13] ));
 sg13g2_a22oi_1 _16373_ (.Y(_09623_),
    .B1(_09493_),
    .B2(\cpu.dcache.r_tag[4][13] ),
    .A2(_09547_),
    .A1(\cpu.dcache.r_tag[3][13] ));
 sg13g2_nand4_1 _16374_ (.B(_09621_),
    .C(_09622_),
    .A(_09619_),
    .Y(_09624_),
    .D(_09623_));
 sg13g2_buf_8 _16375_ (.A(_09406_),
    .X(_09625_));
 sg13g2_mux4_1 _16376_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net908),
    .X(_09626_));
 sg13g2_mux4_1 _16377_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net908),
    .X(_09627_));
 sg13g2_buf_8 _16378_ (.A(_09406_),
    .X(_09628_));
 sg13g2_buf_2 _16379_ (.A(_08298_),
    .X(_09629_));
 sg13g2_mux4_1 _16380_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net906),
    .X(_09630_));
 sg13g2_mux4_1 _16381_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net906),
    .X(_09631_));
 sg13g2_mux4_1 _16382_ (.S0(net781),
    .A0(_09626_),
    .A1(_09627_),
    .A2(_09630_),
    .A3(_09631_),
    .S1(net686),
    .X(_09632_));
 sg13g2_mux4_1 _16383_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(_09537_),
    .X(_09633_));
 sg13g2_mux4_1 _16384_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net908),
    .X(_09634_));
 sg13g2_buf_2 _16385_ (.A(_08298_),
    .X(_09635_));
 sg13g2_mux4_1 _16386_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net905),
    .X(_09636_));
 sg13g2_mux4_1 _16387_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net905),
    .X(_09637_));
 sg13g2_mux4_1 _16388_ (.S0(net781),
    .A0(_09633_),
    .A1(_09634_),
    .A2(_09636_),
    .A3(_09637_),
    .S1(net823),
    .X(_09638_));
 sg13g2_mux2_1 _16389_ (.A0(_09632_),
    .A1(_09638_),
    .S(net687),
    .X(_09639_));
 sg13g2_nand2_1 _16390_ (.Y(_09640_),
    .A(_08540_),
    .B(_09639_));
 sg13g2_o21ai_1 _16391_ (.B1(_09640_),
    .Y(_09641_),
    .A1(_08540_),
    .A2(net1093));
 sg13g2_buf_1 _16392_ (.A(_09641_),
    .X(_09642_));
 sg13g2_xnor2_1 _16393_ (.Y(_09643_),
    .A(_09624_),
    .B(net386));
 sg13g2_mux4_1 _16394_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net905),
    .X(_09644_));
 sg13g2_mux4_1 _16395_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net906),
    .X(_09645_));
 sg13g2_mux4_1 _16396_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net913),
    .X(_09646_));
 sg13g2_mux4_1 _16397_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net913),
    .X(_09647_));
 sg13g2_mux4_1 _16398_ (.S0(net781),
    .A0(_09644_),
    .A1(_09645_),
    .A2(_09646_),
    .A3(_09647_),
    .S1(net823),
    .X(_09648_));
 sg13g2_mux4_1 _16399_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net905),
    .X(_09649_));
 sg13g2_mux4_1 _16400_ (.S0(_09628_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(_09635_),
    .X(_09650_));
 sg13g2_mux4_1 _16401_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(net913),
    .X(_09651_));
 sg13g2_mux4_1 _16402_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(_09402_),
    .X(_09652_));
 sg13g2_mux4_1 _16403_ (.S0(_08425_),
    .A0(_09649_),
    .A1(_09650_),
    .A2(_09651_),
    .A3(_09652_),
    .S1(net823),
    .X(_09653_));
 sg13g2_mux2_1 _16404_ (.A0(_09648_),
    .A1(_09653_),
    .S(_08314_),
    .X(_09654_));
 sg13g2_nand2_1 _16405_ (.Y(_09655_),
    .A(net1155),
    .B(_09654_));
 sg13g2_o21ai_1 _16406_ (.B1(_09655_),
    .Y(_09656_),
    .A1(net1083),
    .A2(_08428_));
 sg13g2_buf_1 _16407_ (.A(_09656_),
    .X(_09657_));
 sg13g2_a22oi_1 _16408_ (.Y(_09658_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[3][12] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][12] ));
 sg13g2_a22oi_1 _16409_ (.Y(_09659_),
    .B1(_09446_),
    .B2(\cpu.dcache.r_tag[2][12] ),
    .A2(_09456_),
    .A1(\cpu.dcache.r_tag[1][12] ));
 sg13g2_mux2_1 _16410_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(\cpu.dcache.r_tag[7][12] ),
    .S(net1063),
    .X(_09660_));
 sg13g2_a22oi_1 _16411_ (.Y(_09661_),
    .B1(_09660_),
    .B2(net918),
    .A2(_09521_),
    .A1(\cpu.dcache.r_tag[4][12] ));
 sg13g2_nand2b_1 _16412_ (.Y(_09662_),
    .B(net909),
    .A_N(_09661_));
 sg13g2_and4_1 _16413_ (.A(net616),
    .B(_09658_),
    .C(_09659_),
    .D(_09662_),
    .X(_09663_));
 sg13g2_a21oi_1 _16414_ (.A1(_00245_),
    .A2(net621),
    .Y(_09664_),
    .B1(_09663_));
 sg13g2_xnor2_1 _16415_ (.Y(_09665_),
    .A(net385),
    .B(_09664_));
 sg13g2_nand2_1 _16416_ (.Y(_09666_),
    .A(_09643_),
    .B(_09665_));
 sg13g2_mux4_1 _16417_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net906),
    .X(_09667_));
 sg13g2_mux4_1 _16418_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net906),
    .X(_09668_));
 sg13g2_mux4_1 _16419_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net905),
    .X(_09669_));
 sg13g2_mux4_1 _16420_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net905),
    .X(_09670_));
 sg13g2_mux4_1 _16421_ (.S0(net781),
    .A0(_09667_),
    .A1(_09668_),
    .A2(_09669_),
    .A3(_09670_),
    .S1(net823),
    .X(_09671_));
 sg13g2_nand2_1 _16422_ (.Y(_09672_),
    .A(net822),
    .B(_09671_));
 sg13g2_mux4_1 _16423_ (.S0(_09625_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(_09629_),
    .X(_09673_));
 sg13g2_mux4_1 _16424_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net906),
    .X(_09674_));
 sg13g2_mux4_1 _16425_ (.S0(_09400_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net905),
    .X(_09675_));
 sg13g2_mux4_1 _16426_ (.S0(_09400_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09635_),
    .X(_09676_));
 sg13g2_mux4_1 _16427_ (.S0(net781),
    .A0(_09673_),
    .A1(_09674_),
    .A2(_09675_),
    .A3(_09676_),
    .S1(_08411_),
    .X(_09677_));
 sg13g2_nand2_1 _16428_ (.Y(_09678_),
    .A(_09416_),
    .B(_09677_));
 sg13g2_a21oi_2 _16429_ (.B1(_08459_),
    .Y(_09679_),
    .A2(_09678_),
    .A1(_09672_));
 sg13g2_buf_1 _16430_ (.A(_09679_),
    .X(_09680_));
 sg13g2_inv_1 _16431_ (.Y(_09681_),
    .A(_00249_));
 sg13g2_a22oi_1 _16432_ (.Y(_09682_),
    .B1(_09489_),
    .B2(\cpu.dcache.r_tag[5][16] ),
    .A2(_09437_),
    .A1(_09681_));
 sg13g2_a22oi_1 _16433_ (.Y(_09683_),
    .B1(net684),
    .B2(\cpu.dcache.r_tag[2][16] ),
    .A2(_09429_),
    .A1(\cpu.dcache.r_tag[7][16] ));
 sg13g2_a22oi_1 _16434_ (.Y(_09684_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[3][16] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][16] ));
 sg13g2_a22oi_1 _16435_ (.Y(_09685_),
    .B1(_09492_),
    .B2(\cpu.dcache.r_tag[4][16] ),
    .A2(_09456_),
    .A1(\cpu.dcache.r_tag[1][16] ));
 sg13g2_nand4_1 _16436_ (.B(_09683_),
    .C(_09684_),
    .A(_09682_),
    .Y(_09686_),
    .D(_09685_));
 sg13g2_xor2_1 _16437_ (.B(_09686_),
    .A(net429),
    .X(_09687_));
 sg13g2_mux4_1 _16438_ (.S0(net782),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net908),
    .X(_09688_));
 sg13g2_mux4_1 _16439_ (.S0(_09506_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net908),
    .X(_09689_));
 sg13g2_mux4_1 _16440_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net906),
    .X(_09690_));
 sg13g2_mux4_1 _16441_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net906),
    .X(_09691_));
 sg13g2_mux4_1 _16442_ (.S0(_09509_),
    .A0(_09688_),
    .A1(_09689_),
    .A2(_09690_),
    .A3(_09691_),
    .S1(net686),
    .X(_09692_));
 sg13g2_nand2_1 _16443_ (.Y(_09693_),
    .A(_08443_),
    .B(_09692_));
 sg13g2_mux4_1 _16444_ (.S0(_09625_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(_09537_),
    .X(_09694_));
 sg13g2_mux4_1 _16445_ (.S0(_09506_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(net908),
    .X(_09695_));
 sg13g2_mux4_1 _16446_ (.S0(_09628_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(net905),
    .X(_09696_));
 sg13g2_mux4_1 _16447_ (.S0(net777),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09629_),
    .X(_09697_));
 sg13g2_mux4_1 _16448_ (.S0(net781),
    .A0(_09694_),
    .A1(_09695_),
    .A2(_09696_),
    .A3(_09697_),
    .S1(_08411_),
    .X(_09698_));
 sg13g2_nand2_1 _16449_ (.Y(_09699_),
    .A(net687),
    .B(_09698_));
 sg13g2_a21oi_2 _16450_ (.B1(_08459_),
    .Y(_09700_),
    .A2(_09699_),
    .A1(_09693_));
 sg13g2_buf_1 _16451_ (.A(_09700_),
    .X(_09701_));
 sg13g2_a22oi_1 _16452_ (.Y(_09702_),
    .B1(net684),
    .B2(\cpu.dcache.r_tag[2][18] ),
    .A2(_09456_),
    .A1(\cpu.dcache.r_tag[1][18] ));
 sg13g2_inv_1 _16453_ (.Y(_09703_),
    .A(_00251_));
 sg13g2_a22oi_1 _16454_ (.Y(_09704_),
    .B1(_09492_),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(_09437_),
    .A1(_09703_));
 sg13g2_a22oi_1 _16455_ (.Y(_09705_),
    .B1(net683),
    .B2(\cpu.dcache.r_tag[5][18] ),
    .A2(_09442_),
    .A1(\cpu.dcache.r_tag[3][18] ));
 sg13g2_a22oi_1 _16456_ (.Y(_09706_),
    .B1(_09453_),
    .B2(\cpu.dcache.r_tag[6][18] ),
    .A2(_09429_),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_nand4_1 _16457_ (.B(_09704_),
    .C(_09705_),
    .A(_09702_),
    .Y(_09707_),
    .D(_09706_));
 sg13g2_xor2_1 _16458_ (.B(_09707_),
    .A(net428),
    .X(_09708_));
 sg13g2_nor2_1 _16459_ (.A(_09687_),
    .B(_09708_),
    .Y(_09709_));
 sg13g2_buf_1 _16460_ (.A(net913),
    .X(_09710_));
 sg13g2_mux4_1 _16461_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net776),
    .X(_09711_));
 sg13g2_mux4_1 _16462_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net776),
    .X(_09712_));
 sg13g2_mux4_1 _16463_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net779),
    .X(_09713_));
 sg13g2_mux4_1 _16464_ (.S0(_09565_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net779),
    .X(_09714_));
 sg13g2_mux4_1 _16465_ (.S0(net788),
    .A0(_09711_),
    .A1(_09712_),
    .A2(_09713_),
    .A3(_09714_),
    .S1(_09413_),
    .X(_09715_));
 sg13g2_nand2_1 _16466_ (.Y(_09716_),
    .A(net822),
    .B(_09715_));
 sg13g2_mux4_1 _16467_ (.S0(net780),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net779),
    .X(_09717_));
 sg13g2_mux4_1 _16468_ (.S0(_09565_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(_09566_),
    .X(_09718_));
 sg13g2_mux4_1 _16469_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net792),
    .X(_09719_));
 sg13g2_mux4_1 _16470_ (.S0(_09401_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net779),
    .X(_09720_));
 sg13g2_mux4_1 _16471_ (.S0(net788),
    .A0(_09717_),
    .A1(_09718_),
    .A2(_09719_),
    .A3(_09720_),
    .S1(net688),
    .X(_09721_));
 sg13g2_nand2_1 _16472_ (.Y(_09722_),
    .A(net687),
    .B(_09721_));
 sg13g2_a21oi_1 _16473_ (.A1(_09716_),
    .A2(_09722_),
    .Y(_09723_),
    .B1(_08460_));
 sg13g2_buf_1 _16474_ (.A(_09723_),
    .X(_09724_));
 sg13g2_nand2_1 _16475_ (.Y(_09725_),
    .A(\cpu.dcache.r_tag[0][21] ),
    .B(net621));
 sg13g2_a22oi_1 _16476_ (.Y(_09726_),
    .B1(net617),
    .B2(\cpu.dcache.r_tag[4][21] ),
    .A2(net615),
    .A1(\cpu.dcache.r_tag[3][21] ));
 sg13g2_a22oi_1 _16477_ (.Y(_09727_),
    .B1(net620),
    .B2(\cpu.dcache.r_tag[2][21] ),
    .A2(_09457_),
    .A1(\cpu.dcache.r_tag[1][21] ));
 sg13g2_buf_1 _16478_ (.A(_09444_),
    .X(_09728_));
 sg13g2_mux2_1 _16479_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(\cpu.dcache.r_tag[7][21] ),
    .S(net1072),
    .X(_09729_));
 sg13g2_a22oi_1 _16480_ (.Y(_09730_),
    .B1(_09729_),
    .B2(net918),
    .A2(net775),
    .A1(\cpu.dcache.r_tag[6][21] ));
 sg13g2_nand2b_1 _16481_ (.Y(_09731_),
    .B(net909),
    .A_N(_09730_));
 sg13g2_nand4_1 _16482_ (.B(_09726_),
    .C(_09727_),
    .A(_09725_),
    .Y(_09732_),
    .D(_09731_));
 sg13g2_xnor2_1 _16483_ (.Y(_09733_),
    .A(net427),
    .B(_09732_));
 sg13g2_nor2_1 _16484_ (.A(_00240_),
    .B(_09515_),
    .Y(_09734_));
 sg13g2_and2_1 _16485_ (.A(net1072),
    .B(\cpu.dcache.r_tag[3][9] ),
    .X(_09735_));
 sg13g2_a21oi_1 _16486_ (.A1(net915),
    .A2(\cpu.dcache.r_tag[1][9] ),
    .Y(_09736_),
    .B1(_09735_));
 sg13g2_buf_1 _16487_ (.A(net1140),
    .X(_09737_));
 sg13g2_a22oi_1 _16488_ (.Y(_09738_),
    .B1(\cpu.dcache.r_tag[2][9] ),
    .B2(net1061),
    .A2(\cpu.dcache.r_tag[6][9] ),
    .A1(_09523_));
 sg13g2_nand2b_1 _16489_ (.Y(_09739_),
    .B(net775),
    .A_N(_09738_));
 sg13g2_o21ai_1 _16490_ (.B1(_09739_),
    .Y(_09740_),
    .A1(_09433_),
    .A2(_09736_));
 sg13g2_inv_1 _16491_ (.Y(_09741_),
    .A(_09427_));
 sg13g2_buf_1 _16492_ (.A(_09741_),
    .X(_09742_));
 sg13g2_mux2_1 _16493_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(net1072),
    .X(_09743_));
 sg13g2_a22oi_1 _16494_ (.Y(_09744_),
    .B1(_09743_),
    .B2(_09235_),
    .A2(_09521_),
    .A1(\cpu.dcache.r_tag[4][9] ));
 sg13g2_nor2_1 _16495_ (.A(net904),
    .B(_09744_),
    .Y(_09745_));
 sg13g2_nor3_1 _16496_ (.A(_09734_),
    .B(_09740_),
    .C(_09745_),
    .Y(_09746_));
 sg13g2_xor2_1 _16497_ (.B(_09746_),
    .A(_00239_),
    .X(_09747_));
 sg13g2_mux2_1 _16498_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(\cpu.dcache.r_tag[3][8] ),
    .S(net1063),
    .X(_09748_));
 sg13g2_mux2_1 _16499_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(\cpu.dcache.r_tag[7][8] ),
    .S(net1063),
    .X(_09749_));
 sg13g2_a22oi_1 _16500_ (.Y(_09750_),
    .B1(_09749_),
    .B2(net1062),
    .A2(_09748_),
    .A1(net1061));
 sg13g2_nand2b_1 _16501_ (.Y(_09751_),
    .B(_09235_),
    .A_N(_09750_));
 sg13g2_a22oi_1 _16502_ (.Y(_09752_),
    .B1(_09492_),
    .B2(\cpu.dcache.r_tag[4][8] ),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[6][8] ));
 sg13g2_nand2b_1 _16503_ (.Y(_09753_),
    .B(_09437_),
    .A_N(_00238_));
 sg13g2_and2_1 _16504_ (.A(net1072),
    .B(net1061),
    .X(_09754_));
 sg13g2_nand3_1 _16505_ (.B(\cpu.dcache.r_tag[2][8] ),
    .C(_09754_),
    .A(net785),
    .Y(_09755_));
 sg13g2_and4_1 _16506_ (.A(_09751_),
    .B(_09752_),
    .C(_09753_),
    .D(_09755_),
    .X(_09756_));
 sg13g2_xor2_1 _16507_ (.B(_09756_),
    .A(_00237_),
    .X(_09757_));
 sg13g2_buf_1 _16508_ (.A(_00231_),
    .X(_09758_));
 sg13g2_inv_1 _16509_ (.Y(_09759_),
    .A(_00232_));
 sg13g2_a22oi_1 _16510_ (.Y(_09760_),
    .B1(_09492_),
    .B2(\cpu.dcache.r_tag[4][5] ),
    .A2(_09437_),
    .A1(_09759_));
 sg13g2_mux2_1 _16511_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(\cpu.dcache.r_tag[7][5] ),
    .S(net918),
    .X(_09761_));
 sg13g2_nor2_2 _16512_ (.A(net904),
    .B(_09313_),
    .Y(_09762_));
 sg13g2_a22oi_1 _16513_ (.Y(_09763_),
    .B1(_09761_),
    .B2(_09762_),
    .A2(net684),
    .A1(\cpu.dcache.r_tag[2][5] ));
 sg13g2_a22oi_1 _16514_ (.Y(_09764_),
    .B1(\cpu.dcache.r_tag[1][5] ),
    .B2(net1061),
    .A2(\cpu.dcache.r_tag[5][5] ),
    .A1(net1062));
 sg13g2_nand3_1 _16515_ (.B(net1061),
    .C(\cpu.dcache.r_tag[3][5] ),
    .A(net1072),
    .Y(_09765_));
 sg13g2_o21ai_1 _16516_ (.B1(_09765_),
    .Y(_09766_),
    .A1(net919),
    .A2(_09764_));
 sg13g2_nand2_1 _16517_ (.Y(_09767_),
    .A(net918),
    .B(_09766_));
 sg13g2_nand3_1 _16518_ (.B(_09763_),
    .C(_09767_),
    .A(_09760_),
    .Y(_09768_));
 sg13g2_xnor2_1 _16519_ (.Y(_09769_),
    .A(_09758_),
    .B(_09768_));
 sg13g2_nor3_1 _16520_ (.A(_09747_),
    .B(_09757_),
    .C(_09769_),
    .Y(_09770_));
 sg13g2_nand2_1 _16521_ (.Y(_09771_),
    .A(_09737_),
    .B(\cpu.dcache.r_tag[2][11] ));
 sg13g2_nand3_1 _16522_ (.B(net1062),
    .C(\cpu.dcache.r_tag[7][11] ),
    .A(net1068),
    .Y(_09772_));
 sg13g2_o21ai_1 _16523_ (.B1(_09772_),
    .Y(_09773_),
    .A1(net1068),
    .A2(_09771_));
 sg13g2_and2_1 _16524_ (.A(net1140),
    .B(\cpu.dcache.r_tag[1][11] ),
    .X(_09774_));
 sg13g2_and2_1 _16525_ (.A(_09427_),
    .B(\cpu.dcache.r_tag[4][11] ),
    .X(_09775_));
 sg13g2_and2_1 _16526_ (.A(net1140),
    .B(\cpu.dcache.r_tag[3][11] ),
    .X(_09776_));
 sg13g2_and2_1 _16527_ (.A(_09427_),
    .B(\cpu.dcache.r_tag[6][11] ),
    .X(_09777_));
 sg13g2_mux4_1 _16528_ (.S0(_09459_),
    .A0(_09774_),
    .A1(_09775_),
    .A2(_09776_),
    .A3(_09777_),
    .S1(net1072),
    .X(_09778_));
 sg13g2_a221oi_1 _16529_ (.B2(net919),
    .C1(_09778_),
    .B1(_09773_),
    .A1(\cpu.dcache.r_tag[5][11] ),
    .Y(_09779_),
    .A2(_09488_));
 sg13g2_mux2_1 _16530_ (.A0(_00244_),
    .A1(_09779_),
    .S(_09515_),
    .X(_09780_));
 sg13g2_xor2_1 _16531_ (.B(_09780_),
    .A(_00243_),
    .X(_09781_));
 sg13g2_mux2_1 _16532_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(\cpu.dcache.r_tag[3][10] ),
    .S(net1068),
    .X(_09782_));
 sg13g2_mux2_1 _16533_ (.A0(\cpu.dcache.r_tag[4][10] ),
    .A1(\cpu.dcache.r_tag[6][10] ),
    .S(net1146),
    .X(_09783_));
 sg13g2_nor2b_1 _16534_ (.A(net1063),
    .B_N(\cpu.dcache.r_tag[5][10] ),
    .Y(_09784_));
 sg13g2_mux2_1 _16535_ (.A0(_09783_),
    .A1(_09784_),
    .S(net1068),
    .X(_09785_));
 sg13g2_inv_1 _16536_ (.Y(_09786_),
    .A(\cpu.dcache.r_tag[1][10] ));
 sg13g2_nand3b_1 _16537_ (.B(net1140),
    .C(_09233_),
    .Y(_09787_),
    .A_N(net1146));
 sg13g2_buf_1 _16538_ (.A(_09787_),
    .X(_09788_));
 sg13g2_nand4_1 _16539_ (.B(net1062),
    .C(net1072),
    .A(net1068),
    .Y(_09789_),
    .D(\cpu.dcache.r_tag[7][10] ));
 sg13g2_o21ai_1 _16540_ (.B1(_09789_),
    .Y(_09790_),
    .A1(_09786_),
    .A2(_09788_));
 sg13g2_a221oi_1 _16541_ (.B2(net1062),
    .C1(_09790_),
    .B1(_09785_),
    .A1(_09754_),
    .Y(_09791_),
    .A2(_09782_));
 sg13g2_mux2_1 _16542_ (.A0(_00242_),
    .A1(_09791_),
    .S(_09515_),
    .X(_09792_));
 sg13g2_xor2_1 _16543_ (.B(_09792_),
    .A(_00241_),
    .X(_09793_));
 sg13g2_inv_1 _16544_ (.Y(_09794_),
    .A(_09433_));
 sg13g2_mux2_1 _16545_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(\cpu.dcache.r_tag[3][7] ),
    .S(net1072),
    .X(_09795_));
 sg13g2_mux2_1 _16546_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(\cpu.dcache.r_tag[7][7] ),
    .S(net1063),
    .X(_09796_));
 sg13g2_nor2b_1 _16547_ (.A(net1063),
    .B_N(\cpu.dcache.r_tag[4][7] ),
    .Y(_09797_));
 sg13g2_mux2_1 _16548_ (.A0(_09796_),
    .A1(_09797_),
    .S(_09459_),
    .X(_09798_));
 sg13g2_a22oi_1 _16549_ (.Y(_09799_),
    .B1(\cpu.dcache.r_tag[2][7] ),
    .B2(_09737_),
    .A2(\cpu.dcache.r_tag[6][7] ),
    .A1(net1062));
 sg13g2_nor2b_1 _16550_ (.A(_09799_),
    .B_N(_09728_),
    .Y(_09800_));
 sg13g2_a221oi_1 _16551_ (.B2(_09524_),
    .C1(_09800_),
    .B1(_09798_),
    .A1(_09794_),
    .Y(_09801_),
    .A2(_09795_));
 sg13g2_mux2_1 _16552_ (.A0(_00236_),
    .A1(_09801_),
    .S(_09515_),
    .X(_09802_));
 sg13g2_xor2_1 _16553_ (.B(_09802_),
    .A(_00235_),
    .X(_09803_));
 sg13g2_nor2b_1 _16554_ (.A(_09449_),
    .B_N(net1068),
    .Y(_09804_));
 sg13g2_buf_2 _16555_ (.A(_09804_),
    .X(_09805_));
 sg13g2_a22oi_1 _16556_ (.Y(_09806_),
    .B1(_09805_),
    .B2(\cpu.dcache.r_tag[5][6] ),
    .A2(_09444_),
    .A1(\cpu.dcache.r_tag[6][6] ));
 sg13g2_nand2_1 _16557_ (.Y(_09807_),
    .A(net1140),
    .B(\cpu.dcache.r_tag[2][6] ));
 sg13g2_nand2_1 _16558_ (.Y(_09808_),
    .A(net1062),
    .B(\cpu.dcache.r_tag[4][6] ));
 sg13g2_a22oi_1 _16559_ (.Y(_09809_),
    .B1(\cpu.dcache.r_tag[3][6] ),
    .B2(net1140),
    .A2(\cpu.dcache.r_tag[7][6] ),
    .A1(net1062));
 sg13g2_nand2_1 _16560_ (.Y(_09810_),
    .A(net1140),
    .B(\cpu.dcache.r_tag[1][6] ));
 sg13g2_mux4_1 _16561_ (.S0(net915),
    .A0(_09807_),
    .A1(_09808_),
    .A2(_09809_),
    .A3(_09810_),
    .S1(net918),
    .X(_09811_));
 sg13g2_o21ai_1 _16562_ (.B1(_09811_),
    .Y(_09812_),
    .A1(net904),
    .A2(_09806_));
 sg13g2_nand2_1 _16563_ (.Y(_09813_),
    .A(_00234_),
    .B(_09437_));
 sg13g2_o21ai_1 _16564_ (.B1(_09813_),
    .Y(_09814_),
    .A1(_09438_),
    .A2(_09812_));
 sg13g2_xor2_1 _16565_ (.B(_09814_),
    .A(_00233_),
    .X(_09815_));
 sg13g2_nor4_1 _16566_ (.A(_09781_),
    .B(_09793_),
    .C(_09803_),
    .D(_09815_),
    .Y(_09816_));
 sg13g2_nand4_1 _16567_ (.B(_09733_),
    .C(_09770_),
    .A(_09709_),
    .Y(_09817_),
    .D(_09816_));
 sg13g2_nor4_1 _16568_ (.A(_09551_),
    .B(_09618_),
    .C(_09666_),
    .D(_09817_),
    .Y(_09818_));
 sg13g2_mux4_1 _16569_ (.S0(net798),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net919),
    .X(_09819_));
 sg13g2_mux4_1 _16570_ (.S0(net918),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net919),
    .X(_09820_));
 sg13g2_mux2_1 _16571_ (.A0(_09819_),
    .A1(_09820_),
    .S(net904),
    .X(_09821_));
 sg13g2_mux4_1 _16572_ (.S0(_09236_),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(_09221_),
    .X(_09822_));
 sg13g2_mux4_1 _16573_ (.S0(net798),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net919),
    .X(_09823_));
 sg13g2_buf_1 _16574_ (.A(net904),
    .X(_09824_));
 sg13g2_mux2_1 _16575_ (.A0(_09822_),
    .A1(_09823_),
    .S(_09824_),
    .X(_09825_));
 sg13g2_nand3_1 _16576_ (.B(_09821_),
    .C(_09825_),
    .A(_09286_),
    .Y(_09826_));
 sg13g2_buf_1 _16577_ (.A(_09826_),
    .X(_09827_));
 sg13g2_a21oi_1 _16578_ (.A1(_09399_),
    .A2(_09818_),
    .Y(_09828_),
    .B1(_09827_));
 sg13g2_inv_1 _16579_ (.Y(_09829_),
    .A(_09827_));
 sg13g2_and2_1 _16580_ (.A(_09821_),
    .B(_09818_),
    .X(_09830_));
 sg13g2_buf_1 _16581_ (.A(_09830_),
    .X(_09831_));
 sg13g2_nor3_1 _16582_ (.A(_09398_),
    .B(_09829_),
    .C(_09831_),
    .Y(_09832_));
 sg13g2_buf_1 _16583_ (.A(_09832_),
    .X(_09833_));
 sg13g2_nand2b_1 _16584_ (.Y(_09834_),
    .B(_09286_),
    .A_N(_08350_));
 sg13g2_a21oi_1 _16585_ (.A1(_08354_),
    .A2(_08408_),
    .Y(_09835_),
    .B1(_09834_));
 sg13g2_o21ai_1 _16586_ (.B1(_09835_),
    .Y(_09836_),
    .A1(_09828_),
    .A2(_09833_));
 sg13g2_o21ai_1 _16587_ (.B1(_09836_),
    .Y(_09837_),
    .A1(_09397_),
    .A2(_08894_));
 sg13g2_nor2_1 _16588_ (.A(_09396_),
    .B(_09837_),
    .Y(_09838_));
 sg13g2_inv_1 _16589_ (.Y(_09839_),
    .A(_09838_));
 sg13g2_buf_1 _16590_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09840_));
 sg13g2_buf_1 _16591_ (.A(\cpu.qspi.r_ind ),
    .X(_09841_));
 sg13g2_buf_1 _16592_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09842_));
 sg13g2_buf_2 _16593_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09843_));
 sg13g2_nor4_2 _16594_ (.A(_09842_),
    .B(_09843_),
    .C(\cpu.qspi.r_count[3] ),
    .Y(_09844_),
    .D(\cpu.qspi.r_count[2] ));
 sg13g2_and2_1 _16595_ (.A(_00254_),
    .B(_09844_),
    .X(_09845_));
 sg13g2_buf_1 _16596_ (.A(_09845_),
    .X(_09846_));
 sg13g2_buf_1 _16597_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09847_));
 sg13g2_buf_1 _16598_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09848_));
 sg13g2_a221oi_1 _16599_ (.B2(_09847_),
    .C1(_09848_),
    .B1(_09846_),
    .A1(_09840_),
    .Y(_09849_),
    .A2(_09841_));
 sg13g2_a21oi_1 _16600_ (.A1(_09839_),
    .A2(_09849_),
    .Y(_00026_),
    .B1(net623));
 sg13g2_buf_1 _16601_ (.A(_09365_),
    .X(_09850_));
 sg13g2_buf_2 _16602_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09851_));
 sg13g2_nand2_1 _16603_ (.Y(_09852_),
    .A(_00254_),
    .B(_09844_));
 sg13g2_buf_1 _16604_ (.A(_09852_),
    .X(_09853_));
 sg13g2_and2_1 _16605_ (.A(_09397_),
    .B(_09828_),
    .X(_09854_));
 sg13g2_buf_1 _16606_ (.A(_09854_),
    .X(_09855_));
 sg13g2_buf_1 _16607_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09856_));
 sg13g2_a22oi_1 _16608_ (.Y(_09857_),
    .B1(net172),
    .B2(net1138),
    .A2(net773),
    .A1(_09851_));
 sg13g2_nor2_1 _16609_ (.A(net614),
    .B(_09857_),
    .Y(_00025_));
 sg13g2_buf_1 _16610_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09858_));
 sg13g2_buf_1 _16611_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09859_));
 sg13g2_a21oi_1 _16612_ (.A1(_09858_),
    .A2(_09846_),
    .Y(_09860_),
    .B1(_09859_));
 sg13g2_nor2_1 _16613_ (.A(net614),
    .B(_09860_),
    .Y(_00022_));
 sg13g2_buf_1 _16614_ (.A(_00279_),
    .X(_09861_));
 sg13g2_buf_1 _16615_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09862_));
 sg13g2_nand2_1 _16616_ (.Y(_09863_),
    .A(net1137),
    .B(net773));
 sg13g2_a21oi_1 _16617_ (.A1(_09861_),
    .A2(_09863_),
    .Y(_00023_),
    .B1(net623));
 sg13g2_buf_1 _16618_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09864_));
 sg13g2_buf_1 _16619_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09865_));
 sg13g2_buf_1 _16620_ (.A(_08310_),
    .X(_09866_));
 sg13g2_inv_1 _16621_ (.Y(_09867_),
    .A(_09426_));
 sg13g2_or2_1 _16622_ (.X(_09868_),
    .B(_08615_),
    .A(_09397_));
 sg13g2_o21ai_1 _16623_ (.B1(_09868_),
    .Y(_09869_),
    .A1(net1060),
    .A2(_09867_));
 sg13g2_nor2_1 _16624_ (.A(_09865_),
    .B(_09869_),
    .Y(_09870_));
 sg13g2_a21oi_1 _16625_ (.A1(_09865_),
    .A2(net172),
    .Y(_09871_),
    .B1(_09870_));
 sg13g2_and2_1 _16626_ (.A(_09864_),
    .B(_09871_),
    .X(_09872_));
 sg13g2_buf_8 _16627_ (.A(_09872_),
    .X(_09873_));
 sg13g2_inv_1 _16628_ (.Y(_09874_),
    .A(_09869_));
 sg13g2_nor3_1 _16629_ (.A(_09865_),
    .B(_09864_),
    .C(_09874_),
    .Y(_09875_));
 sg13g2_buf_2 _16630_ (.A(_09875_),
    .X(_09876_));
 sg13g2_nor2_1 _16631_ (.A(_09876_),
    .B(_09873_),
    .Y(_09877_));
 sg13g2_buf_2 _16632_ (.A(_09877_),
    .X(_09878_));
 sg13g2_and2_1 _16633_ (.A(\cpu.qspi.r_quad[2] ),
    .B(_09876_),
    .X(_09879_));
 sg13g2_a221oi_1 _16634_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09879_),
    .B1(_09878_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09880_),
    .A2(_09873_));
 sg13g2_buf_2 _16635_ (.A(_09880_),
    .X(_09881_));
 sg13g2_nand2_1 _16636_ (.Y(_09882_),
    .A(\cpu.qspi.r_state[17] ),
    .B(_09837_));
 sg13g2_inv_1 _16637_ (.Y(_09883_),
    .A(_09882_));
 sg13g2_a22oi_1 _16638_ (.Y(_09884_),
    .B1(_09881_),
    .B2(_09883_),
    .A2(net773),
    .A1(_09858_));
 sg13g2_nor2_1 _16639_ (.A(net614),
    .B(_09884_),
    .Y(_00028_));
 sg13g2_nand2_1 _16640_ (.Y(_09885_),
    .A(_09847_),
    .B(_09852_));
 sg13g2_buf_1 _16641_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09886_));
 sg13g2_nand2_1 _16642_ (.Y(_09887_),
    .A(net1136),
    .B(_09846_));
 sg13g2_a21oi_1 _16643_ (.A1(_09885_),
    .A2(_09887_),
    .Y(_00027_),
    .B1(net623));
 sg13g2_inv_1 _16644_ (.Y(_09888_),
    .A(_09841_));
 sg13g2_buf_1 _16645_ (.A(net795),
    .X(_09889_));
 sg13g2_a21o_1 _16646_ (.A2(_09888_),
    .A1(_09840_),
    .B1(_09889_),
    .X(_00021_));
 sg13g2_buf_1 _16647_ (.A(\cpu.dec.r_op[10] ),
    .X(_09890_));
 sg13g2_a21oi_1 _16648_ (.A1(net696),
    .A2(_09005_),
    .Y(_09891_),
    .B1(_09013_));
 sg13g2_buf_2 _16649_ (.A(_09891_),
    .X(_09892_));
 sg13g2_nand2_1 _16650_ (.Y(_09893_),
    .A(_09892_),
    .B(_09035_));
 sg13g2_nor3_1 _16651_ (.A(net141),
    .B(_08998_),
    .C(_09893_),
    .Y(_09894_));
 sg13g2_a21o_1 _16652_ (.A2(_08897_),
    .A1(net1135),
    .B1(_09894_),
    .X(_00011_));
 sg13g2_buf_1 _16653_ (.A(_09107_),
    .X(_09895_));
 sg13g2_nor2_1 _16654_ (.A(_09895_),
    .B(_09126_),
    .Y(_09896_));
 sg13g2_a21oi_1 _16655_ (.A1(net800),
    .A2(_08951_),
    .Y(_09897_),
    .B1(_08959_));
 sg13g2_buf_1 _16656_ (.A(_09897_),
    .X(_09898_));
 sg13g2_a21o_1 _16657_ (.A2(_08967_),
    .A1(_08920_),
    .B1(_08975_),
    .X(_09899_));
 sg13g2_buf_1 _16658_ (.A(_09899_),
    .X(_09900_));
 sg13g2_a21oi_2 _16659_ (.B1(_08991_),
    .Y(_09901_),
    .A2(_08984_),
    .A1(net696));
 sg13g2_nor2_2 _16660_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sg13g2_nand2_1 _16661_ (.Y(_09903_),
    .A(_09898_),
    .B(_09902_));
 sg13g2_buf_2 _16662_ (.A(_09903_),
    .X(_09904_));
 sg13g2_a21o_1 _16663_ (.A2(_09147_),
    .A1(net800),
    .B1(_09155_),
    .X(_09905_));
 sg13g2_buf_1 _16664_ (.A(_09905_),
    .X(_09906_));
 sg13g2_buf_1 _16665_ (.A(_09906_),
    .X(_09907_));
 sg13g2_nor2_1 _16666_ (.A(_09116_),
    .B(_09139_),
    .Y(_09908_));
 sg13g2_nand2_1 _16667_ (.Y(_09909_),
    .A(net272),
    .B(_09908_));
 sg13g2_a21o_1 _16668_ (.A2(_09166_),
    .A1(_09122_),
    .B1(_09173_),
    .X(_09910_));
 sg13g2_buf_2 _16669_ (.A(_09910_),
    .X(_09911_));
 sg13g2_buf_1 _16670_ (.A(_09191_),
    .X(_09912_));
 sg13g2_nand3_1 _16671_ (.B(_09911_),
    .C(net271),
    .A(net194),
    .Y(_09913_));
 sg13g2_nor3_1 _16672_ (.A(_09904_),
    .B(_09909_),
    .C(_09913_),
    .Y(_09914_));
 sg13g2_a21oi_1 _16673_ (.A1(_09118_),
    .A2(_09896_),
    .Y(_09915_),
    .B1(_09914_));
 sg13g2_buf_1 _16674_ (.A(\cpu.dec.r_op[1] ),
    .X(_09916_));
 sg13g2_nand2_1 _16675_ (.Y(_09917_),
    .A(_09916_),
    .B(net140));
 sg13g2_o21ai_1 _16676_ (.B1(_09917_),
    .Y(_00012_),
    .A1(net107),
    .A2(_09915_));
 sg13g2_nand2_1 _16677_ (.Y(_09918_),
    .A(net345),
    .B(_09035_));
 sg13g2_nor2_1 _16678_ (.A(_09114_),
    .B(_09918_),
    .Y(_09919_));
 sg13g2_a21oi_1 _16679_ (.A1(_09135_),
    .A2(_09896_),
    .Y(_09920_),
    .B1(_09919_));
 sg13g2_buf_1 _16680_ (.A(\cpu.dec.r_op[9] ),
    .X(_09921_));
 sg13g2_buf_1 _16681_ (.A(net1134),
    .X(_09922_));
 sg13g2_nand2_1 _16682_ (.Y(_09923_),
    .A(net1059),
    .B(net140));
 sg13g2_o21ai_1 _16683_ (.B1(_09923_),
    .Y(_00020_),
    .A1(net107),
    .A2(_09920_));
 sg13g2_buf_2 _16684_ (.A(\cpu.dec.r_op[8] ),
    .X(_09924_));
 sg13g2_inv_1 _16685_ (.Y(_09925_),
    .A(_09924_));
 sg13g2_buf_1 _16686_ (.A(_09925_),
    .X(_09926_));
 sg13g2_nor2_1 _16687_ (.A(_09898_),
    .B(_08994_),
    .Y(_09927_));
 sg13g2_buf_2 _16688_ (.A(_09927_),
    .X(_09928_));
 sg13g2_a21oi_1 _16689_ (.A1(_09122_),
    .A2(_08929_),
    .Y(_09929_),
    .B1(_08939_));
 sg13g2_buf_1 _16690_ (.A(_09929_),
    .X(_09930_));
 sg13g2_nor2_2 _16691_ (.A(_09111_),
    .B(net270),
    .Y(_09931_));
 sg13g2_nand3_1 _16692_ (.B(_09928_),
    .C(_09931_),
    .A(net142),
    .Y(_09932_));
 sg13g2_o21ai_1 _16693_ (.B1(_09932_),
    .Y(_00019_),
    .A1(net903),
    .A2(net108));
 sg13g2_buf_2 _16694_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09933_));
 sg13g2_inv_1 _16695_ (.Y(_09934_),
    .A(_09933_));
 sg13g2_nand2_1 _16696_ (.Y(_09935_),
    .A(net1136),
    .B(net773));
 sg13g2_a21oi_1 _16697_ (.A1(_09934_),
    .A2(_09935_),
    .Y(_00024_),
    .B1(net623));
 sg13g2_nor2_1 _16698_ (.A(net389),
    .B(_09126_),
    .Y(_09936_));
 sg13g2_nand2b_1 _16699_ (.Y(_09937_),
    .B(net342),
    .A_N(_09191_));
 sg13g2_inv_1 _16700_ (.Y(_09938_),
    .A(_09937_));
 sg13g2_nor2_1 _16701_ (.A(_09114_),
    .B(_09909_),
    .Y(_09939_));
 sg13g2_a22oi_1 _16702_ (.Y(_09940_),
    .B1(_09938_),
    .B2(_09939_),
    .A2(_09936_),
    .A1(_09118_));
 sg13g2_buf_1 _16703_ (.A(net174),
    .X(_09941_));
 sg13g2_nand2_1 _16704_ (.Y(_09942_),
    .A(\cpu.dec.r_op[7] ),
    .B(net138));
 sg13g2_o21ai_1 _16705_ (.B1(_09942_),
    .Y(_00018_),
    .A1(_09121_),
    .A2(_09940_));
 sg13g2_buf_1 _16706_ (.A(\cpu.uart.r_div[11] ),
    .X(_09943_));
 sg13g2_nor3_1 _16707_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09944_));
 sg13g2_nor2b_1 _16708_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09944_),
    .Y(_09945_));
 sg13g2_nor2b_1 _16709_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09945_),
    .Y(_09946_));
 sg13g2_nor2b_1 _16710_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09946_),
    .Y(_09947_));
 sg13g2_nor2b_1 _16711_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09947_),
    .Y(_09948_));
 sg13g2_nand2b_1 _16712_ (.Y(_09949_),
    .B(_09948_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16713_ (.A(\cpu.uart.r_div[8] ),
    .B(_09949_),
    .Y(_09950_));
 sg13g2_nand2b_1 _16714_ (.Y(_09951_),
    .B(_09950_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16715_ (.A(_09951_),
    .X(_09952_));
 sg13g2_nor3_1 _16716_ (.A(_09943_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09952_),
    .Y(_09953_));
 sg13g2_buf_2 _16717_ (.A(_09953_),
    .X(_09954_));
 sg13g2_nor2_1 _16718_ (.A(net917),
    .B(_09954_),
    .Y(_09955_));
 sg13g2_buf_1 _16719_ (.A(_09955_),
    .X(_09956_));
 sg13g2_buf_1 _16720_ (.A(net229),
    .X(_09957_));
 sg13g2_mux2_1 _16721_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00281_),
    .S(net209),
    .X(_00079_));
 sg13g2_xnor2_1 _16722_ (.Y(_09958_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16723_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09958_),
    .S(_09957_),
    .X(_00082_));
 sg13g2_o21ai_1 _16724_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09959_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16725_ (.A(_09944_),
    .B_N(_09959_),
    .Y(_09960_));
 sg13g2_nor2_1 _16726_ (.A(\cpu.uart.r_div_value[2] ),
    .B(_09956_),
    .Y(_09961_));
 sg13g2_a21oi_1 _16727_ (.A1(net209),
    .A2(_09960_),
    .Y(_00083_),
    .B1(_09961_));
 sg13g2_xnor2_1 _16728_ (.Y(_09962_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09944_));
 sg13g2_nor2_1 _16729_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net229),
    .Y(_09963_));
 sg13g2_a21oi_1 _16730_ (.A1(net209),
    .A2(_09962_),
    .Y(_00084_),
    .B1(_09963_));
 sg13g2_xnor2_1 _16731_ (.Y(_09964_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09945_));
 sg13g2_nor2_1 _16732_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net229),
    .Y(_09965_));
 sg13g2_a21oi_1 _16733_ (.A1(net209),
    .A2(_09964_),
    .Y(_00085_),
    .B1(_09965_));
 sg13g2_xnor2_1 _16734_ (.Y(_09966_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09946_));
 sg13g2_nor2_1 _16735_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net229),
    .Y(_09967_));
 sg13g2_a21oi_1 _16736_ (.A1(net209),
    .A2(_09966_),
    .Y(_00086_),
    .B1(_09967_));
 sg13g2_xnor2_1 _16737_ (.Y(_09968_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09947_));
 sg13g2_nor2_1 _16738_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net229),
    .Y(_09969_));
 sg13g2_a21oi_1 _16739_ (.A1(_09957_),
    .A2(_09968_),
    .Y(_00087_),
    .B1(_09969_));
 sg13g2_xnor2_1 _16740_ (.Y(_09970_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09948_));
 sg13g2_nor2_1 _16741_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net229),
    .Y(_09971_));
 sg13g2_a21oi_1 _16742_ (.A1(net209),
    .A2(_09970_),
    .Y(_00088_),
    .B1(_09971_));
 sg13g2_xor2_1 _16743_ (.B(_09949_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09972_));
 sg13g2_nor2_1 _16744_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net229),
    .Y(_09973_));
 sg13g2_a21oi_1 _16745_ (.A1(net209),
    .A2(_09972_),
    .Y(_00089_),
    .B1(_09973_));
 sg13g2_xnor2_1 _16746_ (.Y(_09974_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09950_));
 sg13g2_nor2_1 _16747_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net229),
    .Y(_09975_));
 sg13g2_a21oi_1 _16748_ (.A1(net209),
    .A2(_09974_),
    .Y(_00090_),
    .B1(_09975_));
 sg13g2_buf_1 _16749_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09976_));
 sg13g2_inv_1 _16750_ (.Y(_09977_),
    .A(_09976_));
 sg13g2_nand2_1 _16751_ (.Y(_09978_),
    .A(net916),
    .B(_09952_));
 sg13g2_o21ai_1 _16752_ (.B1(_09978_),
    .Y(_09979_),
    .A1(_09943_),
    .A2(_09976_));
 sg13g2_inv_1 _16753_ (.Y(_09980_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16754_ (.A(_09980_),
    .B(net795),
    .C(_09952_),
    .Y(_09981_));
 sg13g2_a221oi_1 _16755_ (.B2(_09980_),
    .C1(_09981_),
    .B1(_09979_),
    .A1(_09977_),
    .Y(_00080_),
    .A2(net691));
 sg13g2_nor2_1 _16756_ (.A(\cpu.uart.r_div[10] ),
    .B(_09952_),
    .Y(_09982_));
 sg13g2_nand2_1 _16757_ (.Y(_09983_),
    .A(_09943_),
    .B(net797));
 sg13g2_o21ai_1 _16758_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09984_),
    .A1(net795),
    .A2(_09954_));
 sg13g2_o21ai_1 _16759_ (.B1(_09984_),
    .Y(_00081_),
    .A1(_09982_),
    .A2(_09983_));
 sg13g2_inv_1 _16760_ (.Y(_09985_),
    .A(_00287_));
 sg13g2_buf_1 _16761_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09986_));
 sg13g2_buf_1 _16762_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09987_));
 sg13g2_buf_1 _16763_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09988_));
 sg13g2_buf_1 _16764_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09989_));
 sg13g2_buf_1 _16765_ (.A(\cpu.intr.r_timer_count[10] ),
    .X(_09990_));
 sg13g2_buf_1 _16766_ (.A(\cpu.intr.r_timer_count[7] ),
    .X(_09991_));
 sg13g2_buf_2 _16767_ (.A(\cpu.intr.r_timer_count[6] ),
    .X(_09992_));
 sg13g2_buf_2 _16768_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09993_));
 sg13g2_buf_2 _16769_ (.A(\cpu.intr.r_timer_count[0] ),
    .X(_09994_));
 sg13g2_buf_1 _16770_ (.A(\cpu.intr.r_timer_count[2] ),
    .X(_09995_));
 sg13g2_nor4_1 _16771_ (.A(_09993_),
    .B(_09994_),
    .C(\cpu.intr.r_timer_count[3] ),
    .D(_09995_),
    .Y(_09996_));
 sg13g2_nor2b_1 _16772_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09996_),
    .Y(_09997_));
 sg13g2_nor2b_1 _16773_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09997_),
    .Y(_09998_));
 sg13g2_inv_1 _16774_ (.Y(_09999_),
    .A(_09998_));
 sg13g2_nor4_2 _16775_ (.A(_09991_),
    .B(_09992_),
    .C(\cpu.intr.r_timer_count[8] ),
    .Y(_10000_),
    .D(_09999_));
 sg13g2_nand2b_1 _16776_ (.Y(_10001_),
    .B(_10000_),
    .A_N(\cpu.intr.r_timer_count[9] ));
 sg13g2_nor3_1 _16777_ (.A(\cpu.intr.r_timer_count[11] ),
    .B(_09990_),
    .C(_10001_),
    .Y(_10002_));
 sg13g2_nor2b_1 _16778_ (.A(\cpu.intr.r_timer_count[12] ),
    .B_N(_10002_),
    .Y(_10003_));
 sg13g2_nor2b_1 _16779_ (.A(\cpu.intr.r_timer_count[13] ),
    .B_N(_10003_),
    .Y(_10004_));
 sg13g2_nor2b_1 _16780_ (.A(\cpu.intr.r_timer_count[14] ),
    .B_N(_10004_),
    .Y(_10005_));
 sg13g2_nand2b_1 _16781_ (.Y(_10006_),
    .B(_10005_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_nor3_1 _16782_ (.A(_09988_),
    .B(_09989_),
    .C(_10006_),
    .Y(_10007_));
 sg13g2_nor2b_1 _16783_ (.A(_09987_),
    .B_N(_10007_),
    .Y(_10008_));
 sg13g2_nand2b_1 _16784_ (.Y(_10009_),
    .B(_10008_),
    .A_N(_09986_));
 sg13g2_buf_1 _16785_ (.A(_10009_),
    .X(_10010_));
 sg13g2_buf_2 _16786_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_10011_));
 sg13g2_buf_1 _16787_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_10012_));
 sg13g2_buf_1 _16788_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_10013_));
 sg13g2_buf_1 _16789_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_10014_));
 sg13g2_nor4_2 _16790_ (.A(_10011_),
    .B(_10012_),
    .C(_10013_),
    .Y(_10015_),
    .D(_10014_));
 sg13g2_nand2b_1 _16791_ (.Y(_10016_),
    .B(_10015_),
    .A_N(_10010_));
 sg13g2_buf_2 _16792_ (.A(_10016_),
    .X(_10017_));
 sg13g2_buf_1 _16793_ (.A(net1067),
    .X(_10018_));
 sg13g2_buf_1 _16794_ (.A(net902),
    .X(_10019_));
 sg13g2_buf_1 _16795_ (.A(net772),
    .X(_10020_));
 sg13g2_buf_1 _16796_ (.A(net681),
    .X(_10021_));
 sg13g2_buf_1 _16797_ (.A(net786),
    .X(_10022_));
 sg13g2_buf_1 _16798_ (.A(net680),
    .X(_10023_));
 sg13g2_buf_1 _16799_ (.A(net612),
    .X(_10024_));
 sg13g2_buf_1 _16800_ (.A(net545),
    .X(_10025_));
 sg13g2_buf_1 _16801_ (.A(\cpu.addr[5] ),
    .X(_10026_));
 sg13g2_buf_1 _16802_ (.A(_10026_),
    .X(_10027_));
 sg13g2_nor3_2 _16803_ (.A(_10027_),
    .B(net1070),
    .C(_09228_),
    .Y(_10028_));
 sg13g2_nand2_1 _16804_ (.Y(_10029_),
    .A(net1071),
    .B(_10028_));
 sg13g2_buf_1 _16805_ (.A(_10029_),
    .X(_10030_));
 sg13g2_nor2_1 _16806_ (.A(_09292_),
    .B(net679),
    .Y(_10031_));
 sg13g2_buf_1 _16807_ (.A(_10031_),
    .X(_10032_));
 sg13g2_nand3_1 _16808_ (.B(net485),
    .C(net193),
    .A(net613),
    .Y(_10033_));
 sg13g2_buf_1 _16809_ (.A(_10033_),
    .X(_10034_));
 sg13g2_nand2_1 _16810_ (.Y(_10035_),
    .A(_10017_),
    .B(_10034_));
 sg13g2_buf_8 _16811_ (.A(_10035_),
    .X(_10036_));
 sg13g2_buf_8 _16812_ (.A(_10036_),
    .X(_10037_));
 sg13g2_buf_8 _16813_ (.A(_10036_),
    .X(_10038_));
 sg13g2_nand2_1 _16814_ (.Y(_10039_),
    .A(\cpu.intr.r_timer_reload[0] ),
    .B(net67));
 sg13g2_o21ai_1 _16815_ (.B1(_10039_),
    .Y(_00055_),
    .A1(_09985_),
    .A2(net68));
 sg13g2_xor2_1 _16816_ (.B(_09994_),
    .A(_09993_),
    .X(_10040_));
 sg13g2_nand2_1 _16817_ (.Y(_10041_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net67));
 sg13g2_o21ai_1 _16818_ (.B1(_10041_),
    .Y(_00066_),
    .A1(net68),
    .A2(_10040_));
 sg13g2_nor3_1 _16819_ (.A(_09993_),
    .B(_09994_),
    .C(_09995_),
    .Y(_10042_));
 sg13g2_o21ai_1 _16820_ (.B1(_09995_),
    .Y(_10043_),
    .A1(_09993_),
    .A2(_09994_));
 sg13g2_nor2b_1 _16821_ (.A(_10042_),
    .B_N(_10043_),
    .Y(_10044_));
 sg13g2_nand2_1 _16822_ (.Y(_10045_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net67));
 sg13g2_o21ai_1 _16823_ (.B1(_10045_),
    .Y(_00071_),
    .A1(net68),
    .A2(_10044_));
 sg13g2_xnor2_1 _16824_ (.Y(_10046_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_10042_));
 sg13g2_nand2_1 _16825_ (.Y(_10047_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(net67));
 sg13g2_o21ai_1 _16826_ (.B1(_10047_),
    .Y(_00072_),
    .A1(net68),
    .A2(_10046_));
 sg13g2_xnor2_1 _16827_ (.Y(_10048_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09996_));
 sg13g2_buf_8 _16828_ (.A(_10036_),
    .X(_10049_));
 sg13g2_nand2_1 _16829_ (.Y(_10050_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(net66));
 sg13g2_o21ai_1 _16830_ (.B1(_10050_),
    .Y(_00073_),
    .A1(net68),
    .A2(_10048_));
 sg13g2_xnor2_1 _16831_ (.Y(_10051_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09997_));
 sg13g2_nand2_1 _16832_ (.Y(_10052_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(net66));
 sg13g2_o21ai_1 _16833_ (.B1(_10052_),
    .Y(_00074_),
    .A1(net68),
    .A2(_10051_));
 sg13g2_xnor2_1 _16834_ (.Y(_10053_),
    .A(_09992_),
    .B(_09998_));
 sg13g2_nand2_1 _16835_ (.Y(_10054_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(net66));
 sg13g2_o21ai_1 _16836_ (.B1(_10054_),
    .Y(_00075_),
    .A1(_10037_),
    .A2(_10053_));
 sg13g2_nor2_1 _16837_ (.A(_09992_),
    .B(_09999_),
    .Y(_10055_));
 sg13g2_xnor2_1 _16838_ (.Y(_10056_),
    .A(_09991_),
    .B(_10055_));
 sg13g2_nand2_1 _16839_ (.Y(_10057_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(net66));
 sg13g2_o21ai_1 _16840_ (.B1(_10057_),
    .Y(_00076_),
    .A1(net68),
    .A2(_10056_));
 sg13g2_nor3_1 _16841_ (.A(_09991_),
    .B(_09992_),
    .C(_09999_),
    .Y(_10058_));
 sg13g2_xnor2_1 _16842_ (.Y(_10059_),
    .A(\cpu.intr.r_timer_count[8] ),
    .B(_10058_));
 sg13g2_nand2_1 _16843_ (.Y(_10060_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(_10049_));
 sg13g2_o21ai_1 _16844_ (.B1(_10060_),
    .Y(_00077_),
    .A1(_10037_),
    .A2(_10059_));
 sg13g2_xnor2_1 _16845_ (.Y(_10061_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(_10000_));
 sg13g2_nand2_1 _16846_ (.Y(_10062_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net66));
 sg13g2_o21ai_1 _16847_ (.B1(_10062_),
    .Y(_00078_),
    .A1(net68),
    .A2(_10061_));
 sg13g2_xor2_1 _16848_ (.B(_10001_),
    .A(_09990_),
    .X(_10063_));
 sg13g2_nand2_1 _16849_ (.Y(_10064_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net66));
 sg13g2_o21ai_1 _16850_ (.B1(_10064_),
    .Y(_00056_),
    .A1(net67),
    .A2(_10063_));
 sg13g2_o21ai_1 _16851_ (.B1(\cpu.intr.r_timer_count[11] ),
    .Y(_10065_),
    .A1(_09990_),
    .A2(_10001_));
 sg13g2_nor2b_1 _16852_ (.A(_10002_),
    .B_N(_10065_),
    .Y(_10066_));
 sg13g2_nand2_1 _16853_ (.Y(_10067_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net66));
 sg13g2_o21ai_1 _16854_ (.B1(_10067_),
    .Y(_00057_),
    .A1(net67),
    .A2(_10066_));
 sg13g2_xnor2_1 _16855_ (.Y(_10068_),
    .A(\cpu.intr.r_timer_count[12] ),
    .B(_10002_));
 sg13g2_nand2_1 _16856_ (.Y(_10069_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(_10049_));
 sg13g2_o21ai_1 _16857_ (.B1(_10069_),
    .Y(_00058_),
    .A1(net67),
    .A2(_10068_));
 sg13g2_xnor2_1 _16858_ (.Y(_10070_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_10003_));
 sg13g2_nand2_1 _16859_ (.Y(_10071_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net66));
 sg13g2_o21ai_1 _16860_ (.B1(_10071_),
    .Y(_00059_),
    .A1(net67),
    .A2(_10070_));
 sg13g2_xnor2_1 _16861_ (.Y(_10072_),
    .A(\cpu.intr.r_timer_count[14] ),
    .B(_10004_));
 sg13g2_nand2_1 _16862_ (.Y(_10073_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(_10036_));
 sg13g2_o21ai_1 _16863_ (.B1(_10073_),
    .Y(_00060_),
    .A1(_10038_),
    .A2(_10072_));
 sg13g2_xnor2_1 _16864_ (.Y(_10074_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_10005_));
 sg13g2_nand2_1 _16865_ (.Y(_10075_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_10036_));
 sg13g2_o21ai_1 _16866_ (.B1(_10075_),
    .Y(_00061_),
    .A1(_10038_),
    .A2(_10074_));
 sg13g2_nor4_1 _16867_ (.A(_09988_),
    .B(_09987_),
    .C(_09986_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_10076_));
 sg13g2_or2_1 _16868_ (.X(_10077_),
    .B(_10006_),
    .A(_09989_));
 sg13g2_a21oi_1 _16869_ (.A1(_10015_),
    .A2(_10076_),
    .Y(_10078_),
    .B1(_10077_));
 sg13g2_a21oi_1 _16870_ (.A1(_09989_),
    .A2(_10006_),
    .Y(_10079_),
    .B1(_10078_));
 sg13g2_buf_1 _16871_ (.A(\cpu.dcache.wdata[0] ),
    .X(_10080_));
 sg13g2_buf_1 _16872_ (.A(_10080_),
    .X(_10081_));
 sg13g2_buf_1 _16873_ (.A(net1057),
    .X(_10082_));
 sg13g2_nor2_1 _16874_ (.A(net901),
    .B(net137),
    .Y(_10083_));
 sg13g2_a21oi_1 _16875_ (.A1(net137),
    .A2(_10079_),
    .Y(_00062_),
    .B1(_10083_));
 sg13g2_nor2_1 _16876_ (.A(\cpu.intr.r_timer_reload[17] ),
    .B(_10017_),
    .Y(_10084_));
 sg13g2_and2_1 _16877_ (.A(_09988_),
    .B(_10077_),
    .X(_10085_));
 sg13g2_o21ai_1 _16878_ (.B1(net137),
    .Y(_10086_),
    .A1(_10007_),
    .A2(_10085_));
 sg13g2_buf_1 _16879_ (.A(\cpu.dcache.wdata[1] ),
    .X(_10087_));
 sg13g2_buf_1 _16880_ (.A(_10087_),
    .X(_10088_));
 sg13g2_inv_2 _16881_ (.Y(_10089_),
    .A(_09238_));
 sg13g2_buf_1 _16882_ (.A(_10089_),
    .X(_10090_));
 sg13g2_buf_1 _16883_ (.A(net900),
    .X(_10091_));
 sg13g2_buf_1 _16884_ (.A(net771),
    .X(_10092_));
 sg13g2_buf_1 _16885_ (.A(net678),
    .X(_10093_));
 sg13g2_buf_1 _16886_ (.A(net611),
    .X(_10094_));
 sg13g2_nor2_2 _16887_ (.A(_09460_),
    .B(net915),
    .Y(_10095_));
 sg13g2_nand2_1 _16888_ (.Y(_10096_),
    .A(net909),
    .B(_10095_));
 sg13g2_buf_2 _16889_ (.A(_10096_),
    .X(_10097_));
 sg13g2_nor4_1 _16890_ (.A(net544),
    .B(_09292_),
    .C(_10097_),
    .D(net679),
    .Y(_10098_));
 sg13g2_buf_1 _16891_ (.A(_10098_),
    .X(_10099_));
 sg13g2_buf_1 _16892_ (.A(_10099_),
    .X(_10100_));
 sg13g2_nand2_1 _16893_ (.Y(_10101_),
    .A(net1056),
    .B(net171));
 sg13g2_o21ai_1 _16894_ (.B1(_10101_),
    .Y(_00063_),
    .A1(_10084_),
    .A2(_10086_));
 sg13g2_nor2_1 _16895_ (.A(\cpu.intr.r_timer_reload[18] ),
    .B(_10017_),
    .Y(_10102_));
 sg13g2_nor2b_1 _16896_ (.A(_10007_),
    .B_N(_09987_),
    .Y(_10103_));
 sg13g2_o21ai_1 _16897_ (.B1(net137),
    .Y(_10104_),
    .A1(_10008_),
    .A2(_10103_));
 sg13g2_buf_1 _16898_ (.A(\cpu.dcache.wdata[2] ),
    .X(_10105_));
 sg13g2_buf_1 _16899_ (.A(_10105_),
    .X(_10106_));
 sg13g2_nand2_1 _16900_ (.Y(_10107_),
    .A(_10106_),
    .B(_10099_));
 sg13g2_o21ai_1 _16901_ (.B1(_10107_),
    .Y(_00064_),
    .A1(_10102_),
    .A2(_10104_));
 sg13g2_xor2_1 _16902_ (.B(_10008_),
    .A(_09986_),
    .X(_10108_));
 sg13g2_o21ai_1 _16903_ (.B1(_10108_),
    .Y(_10109_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_10017_));
 sg13g2_buf_1 _16904_ (.A(\cpu.dcache.wdata[3] ),
    .X(_10110_));
 sg13g2_buf_1 _16905_ (.A(net1133),
    .X(_10111_));
 sg13g2_nand2_1 _16906_ (.Y(_10112_),
    .A(net1054),
    .B(_10099_));
 sg13g2_o21ai_1 _16907_ (.B1(_10112_),
    .Y(_00065_),
    .A1(net171),
    .A2(_10109_));
 sg13g2_nor2b_1 _16908_ (.A(\cpu.intr.r_timer_reload[20] ),
    .B_N(_10015_),
    .Y(_10113_));
 sg13g2_nor3_1 _16909_ (.A(_10011_),
    .B(_10010_),
    .C(_10113_),
    .Y(_10114_));
 sg13g2_a21oi_1 _16910_ (.A1(_10011_),
    .A2(_10010_),
    .Y(_10115_),
    .B1(_10114_));
 sg13g2_buf_2 _16911_ (.A(\cpu.dcache.wdata[4] ),
    .X(_10116_));
 sg13g2_buf_1 _16912_ (.A(_10116_),
    .X(_10117_));
 sg13g2_nor2_1 _16913_ (.A(net1053),
    .B(net137),
    .Y(_10118_));
 sg13g2_a21oi_1 _16914_ (.A1(net137),
    .A2(_10115_),
    .Y(_00067_),
    .B1(_10118_));
 sg13g2_nor2_1 _16915_ (.A(_10011_),
    .B(_10010_),
    .Y(_10119_));
 sg13g2_xnor2_1 _16916_ (.Y(_10120_),
    .A(_10012_),
    .B(_10119_));
 sg13g2_o21ai_1 _16917_ (.B1(net137),
    .Y(_10121_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_10017_));
 sg13g2_buf_2 _16918_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10122_));
 sg13g2_buf_1 _16919_ (.A(_10122_),
    .X(_10123_));
 sg13g2_nand2_1 _16920_ (.Y(_10124_),
    .A(_10123_),
    .B(_10099_));
 sg13g2_o21ai_1 _16921_ (.B1(_10124_),
    .Y(_00068_),
    .A1(_10120_),
    .A2(_10121_));
 sg13g2_nor3_1 _16922_ (.A(_10011_),
    .B(_10012_),
    .C(_10010_),
    .Y(_10125_));
 sg13g2_xnor2_1 _16923_ (.Y(_10126_),
    .A(_10013_),
    .B(_10125_));
 sg13g2_o21ai_1 _16924_ (.B1(net137),
    .Y(_10127_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_10017_));
 sg13g2_buf_2 _16925_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10128_));
 sg13g2_buf_1 _16926_ (.A(_10128_),
    .X(_10129_));
 sg13g2_nand2_1 _16927_ (.Y(_10130_),
    .A(net1051),
    .B(_10099_));
 sg13g2_o21ai_1 _16928_ (.B1(_10130_),
    .Y(_00069_),
    .A1(_10126_),
    .A2(_10127_));
 sg13g2_buf_2 _16929_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10131_));
 sg13g2_buf_1 _16930_ (.A(_10131_),
    .X(_10132_));
 sg13g2_buf_1 _16931_ (.A(net1050),
    .X(_10133_));
 sg13g2_nor2b_1 _16932_ (.A(_10014_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_10134_));
 sg13g2_nor2b_1 _16933_ (.A(_10013_),
    .B_N(_10125_),
    .Y(_10135_));
 sg13g2_mux2_1 _16934_ (.A0(_10014_),
    .A1(_10134_),
    .S(_10135_),
    .X(_10136_));
 sg13g2_mux2_1 _16935_ (.A0(net899),
    .A1(_10136_),
    .S(_10034_),
    .X(_00070_));
 sg13g2_buf_2 _16936_ (.A(net613),
    .X(_10137_));
 sg13g2_nor2b_1 _16937_ (.A(net543),
    .B_N(net1057),
    .Y(_10138_));
 sg13g2_nand2_1 _16938_ (.Y(_10139_),
    .A(net915),
    .B(_09451_));
 sg13g2_buf_1 _16939_ (.A(_10139_),
    .X(_10140_));
 sg13g2_nor3_1 _16940_ (.A(_09292_),
    .B(_10140_),
    .C(net679),
    .Y(_10141_));
 sg13g2_buf_1 _16941_ (.A(_10141_),
    .X(_10142_));
 sg13g2_buf_1 _16942_ (.A(net192),
    .X(_10143_));
 sg13g2_mux2_1 _16943_ (.A0(_00288_),
    .A1(_10138_),
    .S(_10143_),
    .X(_00036_));
 sg13g2_buf_1 _16944_ (.A(_10087_),
    .X(_10144_));
 sg13g2_buf_1 _16945_ (.A(net1049),
    .X(_10145_));
 sg13g2_and2_1 _16946_ (.A(_10093_),
    .B(_10141_),
    .X(_10146_));
 sg13g2_buf_1 _16947_ (.A(_10146_),
    .X(_10147_));
 sg13g2_buf_1 _16948_ (.A(_10147_),
    .X(_10148_));
 sg13g2_buf_1 _16949_ (.A(net136),
    .X(_10149_));
 sg13g2_buf_1 _16950_ (.A(_10147_),
    .X(_10150_));
 sg13g2_nand2_1 _16951_ (.Y(_10151_),
    .A(net785),
    .B(_09238_));
 sg13g2_buf_1 _16952_ (.A(_10151_),
    .X(_10152_));
 sg13g2_buf_1 _16953_ (.A(_10152_),
    .X(_10153_));
 sg13g2_nor2_1 _16954_ (.A(_09463_),
    .B(net542),
    .Y(_10154_));
 sg13g2_buf_1 _16955_ (.A(_10154_),
    .X(_10155_));
 sg13g2_buf_1 _16956_ (.A(_10155_),
    .X(_10156_));
 sg13g2_and2_1 _16957_ (.A(_10032_),
    .B(net384),
    .X(_10157_));
 sg13g2_buf_1 _16958_ (.A(_10157_),
    .X(_10158_));
 sg13g2_buf_1 _16959_ (.A(net134),
    .X(_10159_));
 sg13g2_buf_2 _16960_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10160_));
 sg13g2_buf_2 _16961_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10161_));
 sg13g2_xnor2_1 _16962_ (.Y(_10162_),
    .A(_10160_),
    .B(_10161_));
 sg13g2_nor3_1 _16963_ (.A(net135),
    .B(net104),
    .C(_10162_),
    .Y(_10163_));
 sg13g2_a21o_1 _16964_ (.A2(net105),
    .A1(net898),
    .B1(_10163_),
    .X(_00043_));
 sg13g2_buf_1 _16965_ (.A(_10105_),
    .X(_10164_));
 sg13g2_buf_1 _16966_ (.A(net1048),
    .X(_10165_));
 sg13g2_buf_1 _16967_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10166_));
 sg13g2_nand2_1 _16968_ (.Y(_10167_),
    .A(_10160_),
    .B(_10161_));
 sg13g2_xor2_1 _16969_ (.B(_10167_),
    .A(_10166_),
    .X(_10168_));
 sg13g2_nor3_1 _16970_ (.A(net136),
    .B(net104),
    .C(_10168_),
    .Y(_10169_));
 sg13g2_a21o_1 _16971_ (.A2(net105),
    .A1(net897),
    .B1(_10169_),
    .X(_00044_));
 sg13g2_buf_1 _16972_ (.A(_10111_),
    .X(_10170_));
 sg13g2_buf_1 _16973_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10171_));
 sg13g2_nand2_1 _16974_ (.Y(_10172_),
    .A(_10161_),
    .B(_10166_));
 sg13g2_nor2_1 _16975_ (.A(_00288_),
    .B(_10172_),
    .Y(_10173_));
 sg13g2_xnor2_1 _16976_ (.Y(_10174_),
    .A(_10171_),
    .B(_10173_));
 sg13g2_nor3_1 _16977_ (.A(net136),
    .B(net104),
    .C(_10174_),
    .Y(_10175_));
 sg13g2_a21o_1 _16978_ (.A2(net105),
    .A1(_10170_),
    .B1(_10175_),
    .X(_00045_));
 sg13g2_buf_1 _16979_ (.A(_10116_),
    .X(_10176_));
 sg13g2_buf_1 _16980_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10177_));
 sg13g2_and4_1 _16981_ (.A(_10160_),
    .B(_10161_),
    .C(_10166_),
    .D(_10171_),
    .X(_10178_));
 sg13g2_xnor2_1 _16982_ (.Y(_10179_),
    .A(_10177_),
    .B(_10178_));
 sg13g2_nor3_1 _16983_ (.A(net136),
    .B(net104),
    .C(_10179_),
    .Y(_10180_));
 sg13g2_a21o_1 _16984_ (.A2(net135),
    .A1(net1047),
    .B1(_10180_),
    .X(_00046_));
 sg13g2_buf_1 _16985_ (.A(net1052),
    .X(_10181_));
 sg13g2_buf_1 _16986_ (.A(net134),
    .X(_10182_));
 sg13g2_buf_2 _16987_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10183_));
 sg13g2_and3_1 _16988_ (.X(_10184_),
    .A(_10171_),
    .B(_10177_),
    .C(_10173_));
 sg13g2_buf_2 _16989_ (.A(_10184_),
    .X(_10185_));
 sg13g2_xnor2_1 _16990_ (.Y(_10186_),
    .A(_10183_),
    .B(_10185_));
 sg13g2_nor3_1 _16991_ (.A(net136),
    .B(net103),
    .C(_10186_),
    .Y(_10187_));
 sg13g2_a21o_1 _16992_ (.A2(net135),
    .A1(_10181_),
    .B1(_10187_),
    .X(_00047_));
 sg13g2_buf_1 _16993_ (.A(net1051),
    .X(_10188_));
 sg13g2_buf_1 _16994_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10189_));
 sg13g2_and2_1 _16995_ (.A(_10177_),
    .B(_10178_),
    .X(_10190_));
 sg13g2_buf_1 _16996_ (.A(_10190_),
    .X(_10191_));
 sg13g2_nand2_1 _16997_ (.Y(_10192_),
    .A(_10183_),
    .B(_10191_));
 sg13g2_xor2_1 _16998_ (.B(_10192_),
    .A(_10189_),
    .X(_10193_));
 sg13g2_nor3_1 _16999_ (.A(net136),
    .B(net103),
    .C(_10193_),
    .Y(_10194_));
 sg13g2_a21o_1 _17000_ (.A2(net135),
    .A1(_10188_),
    .B1(_10194_),
    .X(_00048_));
 sg13g2_buf_1 _17001_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10195_));
 sg13g2_nand3_1 _17002_ (.B(_10189_),
    .C(_10185_),
    .A(_10183_),
    .Y(_10196_));
 sg13g2_xor2_1 _17003_ (.B(_10196_),
    .A(_10195_),
    .X(_10197_));
 sg13g2_nor3_1 _17004_ (.A(net136),
    .B(net103),
    .C(_10197_),
    .Y(_10198_));
 sg13g2_a21o_1 _17005_ (.A2(net135),
    .A1(net899),
    .B1(_10198_),
    .X(_00049_));
 sg13g2_buf_2 _17006_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10199_));
 sg13g2_inv_1 _17007_ (.Y(_10200_),
    .A(_10191_));
 sg13g2_nand3_1 _17008_ (.B(_10189_),
    .C(_10195_),
    .A(_10183_),
    .Y(_10201_));
 sg13g2_nor2_1 _17009_ (.A(_10200_),
    .B(_10201_),
    .Y(_10202_));
 sg13g2_xnor2_1 _17010_ (.Y(_10203_),
    .A(_10199_),
    .B(_10202_));
 sg13g2_buf_1 _17011_ (.A(net544),
    .X(_10204_));
 sg13g2_buf_2 _17012_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10205_));
 sg13g2_nand3_1 _17013_ (.B(_10205_),
    .C(net170),
    .A(net484),
    .Y(_10206_));
 sg13g2_o21ai_1 _17014_ (.B1(_10206_),
    .Y(_00050_),
    .A1(net170),
    .A2(_10203_));
 sg13g2_buf_2 _17015_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10207_));
 sg13g2_nand2_1 _17016_ (.Y(_10208_),
    .A(_10199_),
    .B(_10202_));
 sg13g2_xor2_1 _17017_ (.B(_10208_),
    .A(_10207_),
    .X(_10209_));
 sg13g2_buf_2 _17018_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10210_));
 sg13g2_nand3_1 _17019_ (.B(_10210_),
    .C(net170),
    .A(net484),
    .Y(_10211_));
 sg13g2_o21ai_1 _17020_ (.B1(_10211_),
    .Y(_00051_),
    .A1(net170),
    .A2(_10209_));
 sg13g2_buf_1 _17021_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10212_));
 sg13g2_nand3_1 _17022_ (.B(_10207_),
    .C(_10202_),
    .A(_10199_),
    .Y(_10213_));
 sg13g2_xor2_1 _17023_ (.B(_10213_),
    .A(_10212_),
    .X(_10214_));
 sg13g2_buf_2 _17024_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10215_));
 sg13g2_nand3_1 _17025_ (.B(_10215_),
    .C(net192),
    .A(net484),
    .Y(_10216_));
 sg13g2_o21ai_1 _17026_ (.B1(_10216_),
    .Y(_00037_),
    .A1(net170),
    .A2(_10214_));
 sg13g2_buf_2 _17027_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10217_));
 sg13g2_nand3_1 _17028_ (.B(_10207_),
    .C(_10212_),
    .A(_10199_),
    .Y(_10218_));
 sg13g2_nor2_1 _17029_ (.A(_10201_),
    .B(_10218_),
    .Y(_10219_));
 sg13g2_nand2_1 _17030_ (.Y(_10220_),
    .A(_10185_),
    .B(_10219_));
 sg13g2_xor2_1 _17031_ (.B(_10220_),
    .A(_10217_),
    .X(_10221_));
 sg13g2_buf_2 _17032_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10222_));
 sg13g2_nand3_1 _17033_ (.B(_10222_),
    .C(net192),
    .A(net484),
    .Y(_10223_));
 sg13g2_o21ai_1 _17034_ (.B1(_10223_),
    .Y(_00038_),
    .A1(net170),
    .A2(_10221_));
 sg13g2_buf_1 _17035_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10224_));
 sg13g2_nand3_1 _17036_ (.B(_10191_),
    .C(_10219_),
    .A(_10217_),
    .Y(_10225_));
 sg13g2_xor2_1 _17037_ (.B(_10225_),
    .A(_10224_),
    .X(_10226_));
 sg13g2_buf_2 _17038_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10227_));
 sg13g2_nand3_1 _17039_ (.B(_10227_),
    .C(net192),
    .A(net484),
    .Y(_10228_));
 sg13g2_o21ai_1 _17040_ (.B1(_10228_),
    .Y(_00039_),
    .A1(_10143_),
    .A2(_10226_));
 sg13g2_buf_2 _17041_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10229_));
 sg13g2_buf_1 _17042_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10230_));
 sg13g2_nand4_1 _17043_ (.B(_10224_),
    .C(_10185_),
    .A(_10217_),
    .Y(_10231_),
    .D(_10219_));
 sg13g2_xor2_1 _17044_ (.B(_10231_),
    .A(_10230_),
    .X(_10232_));
 sg13g2_nor3_1 _17045_ (.A(_10148_),
    .B(_10182_),
    .C(_10232_),
    .Y(_10233_));
 sg13g2_a21o_1 _17046_ (.A2(net135),
    .A1(_10229_),
    .B1(_10233_),
    .X(_00040_));
 sg13g2_buf_1 _17047_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10234_));
 sg13g2_and4_1 _17048_ (.A(_10217_),
    .B(_10224_),
    .C(_10230_),
    .D(_10219_),
    .X(_10235_));
 sg13g2_buf_1 _17049_ (.A(_10235_),
    .X(_10236_));
 sg13g2_nand2_1 _17050_ (.Y(_10237_),
    .A(_10191_),
    .B(_10236_));
 sg13g2_xor2_1 _17051_ (.B(_10237_),
    .A(_10234_),
    .X(_10238_));
 sg13g2_buf_1 _17052_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10239_));
 sg13g2_nand3_1 _17053_ (.B(_10239_),
    .C(net192),
    .A(net484),
    .Y(_10240_));
 sg13g2_o21ai_1 _17054_ (.B1(_10240_),
    .Y(_00041_),
    .A1(net170),
    .A2(_10238_));
 sg13g2_buf_1 _17055_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10241_));
 sg13g2_nand3_1 _17056_ (.B(_10185_),
    .C(_10236_),
    .A(_10234_),
    .Y(_10242_));
 sg13g2_xor2_1 _17057_ (.B(_10242_),
    .A(_10241_),
    .X(_10243_));
 sg13g2_buf_2 _17058_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10244_));
 sg13g2_nand3_1 _17059_ (.B(_10244_),
    .C(net192),
    .A(net484),
    .Y(_10245_));
 sg13g2_o21ai_1 _17060_ (.B1(_10245_),
    .Y(_00042_),
    .A1(net170),
    .A2(_10243_));
 sg13g2_buf_1 _17061_ (.A(\cpu.ex.r_mult[0] ),
    .X(_10246_));
 sg13g2_buf_1 _17062_ (.A(net689),
    .X(_10247_));
 sg13g2_buf_1 _17063_ (.A(_09390_),
    .X(_10248_));
 sg13g2_inv_1 _17064_ (.Y(_10249_),
    .A(\cpu.ex.r_div_running ));
 sg13g2_inv_4 _17065_ (.A(net1141),
    .Y(_10250_));
 sg13g2_nand2_1 _17066_ (.Y(_10251_),
    .A(_10249_),
    .B(_10250_));
 sg13g2_nor3_2 _17067_ (.A(net610),
    .B(net609),
    .C(_10251_),
    .Y(_10252_));
 sg13g2_buf_1 _17068_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10253_));
 sg13g2_inv_1 _17069_ (.Y(_10254_),
    .A(net1132));
 sg13g2_buf_8 _17070_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10255_));
 sg13g2_buf_2 _17071_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10256_));
 sg13g2_buf_8 _17072_ (.A(_10256_),
    .X(_10257_));
 sg13g2_nand2_1 _17073_ (.Y(_10258_),
    .A(net1131),
    .B(net1046));
 sg13g2_buf_8 _17074_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10259_));
 sg13g2_buf_8 _17075_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10260_));
 sg13g2_inv_1 _17076_ (.Y(_10261_),
    .A(_10260_));
 sg13g2_nor2_1 _17077_ (.A(net1130),
    .B(_10261_),
    .Y(_10262_));
 sg13g2_inv_1 _17078_ (.Y(_10263_),
    .A(_10262_));
 sg13g2_nor3_1 _17079_ (.A(_10254_),
    .B(_10258_),
    .C(_10263_),
    .Y(_10264_));
 sg13g2_buf_1 _17080_ (.A(_10264_),
    .X(_10265_));
 sg13g2_buf_1 _17081_ (.A(\cpu.ex.r_set_cc ),
    .X(_10266_));
 sg13g2_nand2_2 _17082_ (.Y(_10267_),
    .A(net1132),
    .B(_10266_));
 sg13g2_nor2b_1 _17083_ (.A(_10265_),
    .B_N(_10267_),
    .Y(_10268_));
 sg13g2_buf_1 _17084_ (.A(_10268_),
    .X(_10269_));
 sg13g2_nand2b_1 _17085_ (.Y(_10270_),
    .B(_10269_),
    .A_N(_10252_));
 sg13g2_buf_2 _17086_ (.A(_10270_),
    .X(_10271_));
 sg13g2_buf_1 _17087_ (.A(_10271_),
    .X(_10272_));
 sg13g2_buf_2 _17088_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10273_));
 sg13g2_buf_1 _17089_ (.A(\cpu.dec.r_rs2_inv ),
    .X(_10274_));
 sg13g2_or2_1 _17090_ (.X(_10275_),
    .B(_10274_),
    .A(_10273_));
 sg13g2_buf_2 _17091_ (.A(_10275_),
    .X(_10276_));
 sg13g2_nor4_1 _17092_ (.A(net1131),
    .B(_10256_),
    .C(net1130),
    .D(_10260_),
    .Y(_10277_));
 sg13g2_nand2b_1 _17093_ (.Y(_10278_),
    .B(net1132),
    .A_N(_10277_));
 sg13g2_buf_1 _17094_ (.A(_10278_),
    .X(_10279_));
 sg13g2_buf_8 _17095_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10280_));
 sg13g2_xnor2_1 _17096_ (.Y(_10281_),
    .A(net1130),
    .B(_10280_));
 sg13g2_buf_8 _17097_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10282_));
 sg13g2_xnor2_1 _17098_ (.Y(_10283_),
    .A(_10256_),
    .B(_10282_));
 sg13g2_buf_8 _17099_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10284_));
 sg13g2_xnor2_1 _17100_ (.Y(_10285_),
    .A(_10260_),
    .B(_10284_));
 sg13g2_buf_8 _17101_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10286_));
 sg13g2_xnor2_1 _17102_ (.Y(_10287_),
    .A(net1131),
    .B(_10286_));
 sg13g2_nand4_1 _17103_ (.B(_10283_),
    .C(_10285_),
    .A(_10281_),
    .Y(_10288_),
    .D(_10287_));
 sg13g2_buf_1 _17104_ (.A(_10288_),
    .X(_10289_));
 sg13g2_nor2_1 _17105_ (.A(_10279_),
    .B(_10289_),
    .Y(_10290_));
 sg13g2_buf_8 _17106_ (.A(_10290_),
    .X(_10291_));
 sg13g2_buf_1 _17107_ (.A(_10291_),
    .X(_10292_));
 sg13g2_buf_8 _17108_ (.A(_10282_),
    .X(_10293_));
 sg13g2_buf_8 _17109_ (.A(net1045),
    .X(_10294_));
 sg13g2_buf_1 _17110_ (.A(_10294_),
    .X(_10295_));
 sg13g2_buf_1 _17111_ (.A(net770),
    .X(_10296_));
 sg13g2_buf_8 _17112_ (.A(net677),
    .X(_10297_));
 sg13g2_buf_8 _17113_ (.A(_10280_),
    .X(_10298_));
 sg13g2_buf_8 _17114_ (.A(net1044),
    .X(_10299_));
 sg13g2_buf_8 _17115_ (.A(net892),
    .X(_10300_));
 sg13g2_buf_8 _17116_ (.A(net769),
    .X(_10301_));
 sg13g2_buf_1 _17117_ (.A(net676),
    .X(_10302_));
 sg13g2_buf_8 _17118_ (.A(_10284_),
    .X(_10303_));
 sg13g2_nor2b_1 _17119_ (.A(net1043),
    .B_N(_10286_),
    .Y(_10304_));
 sg13g2_buf_2 _17120_ (.A(_10304_),
    .X(_10305_));
 sg13g2_nor2b_1 _17121_ (.A(_10286_),
    .B_N(net1043),
    .Y(_10306_));
 sg13g2_buf_1 _17122_ (.A(_10306_),
    .X(_10307_));
 sg13g2_buf_2 _17123_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10308_));
 sg13g2_a22oi_1 _17124_ (.Y(_10309_),
    .B1(net768),
    .B2(_10308_),
    .A2(_10305_),
    .A1(\cpu.ex.r_epc[15] ));
 sg13g2_buf_8 _17125_ (.A(_10286_),
    .X(_10310_));
 sg13g2_buf_8 _17126_ (.A(net1042),
    .X(_10311_));
 sg13g2_nor2b_1 _17127_ (.A(_10311_),
    .B_N(net892),
    .Y(_10312_));
 sg13g2_buf_8 _17128_ (.A(_10312_),
    .X(_10313_));
 sg13g2_buf_1 _17129_ (.A(net675),
    .X(_10314_));
 sg13g2_buf_8 _17130_ (.A(net1043),
    .X(_10315_));
 sg13g2_buf_2 _17131_ (.A(net890),
    .X(_10316_));
 sg13g2_buf_1 _17132_ (.A(net767),
    .X(_10317_));
 sg13g2_buf_1 _17133_ (.A(net674),
    .X(_10318_));
 sg13g2_mux2_1 _17134_ (.A0(\cpu.ex.r_9[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .S(net604),
    .X(_10319_));
 sg13g2_nand2_1 _17135_ (.Y(_10320_),
    .A(net605),
    .B(_10319_));
 sg13g2_o21ai_1 _17136_ (.B1(_10320_),
    .Y(_10321_),
    .A1(net606),
    .A2(_10309_));
 sg13g2_buf_1 _17137_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10322_));
 sg13g2_buf_8 _17138_ (.A(net1044),
    .X(_10323_));
 sg13g2_nor2b_1 _17139_ (.A(_10323_),
    .B_N(net1042),
    .Y(_10324_));
 sg13g2_buf_2 _17140_ (.A(_10324_),
    .X(_10325_));
 sg13g2_buf_8 _17141_ (.A(_10325_),
    .X(_10326_));
 sg13g2_a22oi_1 _17142_ (.Y(_10327_),
    .B1(net605),
    .B2(\cpu.ex.r_8[15] ),
    .A2(net603),
    .A1(_10322_));
 sg13g2_or2_1 _17143_ (.X(_10328_),
    .B(_10284_),
    .A(_10282_));
 sg13g2_buf_1 _17144_ (.A(_10328_),
    .X(_10329_));
 sg13g2_nor2_1 _17145_ (.A(_10327_),
    .B(_10329_),
    .Y(_10330_));
 sg13g2_a21oi_1 _17146_ (.A1(_10297_),
    .A2(_10321_),
    .Y(_10331_),
    .B1(_10330_));
 sg13g2_buf_8 _17147_ (.A(net891),
    .X(_10332_));
 sg13g2_inv_2 _17148_ (.Y(_10333_),
    .A(net766));
 sg13g2_buf_8 _17149_ (.A(_10333_),
    .X(_10334_));
 sg13g2_inv_1 _17150_ (.Y(_10335_),
    .A(_10293_));
 sg13g2_buf_8 _17151_ (.A(_10335_),
    .X(_10336_));
 sg13g2_buf_1 _17152_ (.A(net765),
    .X(_10337_));
 sg13g2_nor2b_1 _17153_ (.A(_10303_),
    .B_N(net1044),
    .Y(_10338_));
 sg13g2_buf_1 _17154_ (.A(_10338_),
    .X(_10339_));
 sg13g2_mux2_1 _17155_ (.A0(\cpu.ex.r_stmp[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(net606),
    .X(_10340_));
 sg13g2_a22oi_1 _17156_ (.Y(_10341_),
    .B1(_10340_),
    .B2(net604),
    .A2(net764),
    .A1(\cpu.ex.r_10[15] ));
 sg13g2_mux2_1 _17157_ (.A0(\cpu.ex.r_mult[31] ),
    .A1(\cpu.ex.r_15[15] ),
    .S(net606),
    .X(_10342_));
 sg13g2_a221oi_1 _17158_ (.B2(_10318_),
    .C1(net673),
    .B1(_10342_),
    .A1(\cpu.ex.r_11[15] ),
    .Y(_10343_),
    .A2(net764));
 sg13g2_a21oi_1 _17159_ (.A1(net673),
    .A2(_10341_),
    .Y(_10344_),
    .B1(_10343_));
 sg13g2_and2_1 _17160_ (.A(_10298_),
    .B(net1043),
    .X(_10345_));
 sg13g2_buf_1 _17161_ (.A(_10345_),
    .X(_10346_));
 sg13g2_nand3_1 _17162_ (.B(net673),
    .C(net763),
    .A(\cpu.ex.r_12[15] ),
    .Y(_10347_));
 sg13g2_nor2_1 _17163_ (.A(net1044),
    .B(_10284_),
    .Y(_10348_));
 sg13g2_buf_2 _17164_ (.A(_10348_),
    .X(_10349_));
 sg13g2_buf_1 _17165_ (.A(_10349_),
    .X(_10350_));
 sg13g2_nand3_1 _17166_ (.B(net607),
    .C(net672),
    .A(\cpu.ex.r_lr[15] ),
    .Y(_10351_));
 sg13g2_nand3_1 _17167_ (.B(_10347_),
    .C(_10351_),
    .A(net602),
    .Y(_10352_));
 sg13g2_o21ai_1 _17168_ (.B1(_10352_),
    .Y(_10353_),
    .A1(net602),
    .A2(_10344_));
 sg13g2_nor2_1 _17169_ (.A(_10282_),
    .B(_10286_),
    .Y(_10354_));
 sg13g2_buf_2 _17170_ (.A(_10354_),
    .X(_10355_));
 sg13g2_nand2_1 _17171_ (.Y(_10356_),
    .A(_10355_),
    .B(_10349_));
 sg13g2_o21ai_1 _17172_ (.B1(_10356_),
    .Y(_10357_),
    .A1(_10279_),
    .A2(_10289_));
 sg13g2_buf_1 _17173_ (.A(_10357_),
    .X(_10358_));
 sg13g2_a21oi_1 _17174_ (.A1(_10331_),
    .A2(_10353_),
    .Y(_10359_),
    .B1(net540));
 sg13g2_a21o_1 _17175_ (.A2(net541),
    .A1(net907),
    .B1(_10359_),
    .X(_10360_));
 sg13g2_buf_8 _17176_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10361_));
 sg13g2_buf_1 _17177_ (.A(_10361_),
    .X(_10362_));
 sg13g2_mux2_1 _17178_ (.A0(\cpu.dec.imm[15] ),
    .A1(_10360_),
    .S(net1041),
    .X(_10363_));
 sg13g2_buf_8 _17179_ (.A(_10273_),
    .X(_10364_));
 sg13g2_nand2_1 _17180_ (.Y(_10365_),
    .A(net712),
    .B(net1040));
 sg13g2_o21ai_1 _17181_ (.B1(_10365_),
    .Y(_10366_),
    .A1(_10276_),
    .A2(_10363_));
 sg13g2_buf_2 _17182_ (.A(_10366_),
    .X(_10367_));
 sg13g2_buf_1 _17183_ (.A(\cpu.br ),
    .X(_10368_));
 sg13g2_nand2_1 _17184_ (.Y(_10369_),
    .A(_08354_),
    .B(_08363_));
 sg13g2_nand2_1 _17185_ (.Y(_10370_),
    .A(_10368_),
    .B(_10369_));
 sg13g2_a21o_1 _17186_ (.A2(_08452_),
    .A1(net490),
    .B1(_10370_),
    .X(_10371_));
 sg13g2_buf_8 _17187_ (.A(_10371_),
    .X(_10372_));
 sg13g2_buf_1 _17188_ (.A(_10368_),
    .X(_10373_));
 sg13g2_buf_8 _17189_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10374_));
 sg13g2_buf_1 _17190_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10375_));
 sg13g2_nor2_2 _17191_ (.A(net1129),
    .B(net1128),
    .Y(_10376_));
 sg13g2_buf_2 _17192_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10377_));
 sg13g2_buf_8 _17193_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10378_));
 sg13g2_nor2_2 _17194_ (.A(_10377_),
    .B(_10378_),
    .Y(_10379_));
 sg13g2_a21oi_1 _17195_ (.A1(_10376_),
    .A2(_10379_),
    .Y(_10380_),
    .B1(_00275_));
 sg13g2_inv_1 _17196_ (.Y(_10381_),
    .A(_09244_));
 sg13g2_nor2_1 _17197_ (.A(_10381_),
    .B(_09243_),
    .Y(_10382_));
 sg13g2_o21ai_1 _17198_ (.B1(_10382_),
    .Y(_10383_),
    .A1(_09259_),
    .A2(_09268_));
 sg13g2_a21oi_1 _17199_ (.A1(_09242_),
    .A2(_09282_),
    .Y(_10384_),
    .B1(_09241_));
 sg13g2_nand3_1 _17200_ (.B(_10383_),
    .C(_10384_),
    .A(_10380_),
    .Y(_10385_));
 sg13g2_buf_1 _17201_ (.A(_10385_),
    .X(_10386_));
 sg13g2_a21o_1 _17202_ (.A2(_08358_),
    .A1(_08318_),
    .B1(_10386_),
    .X(_10387_));
 sg13g2_buf_8 _17203_ (.A(_10387_),
    .X(_10388_));
 sg13g2_nand2_1 _17204_ (.Y(_10389_),
    .A(net1039),
    .B(_10388_));
 sg13g2_buf_8 _17205_ (.A(_10389_),
    .X(_10390_));
 sg13g2_a21o_1 _17206_ (.A2(_10390_),
    .A1(_10372_),
    .B1(_00299_),
    .X(_10391_));
 sg13g2_buf_1 _17207_ (.A(_10391_),
    .X(_10392_));
 sg13g2_nor2_1 _17208_ (.A(_10254_),
    .B(_10277_),
    .Y(_10393_));
 sg13g2_xor2_1 _17209_ (.B(net1129),
    .A(net1130),
    .X(_10394_));
 sg13g2_xor2_1 _17210_ (.B(_10378_),
    .A(net1046),
    .X(_10395_));
 sg13g2_xor2_1 _17211_ (.B(net1128),
    .A(_10260_),
    .X(_10396_));
 sg13g2_xor2_1 _17212_ (.B(_10377_),
    .A(net1131),
    .X(_10397_));
 sg13g2_nor4_1 _17213_ (.A(_10394_),
    .B(_10395_),
    .C(_10396_),
    .D(_10397_),
    .Y(_10398_));
 sg13g2_and2_1 _17214_ (.A(_10393_),
    .B(_10398_),
    .X(_10399_));
 sg13g2_buf_8 _17215_ (.A(_10399_),
    .X(_10400_));
 sg13g2_inv_1 _17216_ (.Y(_10401_),
    .A(\cpu.ex.r_13[2] ));
 sg13g2_buf_8 _17217_ (.A(_10377_),
    .X(_10402_));
 sg13g2_buf_1 _17218_ (.A(net1038),
    .X(_10403_));
 sg13g2_buf_1 _17219_ (.A(net1128),
    .X(_10404_));
 sg13g2_nand2b_1 _17220_ (.Y(_10405_),
    .B(net1037),
    .A_N(net888));
 sg13g2_inv_1 _17221_ (.Y(_10406_),
    .A(_00262_));
 sg13g2_and2_1 _17222_ (.A(_10377_),
    .B(net1128),
    .X(_10407_));
 sg13g2_buf_1 _17223_ (.A(_10407_),
    .X(_10408_));
 sg13g2_inv_2 _17224_ (.Y(_10409_),
    .A(_10377_));
 sg13g2_buf_8 _17225_ (.A(net1128),
    .X(_10410_));
 sg13g2_nor2_1 _17226_ (.A(_10409_),
    .B(net1036),
    .Y(_10411_));
 sg13g2_a22oi_1 _17227_ (.Y(_10412_),
    .B1(_10411_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10408_),
    .A1(_10406_));
 sg13g2_o21ai_1 _17228_ (.B1(_10412_),
    .Y(_10413_),
    .A1(_10401_),
    .A2(_10405_));
 sg13g2_buf_8 _17229_ (.A(_10378_),
    .X(_10414_));
 sg13g2_buf_8 _17230_ (.A(net1035),
    .X(_10415_));
 sg13g2_buf_8 _17231_ (.A(net1129),
    .X(_10416_));
 sg13g2_buf_1 _17232_ (.A(net1034),
    .X(_10417_));
 sg13g2_and2_1 _17233_ (.A(net887),
    .B(net886),
    .X(_10418_));
 sg13g2_buf_2 _17234_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10419_));
 sg13g2_inv_2 _17235_ (.Y(_10420_),
    .A(_10419_));
 sg13g2_inv_2 _17236_ (.Y(_10421_),
    .A(_10416_));
 sg13g2_nor2b_1 _17237_ (.A(net1038),
    .B_N(_10378_),
    .Y(_10422_));
 sg13g2_buf_1 _17238_ (.A(_10422_),
    .X(_10423_));
 sg13g2_nand2_1 _17239_ (.Y(_10424_),
    .A(_10421_),
    .B(_10423_));
 sg13g2_buf_1 _17240_ (.A(net1034),
    .X(_10425_));
 sg13g2_nor2b_1 _17241_ (.A(net1035),
    .B_N(_10402_),
    .Y(_10426_));
 sg13g2_buf_2 _17242_ (.A(_10426_),
    .X(_10427_));
 sg13g2_nand3_1 _17243_ (.B(\cpu.ex.r_14[2] ),
    .C(_10427_),
    .A(net885),
    .Y(_10428_));
 sg13g2_o21ai_1 _17244_ (.B1(_10428_),
    .Y(_10429_),
    .A1(_10420_),
    .A2(_10424_));
 sg13g2_buf_1 _17245_ (.A(net1036),
    .X(_10430_));
 sg13g2_buf_1 _17246_ (.A(net884),
    .X(_10431_));
 sg13g2_buf_2 _17247_ (.A(net887),
    .X(_10432_));
 sg13g2_nor3_2 _17248_ (.A(_10409_),
    .B(_10421_),
    .C(_10410_),
    .Y(_10433_));
 sg13g2_nor2b_1 _17249_ (.A(net1129),
    .B_N(net1128),
    .Y(_10434_));
 sg13g2_buf_1 _17250_ (.A(_10434_),
    .X(_10435_));
 sg13g2_and2_1 _17251_ (.A(_10409_),
    .B(net883),
    .X(_10436_));
 sg13g2_a22oi_1 _17252_ (.Y(_10437_),
    .B1(_10436_),
    .B2(_08364_),
    .A2(_10433_),
    .A1(\cpu.ex.r_10[2] ));
 sg13g2_nor2_1 _17253_ (.A(net761),
    .B(_10437_),
    .Y(_10438_));
 sg13g2_a221oi_1 _17254_ (.B2(net762),
    .C1(_10438_),
    .B1(_10429_),
    .A1(_10413_),
    .Y(_10439_),
    .A2(_10418_));
 sg13g2_and2_1 _17255_ (.A(_10378_),
    .B(_10375_),
    .X(_10440_));
 sg13g2_buf_1 _17256_ (.A(_10440_),
    .X(_10441_));
 sg13g2_nor2_2 _17257_ (.A(net887),
    .B(net1036),
    .Y(_10442_));
 sg13g2_buf_1 _17258_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10443_));
 sg13g2_a22oi_1 _17259_ (.Y(_10444_),
    .B1(_10442_),
    .B2(_10443_),
    .A2(_10441_),
    .A1(\cpu.ex.r_mult[18] ));
 sg13g2_nor2b_1 _17260_ (.A(net1129),
    .B_N(_10377_),
    .Y(_10445_));
 sg13g2_buf_1 _17261_ (.A(_10445_),
    .X(_10446_));
 sg13g2_nor2b_1 _17262_ (.A(_10444_),
    .B_N(net882),
    .Y(_10447_));
 sg13g2_nor2_1 _17263_ (.A(net1035),
    .B(net1034),
    .Y(_10448_));
 sg13g2_nand3_1 _17264_ (.B(_10408_),
    .C(_10448_),
    .A(\cpu.ex.r_stmp[2] ),
    .Y(_10449_));
 sg13g2_nor2b_1 _17265_ (.A(net1128),
    .B_N(net1129),
    .Y(_10450_));
 sg13g2_buf_2 _17266_ (.A(_10450_),
    .X(_10451_));
 sg13g2_nand3_1 _17267_ (.B(_10379_),
    .C(_10451_),
    .A(\cpu.ex.r_8[2] ),
    .Y(_10452_));
 sg13g2_or2_1 _17268_ (.X(_10453_),
    .B(\cpu.dec.r_rs1[2] ),
    .A(net1129));
 sg13g2_buf_1 _17269_ (.A(_10453_),
    .X(_10454_));
 sg13g2_nand2_1 _17270_ (.Y(_10455_),
    .A(_10377_),
    .B(_10378_));
 sg13g2_nor2_1 _17271_ (.A(_10454_),
    .B(_10455_),
    .Y(_10456_));
 sg13g2_buf_2 _17272_ (.A(_10456_),
    .X(_10457_));
 sg13g2_nand2b_1 _17273_ (.Y(_10458_),
    .B(_10378_),
    .A_N(_10377_));
 sg13g2_buf_1 _17274_ (.A(_10458_),
    .X(_10459_));
 sg13g2_nor2_1 _17275_ (.A(_10410_),
    .B(_10459_),
    .Y(_10460_));
 sg13g2_mux2_1 _17276_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(\cpu.ex.r_9[2] ),
    .S(net1034),
    .X(_10461_));
 sg13g2_a22oi_1 _17277_ (.Y(_10462_),
    .B1(_10460_),
    .B2(_10461_),
    .A2(_10457_),
    .A1(\cpu.ex.r_epc[2] ));
 sg13g2_nand3_1 _17278_ (.B(_10452_),
    .C(_10462_),
    .A(_10449_),
    .Y(_10463_));
 sg13g2_and2_1 _17279_ (.A(_10374_),
    .B(_10375_),
    .X(_10464_));
 sg13g2_buf_1 _17280_ (.A(_10464_),
    .X(_10465_));
 sg13g2_and2_1 _17281_ (.A(_10379_),
    .B(_10465_),
    .X(_10466_));
 sg13g2_buf_1 _17282_ (.A(_10466_),
    .X(_10467_));
 sg13g2_and2_1 _17283_ (.A(\cpu.ex.r_12[2] ),
    .B(_10467_),
    .X(_10468_));
 sg13g2_nor4_1 _17284_ (.A(_10400_),
    .B(_10447_),
    .C(_10463_),
    .D(_10468_),
    .Y(_10469_));
 sg13g2_a22oi_1 _17285_ (.Y(_10470_),
    .B1(_10439_),
    .B2(_10469_),
    .A2(_10400_),
    .A1(_09459_));
 sg13g2_buf_2 _17286_ (.A(_10470_),
    .X(_10471_));
 sg13g2_nand3_1 _17287_ (.B(_10390_),
    .C(_10471_),
    .A(_10372_),
    .Y(_10472_));
 sg13g2_buf_2 _17288_ (.A(_10472_),
    .X(_10473_));
 sg13g2_nand3_1 _17289_ (.B(_10392_),
    .C(_10473_),
    .A(_09384_),
    .Y(_10474_));
 sg13g2_a21o_1 _17290_ (.A2(_10390_),
    .A1(_10372_),
    .B1(_00191_),
    .X(_10475_));
 sg13g2_buf_2 _17291_ (.A(_10475_),
    .X(_10476_));
 sg13g2_buf_8 _17292_ (.A(_10372_),
    .X(_10477_));
 sg13g2_buf_8 _17293_ (.A(_10390_),
    .X(_10478_));
 sg13g2_nand2_1 _17294_ (.Y(_10479_),
    .A(_10393_),
    .B(_10398_));
 sg13g2_buf_2 _17295_ (.A(_10479_),
    .X(_10480_));
 sg13g2_buf_1 _17296_ (.A(_10480_),
    .X(_10481_));
 sg13g2_nand2b_1 _17297_ (.Y(_10482_),
    .B(net1038),
    .A_N(net1035));
 sg13g2_buf_2 _17298_ (.A(_10482_),
    .X(_10483_));
 sg13g2_buf_1 _17299_ (.A(_10451_),
    .X(_10484_));
 sg13g2_a22oi_1 _17300_ (.Y(_10485_),
    .B1(net760),
    .B2(\cpu.ex.r_10[3] ),
    .A2(net883),
    .A1(\cpu.ex.r_stmp[3] ));
 sg13g2_nor2b_1 _17301_ (.A(net1038),
    .B_N(_10416_),
    .Y(_10486_));
 sg13g2_buf_2 _17302_ (.A(_10486_),
    .X(_10487_));
 sg13g2_a22oi_1 _17303_ (.Y(_10488_),
    .B1(net882),
    .B2(\cpu.ex.r_mult[19] ),
    .A2(_10487_),
    .A1(\cpu.ex.r_13[3] ));
 sg13g2_nand2b_1 _17304_ (.Y(_10489_),
    .B(_10441_),
    .A_N(_10488_));
 sg13g2_o21ai_1 _17305_ (.B1(_10489_),
    .Y(_10490_),
    .A1(_10483_),
    .A2(_10485_));
 sg13g2_nand2_1 _17306_ (.Y(_10491_),
    .A(_10409_),
    .B(net885));
 sg13g2_nor2b_1 _17307_ (.A(net761),
    .B_N(net1037),
    .Y(_10492_));
 sg13g2_nor2b_1 _17308_ (.A(net884),
    .B_N(net761),
    .Y(_10493_));
 sg13g2_a22oi_1 _17309_ (.Y(_10494_),
    .B1(_10493_),
    .B2(\cpu.ex.r_9[3] ),
    .A2(_10492_),
    .A1(\cpu.ex.r_12[3] ));
 sg13g2_nor2_1 _17310_ (.A(net888),
    .B(net1037),
    .Y(_10495_));
 sg13g2_a22oi_1 _17311_ (.Y(_10496_),
    .B1(_10495_),
    .B2(\cpu.ex.r_8[3] ),
    .A2(_10408_),
    .A1(\cpu.ex.r_14[3] ));
 sg13g2_nor2b_1 _17312_ (.A(net1035),
    .B_N(net1129),
    .Y(_10497_));
 sg13g2_buf_1 _17313_ (.A(_10497_),
    .X(_10498_));
 sg13g2_buf_1 _17314_ (.A(_10498_),
    .X(_10499_));
 sg13g2_nand2b_1 _17315_ (.Y(_10500_),
    .B(net671),
    .A_N(_10496_));
 sg13g2_o21ai_1 _17316_ (.B1(_10500_),
    .Y(_10501_),
    .A1(_10491_),
    .A2(_10494_));
 sg13g2_inv_2 _17317_ (.Y(_10502_),
    .A(_10415_));
 sg13g2_buf_1 _17318_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10503_));
 sg13g2_a22oi_1 _17319_ (.Y(_10504_),
    .B1(_10436_),
    .B2(_10503_),
    .A2(_10433_),
    .A1(\cpu.ex.r_11[3] ));
 sg13g2_nor2_1 _17320_ (.A(net759),
    .B(_10504_),
    .Y(_10505_));
 sg13g2_buf_8 _17321_ (.A(_10417_),
    .X(_10506_));
 sg13g2_buf_1 _17322_ (.A(net758),
    .X(_10507_));
 sg13g2_nor2_1 _17323_ (.A(net884),
    .B(_10455_),
    .Y(_10508_));
 sg13g2_buf_1 _17324_ (.A(net888),
    .X(_10509_));
 sg13g2_nor2_1 _17325_ (.A(_08449_),
    .B(net757),
    .Y(_10510_));
 sg13g2_a22oi_1 _17326_ (.Y(_10511_),
    .B1(_10510_),
    .B2(_10492_),
    .A2(_10508_),
    .A1(\cpu.ex.r_epc[3] ));
 sg13g2_nor2_1 _17327_ (.A(_10454_),
    .B(_10459_),
    .Y(_10512_));
 sg13g2_buf_2 _17328_ (.A(_10512_),
    .X(_10513_));
 sg13g2_nor2_2 _17329_ (.A(_10454_),
    .B(_10483_),
    .Y(_10514_));
 sg13g2_buf_1 _17330_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10515_));
 sg13g2_nand4_1 _17331_ (.B(net887),
    .C(net1034),
    .A(_10402_),
    .Y(_10516_),
    .D(net1036));
 sg13g2_buf_1 _17332_ (.A(_10516_),
    .X(_10517_));
 sg13g2_nor2_1 _17333_ (.A(_00263_),
    .B(_10517_),
    .Y(_10518_));
 sg13g2_a221oi_1 _17334_ (.B2(_10515_),
    .C1(_10518_),
    .B1(_10514_),
    .A1(\cpu.ex.r_lr[3] ),
    .Y(_10519_),
    .A2(_10513_));
 sg13g2_o21ai_1 _17335_ (.B1(_10519_),
    .Y(_10520_),
    .A1(net670),
    .A2(_10511_));
 sg13g2_nor4_1 _17336_ (.A(_10490_),
    .B(_10501_),
    .C(_10505_),
    .D(_10520_),
    .Y(_10521_));
 sg13g2_nor2_1 _17337_ (.A(_09220_),
    .B(_10480_),
    .Y(_10522_));
 sg13g2_a21oi_1 _17338_ (.A1(net539),
    .A2(_10521_),
    .Y(_10523_),
    .B1(_10522_));
 sg13g2_nand3_1 _17339_ (.B(net269),
    .C(_10523_),
    .A(net339),
    .Y(_10524_));
 sg13g2_buf_1 _17340_ (.A(_10524_),
    .X(_10525_));
 sg13g2_nor2_1 _17341_ (.A(_09372_),
    .B(_09385_),
    .Y(_10526_));
 sg13g2_nor2b_1 _17342_ (.A(_09386_),
    .B_N(_09385_),
    .Y(_10527_));
 sg13g2_a22oi_1 _17343_ (.Y(_10528_),
    .B1(_10527_),
    .B2(net1142),
    .A2(_10526_),
    .A1(_09386_));
 sg13g2_nand2b_1 _17344_ (.Y(_10529_),
    .B(_09382_),
    .A_N(_10528_));
 sg13g2_a21oi_1 _17345_ (.A1(_10476_),
    .A2(_10525_),
    .Y(_10530_),
    .B1(_10529_));
 sg13g2_inv_1 _17346_ (.Y(_10531_),
    .A(_00298_));
 sg13g2_nand2_1 _17347_ (.Y(_10532_),
    .A(_10372_),
    .B(_10390_));
 sg13g2_buf_8 _17348_ (.A(_10532_),
    .X(_10533_));
 sg13g2_a21oi_1 _17349_ (.A1(net490),
    .A2(_08452_),
    .Y(_10534_),
    .B1(_10370_));
 sg13g2_buf_2 _17350_ (.A(_10534_),
    .X(_10535_));
 sg13g2_and2_1 _17351_ (.A(net1039),
    .B(_10388_),
    .X(_10536_));
 sg13g2_buf_8 _17352_ (.A(_10536_),
    .X(_10537_));
 sg13g2_buf_1 _17353_ (.A(_10400_),
    .X(_10538_));
 sg13g2_mux2_1 _17354_ (.A0(\cpu.ex.r_9[5] ),
    .A1(\cpu.ex.r_11[5] ),
    .S(net757),
    .X(_10539_));
 sg13g2_buf_1 _17355_ (.A(net761),
    .X(_10540_));
 sg13g2_and2_1 _17356_ (.A(net669),
    .B(_10451_),
    .X(_10541_));
 sg13g2_and2_1 _17357_ (.A(_10427_),
    .B(_10451_),
    .X(_10542_));
 sg13g2_buf_1 _17358_ (.A(_10542_),
    .X(_10543_));
 sg13g2_a22oi_1 _17359_ (.Y(_10544_),
    .B1(_10543_),
    .B2(\cpu.ex.r_10[5] ),
    .A2(_10541_),
    .A1(_10539_));
 sg13g2_nor2_1 _17360_ (.A(_00265_),
    .B(_10517_),
    .Y(_10545_));
 sg13g2_a21oi_1 _17361_ (.A1(\cpu.ex.r_lr[5] ),
    .A2(_10513_),
    .Y(_10546_),
    .B1(_10545_));
 sg13g2_buf_1 _17362_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10547_));
 sg13g2_a22oi_1 _17363_ (.Y(_10548_),
    .B1(_10442_),
    .B2(\cpu.ex.r_8[5] ),
    .A2(_10441_),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_nor2_1 _17364_ (.A(_10491_),
    .B(_10548_),
    .Y(_10549_));
 sg13g2_a221oi_1 _17365_ (.B2(_10547_),
    .C1(_10549_),
    .B1(_10514_),
    .A1(\cpu.ex.r_epc[5] ),
    .Y(_10550_),
    .A2(_10457_));
 sg13g2_nor2b_1 _17366_ (.A(net1034),
    .B_N(net1035),
    .Y(_10551_));
 sg13g2_buf_1 _17367_ (.A(_10551_),
    .X(_10552_));
 sg13g2_a22oi_1 _17368_ (.Y(_10553_),
    .B1(_10498_),
    .B2(\cpu.ex.r_14[5] ),
    .A2(_10552_),
    .A1(\cpu.ex.r_mult[21] ));
 sg13g2_nor2_1 _17369_ (.A(_10409_),
    .B(_10553_),
    .Y(_10554_));
 sg13g2_a22oi_1 _17370_ (.Y(_10555_),
    .B1(net882),
    .B2(\cpu.ex.r_stmp[5] ),
    .A2(_10487_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_nor2_1 _17371_ (.A(net669),
    .B(_10555_),
    .Y(_10556_));
 sg13g2_buf_1 _17372_ (.A(net1037),
    .X(_10557_));
 sg13g2_buf_1 _17373_ (.A(net881),
    .X(_10558_));
 sg13g2_o21ai_1 _17374_ (.B1(net756),
    .Y(_10559_),
    .A1(_10554_),
    .A2(_10556_));
 sg13g2_nand4_1 _17375_ (.B(_10546_),
    .C(_10550_),
    .A(_10544_),
    .Y(_10560_),
    .D(_10559_));
 sg13g2_inv_1 _17376_ (.Y(_10561_),
    .A(_10026_));
 sg13g2_nand2_1 _17377_ (.Y(_10562_),
    .A(_10561_),
    .B(net538));
 sg13g2_o21ai_1 _17378_ (.B1(_10562_),
    .Y(_10563_),
    .A1(net538),
    .A2(_10560_));
 sg13g2_nor3_1 _17379_ (.A(_10535_),
    .B(_10537_),
    .C(_10563_),
    .Y(_10564_));
 sg13g2_a21o_1 _17380_ (.A2(net228),
    .A1(_10531_),
    .B1(_10564_),
    .X(_10565_));
 sg13g2_buf_8 _17381_ (.A(_10565_),
    .X(_10566_));
 sg13g2_a21oi_1 _17382_ (.A1(_08318_),
    .A2(_08358_),
    .Y(_10567_),
    .B1(_10386_));
 sg13g2_inv_2 _17383_ (.Y(_10568_),
    .A(net1037));
 sg13g2_mux2_1 _17384_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_9[4] ),
    .S(net1034),
    .X(_10569_));
 sg13g2_nand3_1 _17385_ (.B(_10423_),
    .C(_10569_),
    .A(_10568_),
    .Y(_10570_));
 sg13g2_nand2b_1 _17386_ (.Y(_10571_),
    .B(net1037),
    .A_N(_00264_));
 sg13g2_nand2b_1 _17387_ (.Y(_10572_),
    .B(\cpu.ex.r_11[4] ),
    .A_N(net1036));
 sg13g2_nand3_1 _17388_ (.B(net887),
    .C(net886),
    .A(net1038),
    .Y(_10573_));
 sg13g2_a21o_1 _17389_ (.A2(_10572_),
    .A1(_10571_),
    .B1(_10573_),
    .X(_10574_));
 sg13g2_nand3b_1 _17390_ (.B(net886),
    .C(\cpu.ex.r_12[4] ),
    .Y(_10575_),
    .A_N(net888));
 sg13g2_nand3b_1 _17391_ (.B(\cpu.ex.r_stmp[4] ),
    .C(net888),
    .Y(_10576_),
    .A_N(net886));
 sg13g2_nand2b_1 _17392_ (.Y(_10577_),
    .B(net1037),
    .A_N(net887));
 sg13g2_a21o_1 _17393_ (.A2(_10576_),
    .A1(_10575_),
    .B1(_10577_),
    .X(_10578_));
 sg13g2_nand3_1 _17394_ (.B(_10574_),
    .C(_10578_),
    .A(_10570_),
    .Y(_10579_));
 sg13g2_a22oi_1 _17395_ (.Y(_10580_),
    .B1(_10448_),
    .B2(_08311_),
    .A2(_10418_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_nand3b_1 _17396_ (.B(net886),
    .C(\cpu.ex.r_8[4] ),
    .Y(_10581_),
    .A_N(_10403_));
 sg13g2_buf_1 _17397_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10582_));
 sg13g2_nand3b_1 _17398_ (.B(_10582_),
    .C(net888),
    .Y(_10583_),
    .A_N(net886));
 sg13g2_or2_1 _17399_ (.X(_10584_),
    .B(net1036),
    .A(_10415_));
 sg13g2_a21o_1 _17400_ (.A2(_10583_),
    .A1(_10581_),
    .B1(_10584_),
    .X(_10585_));
 sg13g2_o21ai_1 _17401_ (.B1(_10585_),
    .Y(_10586_),
    .A1(_10405_),
    .A2(_10580_));
 sg13g2_mux2_1 _17402_ (.A0(\cpu.ex.r_10[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(net1036),
    .X(_10587_));
 sg13g2_mux2_1 _17403_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(\cpu.ex.r_mult[20] ),
    .S(net1036),
    .X(_10588_));
 sg13g2_a22oi_1 _17404_ (.Y(_10589_),
    .B1(_10588_),
    .B2(_10552_),
    .A2(_10587_),
    .A1(net671));
 sg13g2_nor2_1 _17405_ (.A(_10409_),
    .B(_10589_),
    .Y(_10590_));
 sg13g2_nor4_1 _17406_ (.A(_10400_),
    .B(_10579_),
    .C(_10586_),
    .D(_10590_),
    .Y(_10591_));
 sg13g2_a21oi_2 _17407_ (.B1(_10591_),
    .Y(_10592_),
    .A2(_10400_),
    .A1(net904));
 sg13g2_nand4_1 _17408_ (.B(_08452_),
    .C(_10567_),
    .A(net490),
    .Y(_10593_),
    .D(_10592_));
 sg13g2_a21o_1 _17409_ (.A2(_08392_),
    .A1(_08378_),
    .B1(_08396_),
    .X(_10594_));
 sg13g2_buf_2 _17410_ (.A(_10594_),
    .X(_10595_));
 sg13g2_and4_1 _17411_ (.A(_08410_),
    .B(_08422_),
    .C(_08439_),
    .D(_08450_),
    .X(_10596_));
 sg13g2_nor2b_1 _17412_ (.A(_08488_),
    .B_N(net1039),
    .Y(_10597_));
 sg13g2_and2_1 _17413_ (.A(_10369_),
    .B(_10597_),
    .X(_10598_));
 sg13g2_o21ai_1 _17414_ (.B1(_10598_),
    .Y(_10599_),
    .A1(_10595_),
    .A2(_10596_));
 sg13g2_o21ai_1 _17415_ (.B1(net1039),
    .Y(_10600_),
    .A1(_10369_),
    .A2(_10386_));
 sg13g2_a22oi_1 _17416_ (.Y(_10601_),
    .B1(_10592_),
    .B2(_10600_),
    .A2(_10597_),
    .A1(_10388_));
 sg13g2_and3_1 _17417_ (.X(_10602_),
    .A(_10593_),
    .B(_10599_),
    .C(_10601_));
 sg13g2_buf_2 _17418_ (.A(_10602_),
    .X(_10603_));
 sg13g2_xor2_1 _17419_ (.B(_09385_),
    .A(net1142),
    .X(_10604_));
 sg13g2_and2_1 _17420_ (.A(net622),
    .B(_10604_),
    .X(_10605_));
 sg13g2_buf_2 _17421_ (.A(_10605_),
    .X(_10606_));
 sg13g2_nand2_1 _17422_ (.Y(_10607_),
    .A(_09386_),
    .B(_10606_));
 sg13g2_a21oi_1 _17423_ (.A1(_09384_),
    .A2(_10603_),
    .Y(_10608_),
    .B1(_10607_));
 sg13g2_a22oi_1 _17424_ (.Y(_10609_),
    .B1(_10566_),
    .B2(_10608_),
    .A2(_10530_),
    .A1(_10474_));
 sg13g2_buf_2 _17425_ (.A(_10609_),
    .X(_10610_));
 sg13g2_nand3_1 _17426_ (.B(net622),
    .C(_10527_),
    .A(net1142),
    .Y(_10611_));
 sg13g2_buf_1 _17427_ (.A(_00297_),
    .X(_10612_));
 sg13g2_and3_1 _17428_ (.X(_10613_),
    .A(net1142),
    .B(_09386_),
    .C(net622));
 sg13g2_buf_1 _17429_ (.A(_10613_),
    .X(_10614_));
 sg13g2_nand3b_1 _17430_ (.B(_10614_),
    .C(_09385_),
    .Y(_10615_),
    .A_N(_10612_));
 sg13g2_o21ai_1 _17431_ (.B1(_10615_),
    .Y(_10616_),
    .A1(_00299_),
    .A2(_10611_));
 sg13g2_inv_1 _17432_ (.Y(_10617_),
    .A(_10616_));
 sg13g2_and2_1 _17433_ (.A(_09385_),
    .B(_10614_),
    .X(_10618_));
 sg13g2_inv_2 _17434_ (.Y(_10619_),
    .A(_09224_));
 sg13g2_buf_2 _17435_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10620_));
 sg13g2_a22oi_1 _17436_ (.Y(_10621_),
    .B1(net882),
    .B2(_10620_),
    .A2(_10487_),
    .A1(\cpu.ex.r_13[6] ));
 sg13g2_nor2b_1 _17437_ (.A(_10621_),
    .B_N(_10441_),
    .Y(_10622_));
 sg13g2_a22oi_1 _17438_ (.Y(_10623_),
    .B1(net760),
    .B2(\cpu.ex.r_10[6] ),
    .A2(net883),
    .A1(\cpu.ex.r_stmp[6] ));
 sg13g2_buf_1 _17439_ (.A(_10427_),
    .X(_10624_));
 sg13g2_nand2b_1 _17440_ (.Y(_10625_),
    .B(net668),
    .A_N(_10623_));
 sg13g2_a22oi_1 _17441_ (.Y(_10626_),
    .B1(_10513_),
    .B2(\cpu.ex.r_lr[6] ),
    .A2(_10467_),
    .A1(\cpu.ex.r_12[6] ));
 sg13g2_inv_1 _17442_ (.Y(_10627_),
    .A(_00266_));
 sg13g2_mux2_1 _17443_ (.A0(_10627_),
    .A1(\cpu.ex.r_14[6] ),
    .S(net759),
    .X(_10628_));
 sg13g2_and3_1 _17444_ (.X(_10629_),
    .A(net1038),
    .B(net1034),
    .C(net1128));
 sg13g2_a22oi_1 _17445_ (.Y(_10630_),
    .B1(_10457_),
    .B2(\cpu.ex.r_epc[6] ),
    .A2(_10629_),
    .A1(_10628_));
 sg13g2_nand2_1 _17446_ (.Y(_10631_),
    .A(\cpu.ex.r_sp[6] ),
    .B(_10514_));
 sg13g2_nand4_1 _17447_ (.B(_10626_),
    .C(_10630_),
    .A(_10625_),
    .Y(_10632_),
    .D(_10631_));
 sg13g2_buf_1 _17448_ (.A(_10409_),
    .X(_10633_));
 sg13g2_mux2_1 _17449_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_9[6] ),
    .S(_10540_),
    .X(_10634_));
 sg13g2_and2_1 _17450_ (.A(net1038),
    .B(net1035),
    .X(_10635_));
 sg13g2_buf_2 _17451_ (.A(_10635_),
    .X(_10636_));
 sg13g2_a22oi_1 _17452_ (.Y(_10637_),
    .B1(_10636_),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10634_),
    .A1(_10633_));
 sg13g2_nor2b_1 _17453_ (.A(_10637_),
    .B_N(net760),
    .Y(_10638_));
 sg13g2_nor4_1 _17454_ (.A(net538),
    .B(_10622_),
    .C(_10632_),
    .D(_10638_),
    .Y(_10639_));
 sg13g2_a21oi_2 _17455_ (.B1(_10639_),
    .Y(_10640_),
    .A2(net538),
    .A1(_10619_));
 sg13g2_inv_1 _17456_ (.Y(_10641_),
    .A(_10611_));
 sg13g2_a22oi_1 _17457_ (.Y(_10642_),
    .B1(_10471_),
    .B2(_10641_),
    .A2(_10640_),
    .A1(_10618_));
 sg13g2_nor2_1 _17458_ (.A(_10535_),
    .B(_10537_),
    .Y(_10643_));
 sg13g2_mux2_1 _17459_ (.A0(_10617_),
    .A1(_10642_),
    .S(_10643_),
    .X(_10644_));
 sg13g2_inv_2 _17460_ (.Y(_10645_),
    .A(net1151));
 sg13g2_nand3_1 _17461_ (.B(\cpu.ex.r_9[0] ),
    .C(_10451_),
    .A(net761),
    .Y(_10646_));
 sg13g2_nand3_1 _17462_ (.B(net759),
    .C(net883),
    .A(_09242_),
    .Y(_10647_));
 sg13g2_a21oi_1 _17463_ (.A1(_10646_),
    .A2(_10647_),
    .Y(_10648_),
    .B1(net757));
 sg13g2_buf_1 _17464_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10649_));
 sg13g2_a22oi_1 _17465_ (.Y(_10650_),
    .B1(_10498_),
    .B2(\cpu.ex.r_10[0] ),
    .A2(_10552_),
    .A1(_10649_));
 sg13g2_nor2b_1 _17466_ (.A(_10650_),
    .B_N(_10411_),
    .Y(_10651_));
 sg13g2_nand4_1 _17467_ (.B(net884),
    .C(\cpu.ex.r_14[0] ),
    .A(net885),
    .Y(_10652_),
    .D(_10427_));
 sg13g2_buf_1 _17468_ (.A(_10379_),
    .X(_10653_));
 sg13g2_nand4_1 _17469_ (.B(_10568_),
    .C(\cpu.ex.r_8[0] ),
    .A(net885),
    .Y(_10654_),
    .D(net879));
 sg13g2_nand2_1 _17470_ (.Y(_10655_),
    .A(_10652_),
    .B(_10654_));
 sg13g2_nand4_1 _17471_ (.B(_10568_),
    .C(\cpu.ex.r_11[0] ),
    .A(net885),
    .Y(_10656_),
    .D(_10636_));
 sg13g2_nand4_1 _17472_ (.B(net884),
    .C(\cpu.ex.r_12[0] ),
    .A(net885),
    .Y(_10657_),
    .D(net879));
 sg13g2_nand2_1 _17473_ (.Y(_10658_),
    .A(_10656_),
    .B(_10657_));
 sg13g2_nor4_1 _17474_ (.A(_10648_),
    .B(_10651_),
    .C(_10655_),
    .D(_10658_),
    .Y(_10659_));
 sg13g2_and2_1 _17475_ (.A(net886),
    .B(\cpu.ex.r_15[0] ),
    .X(_10660_));
 sg13g2_a21oi_1 _17476_ (.A1(_10421_),
    .A2(\cpu.ex.r_mult[16] ),
    .Y(_10661_),
    .B1(_10660_));
 sg13g2_buf_1 _17477_ (.A(_10423_),
    .X(_10662_));
 sg13g2_and2_1 _17478_ (.A(_10417_),
    .B(\cpu.ex.r_13[0] ),
    .X(_10663_));
 sg13g2_nor2b_1 _17479_ (.A(net885),
    .B_N(\cpu.ex.r_stmp[0] ),
    .Y(_10664_));
 sg13g2_a22oi_1 _17480_ (.Y(_10665_),
    .B1(_10664_),
    .B2(net668),
    .A2(_10663_),
    .A1(net667));
 sg13g2_o21ai_1 _17481_ (.B1(_10665_),
    .Y(_10666_),
    .A1(_10455_),
    .A2(_10661_));
 sg13g2_a21oi_1 _17482_ (.A1(net756),
    .A2(_10666_),
    .Y(_10667_),
    .B1(_10400_));
 sg13g2_a22oi_1 _17483_ (.Y(_10668_),
    .B1(_10659_),
    .B2(_10667_),
    .A2(_10400_),
    .A1(_10645_));
 sg13g2_buf_1 _17484_ (.A(_10668_),
    .X(_10669_));
 sg13g2_nand3_1 _17485_ (.B(net269),
    .C(_10669_),
    .A(net339),
    .Y(_10670_));
 sg13g2_nand2_1 _17486_ (.Y(_10671_),
    .A(_08309_),
    .B(net1039));
 sg13g2_a221oi_1 _17487_ (.B2(_08452_),
    .C1(_10671_),
    .B1(net490),
    .A1(_08354_),
    .Y(_10672_),
    .A2(_08363_));
 sg13g2_and2_1 _17488_ (.A(_10383_),
    .B(_10384_),
    .X(_10673_));
 sg13g2_buf_1 _17489_ (.A(_10673_),
    .X(_10674_));
 sg13g2_a21oi_1 _17490_ (.A1(_08359_),
    .A2(_10674_),
    .Y(_10675_),
    .B1(_10671_));
 sg13g2_nor2_1 _17491_ (.A(_10672_),
    .B(_10675_),
    .Y(_10676_));
 sg13g2_a21o_1 _17492_ (.A2(_10676_),
    .A1(_10670_),
    .B1(_09388_),
    .X(_10677_));
 sg13g2_nand3_1 _17493_ (.B(_10599_),
    .C(_10601_),
    .A(_10593_),
    .Y(_10678_));
 sg13g2_buf_2 _17494_ (.A(_10678_),
    .X(_10679_));
 sg13g2_and2_1 _17495_ (.A(_10614_),
    .B(_10606_),
    .X(_10680_));
 sg13g2_nor3_1 _17496_ (.A(net1142),
    .B(_09385_),
    .C(_09386_),
    .Y(_10681_));
 sg13g2_xnor2_1 _17497_ (.Y(_10682_),
    .A(\cpu.ex.r_mult_off[3] ),
    .B(_10681_));
 sg13g2_nand2_1 _17498_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(net622),
    .B(_10682_));
 sg13g2_a21oi_1 _17499_ (.A1(_10679_),
    .A2(_10680_),
    .Y(_10683_),
    .B1(\cpu.ex.c_mult_off[3] ));
 sg13g2_nand3b_1 _17500_ (.B(net622),
    .C(_10527_),
    .Y(_10684_),
    .A_N(net1142));
 sg13g2_inv_1 _17501_ (.Y(_10685_),
    .A(_10684_));
 sg13g2_a22oi_1 _17502_ (.Y(_10686_),
    .B1(_10442_),
    .B2(\cpu.ex.r_8[1] ),
    .A2(_10441_),
    .A1(\cpu.ex.r_13[1] ));
 sg13g2_nor2_1 _17503_ (.A(_10491_),
    .B(_10686_),
    .Y(_10687_));
 sg13g2_mux2_1 _17504_ (.A0(\cpu.ex.r_prev_ie ),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(_10414_),
    .X(_10688_));
 sg13g2_nand3_1 _17505_ (.B(net883),
    .C(_10688_),
    .A(_10409_),
    .Y(_10689_));
 sg13g2_nand3_1 _17506_ (.B(_10427_),
    .C(_10451_),
    .A(\cpu.ex.r_10[1] ),
    .Y(_10690_));
 sg13g2_mux2_1 _17507_ (.A0(\cpu.ex.r_stmp[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(_10414_),
    .X(_10691_));
 sg13g2_nand3_1 _17508_ (.B(net882),
    .C(_10691_),
    .A(net884),
    .Y(_10692_));
 sg13g2_nor2b_1 _17509_ (.A(_00261_),
    .B_N(net1035),
    .Y(_10693_));
 sg13g2_nor2b_1 _17510_ (.A(net887),
    .B_N(\cpu.ex.r_14[1] ),
    .Y(_10694_));
 sg13g2_o21ai_1 _17511_ (.B1(_10629_),
    .Y(_10695_),
    .A1(_10693_),
    .A2(_10694_));
 sg13g2_nand4_1 _17512_ (.B(_10690_),
    .C(_10692_),
    .A(_10689_),
    .Y(_10696_),
    .D(_10695_));
 sg13g2_nand3_1 _17513_ (.B(\cpu.ex.r_12[1] ),
    .C(_10487_),
    .A(net884),
    .Y(_10697_));
 sg13g2_buf_1 _17514_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10698_));
 sg13g2_nand3_1 _17515_ (.B(_10698_),
    .C(_10376_),
    .A(_10403_),
    .Y(_10699_));
 sg13g2_a21oi_1 _17516_ (.A1(_10697_),
    .A2(_10699_),
    .Y(_10700_),
    .B1(net761));
 sg13g2_mux4_1 _17517_ (.S0(net1038),
    .A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_epc[1] ),
    .A2(\cpu.ex.r_9[1] ),
    .A3(\cpu.ex.r_11[1] ),
    .S1(net886),
    .X(_10701_));
 sg13g2_and3_1 _17518_ (.X(_10702_),
    .A(net761),
    .B(_10568_),
    .C(_10701_));
 sg13g2_nor4_1 _17519_ (.A(_10687_),
    .B(_10696_),
    .C(_10700_),
    .D(_10702_),
    .Y(_10703_));
 sg13g2_nor2_1 _17520_ (.A(_09238_),
    .B(_10480_),
    .Y(_10704_));
 sg13g2_a21oi_2 _17521_ (.B1(_10704_),
    .Y(_10705_),
    .A2(_10703_),
    .A1(_10480_));
 sg13g2_nand4_1 _17522_ (.B(_08452_),
    .C(_10567_),
    .A(_08398_),
    .Y(_10706_),
    .D(_10705_));
 sg13g2_nand2_1 _17523_ (.Y(_10707_),
    .A(_10600_),
    .B(_10705_));
 sg13g2_nor2b_1 _17524_ (.A(_00200_),
    .B_N(_10368_),
    .Y(_10708_));
 sg13g2_nand2_1 _17525_ (.Y(_10709_),
    .A(_10388_),
    .B(_10708_));
 sg13g2_and2_1 _17526_ (.A(_10369_),
    .B(_10708_),
    .X(_10710_));
 sg13g2_o21ai_1 _17527_ (.B1(_10710_),
    .Y(_10711_),
    .A1(_10595_),
    .A2(_10596_));
 sg13g2_nand4_1 _17528_ (.B(_10707_),
    .C(_10709_),
    .A(_10706_),
    .Y(_10712_),
    .D(_10711_));
 sg13g2_buf_2 _17529_ (.A(_10712_),
    .X(_10713_));
 sg13g2_buf_1 _17530_ (.A(_00296_),
    .X(_10714_));
 sg13g2_inv_2 _17531_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_10606_));
 sg13g2_xnor2_1 _17532_ (.Y(_10715_),
    .A(_09386_),
    .B(_10526_));
 sg13g2_o21ai_1 _17533_ (.B1(net622),
    .Y(_10716_),
    .A1(net1142),
    .A2(_10715_));
 sg13g2_nand2_1 _17534_ (.Y(_10717_),
    .A(\cpu.ex.c_mult_off[1] ),
    .B(_10716_));
 sg13g2_nor2_1 _17535_ (.A(_10714_),
    .B(_10717_),
    .Y(_10718_));
 sg13g2_nand2_1 _17536_ (.Y(_10719_),
    .A(net758),
    .B(net881));
 sg13g2_nor2_1 _17537_ (.A(_10719_),
    .B(_10459_),
    .Y(_10720_));
 sg13g2_buf_1 _17538_ (.A(\cpu.dec.user_io ),
    .X(_10721_));
 sg13g2_a22oi_1 _17539_ (.Y(_10722_),
    .B1(_10636_),
    .B2(\cpu.ex.r_mult[23] ),
    .A2(net879),
    .A1(_10721_));
 sg13g2_nor2b_1 _17540_ (.A(_10722_),
    .B_N(_10435_),
    .Y(_10723_));
 sg13g2_a221oi_1 _17541_ (.B2(\cpu.ex.r_13[7] ),
    .C1(_10723_),
    .B1(_10720_),
    .A1(\cpu.ex.r_lr[7] ),
    .Y(_10724_),
    .A2(_10513_));
 sg13g2_buf_1 _17542_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10725_));
 sg13g2_mux2_1 _17543_ (.A0(\cpu.ex.r_12[7] ),
    .A1(\cpu.ex.r_14[7] ),
    .S(net888),
    .X(_10726_));
 sg13g2_nand3_1 _17544_ (.B(_10499_),
    .C(_10726_),
    .A(_10431_),
    .Y(_10727_));
 sg13g2_o21ai_1 _17545_ (.B1(_10727_),
    .Y(_10728_),
    .A1(_00267_),
    .A2(_10517_));
 sg13g2_a221oi_1 _17546_ (.B2(_10725_),
    .C1(_10728_),
    .B1(_10514_),
    .A1(\cpu.ex.r_epc[7] ),
    .Y(_10729_),
    .A2(_10457_));
 sg13g2_mux2_1 _17547_ (.A0(\cpu.ex.r_10[7] ),
    .A1(\cpu.ex.r_11[7] ),
    .S(_10432_),
    .X(_10730_));
 sg13g2_a22oi_1 _17548_ (.Y(_10731_),
    .B1(_10730_),
    .B2(_10509_),
    .A2(net667),
    .A1(\cpu.ex.r_9[7] ));
 sg13g2_inv_1 _17549_ (.Y(_10732_),
    .A(_10731_));
 sg13g2_buf_1 _17550_ (.A(_10568_),
    .X(_10733_));
 sg13g2_nand3_1 _17551_ (.B(\cpu.ex.r_8[7] ),
    .C(_10487_),
    .A(net755),
    .Y(_10734_));
 sg13g2_nand3_1 _17552_ (.B(\cpu.ex.r_stmp[7] ),
    .C(net882),
    .A(net762),
    .Y(_10735_));
 sg13g2_nand2_1 _17553_ (.Y(_10736_),
    .A(_10734_),
    .B(_10735_));
 sg13g2_a22oi_1 _17554_ (.Y(_10737_),
    .B1(_10736_),
    .B2(net759),
    .A2(_10732_),
    .A1(net760));
 sg13g2_nand4_1 _17555_ (.B(_10724_),
    .C(_10729_),
    .A(_10480_),
    .Y(_10738_),
    .D(_10737_));
 sg13g2_o21ai_1 _17556_ (.B1(_10738_),
    .Y(_10739_),
    .A1(_09228_),
    .A2(net539));
 sg13g2_buf_1 _17557_ (.A(_10739_),
    .X(_10740_));
 sg13g2_nor4_1 _17558_ (.A(_10535_),
    .B(_10537_),
    .C(_10717_),
    .D(_10740_),
    .Y(_10741_));
 sg13g2_a221oi_1 _17559_ (.B2(net228),
    .C1(_10741_),
    .B1(_10718_),
    .A1(_10685_),
    .Y(_10742_),
    .A2(_10713_));
 sg13g2_and4_1 _17560_ (.A(_10644_),
    .B(_10677_),
    .C(_10683_),
    .D(_10742_),
    .X(_10743_));
 sg13g2_buf_2 _17561_ (.A(_10743_),
    .X(_10744_));
 sg13g2_inv_1 _17562_ (.Y(_10745_),
    .A(_00194_));
 sg13g2_nand2_1 _17563_ (.Y(_10746_),
    .A(_00196_),
    .B(_10606_));
 sg13g2_o21ai_1 _17564_ (.B1(_10746_),
    .Y(_10747_),
    .A1(_10745_),
    .A2(_10606_));
 sg13g2_o21ai_1 _17565_ (.B1(_10747_),
    .Y(_10748_),
    .A1(_10535_),
    .A2(_10537_));
 sg13g2_buf_1 _17566_ (.A(net788),
    .X(_10749_));
 sg13g2_nand3b_1 _17567_ (.B(\cpu.ex.r_epc[15] ),
    .C(net761),
    .Y(_10750_),
    .A_N(net1037));
 sg13g2_nand3b_1 _17568_ (.B(_10430_),
    .C(\cpu.ex.r_stmp[15] ),
    .Y(_10751_),
    .A_N(net887));
 sg13g2_a21o_1 _17569_ (.A2(_10751_),
    .A1(_10750_),
    .B1(_10506_),
    .X(_10752_));
 sg13g2_mux2_1 _17570_ (.A0(\cpu.ex.r_10[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(_10404_),
    .X(_10753_));
 sg13g2_nand2_1 _17571_ (.Y(_10754_),
    .A(net671),
    .B(_10753_));
 sg13g2_nand3_1 _17572_ (.B(_10752_),
    .C(_10754_),
    .A(net757),
    .Y(_10755_));
 sg13g2_nand3_1 _17573_ (.B(\cpu.ex.r_lr[15] ),
    .C(_10376_),
    .A(net669),
    .Y(_10756_));
 sg13g2_nand3_1 _17574_ (.B(\cpu.ex.r_12[15] ),
    .C(net671),
    .A(_10557_),
    .Y(_10757_));
 sg13g2_nand3_1 _17575_ (.B(_10756_),
    .C(_10757_),
    .A(net880),
    .Y(_10758_));
 sg13g2_mux2_1 _17576_ (.A0(\cpu.ex.r_9[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .S(_10404_),
    .X(_10759_));
 sg13g2_a22oi_1 _17577_ (.Y(_10760_),
    .B1(_10759_),
    .B2(_10506_),
    .A2(net883),
    .A1(_10308_));
 sg13g2_nand3_1 _17578_ (.B(\cpu.ex.r_11[15] ),
    .C(net760),
    .A(net757),
    .Y(_10761_));
 sg13g2_o21ai_1 _17579_ (.B1(_10761_),
    .Y(_10762_),
    .A1(_10509_),
    .A2(_10760_));
 sg13g2_a22oi_1 _17580_ (.Y(_10763_),
    .B1(_10446_),
    .B2(_10322_),
    .A2(_10487_),
    .A1(\cpu.ex.r_8[15] ));
 sg13g2_mux2_1 _17581_ (.A0(\cpu.ex.r_mult[31] ),
    .A1(\cpu.ex.r_15[15] ),
    .S(net885),
    .X(_10764_));
 sg13g2_nand3_1 _17582_ (.B(_10636_),
    .C(_10764_),
    .A(net762),
    .Y(_10765_));
 sg13g2_o21ai_1 _17583_ (.B1(_10765_),
    .Y(_10766_),
    .A1(_10584_),
    .A2(_10763_));
 sg13g2_a221oi_1 _17584_ (.B2(net669),
    .C1(_10766_),
    .B1(_10762_),
    .A1(_10755_),
    .Y(_10767_),
    .A2(_10758_));
 sg13g2_mux2_1 _17585_ (.A0(net666),
    .A1(_10767_),
    .S(_10480_),
    .X(_10768_));
 sg13g2_nand2b_1 _17586_ (.Y(_10769_),
    .B(\cpu.ex.c_mult_off[1] ),
    .A_N(_10768_));
 sg13g2_nand2_1 _17587_ (.Y(_10770_),
    .A(net1093),
    .B(net538));
 sg13g2_a22oi_1 _17588_ (.Y(_10771_),
    .B1(_10636_),
    .B2(\cpu.ex.r_11[13] ),
    .A2(_10653_),
    .A1(\cpu.ex.r_8[13] ));
 sg13g2_inv_1 _17589_ (.Y(_10772_),
    .A(_10771_));
 sg13g2_nand2_1 _17590_ (.Y(_10773_),
    .A(_10568_),
    .B(\cpu.ex.r_10[13] ));
 sg13g2_nand3_1 _17591_ (.B(\cpu.ex.r_13[13] ),
    .C(_10662_),
    .A(net762),
    .Y(_10774_));
 sg13g2_o21ai_1 _17592_ (.B1(_10774_),
    .Y(_10775_),
    .A1(_10483_),
    .A2(_10773_));
 sg13g2_inv_1 _17593_ (.Y(_10776_),
    .A(_00273_));
 sg13g2_a22oi_1 _17594_ (.Y(_10777_),
    .B1(_10636_),
    .B2(_10776_),
    .A2(_10653_),
    .A1(\cpu.ex.r_12[13] ));
 sg13g2_nor2_1 _17595_ (.A(_10719_),
    .B(_10777_),
    .Y(_10778_));
 sg13g2_a221oi_1 _17596_ (.B2(net670),
    .C1(_10778_),
    .B1(_10775_),
    .A1(net760),
    .Y(_10779_),
    .A2(_10772_));
 sg13g2_mux2_1 _17597_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(\cpu.ex.r_9[13] ),
    .S(_10425_),
    .X(_10780_));
 sg13g2_a22oi_1 _17598_ (.Y(_10781_),
    .B1(_10780_),
    .B2(net880),
    .A2(_10446_),
    .A1(\cpu.ex.r_epc[13] ));
 sg13g2_nor2_1 _17599_ (.A(net759),
    .B(_10781_),
    .Y(_10782_));
 sg13g2_buf_1 _17600_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10783_));
 sg13g2_nor2_1 _17601_ (.A(net758),
    .B(_10483_),
    .Y(_10784_));
 sg13g2_and2_1 _17602_ (.A(_10783_),
    .B(_10784_),
    .X(_10785_));
 sg13g2_o21ai_1 _17603_ (.B1(net755),
    .Y(_10786_),
    .A1(_10782_),
    .A2(_10785_));
 sg13g2_a22oi_1 _17604_ (.Y(_10787_),
    .B1(net667),
    .B2(\cpu.ex.mmu_read[13] ),
    .A2(net668),
    .A1(\cpu.ex.r_stmp[13] ));
 sg13g2_nor2_1 _17605_ (.A(net670),
    .B(_10787_),
    .Y(_10788_));
 sg13g2_buf_2 _17606_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10789_));
 sg13g2_a22oi_1 _17607_ (.Y(_10790_),
    .B1(net671),
    .B2(\cpu.ex.r_14[13] ),
    .A2(_10552_),
    .A1(_10789_));
 sg13g2_nor2_1 _17608_ (.A(net880),
    .B(_10790_),
    .Y(_10791_));
 sg13g2_o21ai_1 _17609_ (.B1(net756),
    .Y(_10792_),
    .A1(_10788_),
    .A2(_10791_));
 sg13g2_nand4_1 _17610_ (.B(_10779_),
    .C(_10786_),
    .A(net539),
    .Y(_10793_),
    .D(_10792_));
 sg13g2_nand3_1 _17611_ (.B(_10770_),
    .C(_10793_),
    .A(_10606_),
    .Y(_10794_));
 sg13g2_nand4_1 _17612_ (.B(net269),
    .C(_10769_),
    .A(net339),
    .Y(_10795_),
    .D(_10794_));
 sg13g2_and3_1 _17613_ (.X(_10796_),
    .A(_10716_),
    .B(_10748_),
    .C(_10795_));
 sg13g2_buf_1 _17614_ (.A(_10796_),
    .X(_10797_));
 sg13g2_buf_8 _17615_ (.A(_10535_),
    .X(_10798_));
 sg13g2_buf_8 _17616_ (.A(_10537_),
    .X(_10799_));
 sg13g2_nor2_1 _17617_ (.A(_09226_),
    .B(net539),
    .Y(_10800_));
 sg13g2_nor2_1 _17618_ (.A(_10421_),
    .B(_10459_),
    .Y(_10801_));
 sg13g2_buf_1 _17619_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10802_));
 sg13g2_a22oi_1 _17620_ (.Y(_10803_),
    .B1(_10784_),
    .B2(_10802_),
    .A2(_10801_),
    .A1(\cpu.ex.r_9[8] ));
 sg13g2_a221oi_1 _17621_ (.B2(\cpu.ex.r_stmp[8] ),
    .C1(net755),
    .B1(_10784_),
    .A1(\cpu.ex.r_13[8] ),
    .Y(_10804_),
    .A2(_10801_));
 sg13g2_a21oi_1 _17622_ (.A1(_10733_),
    .A2(_10803_),
    .Y(_10805_),
    .B1(_10804_));
 sg13g2_and2_1 _17623_ (.A(net762),
    .B(net879),
    .X(_10806_));
 sg13g2_a22oi_1 _17624_ (.Y(_10807_),
    .B1(_10806_),
    .B2(\cpu.ex.r_12[8] ),
    .A2(_10508_),
    .A1(\cpu.ex.r_11[8] ));
 sg13g2_nand3_1 _17625_ (.B(\cpu.ex.r_14[8] ),
    .C(net671),
    .A(net762),
    .Y(_10808_));
 sg13g2_nand3_1 _17626_ (.B(\cpu.ex.r_epc[8] ),
    .C(_10376_),
    .A(_10540_),
    .Y(_10809_));
 sg13g2_a21o_1 _17627_ (.A2(_10809_),
    .A1(_10808_),
    .B1(_10633_),
    .X(_10810_));
 sg13g2_o21ai_1 _17628_ (.B1(_10810_),
    .Y(_10811_),
    .A1(_10421_),
    .A2(_10807_));
 sg13g2_a22oi_1 _17629_ (.Y(_10812_),
    .B1(_10543_),
    .B2(\cpu.ex.r_10[8] ),
    .A2(_10513_),
    .A1(\cpu.ex.r_lr[8] ));
 sg13g2_nand3_1 _17630_ (.B(net879),
    .C(_10484_),
    .A(\cpu.ex.r_8[8] ),
    .Y(_10813_));
 sg13g2_nand3_1 _17631_ (.B(_10636_),
    .C(net883),
    .A(\cpu.ex.r_mult[24] ),
    .Y(_10814_));
 sg13g2_or2_1 _17632_ (.X(_10815_),
    .B(_10517_),
    .A(_00268_));
 sg13g2_nand4_1 _17633_ (.B(_10813_),
    .C(_10814_),
    .A(_10812_),
    .Y(_10816_),
    .D(_10815_));
 sg13g2_nor4_2 _17634_ (.A(net538),
    .B(_10805_),
    .C(_10811_),
    .Y(_10817_),
    .D(_10816_));
 sg13g2_nor3_1 _17635_ (.A(_09388_),
    .B(_10800_),
    .C(_10817_),
    .Y(_10818_));
 sg13g2_buf_2 _17636_ (.A(\cpu.addr[9] ),
    .X(_10819_));
 sg13g2_a22oi_1 _17637_ (.Y(_10820_),
    .B1(_10484_),
    .B2(\cpu.ex.r_11[9] ),
    .A2(net883),
    .A1(\cpu.ex.r_mult[25] ));
 sg13g2_nand2b_1 _17638_ (.Y(_10821_),
    .B(_10636_),
    .A_N(_10820_));
 sg13g2_inv_1 _17639_ (.Y(_10822_),
    .A(\cpu.ex.r_sp[9] ));
 sg13g2_nand3_1 _17640_ (.B(net881),
    .C(\cpu.ex.r_14[9] ),
    .A(net758),
    .Y(_10823_));
 sg13g2_o21ai_1 _17641_ (.B1(_10823_),
    .Y(_10824_),
    .A1(_10822_),
    .A2(_10454_));
 sg13g2_mux2_1 _17642_ (.A0(\cpu.ex.r_9[9] ),
    .A1(\cpu.ex.r_13[9] ),
    .S(net881),
    .X(_10825_));
 sg13g2_nor2_1 _17643_ (.A(_00269_),
    .B(_10517_),
    .Y(_10826_));
 sg13g2_a221oi_1 _17644_ (.B2(_10801_),
    .C1(_10826_),
    .B1(_10825_),
    .A1(net668),
    .Y(_10827_),
    .A2(_10824_));
 sg13g2_nand3_1 _17645_ (.B(\cpu.ex.r_stmp[9] ),
    .C(_10624_),
    .A(_10431_),
    .Y(_10828_));
 sg13g2_nand3_1 _17646_ (.B(\cpu.ex.r_lr[9] ),
    .C(net667),
    .A(_10733_),
    .Y(_10829_));
 sg13g2_a21o_1 _17647_ (.A2(_10829_),
    .A1(_10828_),
    .B1(_10507_),
    .X(_10830_));
 sg13g2_mux2_1 _17648_ (.A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_12[9] ),
    .S(_10430_),
    .X(_10831_));
 sg13g2_and3_1 _17649_ (.X(_10832_),
    .A(net758),
    .B(net879),
    .C(_10831_));
 sg13g2_a221oi_1 _17650_ (.B2(\cpu.ex.r_10[9] ),
    .C1(_10832_),
    .B1(_10543_),
    .A1(\cpu.ex.r_epc[9] ),
    .Y(_10833_),
    .A2(_10457_));
 sg13g2_nand4_1 _17651_ (.B(_10827_),
    .C(_10830_),
    .A(_10821_),
    .Y(_10834_),
    .D(_10833_));
 sg13g2_mux2_1 _17652_ (.A0(_10819_),
    .A1(_10834_),
    .S(_10481_),
    .X(_10835_));
 sg13g2_and2_1 _17653_ (.A(_10685_),
    .B(_10835_),
    .X(_10836_));
 sg13g2_nor4_1 _17654_ (.A(_10798_),
    .B(_10799_),
    .C(_10818_),
    .D(_10836_),
    .Y(_10837_));
 sg13g2_inv_1 _17655_ (.Y(_10838_),
    .A(_00294_));
 sg13g2_nor2_1 _17656_ (.A(_00295_),
    .B(_09388_),
    .Y(_10839_));
 sg13g2_a221oi_1 _17657_ (.B2(_10838_),
    .C1(_10839_),
    .B1(_10685_),
    .A1(_10477_),
    .Y(_10840_),
    .A2(_10478_));
 sg13g2_o21ai_1 _17658_ (.B1(\cpu.ex.c_mult_off[3] ),
    .Y(_10841_),
    .A1(_10837_),
    .A2(_10840_));
 sg13g2_inv_1 _17659_ (.Y(_10842_),
    .A(_00195_));
 sg13g2_nand2_1 _17660_ (.Y(_10843_),
    .A(_00291_),
    .B(_10606_));
 sg13g2_o21ai_1 _17661_ (.B1(_10843_),
    .Y(_10844_),
    .A1(_10842_),
    .A2(_10606_));
 sg13g2_nor2b_1 _17662_ (.A(_10844_),
    .B_N(_10614_),
    .Y(_10845_));
 sg13g2_inv_1 _17663_ (.Y(_10846_),
    .A(_00272_));
 sg13g2_mux4_1 _17664_ (.S0(_10502_),
    .A0(_10846_),
    .A1(\cpu.ex.r_14[12] ),
    .A2(\cpu.ex.r_13[12] ),
    .A3(\cpu.ex.r_12[12] ),
    .S1(net880),
    .X(_10847_));
 sg13g2_mux4_1 _17665_ (.S0(_10432_),
    .A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .A2(\cpu.ex.r_10[12] ),
    .A3(\cpu.ex.r_11[12] ),
    .S1(net757),
    .X(_10848_));
 sg13g2_or2_1 _17666_ (.X(_10849_),
    .B(_10848_),
    .A(_10558_));
 sg13g2_o21ai_1 _17667_ (.B1(_10849_),
    .Y(_10850_),
    .A1(net755),
    .A2(_10847_));
 sg13g2_buf_2 _17668_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10851_));
 sg13g2_buf_8 _17669_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10852_));
 sg13g2_mux4_1 _17670_ (.S0(net757),
    .A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_epc[12] ),
    .A2(_10851_),
    .A3(_10852_),
    .S1(net756),
    .X(_10853_));
 sg13g2_buf_1 _17671_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10854_));
 sg13g2_mux2_1 _17672_ (.A0(_10854_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net756),
    .X(_10855_));
 sg13g2_a221oi_1 _17673_ (.B2(_10624_),
    .C1(net670),
    .B1(_10855_),
    .A1(net669),
    .Y(_10856_),
    .A2(_10853_));
 sg13g2_a21oi_1 _17674_ (.A1(_10507_),
    .A2(_10850_),
    .Y(_10857_),
    .B1(_10856_));
 sg13g2_nand3_1 _17675_ (.B(\cpu.ex.r_14[14] ),
    .C(net668),
    .A(net756),
    .Y(_10858_));
 sg13g2_nand3_1 _17676_ (.B(\cpu.ex.r_9[14] ),
    .C(_10662_),
    .A(net755),
    .Y(_10859_));
 sg13g2_a21oi_1 _17677_ (.A1(_10858_),
    .A2(_10859_),
    .Y(_10860_),
    .B1(_10421_));
 sg13g2_buf_1 _17678_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10861_));
 sg13g2_mux2_1 _17679_ (.A0(_10861_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(_10557_),
    .X(_10862_));
 sg13g2_a22oi_1 _17680_ (.Y(_10863_),
    .B1(_10862_),
    .B2(net759),
    .A2(_10441_),
    .A1(\cpu.ex.r_mult[30] ));
 sg13g2_nor2b_1 _17681_ (.A(_10863_),
    .B_N(net882),
    .Y(_10864_));
 sg13g2_nand2_1 _17682_ (.Y(_10865_),
    .A(net880),
    .B(net755));
 sg13g2_a22oi_1 _17683_ (.Y(_10866_),
    .B1(_10499_),
    .B2(\cpu.ex.r_8[14] ),
    .A2(_10552_),
    .A1(\cpu.ex.r_lr[14] ));
 sg13g2_mux2_1 _17684_ (.A0(\cpu.ex.r_10[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net669),
    .X(_10867_));
 sg13g2_a22oi_1 _17685_ (.Y(_10868_),
    .B1(_10433_),
    .B2(_10867_),
    .A2(_10467_),
    .A1(\cpu.ex.r_12[14] ));
 sg13g2_o21ai_1 _17686_ (.B1(_10868_),
    .Y(_10869_),
    .A1(_10865_),
    .A2(_10866_));
 sg13g2_inv_1 _17687_ (.Y(_10870_),
    .A(_00274_));
 sg13g2_a22oi_1 _17688_ (.Y(_10871_),
    .B1(_10465_),
    .B2(_10870_),
    .A2(_10376_),
    .A1(\cpu.ex.r_epc[14] ));
 sg13g2_buf_2 _17689_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10872_));
 sg13g2_mux2_1 _17690_ (.A0(_10872_),
    .A1(\cpu.ex.r_13[14] ),
    .S(_10425_),
    .X(_10873_));
 sg13g2_nand2b_1 _17691_ (.Y(_10874_),
    .B(_10873_),
    .A_N(_10405_));
 sg13g2_o21ai_1 _17692_ (.B1(_10874_),
    .Y(_10875_),
    .A1(net880),
    .A2(_10871_));
 sg13g2_and2_1 _17693_ (.A(net669),
    .B(_10875_),
    .X(_10876_));
 sg13g2_or4_1 _17694_ (.A(_10860_),
    .B(_10864_),
    .C(_10869_),
    .D(_10876_),
    .X(_10877_));
 sg13g2_mux4_1 _17695_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(net780),
    .A1(net688),
    .A2(_10857_),
    .A3(_10877_),
    .S1(net539),
    .X(_10878_));
 sg13g2_and2_1 _17696_ (.A(_10614_),
    .B(_10878_),
    .X(_10879_));
 sg13g2_mux2_1 _17697_ (.A0(_10845_),
    .A1(_10879_),
    .S(_10643_),
    .X(_10880_));
 sg13g2_inv_2 _17698_ (.Y(_10881_),
    .A(_00293_));
 sg13g2_nor2_1 _17699_ (.A(_00292_),
    .B(_09384_),
    .Y(_10882_));
 sg13g2_a221oi_1 _17700_ (.B2(_10478_),
    .C1(_10882_),
    .B1(_10477_),
    .A1(_10881_),
    .Y(_10883_),
    .A2(_09384_));
 sg13g2_a22oi_1 _17701_ (.Y(_10884_),
    .B1(_10493_),
    .B2(\cpu.ex.r_epc[10] ),
    .A2(_10492_),
    .A1(\cpu.ex.r_stmp[10] ));
 sg13g2_nand2b_1 _17702_ (.Y(_10885_),
    .B(net882),
    .A_N(_10884_));
 sg13g2_and3_1 _17703_ (.X(_10886_),
    .A(net755),
    .B(\cpu.ex.r_9[10] ),
    .C(_10487_));
 sg13g2_buf_2 _17704_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10887_));
 sg13g2_inv_2 _17705_ (.Y(_10888_),
    .A(_10887_));
 sg13g2_nor4_1 _17706_ (.A(net880),
    .B(net758),
    .C(net755),
    .D(_10888_),
    .Y(_10889_));
 sg13g2_o21ai_1 _17707_ (.B1(net669),
    .Y(_10890_),
    .A1(_10886_),
    .A2(_10889_));
 sg13g2_buf_1 _17708_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10891_));
 sg13g2_mux2_1 _17709_ (.A0(\cpu.ex.r_12[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net888),
    .X(_10892_));
 sg13g2_and3_1 _17710_ (.X(_10893_),
    .A(net762),
    .B(net671),
    .C(_10892_));
 sg13g2_a221oi_1 _17711_ (.B2(_10891_),
    .C1(_10893_),
    .B1(_10514_),
    .A1(\cpu.ex.r_lr[10] ),
    .Y(_10894_),
    .A2(_10513_));
 sg13g2_nand2b_1 _17712_ (.Y(_10895_),
    .B(net881),
    .A_N(_00270_));
 sg13g2_nand2b_1 _17713_ (.Y(_10896_),
    .B(\cpu.ex.r_11[10] ),
    .A_N(net884));
 sg13g2_a21o_1 _17714_ (.A2(_10896_),
    .A1(_10895_),
    .B1(_10573_),
    .X(_10897_));
 sg13g2_nand3_1 _17715_ (.B(net879),
    .C(net760),
    .A(\cpu.ex.r_8[10] ),
    .Y(_10898_));
 sg13g2_nand3_1 _17716_ (.B(_10465_),
    .C(net667),
    .A(\cpu.ex.r_13[10] ),
    .Y(_10899_));
 sg13g2_nand3_1 _17717_ (.B(net668),
    .C(net760),
    .A(\cpu.ex.r_10[10] ),
    .Y(_10900_));
 sg13g2_and4_1 _17718_ (.A(_10897_),
    .B(_10898_),
    .C(_10899_),
    .D(_10900_),
    .X(_10901_));
 sg13g2_nand4_1 _17719_ (.B(_10890_),
    .C(_10894_),
    .A(_10885_),
    .Y(_10902_),
    .D(_10901_));
 sg13g2_buf_2 _17720_ (.A(\cpu.addr[10] ),
    .X(_10903_));
 sg13g2_nand2b_1 _17721_ (.Y(_10904_),
    .B(net538),
    .A_N(_10903_));
 sg13g2_o21ai_1 _17722_ (.B1(_10904_),
    .Y(_10905_),
    .A1(net538),
    .A2(_10902_));
 sg13g2_nor2_1 _17723_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_10905_),
    .Y(_10906_));
 sg13g2_buf_1 _17724_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10907_));
 sg13g2_a221oi_1 _17725_ (.B2(\cpu.ex.r_lr[11] ),
    .C1(net670),
    .B1(net667),
    .A1(_10907_),
    .Y(_10908_),
    .A2(net668));
 sg13g2_a221oi_1 _17726_ (.B2(\cpu.ex.r_9[11] ),
    .C1(_10421_),
    .B1(net667),
    .A1(\cpu.ex.r_10[11] ),
    .Y(_10909_),
    .A2(net668));
 sg13g2_or3_1 _17727_ (.A(net756),
    .B(_10908_),
    .C(_10909_),
    .X(_10910_));
 sg13g2_nand3b_1 _17728_ (.B(net881),
    .C(\cpu.ex.r_mult[27] ),
    .Y(_10911_),
    .A_N(net758));
 sg13g2_nand3b_1 _17729_ (.B(\cpu.ex.r_11[11] ),
    .C(net758),
    .Y(_10912_),
    .A_N(net881));
 sg13g2_a21oi_1 _17730_ (.A1(_10911_),
    .A2(_10912_),
    .Y(_10913_),
    .B1(net759));
 sg13g2_and3_1 _17731_ (.X(_10914_),
    .A(net762),
    .B(\cpu.ex.r_14[11] ),
    .C(net671));
 sg13g2_o21ai_1 _17732_ (.B1(net757),
    .Y(_10915_),
    .A1(_10913_),
    .A2(_10914_));
 sg13g2_and3_1 _17733_ (.X(_10916_),
    .A(net670),
    .B(\cpu.ex.r_13[11] ),
    .C(net667));
 sg13g2_inv_1 _17734_ (.Y(_10917_),
    .A(\cpu.ex.r_stmp[11] ));
 sg13g2_nor3_1 _17735_ (.A(net670),
    .B(_10917_),
    .C(_10483_),
    .Y(_10918_));
 sg13g2_o21ai_1 _17736_ (.B1(net756),
    .Y(_10919_),
    .A1(_10916_),
    .A2(_10918_));
 sg13g2_and2_1 _17737_ (.A(net670),
    .B(net879),
    .X(_10920_));
 sg13g2_mux2_1 _17738_ (.A0(\cpu.ex.r_8[11] ),
    .A1(\cpu.ex.r_12[11] ),
    .S(net881),
    .X(_10921_));
 sg13g2_nor2_1 _17739_ (.A(_00271_),
    .B(_10517_),
    .Y(_10922_));
 sg13g2_a221oi_1 _17740_ (.B2(_10921_),
    .C1(_10922_),
    .B1(_10920_),
    .A1(\cpu.ex.r_epc[11] ),
    .Y(_10923_),
    .A2(_10457_));
 sg13g2_nand4_1 _17741_ (.B(_10915_),
    .C(_10919_),
    .A(_10910_),
    .Y(_10924_),
    .D(_10923_));
 sg13g2_buf_2 _17742_ (.A(\cpu.addr[11] ),
    .X(_10925_));
 sg13g2_nand2b_1 _17743_ (.Y(_10926_),
    .B(_10538_),
    .A_N(_10925_));
 sg13g2_o21ai_1 _17744_ (.B1(_10926_),
    .Y(_10927_),
    .A1(_10538_),
    .A2(_10924_));
 sg13g2_nor2_1 _17745_ (.A(_09384_),
    .B(_10927_),
    .Y(_10928_));
 sg13g2_nor4_1 _17746_ (.A(net338),
    .B(net268),
    .C(_10906_),
    .D(_10928_),
    .Y(_10929_));
 sg13g2_nor3_1 _17747_ (.A(_10529_),
    .B(_10883_),
    .C(_10929_),
    .Y(_10930_));
 sg13g2_nor4_2 _17748_ (.A(_10797_),
    .B(_10841_),
    .C(_10880_),
    .Y(_10931_),
    .D(_10930_));
 sg13g2_a21o_1 _17749_ (.A2(_10744_),
    .A1(_10610_),
    .B1(_10931_),
    .X(_10932_));
 sg13g2_buf_1 _17750_ (.A(_10932_),
    .X(_10933_));
 sg13g2_nand2b_1 _17751_ (.Y(_10934_),
    .B(_10364_),
    .A_N(_08492_));
 sg13g2_and4_1 _17752_ (.A(_10281_),
    .B(_10283_),
    .C(_10285_),
    .D(_10287_),
    .X(_10935_));
 sg13g2_a22oi_1 _17753_ (.Y(_10936_),
    .B1(_10355_),
    .B2(_10349_),
    .A2(_10935_),
    .A1(_10393_));
 sg13g2_buf_2 _17754_ (.A(_10936_),
    .X(_10937_));
 sg13g2_nand2_1 _17755_ (.Y(_10938_),
    .A(_10361_),
    .B(net601));
 sg13g2_nand3b_1 _17756_ (.B(net889),
    .C(\cpu.ex.r_8[3] ),
    .Y(_10939_),
    .A_N(net891));
 sg13g2_nand3b_1 _17757_ (.B(net891),
    .C(_10515_),
    .Y(_10940_),
    .A_N(net889));
 sg13g2_a21o_1 _17758_ (.A2(_10940_),
    .A1(_10939_),
    .B1(_10329_),
    .X(_10941_));
 sg13g2_buf_8 _17759_ (.A(_10282_),
    .X(_10942_));
 sg13g2_nor2b_1 _17760_ (.A(net1033),
    .B_N(net1042),
    .Y(_10943_));
 sg13g2_buf_1 _17761_ (.A(_10943_),
    .X(_10944_));
 sg13g2_buf_8 _17762_ (.A(_10284_),
    .X(_10945_));
 sg13g2_mux2_1 _17763_ (.A0(\cpu.ex.r_10[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net1032),
    .X(_10946_));
 sg13g2_nand3_1 _17764_ (.B(_10944_),
    .C(_10946_),
    .A(net769),
    .Y(_10947_));
 sg13g2_mux2_1 _17765_ (.A0(_10503_),
    .A1(\cpu.ex.r_13[3] ),
    .S(net889),
    .X(_10948_));
 sg13g2_nand3_1 _17766_ (.B(net768),
    .C(_10948_),
    .A(net893),
    .Y(_10949_));
 sg13g2_nand3_1 _17767_ (.B(_10947_),
    .C(_10949_),
    .A(_10941_),
    .Y(_10950_));
 sg13g2_nor2b_1 _17768_ (.A(_10282_),
    .B_N(_10303_),
    .Y(_10951_));
 sg13g2_buf_1 _17769_ (.A(_10951_),
    .X(_10952_));
 sg13g2_nor2b_1 _17770_ (.A(net1032),
    .B_N(net1033),
    .Y(_10953_));
 sg13g2_a221oi_1 _17771_ (.B2(\cpu.ex.r_lr[3] ),
    .C1(net769),
    .B1(_10953_),
    .A1(net1155),
    .Y(_10954_),
    .A2(_10952_));
 sg13g2_inv_4 _17772_ (.A(net889),
    .Y(_10955_));
 sg13g2_a221oi_1 _17773_ (.B2(\cpu.ex.r_9[3] ),
    .C1(net754),
    .B1(_10953_),
    .A1(\cpu.ex.r_12[3] ),
    .Y(_10956_),
    .A2(_10952_));
 sg13g2_nor3_1 _17774_ (.A(net766),
    .B(_10954_),
    .C(_10956_),
    .Y(_10957_));
 sg13g2_nor2_1 _17775_ (.A(net1033),
    .B(_10299_),
    .Y(_10958_));
 sg13g2_buf_2 _17776_ (.A(_10958_),
    .X(_10959_));
 sg13g2_nand2_1 _17777_ (.Y(_10960_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(_10959_));
 sg13g2_nor2b_1 _17778_ (.A(_00263_),
    .B_N(net889),
    .Y(_10961_));
 sg13g2_nor2b_1 _17779_ (.A(net769),
    .B_N(\cpu.ex.r_mult[19] ),
    .Y(_10962_));
 sg13g2_o21ai_1 _17780_ (.B1(net893),
    .Y(_10963_),
    .A1(_10961_),
    .A2(_10962_));
 sg13g2_nand2_1 _17781_ (.Y(_10964_),
    .A(_10332_),
    .B(net890));
 sg13g2_a21oi_1 _17782_ (.A1(_10960_),
    .A2(_10963_),
    .Y(_10965_),
    .B1(_10964_));
 sg13g2_buf_8 _17783_ (.A(net890),
    .X(_10966_));
 sg13g2_and2_1 _17784_ (.A(\cpu.ex.r_11[3] ),
    .B(net889),
    .X(_10967_));
 sg13g2_a21oi_1 _17785_ (.A1(\cpu.ex.r_epc[3] ),
    .A2(net754),
    .Y(_10968_),
    .B1(_10967_));
 sg13g2_nor4_1 _17786_ (.A(net765),
    .B(_10333_),
    .C(net753),
    .D(_10968_),
    .Y(_10969_));
 sg13g2_nor4_2 _17787_ (.A(_10950_),
    .B(_10957_),
    .C(_10965_),
    .Y(_10970_),
    .D(_10969_));
 sg13g2_inv_1 _17788_ (.Y(_10971_),
    .A(_10361_));
 sg13g2_nor3_1 _17789_ (.A(_10971_),
    .B(_10279_),
    .C(_10289_),
    .Y(_10972_));
 sg13g2_inv_1 _17790_ (.Y(_10973_),
    .A(\cpu.dec.imm[3] ));
 sg13g2_nor2_1 _17791_ (.A(_10273_),
    .B(_10274_),
    .Y(_10974_));
 sg13g2_o21ai_1 _17792_ (.B1(_10974_),
    .Y(_10975_),
    .A1(_10973_),
    .A2(_10361_));
 sg13g2_a21oi_1 _17793_ (.A1(_09219_),
    .A2(_10972_),
    .Y(_10976_),
    .B1(_10975_));
 sg13g2_o21ai_1 _17794_ (.B1(_10976_),
    .Y(_10977_),
    .A1(_10938_),
    .A2(_10970_));
 sg13g2_buf_1 _17795_ (.A(_10977_),
    .X(_10978_));
 sg13g2_nand2_2 _17796_ (.Y(_10979_),
    .A(_10934_),
    .B(_10978_));
 sg13g2_buf_8 _17797_ (.A(_10979_),
    .X(_10980_));
 sg13g2_nand2_1 _17798_ (.Y(_10981_),
    .A(_08501_),
    .B(_10273_));
 sg13g2_nand3_1 _17799_ (.B(net893),
    .C(net764),
    .A(\cpu.ex.r_9[2] ),
    .Y(_10982_));
 sg13g2_nor2b_2 _17800_ (.A(_10323_),
    .B_N(net1032),
    .Y(_10983_));
 sg13g2_nor2b_1 _17801_ (.A(net1045),
    .B_N(_08364_),
    .Y(_10984_));
 sg13g2_a21oi_1 _17802_ (.A1(_10983_),
    .A2(_10984_),
    .Y(_10985_),
    .B1(net766));
 sg13g2_nand3_1 _17803_ (.B(_10335_),
    .C(net763),
    .A(\cpu.ex.r_12[2] ),
    .Y(_10986_));
 sg13g2_nand3_1 _17804_ (.B(net1045),
    .C(_10349_),
    .A(\cpu.ex.r_lr[2] ),
    .Y(_10987_));
 sg13g2_nand4_1 _17805_ (.B(_10985_),
    .C(_10986_),
    .A(_10982_),
    .Y(_10988_),
    .D(_10987_));
 sg13g2_buf_8 _17806_ (.A(net766),
    .X(_10989_));
 sg13g2_nor2b_2 _17807_ (.A(net1045),
    .B_N(_10299_),
    .Y(_10990_));
 sg13g2_mux2_1 _17808_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net1032),
    .X(_10991_));
 sg13g2_mux2_1 _17809_ (.A0(_10443_),
    .A1(\cpu.ex.r_stmp[2] ),
    .S(net1032),
    .X(_10992_));
 sg13g2_a22oi_1 _17810_ (.Y(_10993_),
    .B1(_10992_),
    .B2(_10959_),
    .A2(_10991_),
    .A1(_10990_));
 sg13g2_nand2_1 _17811_ (.Y(_10994_),
    .A(net665),
    .B(_10993_));
 sg13g2_and2_1 _17812_ (.A(\cpu.ex.r_11[2] ),
    .B(_10305_),
    .X(_10995_));
 sg13g2_a21o_1 _17813_ (.A2(net768),
    .A1(\cpu.ex.r_13[2] ),
    .B1(_10995_),
    .X(_10996_));
 sg13g2_and2_1 _17814_ (.A(net1045),
    .B(net769),
    .X(_10997_));
 sg13g2_buf_2 _17815_ (.A(_10997_),
    .X(_10998_));
 sg13g2_nor2b_1 _17816_ (.A(_00262_),
    .B_N(net889),
    .Y(_10999_));
 sg13g2_nor2b_1 _17817_ (.A(net769),
    .B_N(\cpu.ex.r_mult[18] ),
    .Y(_11000_));
 sg13g2_and3_1 _17818_ (.X(_11001_),
    .A(net1045),
    .B(net891),
    .C(net890));
 sg13g2_o21ai_1 _17819_ (.B1(_11001_),
    .Y(_11002_),
    .A1(_10999_),
    .A2(_11000_));
 sg13g2_nand3b_1 _17820_ (.B(net891),
    .C(\cpu.ex.r_epc[2] ),
    .Y(_11003_),
    .A_N(net890));
 sg13g2_nand3b_1 _17821_ (.B(net890),
    .C(_10419_),
    .Y(_11004_),
    .A_N(net891));
 sg13g2_nand2b_1 _17822_ (.Y(_11005_),
    .B(net1045),
    .A_N(net889));
 sg13g2_a21o_1 _17823_ (.A2(_11004_),
    .A1(_11003_),
    .B1(_11005_),
    .X(_11006_));
 sg13g2_nand3_1 _17824_ (.B(_10355_),
    .C(net764),
    .A(\cpu.ex.r_8[2] ),
    .Y(_11007_));
 sg13g2_nand3_1 _17825_ (.B(_11006_),
    .C(_11007_),
    .A(_11002_),
    .Y(_11008_));
 sg13g2_a221oi_1 _17826_ (.B2(_10998_),
    .C1(_11008_),
    .B1(_10996_),
    .A1(_10988_),
    .Y(_11009_),
    .A2(_10994_));
 sg13g2_buf_1 _17827_ (.A(\cpu.dec.imm[2] ),
    .X(_11010_));
 sg13g2_a221oi_1 _17828_ (.B2(_09234_),
    .C1(_10276_),
    .B1(_10972_),
    .A1(_11010_),
    .Y(_11011_),
    .A2(_10971_));
 sg13g2_o21ai_1 _17829_ (.B1(_11011_),
    .Y(_11012_),
    .A1(_10938_),
    .A2(_11009_));
 sg13g2_buf_1 _17830_ (.A(_11012_),
    .X(_11013_));
 sg13g2_nand2_1 _17831_ (.Y(_11014_),
    .A(_10981_),
    .B(_11013_));
 sg13g2_buf_1 _17832_ (.A(_11014_),
    .X(_11015_));
 sg13g2_and2_1 _17833_ (.A(_10942_),
    .B(_10310_),
    .X(_11016_));
 sg13g2_buf_1 _17834_ (.A(_11016_),
    .X(_11017_));
 sg13g2_inv_1 _17835_ (.Y(_11018_),
    .A(\cpu.ex.r_epc[1] ));
 sg13g2_or2_1 _17836_ (.X(_11019_),
    .B(net1043),
    .A(net1044));
 sg13g2_nand3b_1 _17837_ (.B(net892),
    .C(_10945_),
    .Y(_11020_),
    .A_N(_00261_));
 sg13g2_o21ai_1 _17838_ (.B1(_11020_),
    .Y(_11021_),
    .A1(_11018_),
    .A2(_11019_));
 sg13g2_inv_1 _17839_ (.Y(_11022_),
    .A(\cpu.ex.r_prev_ie ));
 sg13g2_or2_1 _17840_ (.X(_11023_),
    .B(net1044),
    .A(net1033));
 sg13g2_nand3_1 _17841_ (.B(net1033),
    .C(net892),
    .A(\cpu.ex.r_13[1] ),
    .Y(_11024_));
 sg13g2_o21ai_1 _17842_ (.B1(_11024_),
    .Y(_11025_),
    .A1(_11022_),
    .A2(_11023_));
 sg13g2_a22oi_1 _17843_ (.Y(_11026_),
    .B1(_11025_),
    .B2(net768),
    .A2(_11021_),
    .A1(_11017_));
 sg13g2_nand3b_1 _17844_ (.B(net1032),
    .C(\cpu.ex.r_14[1] ),
    .Y(_11027_),
    .A_N(net1033));
 sg13g2_nand3b_1 _17845_ (.B(_10942_),
    .C(\cpu.ex.r_11[1] ),
    .Y(_11028_),
    .A_N(net1043));
 sg13g2_nand2_1 _17846_ (.Y(_11029_),
    .A(net1042),
    .B(net892));
 sg13g2_a21oi_1 _17847_ (.A1(_11027_),
    .A2(_11028_),
    .Y(_11030_),
    .B1(_11029_));
 sg13g2_nand3b_1 _17848_ (.B(net892),
    .C(\cpu.ex.r_8[1] ),
    .Y(_11031_),
    .A_N(net1042));
 sg13g2_nand3b_1 _17849_ (.B(net1042),
    .C(_10698_),
    .Y(_11032_),
    .A_N(net1044));
 sg13g2_a21oi_1 _17850_ (.A1(_11031_),
    .A2(_11032_),
    .Y(_11033_),
    .B1(_10329_));
 sg13g2_nand3b_1 _17851_ (.B(net1042),
    .C(\cpu.ex.r_10[1] ),
    .Y(_11034_),
    .A_N(net1043));
 sg13g2_nand3b_1 _17852_ (.B(net1032),
    .C(\cpu.ex.r_12[1] ),
    .Y(_11035_),
    .A_N(net1042));
 sg13g2_nand2b_1 _17853_ (.Y(_11036_),
    .B(net892),
    .A_N(net1033));
 sg13g2_a21oi_1 _17854_ (.A1(_11034_),
    .A2(_11035_),
    .Y(_11037_),
    .B1(_11036_));
 sg13g2_nor3_1 _17855_ (.A(_11030_),
    .B(_11033_),
    .C(_11037_),
    .Y(_11038_));
 sg13g2_mux2_1 _17856_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_9[1] ),
    .S(net892),
    .X(_11039_));
 sg13g2_nand2b_1 _17857_ (.Y(_11040_),
    .B(_10282_),
    .A_N(_10286_));
 sg13g2_buf_1 _17858_ (.A(_11040_),
    .X(_11041_));
 sg13g2_nor2_1 _17859_ (.A(_10945_),
    .B(_11041_),
    .Y(_11042_));
 sg13g2_mux2_1 _17860_ (.A0(\cpu.ex.r_stmp[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(net1033),
    .X(_11043_));
 sg13g2_inv_1 _17861_ (.Y(_11044_),
    .A(net1043));
 sg13g2_nand2b_1 _17862_ (.Y(_11045_),
    .B(_10310_),
    .A_N(net1044));
 sg13g2_nor2_1 _17863_ (.A(_11044_),
    .B(_11045_),
    .Y(_11046_));
 sg13g2_nor2b_1 _17864_ (.A(_10298_),
    .B_N(_10282_),
    .Y(_11047_));
 sg13g2_and3_1 _17865_ (.X(_11048_),
    .A(\cpu.ex.mmu_read[1] ),
    .B(_10306_),
    .C(_11047_));
 sg13g2_a221oi_1 _17866_ (.B2(_11046_),
    .C1(_11048_),
    .B1(_11043_),
    .A1(_11039_),
    .Y(_11049_),
    .A2(_11042_));
 sg13g2_and3_1 _17867_ (.X(_11050_),
    .A(_11026_),
    .B(_11038_),
    .C(_11049_));
 sg13g2_buf_2 _17868_ (.A(\cpu.dec.imm[1] ),
    .X(_11051_));
 sg13g2_nor2_1 _17869_ (.A(_10089_),
    .B(_10971_),
    .Y(_11052_));
 sg13g2_a221oi_1 _17870_ (.B2(_11052_),
    .C1(_10276_),
    .B1(net608),
    .A1(_11051_),
    .Y(_11053_),
    .A2(_10971_));
 sg13g2_o21ai_1 _17871_ (.B1(_11053_),
    .Y(_11054_),
    .A1(_10938_),
    .A2(_11050_));
 sg13g2_buf_2 _17872_ (.A(_11054_),
    .X(_11055_));
 sg13g2_nand2_1 _17873_ (.Y(_11056_),
    .A(net1077),
    .B(_10273_));
 sg13g2_buf_2 _17874_ (.A(_11056_),
    .X(_11057_));
 sg13g2_buf_1 _17875_ (.A(_00311_),
    .X(_11058_));
 sg13g2_a21oi_1 _17876_ (.A1(_11055_),
    .A2(_11057_),
    .Y(_11059_),
    .B1(_11058_));
 sg13g2_and2_1 _17877_ (.A(net266),
    .B(_11059_),
    .X(_11060_));
 sg13g2_buf_2 _17878_ (.A(_00309_),
    .X(_11061_));
 sg13g2_inv_2 _17879_ (.Y(_11062_),
    .A(_11061_));
 sg13g2_o21ai_1 _17880_ (.B1(_11062_),
    .Y(_11063_),
    .A1(net267),
    .A2(_11060_));
 sg13g2_buf_1 _17881_ (.A(net267),
    .X(_11064_));
 sg13g2_nand2_1 _17882_ (.Y(_11065_),
    .A(net227),
    .B(_11060_));
 sg13g2_a21oi_1 _17883_ (.A1(_11063_),
    .A2(_11065_),
    .Y(_11066_),
    .B1(net690));
 sg13g2_nand3_1 _17884_ (.B(net676),
    .C(net767),
    .A(net665),
    .Y(_11067_));
 sg13g2_buf_1 _17885_ (.A(net1045),
    .X(_11068_));
 sg13g2_and2_1 _17886_ (.A(\cpu.ex.r_15[0] ),
    .B(net878),
    .X(_11069_));
 sg13g2_a21oi_1 _17887_ (.A1(\cpu.ex.r_14[0] ),
    .A2(net765),
    .Y(_11070_),
    .B1(_11069_));
 sg13g2_mux2_1 _17888_ (.A0(\cpu.ex.r_8[0] ),
    .A1(\cpu.ex.r_12[0] ),
    .S(net753),
    .X(_11071_));
 sg13g2_nand3_1 _17889_ (.B(net675),
    .C(_11071_),
    .A(net765),
    .Y(_11072_));
 sg13g2_o21ai_1 _17890_ (.B1(_11072_),
    .Y(_11073_),
    .A1(_11067_),
    .A2(_11070_));
 sg13g2_nand3b_1 _17891_ (.B(net676),
    .C(_11068_),
    .Y(_11074_),
    .A_N(net767));
 sg13g2_and2_1 _17892_ (.A(\cpu.ex.r_11[0] ),
    .B(net766),
    .X(_11075_));
 sg13g2_a21oi_1 _17893_ (.A1(\cpu.ex.r_9[0] ),
    .A2(_10333_),
    .Y(_11076_),
    .B1(_11075_));
 sg13g2_mux2_1 _17894_ (.A0(_10649_),
    .A1(\cpu.ex.r_mult[16] ),
    .S(net753),
    .X(_11077_));
 sg13g2_nand3_1 _17895_ (.B(_10325_),
    .C(_11077_),
    .A(net770),
    .Y(_11078_));
 sg13g2_o21ai_1 _17896_ (.B1(_11078_),
    .Y(_11079_),
    .A1(_11074_),
    .A2(_11076_));
 sg13g2_a22oi_1 _17897_ (.Y(_11080_),
    .B1(_10959_),
    .B2(_09242_),
    .A2(_10998_),
    .A1(\cpu.ex.r_13[0] ));
 sg13g2_nor2b_1 _17898_ (.A(_11080_),
    .B_N(net768),
    .Y(_11081_));
 sg13g2_a22oi_1 _17899_ (.Y(_11082_),
    .B1(net764),
    .B2(\cpu.ex.r_10[0] ),
    .A2(_10983_),
    .A1(\cpu.ex.r_stmp[0] ));
 sg13g2_nor2b_1 _17900_ (.A(_11082_),
    .B_N(_10944_),
    .Y(_11083_));
 sg13g2_nor4_1 _17901_ (.A(_11073_),
    .B(_11079_),
    .C(_11081_),
    .D(_11083_),
    .Y(_11084_));
 sg13g2_nand2_1 _17902_ (.Y(_11085_),
    .A(net1151),
    .B(net608));
 sg13g2_o21ai_1 _17903_ (.B1(_11085_),
    .Y(_11086_),
    .A1(net540),
    .A2(_11084_));
 sg13g2_nand2b_1 _17904_ (.Y(_11087_),
    .B(_10362_),
    .A_N(_10274_));
 sg13g2_buf_1 _17905_ (.A(\cpu.dec.imm[0] ),
    .X(_11088_));
 sg13g2_nor3_1 _17906_ (.A(_11088_),
    .B(net1041),
    .C(_10274_),
    .Y(_11089_));
 sg13g2_nor2_1 _17907_ (.A(net1040),
    .B(_11089_),
    .Y(_11090_));
 sg13g2_o21ai_1 _17908_ (.B1(_11090_),
    .Y(_11091_),
    .A1(_11086_),
    .A2(_11087_));
 sg13g2_buf_2 _17909_ (.A(_11091_),
    .X(_11092_));
 sg13g2_buf_1 _17910_ (.A(_11092_),
    .X(_11093_));
 sg13g2_nor2_1 _17911_ (.A(_11066_),
    .B(net226),
    .Y(_11094_));
 sg13g2_buf_1 _17912_ (.A(_10971_),
    .X(_11095_));
 sg13g2_nor2_1 _17913_ (.A(net877),
    .B(_10276_),
    .Y(_11096_));
 sg13g2_buf_1 _17914_ (.A(_11096_),
    .X(_11097_));
 sg13g2_a22oi_1 _17915_ (.Y(_11098_),
    .B1(_10313_),
    .B2(\cpu.ex.r_9[5] ),
    .A2(_10325_),
    .A1(\cpu.ex.r_epc[5] ));
 sg13g2_nor2_1 _17916_ (.A(net767),
    .B(_11098_),
    .Y(_11099_));
 sg13g2_buf_8 _17917_ (.A(net665),
    .X(_11100_));
 sg13g2_a22oi_1 _17918_ (.Y(_11101_),
    .B1(net763),
    .B2(\cpu.ex.r_13[5] ),
    .A2(net672),
    .A1(\cpu.ex.r_lr[5] ));
 sg13g2_nor2_1 _17919_ (.A(net600),
    .B(_11101_),
    .Y(_11102_));
 sg13g2_o21ai_1 _17920_ (.B1(net677),
    .Y(_11103_),
    .A1(_11099_),
    .A2(_11102_));
 sg13g2_a22oi_1 _17921_ (.Y(_11104_),
    .B1(_10313_),
    .B2(\cpu.ex.r_12[5] ),
    .A2(_10326_),
    .A1(\cpu.ex.r_stmp[5] ));
 sg13g2_nand2b_1 _17922_ (.Y(_11105_),
    .B(_10952_),
    .A_N(_11104_));
 sg13g2_a22oi_1 _17923_ (.Y(_11106_),
    .B1(_10959_),
    .B2(_10547_),
    .A2(_10998_),
    .A1(\cpu.ex.r_11[5] ));
 sg13g2_nand2b_1 _17924_ (.Y(_11107_),
    .B(_10305_),
    .A_N(_11106_));
 sg13g2_and2_1 _17925_ (.A(_10355_),
    .B(_10339_),
    .X(_11108_));
 sg13g2_nand2_1 _17926_ (.Y(_11109_),
    .A(net893),
    .B(net890));
 sg13g2_nor2_1 _17927_ (.A(net893),
    .B(_10315_),
    .Y(_11110_));
 sg13g2_nand2_1 _17928_ (.Y(_11111_),
    .A(\cpu.ex.r_10[5] ),
    .B(_11110_));
 sg13g2_o21ai_1 _17929_ (.B1(_11111_),
    .Y(_11112_),
    .A1(_00265_),
    .A2(_11109_));
 sg13g2_and2_1 _17930_ (.A(_10332_),
    .B(net769),
    .X(_11113_));
 sg13g2_a22oi_1 _17931_ (.Y(_11114_),
    .B1(_10990_),
    .B2(\cpu.ex.r_14[5] ),
    .A2(_11047_),
    .A1(\cpu.ex.r_mult[21] ));
 sg13g2_nor2_1 _17932_ (.A(_10964_),
    .B(_11114_),
    .Y(_11115_));
 sg13g2_a221oi_1 _17933_ (.B2(_11113_),
    .C1(_11115_),
    .B1(_11112_),
    .A1(\cpu.ex.r_8[5] ),
    .Y(_11116_),
    .A2(_11108_));
 sg13g2_nand4_1 _17934_ (.B(_11105_),
    .C(_11107_),
    .A(_11103_),
    .Y(_11117_),
    .D(_11116_));
 sg13g2_a22oi_1 _17935_ (.Y(_11118_),
    .B1(net601),
    .B2(_11117_),
    .A2(net608),
    .A1(_10027_));
 sg13g2_buf_2 _17936_ (.A(_11118_),
    .X(_11119_));
 sg13g2_inv_1 _17937_ (.Y(_11120_),
    .A(_10273_));
 sg13g2_inv_1 _17938_ (.Y(_11121_),
    .A(\cpu.dec.imm[5] ));
 sg13g2_buf_1 _17939_ (.A(_10974_),
    .X(_11122_));
 sg13g2_nand3_1 _17940_ (.B(_11121_),
    .C(net876),
    .A(net877),
    .Y(_11123_));
 sg13g2_o21ai_1 _17941_ (.B1(_11123_),
    .Y(_11124_),
    .A1(_08815_),
    .A2(net1031));
 sg13g2_a21oi_1 _17942_ (.A1(_11097_),
    .A2(_11119_),
    .Y(_11125_),
    .B1(_11124_));
 sg13g2_buf_1 _17943_ (.A(_11125_),
    .X(_11126_));
 sg13g2_a22oi_1 _17944_ (.Y(_11127_),
    .B1(net764),
    .B2(\cpu.ex.r_10[4] ),
    .A2(_10983_),
    .A1(\cpu.ex.r_stmp[4] ));
 sg13g2_nand2b_1 _17945_ (.Y(_11128_),
    .B(_11100_),
    .A_N(_11127_));
 sg13g2_nor2_1 _17946_ (.A(net891),
    .B(net890),
    .Y(_11129_));
 sg13g2_buf_2 _17947_ (.A(_11129_),
    .X(_11130_));
 sg13g2_and2_1 _17948_ (.A(_10311_),
    .B(net1032),
    .X(_11131_));
 sg13g2_buf_2 _17949_ (.A(_11131_),
    .X(_11132_));
 sg13g2_a22oi_1 _17950_ (.Y(_11133_),
    .B1(_11132_),
    .B2(\cpu.ex.r_14[4] ),
    .A2(_11130_),
    .A1(\cpu.ex.r_8[4] ));
 sg13g2_nand2b_1 _17951_ (.Y(_11134_),
    .B(_10301_),
    .A_N(_11133_));
 sg13g2_a21oi_1 _17952_ (.A1(_11128_),
    .A2(_11134_),
    .Y(_11135_),
    .B1(_10296_));
 sg13g2_nand3b_1 _17953_ (.B(_11068_),
    .C(_10346_),
    .Y(_11136_),
    .A_N(_00264_));
 sg13g2_nand3_1 _17954_ (.B(_10336_),
    .C(net672),
    .A(_10582_),
    .Y(_11137_));
 sg13g2_a21oi_1 _17955_ (.A1(_11136_),
    .A2(_11137_),
    .Y(_11138_),
    .B1(net602));
 sg13g2_a22oi_1 _17956_ (.Y(_11139_),
    .B1(_10953_),
    .B2(\cpu.ex.r_9[4] ),
    .A2(_10952_),
    .A1(\cpu.ex.r_12[4] ));
 sg13g2_nor2b_1 _17957_ (.A(_11139_),
    .B_N(net675),
    .Y(_11140_));
 sg13g2_a22oi_1 _17958_ (.Y(_11141_),
    .B1(_10959_),
    .B2(_08311_),
    .A2(_10998_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_nor2b_1 _17959_ (.A(_11141_),
    .B_N(net768),
    .Y(_11142_));
 sg13g2_a22oi_1 _17960_ (.Y(_11143_),
    .B1(_11132_),
    .B2(\cpu.ex.r_mult[20] ),
    .A2(_11130_),
    .A1(\cpu.ex.r_lr[4] ));
 sg13g2_buf_1 _17961_ (.A(_11044_),
    .X(_11144_));
 sg13g2_mux2_1 _17962_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(\cpu.ex.r_11[4] ),
    .S(net676),
    .X(_11145_));
 sg13g2_nand3_1 _17963_ (.B(_11017_),
    .C(_11145_),
    .A(net752),
    .Y(_11146_));
 sg13g2_o21ai_1 _17964_ (.B1(_11146_),
    .Y(_11147_),
    .A1(_11005_),
    .A2(_11143_));
 sg13g2_or4_1 _17965_ (.A(_11138_),
    .B(_11140_),
    .C(_11142_),
    .D(_11147_),
    .X(_11148_));
 sg13g2_nor2_1 _17966_ (.A(net877),
    .B(net540),
    .Y(_11149_));
 sg13g2_o21ai_1 _17967_ (.B1(_11149_),
    .Y(_11150_),
    .A1(_11135_),
    .A2(_11148_));
 sg13g2_nor2_1 _17968_ (.A(_09742_),
    .B(_11095_),
    .Y(_11151_));
 sg13g2_a221oi_1 _17969_ (.B2(_11151_),
    .C1(_10276_),
    .B1(net608),
    .A1(_11095_),
    .Y(_11152_),
    .A2(\cpu.dec.imm[4] ));
 sg13g2_nor2_1 _17970_ (.A(net1150),
    .B(net1031),
    .Y(_11153_));
 sg13g2_a21oi_1 _17971_ (.A1(_11150_),
    .A2(_11152_),
    .Y(_11154_),
    .B1(_11153_));
 sg13g2_buf_1 _17972_ (.A(_11154_),
    .X(_11155_));
 sg13g2_o21ai_1 _17973_ (.B1(net690),
    .Y(_11156_),
    .A1(net225),
    .A2(net265));
 sg13g2_buf_1 _17974_ (.A(_00307_),
    .X(_11157_));
 sg13g2_buf_1 _17975_ (.A(_00308_),
    .X(_11158_));
 sg13g2_inv_2 _17976_ (.Y(_11159_),
    .A(_11158_));
 sg13g2_a21o_1 _17977_ (.A2(_11152_),
    .A1(_11150_),
    .B1(_11153_),
    .X(_11160_));
 sg13g2_buf_1 _17978_ (.A(_11160_),
    .X(_11161_));
 sg13g2_nor2_1 _17979_ (.A(_11159_),
    .B(net264),
    .Y(_11162_));
 sg13g2_a21oi_1 _17980_ (.A1(_11157_),
    .A2(net225),
    .Y(_11163_),
    .B1(_11162_));
 sg13g2_inv_1 _17981_ (.Y(_11164_),
    .A(_10620_));
 sg13g2_nand2_1 _17982_ (.Y(_11165_),
    .A(net1041),
    .B(net876));
 sg13g2_a221oi_1 _17983_ (.B2(\cpu.ex.r_12[7] ),
    .C1(net878),
    .B1(net768),
    .A1(\cpu.ex.r_10[7] ),
    .Y(_11166_),
    .A2(_10305_));
 sg13g2_a221oi_1 _17984_ (.B2(\cpu.ex.r_13[7] ),
    .C1(net765),
    .B1(_10307_),
    .A1(\cpu.ex.r_11[7] ),
    .Y(_11167_),
    .A2(_10305_));
 sg13g2_nor2b_1 _17985_ (.A(net893),
    .B_N(\cpu.ex.r_14[7] ),
    .Y(_11168_));
 sg13g2_and2_1 _17986_ (.A(\cpu.ex.r_9[7] ),
    .B(net893),
    .X(_11169_));
 sg13g2_a22oi_1 _17987_ (.Y(_11170_),
    .B1(_11169_),
    .B2(_11130_),
    .A2(_11168_),
    .A1(_11132_));
 sg13g2_o21ai_1 _17988_ (.B1(_11170_),
    .Y(_11171_),
    .A1(_11166_),
    .A2(_11167_));
 sg13g2_nand3_1 _17989_ (.B(net754),
    .C(_10355_),
    .A(_10721_),
    .Y(_11172_));
 sg13g2_nand3b_1 _17990_ (.B(net770),
    .C(_11113_),
    .Y(_11173_),
    .A_N(_00267_));
 sg13g2_nand3_1 _17991_ (.B(_11172_),
    .C(_11173_),
    .A(net674),
    .Y(_11174_));
 sg13g2_a22oi_1 _17992_ (.Y(_11175_),
    .B1(net675),
    .B2(\cpu.ex.r_8[7] ),
    .A2(_10325_),
    .A1(_10725_));
 sg13g2_o21ai_1 _17993_ (.B1(net752),
    .Y(_11176_),
    .A1(net770),
    .A2(_11175_));
 sg13g2_a22oi_1 _17994_ (.Y(_11177_),
    .B1(_11132_),
    .B2(\cpu.ex.r_mult[23] ),
    .A2(_11130_),
    .A1(\cpu.ex.r_lr[7] ));
 sg13g2_nand3b_1 _17995_ (.B(net753),
    .C(\cpu.ex.r_stmp[7] ),
    .Y(_11178_),
    .A_N(_10294_));
 sg13g2_nand3b_1 _17996_ (.B(net878),
    .C(\cpu.ex.r_epc[7] ),
    .Y(_11179_),
    .A_N(_10966_));
 sg13g2_a21o_1 _17997_ (.A2(_11179_),
    .A1(_11178_),
    .B1(_11045_),
    .X(_11180_));
 sg13g2_o21ai_1 _17998_ (.B1(_11180_),
    .Y(_11181_),
    .A1(_11005_),
    .A2(_11177_));
 sg13g2_a221oi_1 _17999_ (.B2(_11176_),
    .C1(_11181_),
    .B1(_11174_),
    .A1(_10302_),
    .Y(_11182_),
    .A2(_11171_));
 sg13g2_nand2_1 _18000_ (.Y(_11183_),
    .A(_09228_),
    .B(net608));
 sg13g2_o21ai_1 _18001_ (.B1(_11183_),
    .Y(_11184_),
    .A1(net540),
    .A2(_11182_));
 sg13g2_nor2_1 _18002_ (.A(_10361_),
    .B(\cpu.dec.imm[7] ),
    .Y(_11185_));
 sg13g2_a22oi_1 _18003_ (.Y(_11186_),
    .B1(net876),
    .B2(_11185_),
    .A2(net1040),
    .A1(_08872_));
 sg13g2_o21ai_1 _18004_ (.B1(_11186_),
    .Y(_11187_),
    .A1(_11165_),
    .A2(_11184_));
 sg13g2_buf_2 _18005_ (.A(_11187_),
    .X(_11188_));
 sg13g2_inv_1 _18006_ (.Y(_11189_),
    .A(_11188_));
 sg13g2_buf_1 _18007_ (.A(_11189_),
    .X(_11190_));
 sg13g2_nand3_1 _18008_ (.B(_10966_),
    .C(_10325_),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_11191_));
 sg13g2_nand3_1 _18009_ (.B(_11044_),
    .C(_10312_),
    .A(\cpu.ex.r_8[6] ),
    .Y(_11192_));
 sg13g2_a21o_1 _18010_ (.A2(_11192_),
    .A1(_11191_),
    .B1(net770),
    .X(_11193_));
 sg13g2_and3_1 _18011_ (.X(_11194_),
    .A(\cpu.ex.r_epc[6] ),
    .B(net878),
    .C(_10349_));
 sg13g2_and3_1 _18012_ (.X(_11195_),
    .A(\cpu.ex.r_14[6] ),
    .B(_10335_),
    .C(net763));
 sg13g2_o21ai_1 _18013_ (.B1(_10989_),
    .Y(_11196_),
    .A1(_11194_),
    .A2(_11195_));
 sg13g2_nor2_1 _18014_ (.A(_11019_),
    .B(_11041_),
    .Y(_11197_));
 sg13g2_inv_1 _18015_ (.Y(_11198_),
    .A(\cpu.ex.r_sp[6] ));
 sg13g2_nand3_1 _18016_ (.B(net893),
    .C(_10300_),
    .A(\cpu.ex.r_11[6] ),
    .Y(_11199_));
 sg13g2_o21ai_1 _18017_ (.B1(_11199_),
    .Y(_11200_),
    .A1(_11198_),
    .A2(_11023_));
 sg13g2_nand3b_1 _18018_ (.B(_10300_),
    .C(\cpu.ex.r_13[6] ),
    .Y(_11201_),
    .A_N(net766));
 sg13g2_nand3b_1 _18019_ (.B(net766),
    .C(_10620_),
    .Y(_11202_),
    .A_N(net769));
 sg13g2_a21oi_1 _18020_ (.A1(_11201_),
    .A2(_11202_),
    .Y(_11203_),
    .B1(_11109_));
 sg13g2_a221oi_1 _18021_ (.B2(_10305_),
    .C1(_11203_),
    .B1(_11200_),
    .A1(\cpu.ex.r_lr[6] ),
    .Y(_11204_),
    .A2(_11197_));
 sg13g2_nor2b_1 _18022_ (.A(net891),
    .B_N(_10293_),
    .Y(_11205_));
 sg13g2_a221oi_1 _18023_ (.B2(\cpu.ex.r_10[6] ),
    .C1(net753),
    .B1(_10944_),
    .A1(\cpu.ex.r_9[6] ),
    .Y(_11206_),
    .A2(_11205_));
 sg13g2_a221oi_1 _18024_ (.B2(_10627_),
    .C1(_11044_),
    .B1(_11017_),
    .A1(\cpu.ex.r_12[6] ),
    .Y(_11207_),
    .A2(_10355_));
 sg13g2_or3_1 _18025_ (.A(net754),
    .B(_11206_),
    .C(_11207_),
    .X(_11208_));
 sg13g2_and4_1 _18026_ (.A(_11193_),
    .B(_11196_),
    .C(_11204_),
    .D(_11208_),
    .X(_11209_));
 sg13g2_nand2_1 _18027_ (.Y(_11210_),
    .A(_09224_),
    .B(net608));
 sg13g2_o21ai_1 _18028_ (.B1(_11210_),
    .Y(_11211_),
    .A1(_10358_),
    .A2(_11209_));
 sg13g2_inv_1 _18029_ (.Y(_11212_),
    .A(_11211_));
 sg13g2_inv_1 _18030_ (.Y(_11213_),
    .A(\cpu.dec.imm[6] ));
 sg13g2_nand3_1 _18031_ (.B(_11213_),
    .C(net876),
    .A(_10971_),
    .Y(_11214_));
 sg13g2_o21ai_1 _18032_ (.B1(_11214_),
    .Y(_11215_),
    .A1(_08863_),
    .A2(net1031));
 sg13g2_a21oi_1 _18033_ (.A1(_11097_),
    .A2(_11212_),
    .Y(_11216_),
    .B1(_11215_));
 sg13g2_buf_8 _18034_ (.A(_11216_),
    .X(_11217_));
 sg13g2_buf_1 _18035_ (.A(_00306_),
    .X(_11218_));
 sg13g2_buf_1 _18036_ (.A(_11188_),
    .X(_11219_));
 sg13g2_inv_1 _18037_ (.Y(_11220_),
    .A(_11215_));
 sg13g2_o21ai_1 _18038_ (.B1(_11220_),
    .Y(_11221_),
    .A1(_11165_),
    .A2(_11211_));
 sg13g2_buf_1 _18039_ (.A(_11221_),
    .X(_11222_));
 sg13g2_nor2_1 _18040_ (.A(_09303_),
    .B(_09376_),
    .Y(_11223_));
 sg13g2_nand2_1 _18041_ (.Y(_11224_),
    .A(\cpu.dec.div ),
    .B(_11223_));
 sg13g2_buf_1 _18042_ (.A(_11224_),
    .X(_11225_));
 sg13g2_a21oi_1 _18043_ (.A1(net263),
    .A2(net337),
    .Y(_11226_),
    .B1(_11225_));
 sg13g2_a221oi_1 _18044_ (.B2(net1127),
    .C1(_11226_),
    .B1(_11217_),
    .A1(_11164_),
    .Y(_11227_),
    .A2(net224));
 sg13g2_and3_1 _18045_ (.X(_11228_),
    .A(_11156_),
    .B(_11163_),
    .C(_11227_));
 sg13g2_buf_1 _18046_ (.A(_11015_),
    .X(_11229_));
 sg13g2_nand3_1 _18047_ (.B(_11055_),
    .C(_11057_),
    .A(_11058_),
    .Y(_11230_));
 sg13g2_a21oi_1 _18048_ (.A1(_10934_),
    .A2(_10978_),
    .Y(_11231_),
    .B1(_11058_));
 sg13g2_a21o_1 _18049_ (.A2(_11230_),
    .A1(_11062_),
    .B1(_11231_),
    .X(_11232_));
 sg13g2_a22oi_1 _18050_ (.Y(_11233_),
    .B1(net223),
    .B2(_11232_),
    .A2(net227),
    .A1(_11062_));
 sg13g2_buf_8 _18051_ (.A(_00310_),
    .X(_11234_));
 sg13g2_inv_1 _18052_ (.Y(_11235_),
    .A(_11234_));
 sg13g2_nand2_1 _18053_ (.Y(_11236_),
    .A(_11235_),
    .B(_11225_));
 sg13g2_nor2_1 _18054_ (.A(_08529_),
    .B(net1031),
    .Y(_11237_));
 sg13g2_or4_1 _18055_ (.A(_10950_),
    .B(_10957_),
    .C(_10965_),
    .D(_10969_),
    .X(_11238_));
 sg13g2_a221oi_1 _18056_ (.B2(_09220_),
    .C1(_10975_),
    .B1(_10972_),
    .A1(_11149_),
    .Y(_11239_),
    .A2(_11238_));
 sg13g2_buf_1 _18057_ (.A(_11239_),
    .X(_11240_));
 sg13g2_nor2_1 _18058_ (.A(_11237_),
    .B(_11240_),
    .Y(_11241_));
 sg13g2_buf_1 _18059_ (.A(_11241_),
    .X(_11242_));
 sg13g2_o21ai_1 _18060_ (.B1(_11242_),
    .Y(_11243_),
    .A1(_11061_),
    .A2(_11236_));
 sg13g2_or2_1 _18061_ (.X(_11244_),
    .B(_11230_),
    .A(net266));
 sg13g2_and2_1 _18062_ (.A(_10981_),
    .B(_11013_),
    .X(_11245_));
 sg13g2_buf_1 _18063_ (.A(_11245_),
    .X(_11246_));
 sg13g2_and2_1 _18064_ (.A(_11055_),
    .B(_11057_),
    .X(_11247_));
 sg13g2_buf_1 _18065_ (.A(_11247_),
    .X(_11248_));
 sg13g2_buf_1 _18066_ (.A(_11248_),
    .X(_11249_));
 sg13g2_o21ai_1 _18067_ (.B1(_11236_),
    .Y(_11250_),
    .A1(net261),
    .A2(net260));
 sg13g2_nand3_1 _18068_ (.B(_11244_),
    .C(_11250_),
    .A(_11243_),
    .Y(_11251_));
 sg13g2_o21ai_1 _18069_ (.B1(_11251_),
    .Y(_11252_),
    .A1(net690),
    .A2(_11233_));
 sg13g2_nand2_1 _18070_ (.Y(_11253_),
    .A(_11228_),
    .B(_11252_));
 sg13g2_a21o_1 _18071_ (.A2(_11094_),
    .A1(_10933_),
    .B1(_11253_),
    .X(_11254_));
 sg13g2_buf_1 _18072_ (.A(_11217_),
    .X(_11255_));
 sg13g2_nor2_1 _18073_ (.A(net224),
    .B(net222),
    .Y(_11256_));
 sg13g2_buf_1 _18074_ (.A(_11225_),
    .X(_11257_));
 sg13g2_nand2_2 _18075_ (.Y(_11258_),
    .A(_10620_),
    .B(net599));
 sg13g2_nor2_1 _18076_ (.A(net222),
    .B(_11258_),
    .Y(_11259_));
 sg13g2_a21o_1 _18077_ (.A2(_11119_),
    .A1(_11097_),
    .B1(_11124_),
    .X(_11260_));
 sg13g2_buf_1 _18078_ (.A(_11260_),
    .X(_11261_));
 sg13g2_nor2_1 _18079_ (.A(_11158_),
    .B(net265),
    .Y(_11262_));
 sg13g2_nand3_1 _18080_ (.B(_11261_),
    .C(_11262_),
    .A(net599),
    .Y(_11263_));
 sg13g2_nor2_1 _18081_ (.A(_11157_),
    .B(net690),
    .Y(_11264_));
 sg13g2_o21ai_1 _18082_ (.B1(_11264_),
    .Y(_11265_),
    .A1(_11261_),
    .A2(_11262_));
 sg13g2_nand2_1 _18083_ (.Y(_11266_),
    .A(_11263_),
    .B(_11265_));
 sg13g2_o21ai_1 _18084_ (.B1(_11266_),
    .Y(_11267_),
    .A1(_11256_),
    .A2(_11259_));
 sg13g2_nor2_1 _18085_ (.A(net1127),
    .B(net690),
    .Y(_11268_));
 sg13g2_and2_1 _18086_ (.A(net263),
    .B(_11268_),
    .X(_11269_));
 sg13g2_nor3_1 _18087_ (.A(_11164_),
    .B(net1127),
    .C(net690),
    .Y(_11270_));
 sg13g2_o21ai_1 _18088_ (.B1(_11266_),
    .Y(_11271_),
    .A1(_11269_),
    .A2(_11270_));
 sg13g2_nor2_1 _18089_ (.A(net224),
    .B(_11258_),
    .Y(_11272_));
 sg13g2_a221oi_1 _18090_ (.B2(net337),
    .C1(_11272_),
    .B1(_11270_),
    .A1(_11256_),
    .Y(_11273_),
    .A2(_11268_));
 sg13g2_nor2_1 _18091_ (.A(net266),
    .B(_11059_),
    .Y(_11274_));
 sg13g2_nor2_1 _18092_ (.A(_11062_),
    .B(net267),
    .Y(_11275_));
 sg13g2_nor3_1 _18093_ (.A(_11236_),
    .B(_11274_),
    .C(_11275_),
    .Y(_11276_));
 sg13g2_nand2_1 _18094_ (.Y(_11277_),
    .A(_11228_),
    .B(_11276_));
 sg13g2_and4_1 _18095_ (.A(_11267_),
    .B(_11271_),
    .C(_11273_),
    .D(_11277_),
    .X(_11278_));
 sg13g2_nand2b_1 _18096_ (.Y(_11279_),
    .B(net1040),
    .A_N(_08841_));
 sg13g2_buf_1 _18097_ (.A(_11279_),
    .X(_11280_));
 sg13g2_and3_1 _18098_ (.X(_11281_),
    .A(\cpu.ex.r_11[10] ),
    .B(net770),
    .C(net676));
 sg13g2_a221oi_1 _18099_ (.B2(_10891_),
    .C1(_11281_),
    .B1(_10959_),
    .A1(\cpu.ex.r_10[10] ),
    .Y(_11282_),
    .A2(_10990_));
 sg13g2_nand2_1 _18100_ (.Y(_11283_),
    .A(\cpu.ex.r_lr[10] ),
    .B(_11047_));
 sg13g2_mux2_1 _18101_ (.A0(_11282_),
    .A1(_11283_),
    .S(net602),
    .X(_11284_));
 sg13g2_nor2_1 _18102_ (.A(net604),
    .B(_11284_),
    .Y(_11285_));
 sg13g2_nand3_1 _18103_ (.B(net674),
    .C(net603),
    .A(_10887_),
    .Y(_11286_));
 sg13g2_nand3_1 _18104_ (.B(_11144_),
    .C(net605),
    .A(\cpu.ex.r_9[10] ),
    .Y(_11287_));
 sg13g2_a21oi_1 _18105_ (.A1(_11286_),
    .A2(_11287_),
    .Y(_11288_),
    .B1(net673));
 sg13g2_nand3_1 _18106_ (.B(net677),
    .C(net603),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_11289_));
 sg13g2_nand3_1 _18107_ (.B(net765),
    .C(net605),
    .A(\cpu.ex.r_8[10] ),
    .Y(_11290_));
 sg13g2_a21oi_1 _18108_ (.A1(_11289_),
    .A2(_11290_),
    .Y(_11291_),
    .B1(net674));
 sg13g2_nand2_1 _18109_ (.Y(_11292_),
    .A(\cpu.ex.r_12[10] ),
    .B(_10355_));
 sg13g2_nor2b_1 _18110_ (.A(_00270_),
    .B_N(net665),
    .Y(_11293_));
 sg13g2_nor2b_1 _18111_ (.A(net600),
    .B_N(\cpu.ex.r_13[10] ),
    .Y(_11294_));
 sg13g2_o21ai_1 _18112_ (.B1(net677),
    .Y(_11295_),
    .A1(_11293_),
    .A2(_11294_));
 sg13g2_nand2_1 _18113_ (.Y(_11296_),
    .A(net606),
    .B(net674));
 sg13g2_a21oi_1 _18114_ (.A1(_11292_),
    .A2(_11295_),
    .Y(_11297_),
    .B1(_11296_));
 sg13g2_and2_1 _18115_ (.A(\cpu.ex.r_14[10] ),
    .B(net676),
    .X(_11298_));
 sg13g2_a21oi_1 _18116_ (.A1(\cpu.ex.r_stmp[10] ),
    .A2(net754),
    .Y(_11299_),
    .B1(_11298_));
 sg13g2_nor4_1 _18117_ (.A(net607),
    .B(net602),
    .C(net752),
    .D(_11299_),
    .Y(_11300_));
 sg13g2_or4_1 _18118_ (.A(_11288_),
    .B(_11291_),
    .C(_11297_),
    .D(_11300_),
    .X(_11301_));
 sg13g2_o21ai_1 _18119_ (.B1(net601),
    .Y(_11302_),
    .A1(_11285_),
    .A2(_11301_));
 sg13g2_nand2_1 _18120_ (.Y(_11303_),
    .A(_10903_),
    .B(_10292_));
 sg13g2_a21oi_1 _18121_ (.A1(_11302_),
    .A2(_11303_),
    .Y(_11304_),
    .B1(net877));
 sg13g2_nand2_1 _18122_ (.Y(_11305_),
    .A(net877),
    .B(\cpu.dec.imm[10] ));
 sg13g2_nand3b_1 _18123_ (.B(_11305_),
    .C(net876),
    .Y(_11306_),
    .A_N(_11304_));
 sg13g2_buf_2 _18124_ (.A(_11306_),
    .X(_11307_));
 sg13g2_and2_1 _18125_ (.A(_11280_),
    .B(_11307_),
    .X(_11308_));
 sg13g2_buf_2 _18126_ (.A(_11308_),
    .X(_11309_));
 sg13g2_buf_1 _18127_ (.A(_00303_),
    .X(_11310_));
 sg13g2_nor2_1 _18128_ (.A(_11310_),
    .B(net690),
    .Y(_11311_));
 sg13g2_buf_2 _18129_ (.A(_00304_),
    .X(_11312_));
 sg13g2_nor2_1 _18130_ (.A(_10361_),
    .B(\cpu.dec.imm[9] ),
    .Y(_11313_));
 sg13g2_nor2_1 _18131_ (.A(_08824_),
    .B(_11120_),
    .Y(_11314_));
 sg13g2_a21oi_2 _18132_ (.B1(_11314_),
    .Y(_11315_),
    .A2(_11313_),
    .A1(_11122_));
 sg13g2_nor2b_1 _18133_ (.A(_00269_),
    .B_N(_10315_),
    .Y(_11316_));
 sg13g2_a21oi_1 _18134_ (.A1(\cpu.ex.r_11[9] ),
    .A2(net752),
    .Y(_11317_),
    .B1(_11316_));
 sg13g2_nand3_1 _18135_ (.B(_10989_),
    .C(net672),
    .A(\cpu.ex.r_epc[9] ),
    .Y(_11318_));
 sg13g2_o21ai_1 _18136_ (.B1(_11318_),
    .Y(_11319_),
    .A1(_11029_),
    .A2(_11317_));
 sg13g2_a22oi_1 _18137_ (.Y(_11320_),
    .B1(net763),
    .B2(\cpu.ex.r_13[9] ),
    .A2(net672),
    .A1(\cpu.ex.r_lr[9] ));
 sg13g2_nor2_1 _18138_ (.A(_11100_),
    .B(_11320_),
    .Y(_11321_));
 sg13g2_o21ai_1 _18139_ (.B1(_10296_),
    .Y(_11322_),
    .A1(_11319_),
    .A2(_11321_));
 sg13g2_nand3_1 _18140_ (.B(net878),
    .C(_10983_),
    .A(\cpu.ex.r_mult[25] ),
    .Y(_11323_));
 sg13g2_nand3_1 _18141_ (.B(net765),
    .C(net764),
    .A(\cpu.ex.r_10[9] ),
    .Y(_11324_));
 sg13g2_a21oi_1 _18142_ (.A1(_11323_),
    .A2(_11324_),
    .Y(_11325_),
    .B1(net602));
 sg13g2_a22oi_1 _18143_ (.Y(_11326_),
    .B1(_11132_),
    .B2(\cpu.ex.r_14[9] ),
    .A2(_11130_),
    .A1(\cpu.ex.r_8[9] ));
 sg13g2_nor2_1 _18144_ (.A(_11036_),
    .B(_11326_),
    .Y(_11327_));
 sg13g2_nand3_1 _18145_ (.B(net878),
    .C(net675),
    .A(\cpu.ex.r_9[9] ),
    .Y(_11328_));
 sg13g2_nand3_1 _18146_ (.B(_10336_),
    .C(_10325_),
    .A(\cpu.ex.r_sp[9] ),
    .Y(_11329_));
 sg13g2_a21oi_1 _18147_ (.A1(_11328_),
    .A2(_11329_),
    .Y(_11330_),
    .B1(_10316_));
 sg13g2_a22oi_1 _18148_ (.Y(_11331_),
    .B1(net675),
    .B2(\cpu.ex.r_12[9] ),
    .A2(_10325_),
    .A1(\cpu.ex.r_stmp[9] ));
 sg13g2_nor2b_1 _18149_ (.A(_11331_),
    .B_N(_10952_),
    .Y(_11332_));
 sg13g2_nor4_1 _18150_ (.A(_11325_),
    .B(_11327_),
    .C(_11330_),
    .D(_11332_),
    .Y(_11333_));
 sg13g2_a21o_1 _18151_ (.A2(_11333_),
    .A1(_11322_),
    .B1(net540),
    .X(_11334_));
 sg13g2_buf_1 _18152_ (.A(_11334_),
    .X(_11335_));
 sg13g2_nand2_1 _18153_ (.Y(_11336_),
    .A(_10819_),
    .B(net608));
 sg13g2_nand3_1 _18154_ (.B(_11335_),
    .C(_11336_),
    .A(_11097_),
    .Y(_11337_));
 sg13g2_buf_1 _18155_ (.A(_11337_),
    .X(_11338_));
 sg13g2_nand2_1 _18156_ (.Y(_11339_),
    .A(_11315_),
    .B(_11338_));
 sg13g2_buf_1 _18157_ (.A(_11339_),
    .X(_11340_));
 sg13g2_xnor2_1 _18158_ (.Y(_11341_),
    .A(_11312_),
    .B(_11340_));
 sg13g2_nand3_1 _18159_ (.B(_11311_),
    .C(_11341_),
    .A(_11309_),
    .Y(_11342_));
 sg13g2_a21o_1 _18160_ (.A2(_11313_),
    .A1(net876),
    .B1(_11314_),
    .X(_11343_));
 sg13g2_buf_1 _18161_ (.A(_11343_),
    .X(_11344_));
 sg13g2_and3_1 _18162_ (.X(_11345_),
    .A(_11097_),
    .B(_11335_),
    .C(_11336_));
 sg13g2_buf_2 _18163_ (.A(_11345_),
    .X(_11346_));
 sg13g2_o21ai_1 _18164_ (.B1(_11312_),
    .Y(_11347_),
    .A1(_11344_),
    .A2(_11346_));
 sg13g2_nor2_1 _18165_ (.A(_11312_),
    .B(_09380_),
    .Y(_11348_));
 sg13g2_nand3_1 _18166_ (.B(_11338_),
    .C(_11348_),
    .A(_11315_),
    .Y(_11349_));
 sg13g2_inv_1 _18167_ (.Y(_11350_),
    .A(_11310_));
 sg13g2_a21oi_1 _18168_ (.A1(_11347_),
    .A2(_11349_),
    .Y(_11351_),
    .B1(_11350_));
 sg13g2_nor2_1 _18169_ (.A(_11344_),
    .B(_11346_),
    .Y(_11352_));
 sg13g2_buf_2 _18170_ (.A(_11352_),
    .X(_11353_));
 sg13g2_nor2_1 _18171_ (.A(_11257_),
    .B(_11353_),
    .Y(_11354_));
 sg13g2_nand2_1 _18172_ (.Y(_11355_),
    .A(_11280_),
    .B(_11307_));
 sg13g2_buf_1 _18173_ (.A(_11355_),
    .X(_11356_));
 sg13g2_o21ai_1 _18174_ (.B1(net169),
    .Y(_11357_),
    .A1(_11351_),
    .A2(_11354_));
 sg13g2_a22oi_1 _18175_ (.Y(_11358_),
    .B1(net763),
    .B2(\cpu.ex.r_13[8] ),
    .A2(_10350_),
    .A1(\cpu.ex.r_lr[8] ));
 sg13g2_nand2b_1 _18176_ (.Y(_11359_),
    .B(_11205_),
    .A_N(_11358_));
 sg13g2_nor2_1 _18177_ (.A(_10329_),
    .B(_11029_),
    .Y(_11360_));
 sg13g2_and2_1 _18178_ (.A(_10350_),
    .B(_11017_),
    .X(_11361_));
 sg13g2_nand2b_1 _18179_ (.Y(_11362_),
    .B(_10295_),
    .A_N(_00268_));
 sg13g2_nand2b_1 _18180_ (.Y(_11363_),
    .B(\cpu.ex.r_14[8] ),
    .A_N(_10295_));
 sg13g2_a21oi_1 _18181_ (.A1(_11362_),
    .A2(_11363_),
    .Y(_11364_),
    .B1(_11067_));
 sg13g2_a221oi_1 _18182_ (.B2(\cpu.ex.r_epc[8] ),
    .C1(_11364_),
    .B1(_11361_),
    .A1(\cpu.ex.r_10[8] ),
    .Y(_11365_),
    .A2(_11360_));
 sg13g2_mux2_1 _18183_ (.A0(\cpu.ex.r_8[8] ),
    .A1(\cpu.ex.r_12[8] ),
    .S(net753),
    .X(_11366_));
 sg13g2_mux2_1 _18184_ (.A0(_10802_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net753),
    .X(_11367_));
 sg13g2_a22oi_1 _18185_ (.Y(_11368_),
    .B1(_11367_),
    .B2(_10326_),
    .A2(_11366_),
    .A1(_10314_));
 sg13g2_or2_1 _18186_ (.X(_11369_),
    .B(_11368_),
    .A(net677));
 sg13g2_nand3b_1 _18187_ (.B(_10301_),
    .C(\cpu.ex.r_11[8] ),
    .Y(_11370_),
    .A_N(_10316_));
 sg13g2_nand3b_1 _18188_ (.B(net767),
    .C(\cpu.ex.r_mult[24] ),
    .Y(_11371_),
    .A_N(net676));
 sg13g2_a21oi_1 _18189_ (.A1(_11370_),
    .A2(_11371_),
    .Y(_11372_),
    .B1(_10334_));
 sg13g2_and3_1 _18190_ (.X(_11373_),
    .A(\cpu.ex.r_9[8] ),
    .B(net752),
    .C(net675));
 sg13g2_o21ai_1 _18191_ (.B1(net677),
    .Y(_11374_),
    .A1(_11372_),
    .A2(_11373_));
 sg13g2_nand4_1 _18192_ (.B(_11365_),
    .C(_11369_),
    .A(_11359_),
    .Y(_11375_),
    .D(_11374_));
 sg13g2_a221oi_1 _18193_ (.B2(_11375_),
    .C1(_11165_),
    .B1(net601),
    .A1(_09226_),
    .Y(_11376_),
    .A2(_10291_));
 sg13g2_buf_1 _18194_ (.A(_11376_),
    .X(_11377_));
 sg13g2_or4_1 _18195_ (.A(_10361_),
    .B(net1040),
    .C(_10274_),
    .D(\cpu.dec.imm[8] ),
    .X(_11378_));
 sg13g2_o21ai_1 _18196_ (.B1(_11378_),
    .Y(_11379_),
    .A1(_08850_),
    .A2(net1031));
 sg13g2_buf_1 _18197_ (.A(_11379_),
    .X(_11380_));
 sg13g2_or2_1 _18198_ (.X(_11381_),
    .B(_11380_),
    .A(_11377_));
 sg13g2_buf_2 _18199_ (.A(_11381_),
    .X(_11382_));
 sg13g2_buf_8 _18200_ (.A(_11382_),
    .X(_11383_));
 sg13g2_buf_1 _18201_ (.A(_00305_),
    .X(_11384_));
 sg13g2_nor2_1 _18202_ (.A(_11384_),
    .B(_09390_),
    .Y(_11385_));
 sg13g2_xnor2_1 _18203_ (.Y(_11386_),
    .A(net208),
    .B(_11385_));
 sg13g2_a21oi_2 _18204_ (.B1(_11386_),
    .Y(_11387_),
    .A2(_11357_),
    .A1(_11342_));
 sg13g2_inv_1 _18205_ (.Y(_11388_),
    .A(_11387_));
 sg13g2_a21oi_1 _18206_ (.A1(_11254_),
    .A2(_11278_),
    .Y(_11389_),
    .B1(_11388_));
 sg13g2_nor2_1 _18207_ (.A(net821),
    .B(net1031),
    .Y(_11390_));
 sg13g2_nand3_1 _18208_ (.B(net607),
    .C(net603),
    .A(\cpu.ex.r_epc[12] ),
    .Y(_11391_));
 sg13g2_nand3_1 _18209_ (.B(net673),
    .C(net605),
    .A(\cpu.ex.r_8[12] ),
    .Y(_11392_));
 sg13g2_a21o_1 _18210_ (.A2(_11392_),
    .A1(_11391_),
    .B1(net604),
    .X(_11393_));
 sg13g2_a22oi_1 _18211_ (.Y(_11394_),
    .B1(_10314_),
    .B2(\cpu.ex.r_13[12] ),
    .A2(net603),
    .A1(_10852_));
 sg13g2_and2_1 _18212_ (.A(net677),
    .B(_10317_),
    .X(_11395_));
 sg13g2_buf_1 _18213_ (.A(_11395_),
    .X(_11396_));
 sg13g2_nand2b_1 _18214_ (.Y(_11397_),
    .B(_11396_),
    .A_N(_11394_));
 sg13g2_nand2_1 _18215_ (.Y(_11398_),
    .A(\cpu.ex.r_11[12] ),
    .B(net600));
 sg13g2_nand2b_1 _18216_ (.Y(_11399_),
    .B(\cpu.ex.r_9[12] ),
    .A_N(net600));
 sg13g2_a21oi_1 _18217_ (.A1(_11398_),
    .A2(_11399_),
    .Y(_11400_),
    .B1(_11074_));
 sg13g2_a21oi_1 _18218_ (.A1(\cpu.ex.r_lr[12] ),
    .A2(_11197_),
    .Y(_11401_),
    .B1(_11400_));
 sg13g2_a22oi_1 _18219_ (.Y(_11402_),
    .B1(_10959_),
    .B2(\cpu.ex.r_stmp[12] ),
    .A2(_10998_),
    .A1(_10846_));
 sg13g2_nand2b_1 _18220_ (.Y(_11403_),
    .B(_11132_),
    .A_N(_11402_));
 sg13g2_nand4_1 _18221_ (.B(_11397_),
    .C(_11401_),
    .A(_11393_),
    .Y(_11404_),
    .D(_11403_));
 sg13g2_nor2_1 _18222_ (.A(net752),
    .B(_11041_),
    .Y(_11405_));
 sg13g2_and2_1 _18223_ (.A(net673),
    .B(_10305_),
    .X(_11406_));
 sg13g2_a22oi_1 _18224_ (.Y(_11407_),
    .B1(_11406_),
    .B2(_10854_),
    .A2(_11405_),
    .A1(_10851_));
 sg13g2_mux2_1 _18225_ (.A0(\cpu.ex.r_10[12] ),
    .A1(\cpu.ex.r_14[12] ),
    .S(net674),
    .X(_11408_));
 sg13g2_a22oi_1 _18226_ (.Y(_11409_),
    .B1(_11408_),
    .B2(net600),
    .A2(_10307_),
    .A1(\cpu.ex.r_12[12] ));
 sg13g2_nand2b_1 _18227_ (.Y(_11410_),
    .B(_10990_),
    .A_N(_11409_));
 sg13g2_o21ai_1 _18228_ (.B1(_11410_),
    .Y(_11411_),
    .A1(net606),
    .A2(_11407_));
 sg13g2_o21ai_1 _18229_ (.B1(net601),
    .Y(_11412_),
    .A1(_11404_),
    .A2(_11411_));
 sg13g2_buf_1 _18230_ (.A(net780),
    .X(_11413_));
 sg13g2_nand2_1 _18231_ (.Y(_11414_),
    .A(net664),
    .B(net541));
 sg13g2_a21oi_1 _18232_ (.A1(_11412_),
    .A2(_11414_),
    .Y(_11415_),
    .B1(net877));
 sg13g2_inv_1 _18233_ (.Y(_11416_),
    .A(\cpu.dec.imm[12] ));
 sg13g2_nor2_1 _18234_ (.A(net1041),
    .B(_11416_),
    .Y(_11417_));
 sg13g2_nor3_2 _18235_ (.A(_10276_),
    .B(_11415_),
    .C(_11417_),
    .Y(_11418_));
 sg13g2_buf_2 _18236_ (.A(_00302_),
    .X(_11419_));
 sg13g2_o21ai_1 _18237_ (.B1(_11419_),
    .Y(_11420_),
    .A1(_11390_),
    .A2(_11418_));
 sg13g2_or3_1 _18238_ (.A(_11419_),
    .B(_11390_),
    .C(_11418_),
    .X(_11421_));
 sg13g2_nand2b_1 _18239_ (.Y(_11422_),
    .B(_10364_),
    .A_N(net714));
 sg13g2_buf_1 _18240_ (.A(_11422_),
    .X(_11423_));
 sg13g2_nand3_1 _18241_ (.B(net600),
    .C(net672),
    .A(\cpu.ex.r_epc[13] ),
    .Y(_11424_));
 sg13g2_nand3_1 _18242_ (.B(net602),
    .C(net763),
    .A(\cpu.ex.r_13[13] ),
    .Y(_11425_));
 sg13g2_nand3_1 _18243_ (.B(_11424_),
    .C(_11425_),
    .A(_10297_),
    .Y(_11426_));
 sg13g2_nand3_1 _18244_ (.B(net604),
    .C(net603),
    .A(\cpu.ex.r_stmp[13] ),
    .Y(_11427_));
 sg13g2_nand3_1 _18245_ (.B(_11144_),
    .C(net605),
    .A(\cpu.ex.r_8[13] ),
    .Y(_11428_));
 sg13g2_nand3_1 _18246_ (.B(_11427_),
    .C(_11428_),
    .A(_10337_),
    .Y(_11429_));
 sg13g2_nand2_1 _18247_ (.Y(_11430_),
    .A(\cpu.ex.r_12[13] ),
    .B(net768));
 sg13g2_nand3_1 _18248_ (.B(net607),
    .C(_10305_),
    .A(\cpu.ex.r_11[13] ),
    .Y(_11431_));
 sg13g2_o21ai_1 _18249_ (.B1(_11431_),
    .Y(_11432_),
    .A1(net607),
    .A2(_11430_));
 sg13g2_buf_1 _18250_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_11433_));
 sg13g2_mux2_1 _18251_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(_11433_),
    .S(net674),
    .X(_11434_));
 sg13g2_a22oi_1 _18252_ (.Y(_11435_),
    .B1(_11434_),
    .B2(net754),
    .A2(net764),
    .A1(\cpu.ex.r_9[13] ));
 sg13g2_nor2_1 _18253_ (.A(_11041_),
    .B(_11435_),
    .Y(_11436_));
 sg13g2_a221oi_1 _18254_ (.B2(net606),
    .C1(_11436_),
    .B1(_11432_),
    .A1(_11426_),
    .Y(_11437_),
    .A2(_11429_));
 sg13g2_mux2_1 _18255_ (.A0(\cpu.ex.r_10[13] ),
    .A1(\cpu.ex.r_14[13] ),
    .S(_10317_),
    .X(_11438_));
 sg13g2_a22oi_1 _18256_ (.Y(_11439_),
    .B1(_11438_),
    .B2(net673),
    .A2(_11396_),
    .A1(_10776_));
 sg13g2_a221oi_1 _18257_ (.B2(_10789_),
    .C1(_10302_),
    .B1(_11396_),
    .A1(_10783_),
    .Y(_11440_),
    .A2(_11110_));
 sg13g2_a21oi_1 _18258_ (.A1(net606),
    .A2(_11439_),
    .Y(_11441_),
    .B1(_11440_));
 sg13g2_nand2_1 _18259_ (.Y(_11442_),
    .A(net600),
    .B(_11441_));
 sg13g2_a21oi_1 _18260_ (.A1(_11437_),
    .A2(_11442_),
    .Y(_11443_),
    .B1(net540));
 sg13g2_buf_1 _18261_ (.A(net1093),
    .X(_11444_));
 sg13g2_nor3_1 _18262_ (.A(net875),
    .B(_10279_),
    .C(_10289_),
    .Y(_11445_));
 sg13g2_nor3_1 _18263_ (.A(net877),
    .B(_11443_),
    .C(_11445_),
    .Y(_11446_));
 sg13g2_nor2_1 _18264_ (.A(net1041),
    .B(\cpu.dec.imm[13] ),
    .Y(_11447_));
 sg13g2_o21ai_1 _18265_ (.B1(net876),
    .Y(_11448_),
    .A1(_11446_),
    .A2(_11447_));
 sg13g2_buf_2 _18266_ (.A(_11448_),
    .X(_11449_));
 sg13g2_nand3_1 _18267_ (.B(_11423_),
    .C(_11449_),
    .A(_10852_),
    .Y(_11450_));
 sg13g2_a21oi_1 _18268_ (.A1(_11420_),
    .A2(_11421_),
    .Y(_11451_),
    .B1(_11450_));
 sg13g2_and2_1 _18269_ (.A(_11423_),
    .B(_11449_),
    .X(_11452_));
 sg13g2_buf_2 _18270_ (.A(_11452_),
    .X(_11453_));
 sg13g2_or2_1 _18271_ (.X(_11454_),
    .B(_11418_),
    .A(_11390_));
 sg13g2_buf_2 _18272_ (.A(_11454_),
    .X(_11455_));
 sg13g2_nor4_1 _18273_ (.A(_10852_),
    .B(_11419_),
    .C(_11453_),
    .D(_11455_),
    .Y(_11456_));
 sg13g2_o21ai_1 _18274_ (.B1(net599),
    .Y(_11457_),
    .A1(_11451_),
    .A2(_11456_));
 sg13g2_buf_1 _18275_ (.A(_11453_),
    .X(_11458_));
 sg13g2_nor2_1 _18276_ (.A(_11390_),
    .B(_11418_),
    .Y(_11459_));
 sg13g2_buf_1 _18277_ (.A(_11459_),
    .X(_11460_));
 sg13g2_inv_4 _18278_ (.A(_10852_),
    .Y(_11461_));
 sg13g2_a21oi_1 _18279_ (.A1(_11461_),
    .A2(_11419_),
    .Y(_11462_),
    .B1(net609));
 sg13g2_or3_1 _18280_ (.A(net133),
    .B(net191),
    .C(_11462_),
    .X(_11463_));
 sg13g2_nand2_1 _18281_ (.Y(_11464_),
    .A(_10925_),
    .B(net608));
 sg13g2_nand3_1 _18282_ (.B(net767),
    .C(_10325_),
    .A(\cpu.ex.r_mult[27] ),
    .Y(_11465_));
 sg13g2_nand3_1 _18283_ (.B(net752),
    .C(net675),
    .A(\cpu.ex.r_9[11] ),
    .Y(_11466_));
 sg13g2_and2_1 _18284_ (.A(_11465_),
    .B(_11466_),
    .X(_11467_));
 sg13g2_mux4_1 _18285_ (.S0(net767),
    .A0(_10907_),
    .A1(\cpu.ex.r_stmp[11] ),
    .A2(\cpu.ex.r_10[11] ),
    .A3(\cpu.ex.r_14[11] ),
    .S1(net676),
    .X(_11468_));
 sg13g2_nand2_1 _18286_ (.Y(_11469_),
    .A(_10944_),
    .B(_11468_));
 sg13g2_o21ai_1 _18287_ (.B1(_11469_),
    .Y(_11470_),
    .A1(net765),
    .A2(_11467_));
 sg13g2_inv_1 _18288_ (.Y(_11471_),
    .A(\cpu.ex.r_12[11] ));
 sg13g2_or2_1 _18289_ (.X(_11472_),
    .B(net766),
    .A(net878));
 sg13g2_nand3b_1 _18290_ (.B(net878),
    .C(net665),
    .Y(_11473_),
    .A_N(_00271_));
 sg13g2_o21ai_1 _18291_ (.B1(_11473_),
    .Y(_11474_),
    .A1(_11471_),
    .A2(_11472_));
 sg13g2_nand3b_1 _18292_ (.B(net665),
    .C(\cpu.ex.r_11[11] ),
    .Y(_11475_),
    .A_N(net753));
 sg13g2_nand3b_1 _18293_ (.B(net767),
    .C(\cpu.ex.r_13[11] ),
    .Y(_11476_),
    .A_N(net665));
 sg13g2_nand3_1 _18294_ (.B(_11475_),
    .C(_11476_),
    .A(net770),
    .Y(_11477_));
 sg13g2_a21o_1 _18295_ (.A2(_11130_),
    .A1(\cpu.ex.r_8[11] ),
    .B1(net770),
    .X(_11478_));
 sg13g2_a22oi_1 _18296_ (.Y(_11479_),
    .B1(_11477_),
    .B2(_11478_),
    .A2(_11474_),
    .A1(net674));
 sg13g2_mux2_1 _18297_ (.A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net665),
    .X(_11480_));
 sg13g2_nand3_1 _18298_ (.B(net672),
    .C(_11480_),
    .A(net677),
    .Y(_11481_));
 sg13g2_o21ai_1 _18299_ (.B1(_11481_),
    .Y(_11482_),
    .A1(net754),
    .A2(_11479_));
 sg13g2_o21ai_1 _18300_ (.B1(net601),
    .Y(_11483_),
    .A1(_11470_),
    .A2(_11482_));
 sg13g2_nand3_1 _18301_ (.B(_11464_),
    .C(_11483_),
    .A(_11097_),
    .Y(_11484_));
 sg13g2_buf_1 _18302_ (.A(_11484_),
    .X(_11485_));
 sg13g2_nor2_1 _18303_ (.A(_10362_),
    .B(\cpu.dec.imm[11] ),
    .Y(_11486_));
 sg13g2_a22oi_1 _18304_ (.Y(_11487_),
    .B1(_11122_),
    .B2(_11486_),
    .A2(net1040),
    .A1(_08882_));
 sg13g2_buf_1 _18305_ (.A(_11487_),
    .X(_11488_));
 sg13g2_and2_1 _18306_ (.A(_11485_),
    .B(_11488_),
    .X(_11489_));
 sg13g2_buf_2 _18307_ (.A(_11489_),
    .X(_11490_));
 sg13g2_buf_1 _18308_ (.A(_11490_),
    .X(_11491_));
 sg13g2_nand2_1 _18309_ (.Y(_11492_),
    .A(_10887_),
    .B(net599));
 sg13g2_xnor2_1 _18310_ (.Y(_11493_),
    .A(net190),
    .B(_11492_));
 sg13g2_a21oi_1 _18311_ (.A1(_11457_),
    .A2(_11463_),
    .Y(_11494_),
    .B1(_11493_));
 sg13g2_inv_1 _18312_ (.Y(_11495_),
    .A(_11384_));
 sg13g2_o21ai_1 _18313_ (.B1(_11495_),
    .Y(_11496_),
    .A1(_11377_),
    .A2(_11380_));
 sg13g2_a21o_1 _18314_ (.A2(_11338_),
    .A1(_11315_),
    .B1(_11496_),
    .X(_11497_));
 sg13g2_inv_1 _18315_ (.Y(_11498_),
    .A(_11312_));
 sg13g2_nand3_1 _18316_ (.B(_11495_),
    .C(net208),
    .A(_11498_),
    .Y(_11499_));
 sg13g2_o21ai_1 _18317_ (.B1(_11498_),
    .Y(_11500_),
    .A1(_11344_),
    .A2(_11346_));
 sg13g2_nand3_1 _18318_ (.B(_11499_),
    .C(_11500_),
    .A(_11497_),
    .Y(_11501_));
 sg13g2_and2_1 _18319_ (.A(_11310_),
    .B(_11280_),
    .X(_11502_));
 sg13g2_a21oi_1 _18320_ (.A1(_11307_),
    .A2(_11502_),
    .Y(_11503_),
    .B1(_11490_));
 sg13g2_a221oi_1 _18321_ (.B2(_10888_),
    .C1(_11310_),
    .B1(_11490_),
    .A1(_11280_),
    .Y(_11504_),
    .A2(_11307_));
 sg13g2_a21oi_1 _18322_ (.A1(_11501_),
    .A2(_11503_),
    .Y(_11505_),
    .B1(_11504_));
 sg13g2_nand2_1 _18323_ (.Y(_11506_),
    .A(_11485_),
    .B(_11488_));
 sg13g2_buf_1 _18324_ (.A(_11506_),
    .X(_11507_));
 sg13g2_a21oi_1 _18325_ (.A1(_11307_),
    .A2(_11502_),
    .Y(_11508_),
    .B1(_10888_));
 sg13g2_a22oi_1 _18326_ (.Y(_11509_),
    .B1(_11501_),
    .B2(_11508_),
    .A2(net207),
    .A1(_10887_));
 sg13g2_nand3_1 _18327_ (.B(_11423_),
    .C(_11449_),
    .A(_11461_),
    .Y(_11510_));
 sg13g2_buf_1 _18328_ (.A(_11510_),
    .X(_11511_));
 sg13g2_nand3_1 _18329_ (.B(_11455_),
    .C(_11511_),
    .A(net599),
    .Y(_11512_));
 sg13g2_nor2_2 _18330_ (.A(_11419_),
    .B(net609),
    .Y(_11513_));
 sg13g2_nand2_1 _18331_ (.Y(_11514_),
    .A(_11511_),
    .B(_11513_));
 sg13g2_a22oi_1 _18332_ (.Y(_11515_),
    .B1(_11512_),
    .B2(_11514_),
    .A2(_11509_),
    .A1(_11505_));
 sg13g2_buf_1 _18333_ (.A(net599),
    .X(_11516_));
 sg13g2_nor2_1 _18334_ (.A(_11461_),
    .B(net133),
    .Y(_11517_));
 sg13g2_and2_1 _18335_ (.A(_11455_),
    .B(_11513_),
    .X(_11518_));
 sg13g2_a22oi_1 _18336_ (.Y(_11519_),
    .B1(_11511_),
    .B2(_11518_),
    .A2(_11517_),
    .A1(net537));
 sg13g2_nand2b_1 _18337_ (.Y(_11520_),
    .B(_11519_),
    .A_N(_11515_));
 sg13g2_a21o_1 _18338_ (.A2(_11494_),
    .A1(_11389_),
    .B1(_11520_),
    .X(_11521_));
 sg13g2_buf_1 _18339_ (.A(_11521_),
    .X(_11522_));
 sg13g2_buf_1 _18340_ (.A(net688),
    .X(_11523_));
 sg13g2_a221oi_1 _18341_ (.B2(_10861_),
    .C1(net606),
    .B1(_11406_),
    .A1(_10872_),
    .Y(_11524_),
    .A2(_11405_));
 sg13g2_a22oi_1 _18342_ (.Y(_11525_),
    .B1(_11017_),
    .B2(_10870_),
    .A2(_10355_),
    .A1(\cpu.ex.r_12[14] ));
 sg13g2_mux2_1 _18343_ (.A0(\cpu.ex.r_9[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net600),
    .X(_11526_));
 sg13g2_a221oi_1 _18344_ (.B2(net607),
    .C1(net604),
    .B1(_11526_),
    .A1(\cpu.ex.r_10[14] ),
    .Y(_11527_),
    .A2(_10944_));
 sg13g2_a21oi_1 _18345_ (.A1(net604),
    .A2(_11525_),
    .Y(_11528_),
    .B1(_11527_));
 sg13g2_nor2_1 _18346_ (.A(net754),
    .B(_11528_),
    .Y(_11529_));
 sg13g2_a22oi_1 _18347_ (.Y(_11530_),
    .B1(net605),
    .B2(\cpu.ex.r_13[14] ),
    .A2(net603),
    .A1(\cpu.ex.r_mult[30] ));
 sg13g2_nor2_1 _18348_ (.A(_11109_),
    .B(_11530_),
    .Y(_11531_));
 sg13g2_and2_1 _18349_ (.A(\cpu.ex.r_lr[14] ),
    .B(_11197_),
    .X(_11532_));
 sg13g2_nand3_1 _18350_ (.B(net604),
    .C(net603),
    .A(\cpu.ex.r_stmp[14] ),
    .Y(_11533_));
 sg13g2_nand3_1 _18351_ (.B(net752),
    .C(net605),
    .A(\cpu.ex.r_8[14] ),
    .Y(_11534_));
 sg13g2_a21oi_1 _18352_ (.A1(_11533_),
    .A2(_11534_),
    .Y(_11535_),
    .B1(net607));
 sg13g2_nand3_1 _18353_ (.B(net607),
    .C(net672),
    .A(\cpu.ex.r_epc[14] ),
    .Y(_11536_));
 sg13g2_nand3_1 _18354_ (.B(net673),
    .C(net763),
    .A(\cpu.ex.r_14[14] ),
    .Y(_11537_));
 sg13g2_a21oi_1 _18355_ (.A1(_11536_),
    .A2(_11537_),
    .Y(_11538_),
    .B1(net602));
 sg13g2_nor4_1 _18356_ (.A(_11531_),
    .B(_11532_),
    .C(_11535_),
    .D(_11538_),
    .Y(_11539_));
 sg13g2_o21ai_1 _18357_ (.B1(_11539_),
    .Y(_11540_),
    .A1(_11524_),
    .A2(_11529_));
 sg13g2_a22oi_1 _18358_ (.Y(_11541_),
    .B1(_10937_),
    .B2(_11540_),
    .A2(net541),
    .A1(net598));
 sg13g2_nor2_1 _18359_ (.A(net1041),
    .B(\cpu.dec.imm[14] ),
    .Y(_11542_));
 sg13g2_a21oi_1 _18360_ (.A1(net1041),
    .A2(_11541_),
    .Y(_11543_),
    .B1(_11542_));
 sg13g2_nand2b_1 _18361_ (.Y(_11544_),
    .B(net1040),
    .A_N(_08637_));
 sg13g2_o21ai_1 _18362_ (.B1(_11544_),
    .Y(_11545_),
    .A1(_10276_),
    .A2(_11543_));
 sg13g2_buf_1 _18363_ (.A(_11545_),
    .X(_11546_));
 sg13g2_buf_1 _18364_ (.A(_11546_),
    .X(_11547_));
 sg13g2_nand3_1 _18365_ (.B(_11522_),
    .C(net168),
    .A(_10367_),
    .Y(_11548_));
 sg13g2_buf_8 _18366_ (.A(_11548_),
    .X(_11549_));
 sg13g2_and2_1 _18367_ (.A(_11254_),
    .B(_11278_),
    .X(_11550_));
 sg13g2_buf_2 _18368_ (.A(_11550_),
    .X(_11551_));
 sg13g2_nand3_1 _18369_ (.B(_11494_),
    .C(net168),
    .A(_11387_),
    .Y(_11552_));
 sg13g2_a21oi_1 _18370_ (.A1(_11520_),
    .A2(net168),
    .Y(_11553_),
    .B1(_10367_));
 sg13g2_o21ai_1 _18371_ (.B1(_11553_),
    .Y(_11554_),
    .A1(_11551_),
    .A2(_11552_));
 sg13g2_buf_1 _18372_ (.A(_00301_),
    .X(_11555_));
 sg13g2_nor2_1 _18373_ (.A(_11555_),
    .B(net609),
    .Y(_11556_));
 sg13g2_nand3_1 _18374_ (.B(_11387_),
    .C(_11494_),
    .A(_10789_),
    .Y(_11557_));
 sg13g2_o21ai_1 _18375_ (.B1(_10789_),
    .Y(_11558_),
    .A1(_11520_),
    .A2(net168));
 sg13g2_o21ai_1 _18376_ (.B1(_11558_),
    .Y(_11559_),
    .A1(_11551_),
    .A2(_11557_));
 sg13g2_inv_1 _18377_ (.Y(_11560_),
    .A(_10363_));
 sg13g2_a22oi_1 _18378_ (.Y(_11561_),
    .B1(net876),
    .B2(_11560_),
    .A2(net1040),
    .A1(net712));
 sg13g2_buf_2 _18379_ (.A(_11561_),
    .X(_11562_));
 sg13g2_a21oi_1 _18380_ (.A1(_11555_),
    .A2(_11562_),
    .Y(_11563_),
    .B1(net609));
 sg13g2_a22oi_1 _18381_ (.Y(_11564_),
    .B1(_11559_),
    .B2(_11563_),
    .A2(_11556_),
    .A1(_11554_));
 sg13g2_buf_8 _18382_ (.A(_11564_),
    .X(_11565_));
 sg13g2_nor2_1 _18383_ (.A(_11377_),
    .B(_11380_),
    .Y(_11566_));
 sg13g2_buf_1 _18384_ (.A(_11566_),
    .X(_11567_));
 sg13g2_nor4_1 _18385_ (.A(_11567_),
    .B(net225),
    .C(net265),
    .D(net190),
    .Y(_11568_));
 sg13g2_nand4_1 _18386_ (.B(_11256_),
    .C(_11546_),
    .A(_10367_),
    .Y(_11569_),
    .D(_11568_));
 sg13g2_buf_1 _18387_ (.A(_11353_),
    .X(_11570_));
 sg13g2_a21o_1 _18388_ (.A2(_11307_),
    .A1(_11280_),
    .B1(net189),
    .X(_11571_));
 sg13g2_nand2_1 _18389_ (.Y(_11572_),
    .A(net267),
    .B(net266));
 sg13g2_nand2_1 _18390_ (.Y(_11573_),
    .A(_11055_),
    .B(_11057_));
 sg13g2_buf_1 _18391_ (.A(_11573_),
    .X(_11574_));
 sg13g2_nand2_1 _18392_ (.Y(_11575_),
    .A(net336),
    .B(_11092_));
 sg13g2_buf_1 _18393_ (.A(_11575_),
    .X(_11576_));
 sg13g2_or2_1 _18394_ (.X(_11577_),
    .B(_11576_),
    .A(_11572_));
 sg13g2_buf_1 _18395_ (.A(_11577_),
    .X(_11578_));
 sg13g2_or4_1 _18396_ (.A(_11453_),
    .B(_11459_),
    .C(_11571_),
    .D(_11578_),
    .X(_11579_));
 sg13g2_buf_1 _18397_ (.A(_11223_),
    .X(_11580_));
 sg13g2_a221oi_1 _18398_ (.B2(_10249_),
    .C1(net1141),
    .B1(net599),
    .A1(_09373_),
    .Y(_11581_),
    .A2(net751));
 sg13g2_o21ai_1 _18399_ (.B1(_11581_),
    .Y(_11582_),
    .A1(_11569_),
    .A2(_11579_));
 sg13g2_buf_1 _18400_ (.A(_11582_),
    .X(_11583_));
 sg13g2_a21o_1 _18401_ (.A2(_11565_),
    .A1(_11549_),
    .B1(net86),
    .X(_11584_));
 sg13g2_nor2_1 _18402_ (.A(_09392_),
    .B(net689),
    .Y(_11585_));
 sg13g2_a21oi_1 _18403_ (.A1(_10610_),
    .A2(_10744_),
    .Y(_11586_),
    .B1(_10931_));
 sg13g2_buf_2 _18404_ (.A(_11586_),
    .X(_11587_));
 sg13g2_buf_1 _18405_ (.A(_11587_),
    .X(_11588_));
 sg13g2_inv_4 _18406_ (.A(_11092_),
    .Y(_11589_));
 sg13g2_nand3b_1 _18407_ (.B(net78),
    .C(_11589_),
    .Y(_11590_),
    .A_N(_11585_));
 sg13g2_nand2b_1 _18408_ (.Y(_11591_),
    .B(_10267_),
    .A_N(_10265_));
 sg13g2_buf_1 _18409_ (.A(_11591_),
    .X(_11592_));
 sg13g2_buf_1 _18410_ (.A(_11592_),
    .X(_11593_));
 sg13g2_a21oi_1 _18411_ (.A1(_11584_),
    .A2(_11590_),
    .Y(_11594_),
    .B1(net425));
 sg13g2_a21o_1 _18412_ (.A2(net340),
    .A1(_10246_),
    .B1(_11594_),
    .X(\cpu.ex.c_mult[0] ));
 sg13g2_buf_1 _18413_ (.A(\cpu.dec.load ),
    .X(_11595_));
 sg13g2_nand2_1 _18414_ (.Y(_11596_),
    .A(net1060),
    .B(_08457_));
 sg13g2_nor2_1 _18415_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11597_));
 sg13g2_nand2_1 _18416_ (.Y(_11598_),
    .A(net1039),
    .B(\cpu.cond[2] ));
 sg13g2_inv_1 _18417_ (.Y(_11599_),
    .A(_08402_));
 sg13g2_a21o_1 _18418_ (.A2(_11598_),
    .A1(_00260_),
    .B1(_11599_),
    .X(_11600_));
 sg13g2_buf_1 _18419_ (.A(_11600_),
    .X(_11601_));
 sg13g2_o21ai_1 _18420_ (.B1(_11601_),
    .Y(_11602_),
    .A1(net1039),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand3b_1 _18421_ (.B(net751),
    .C(_11602_),
    .Y(_11603_),
    .A_N(net1092));
 sg13g2_a21oi_1 _18422_ (.A1(_10649_),
    .A2(\cpu.dec.r_swapsp ),
    .Y(_11604_),
    .B1(_11603_));
 sg13g2_nor2_1 _18423_ (.A(_09303_),
    .B(_09389_),
    .Y(_11605_));
 sg13g2_a21oi_1 _18424_ (.A1(_10249_),
    .A2(_10250_),
    .Y(_11606_),
    .B1(_11605_));
 sg13g2_buf_1 _18425_ (.A(_11606_),
    .X(_11607_));
 sg13g2_a21oi_1 _18426_ (.A1(_11597_),
    .A2(_11604_),
    .Y(_11608_),
    .B1(net188));
 sg13g2_a21oi_1 _18427_ (.A1(_11596_),
    .A2(_11608_),
    .Y(_11609_),
    .B1(_09303_));
 sg13g2_buf_1 _18428_ (.A(_11609_),
    .X(_11610_));
 sg13g2_nand2_1 _18429_ (.Y(_11611_),
    .A(_00312_),
    .B(_11610_));
 sg13g2_buf_1 _18430_ (.A(_11610_),
    .X(_11612_));
 sg13g2_nand2_1 _18431_ (.Y(_11613_),
    .A(_09398_),
    .B(_09829_));
 sg13g2_a21oi_1 _18432_ (.A1(_09831_),
    .A2(_11613_),
    .Y(_11614_),
    .B1(_09834_));
 sg13g2_or2_1 _18433_ (.X(_11615_),
    .B(_11614_),
    .A(_08408_));
 sg13g2_o21ai_1 _18434_ (.B1(_11611_),
    .Y(_11616_),
    .A1(net85),
    .A2(_11615_));
 sg13g2_nand2_1 _18435_ (.Y(_11617_),
    .A(net1092),
    .B(_11616_));
 sg13g2_o21ai_1 _18436_ (.B1(_11617_),
    .Y(_00054_),
    .A1(_11595_),
    .A2(_11611_));
 sg13g2_buf_1 _18437_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11618_));
 sg13g2_nand2_1 _18438_ (.Y(_11619_),
    .A(_09373_),
    .B(_11223_));
 sg13g2_buf_2 _18439_ (.A(_11619_),
    .X(_11620_));
 sg13g2_buf_1 _18440_ (.A(_11620_),
    .X(_11621_));
 sg13g2_buf_8 _18441_ (.A(_11621_),
    .X(_11622_));
 sg13g2_nand2_1 _18442_ (.Y(_11623_),
    .A(_10246_),
    .B(_11622_));
 sg13g2_buf_1 _18443_ (.A(_10933_),
    .X(_11624_));
 sg13g2_nor2_1 _18444_ (.A(net336),
    .B(net77),
    .Y(_11625_));
 sg13g2_mux2_1 _18445_ (.A0(_11623_),
    .A1(_10246_),
    .S(_11625_),
    .X(_11626_));
 sg13g2_nor2_1 _18446_ (.A(_11569_),
    .B(_11579_),
    .Y(_11627_));
 sg13g2_nor2b_1 _18447_ (.A(_11627_),
    .B_N(_11581_),
    .Y(_11628_));
 sg13g2_buf_8 _18448_ (.A(_11628_),
    .X(_11629_));
 sg13g2_buf_1 _18449_ (.A(_10247_),
    .X(_11630_));
 sg13g2_a22oi_1 _18450_ (.Y(_11631_),
    .B1(_11625_),
    .B2(net535),
    .A2(_11629_),
    .A1(_10246_));
 sg13g2_o21ai_1 _18451_ (.B1(_11631_),
    .Y(_11632_),
    .A1(_10250_),
    .A2(_11626_));
 sg13g2_a22oi_1 _18452_ (.Y(_11633_),
    .B1(_11632_),
    .B2(net483),
    .A2(_10271_),
    .A1(_11618_));
 sg13g2_inv_1 _18453_ (.Y(\cpu.ex.c_mult[1] ),
    .A(_11633_));
 sg13g2_nor2_2 _18454_ (.A(_10250_),
    .B(net535),
    .Y(_11634_));
 sg13g2_nand3_1 _18455_ (.B(_11055_),
    .C(_11057_),
    .A(_10246_),
    .Y(_11635_));
 sg13g2_buf_1 _18456_ (.A(_11635_),
    .X(_11636_));
 sg13g2_a21oi_1 _18457_ (.A1(_10981_),
    .A2(_11013_),
    .Y(_11637_),
    .B1(_11618_));
 sg13g2_buf_1 _18458_ (.A(net261),
    .X(_11638_));
 sg13g2_and2_1 _18459_ (.A(_11618_),
    .B(net221),
    .X(_11639_));
 sg13g2_a21oi_1 _18460_ (.A1(_11587_),
    .A2(_11637_),
    .Y(_11640_),
    .B1(_11639_));
 sg13g2_and2_1 _18461_ (.A(net223),
    .B(_11636_),
    .X(_11641_));
 sg13g2_o21ai_1 _18462_ (.B1(_11618_),
    .Y(_11642_),
    .A1(net77),
    .A2(_11641_));
 sg13g2_o21ai_1 _18463_ (.B1(_11642_),
    .Y(_11643_),
    .A1(_11636_),
    .A2(_11640_));
 sg13g2_nor2_1 _18464_ (.A(_10250_),
    .B(_11618_),
    .Y(_11644_));
 sg13g2_a21oi_1 _18465_ (.A1(_11636_),
    .A2(_11644_),
    .Y(_11645_),
    .B1(net610));
 sg13g2_nor3_1 _18466_ (.A(net223),
    .B(net77),
    .C(_11645_),
    .Y(_11646_));
 sg13g2_a221oi_1 _18467_ (.B2(_11643_),
    .C1(_11646_),
    .B1(_11634_),
    .A1(_11618_),
    .Y(_11647_),
    .A2(_11629_));
 sg13g2_nand2_1 _18468_ (.Y(_11648_),
    .A(\cpu.ex.r_mult[2] ),
    .B(_10271_));
 sg13g2_o21ai_1 _18469_ (.B1(_11648_),
    .Y(\cpu.ex.c_mult[2] ),
    .A1(net425),
    .A2(_11647_));
 sg13g2_nand3_1 _18470_ (.B(_10981_),
    .C(_11013_),
    .A(_11618_),
    .Y(_11649_));
 sg13g2_a21oi_1 _18471_ (.A1(_11636_),
    .A2(_11649_),
    .Y(_11650_),
    .B1(_11637_));
 sg13g2_a21o_1 _18472_ (.A2(_11650_),
    .A1(net597),
    .B1(net227),
    .X(_11651_));
 sg13g2_nand3_1 _18473_ (.B(net227),
    .C(_11650_),
    .A(net597),
    .Y(_11652_));
 sg13g2_a21oi_1 _18474_ (.A1(_11651_),
    .A2(_11652_),
    .Y(_11653_),
    .B1(_10933_));
 sg13g2_buf_1 _18475_ (.A(_00120_),
    .X(_11654_));
 sg13g2_nor2_1 _18476_ (.A(_11654_),
    .B(net610),
    .Y(_11655_));
 sg13g2_mux2_1 _18477_ (.A0(_11655_),
    .A1(_11654_),
    .S(_11653_),
    .X(_11656_));
 sg13g2_nor2_1 _18478_ (.A(_11654_),
    .B(net86),
    .Y(_11657_));
 sg13g2_a221oi_1 _18479_ (.B2(net1141),
    .C1(_11657_),
    .B1(_11656_),
    .A1(net535),
    .Y(_11658_),
    .A2(_11653_));
 sg13g2_nand2_1 _18480_ (.Y(_11659_),
    .A(\cpu.ex.r_mult[3] ),
    .B(_10271_));
 sg13g2_o21ai_1 _18481_ (.B1(_11659_),
    .Y(\cpu.ex.c_mult[3] ),
    .A1(net425),
    .A2(_11658_));
 sg13g2_nor2_1 _18482_ (.A(_11654_),
    .B(_10979_),
    .Y(_11660_));
 sg13g2_nand2_1 _18483_ (.Y(_11661_),
    .A(_11654_),
    .B(_10979_));
 sg13g2_o21ai_1 _18484_ (.B1(_11661_),
    .Y(_11662_),
    .A1(_11650_),
    .A2(_11660_));
 sg13g2_buf_1 _18485_ (.A(_11662_),
    .X(_11663_));
 sg13g2_o21ai_1 _18486_ (.B1(net265),
    .Y(_11664_),
    .A1(net610),
    .A2(_11663_));
 sg13g2_nand3b_1 _18487_ (.B(net264),
    .C(net597),
    .Y(_11665_),
    .A_N(_11663_));
 sg13g2_a221oi_1 _18488_ (.B2(_11665_),
    .C1(_10931_),
    .B1(_11664_),
    .A1(_10610_),
    .Y(_11666_),
    .A2(_10744_));
 sg13g2_buf_1 _18489_ (.A(_00127_),
    .X(_11667_));
 sg13g2_nor2_1 _18490_ (.A(_11667_),
    .B(net794),
    .Y(_11668_));
 sg13g2_mux2_1 _18491_ (.A0(_11668_),
    .A1(_11667_),
    .S(_11666_),
    .X(_11669_));
 sg13g2_nor2_1 _18492_ (.A(_11667_),
    .B(net86),
    .Y(_11670_));
 sg13g2_a221oi_1 _18493_ (.B2(net1141),
    .C1(_11670_),
    .B1(_11669_),
    .A1(net535),
    .Y(_11671_),
    .A2(_11666_));
 sg13g2_nand2_1 _18494_ (.Y(_11672_),
    .A(\cpu.ex.r_mult[4] ),
    .B(_10271_));
 sg13g2_o21ai_1 _18495_ (.B1(_11672_),
    .Y(\cpu.ex.c_mult[4] ),
    .A1(net425),
    .A2(_11671_));
 sg13g2_buf_1 _18496_ (.A(_11261_),
    .X(_11673_));
 sg13g2_a21oi_1 _18497_ (.A1(net264),
    .A2(_11663_),
    .Y(_11674_),
    .B1(_11667_));
 sg13g2_nor2_1 _18498_ (.A(net264),
    .B(_11663_),
    .Y(_11675_));
 sg13g2_o21ai_1 _18499_ (.B1(net597),
    .Y(_11676_),
    .A1(_11674_),
    .A2(_11675_));
 sg13g2_xnor2_1 _18500_ (.Y(_11677_),
    .A(net206),
    .B(_11676_));
 sg13g2_nor2_1 _18501_ (.A(net77),
    .B(_11677_),
    .Y(_11678_));
 sg13g2_buf_1 _18502_ (.A(_00139_),
    .X(_11679_));
 sg13g2_nor2_1 _18503_ (.A(_11679_),
    .B(net535),
    .Y(_11680_));
 sg13g2_mux2_1 _18504_ (.A0(_11680_),
    .A1(_11679_),
    .S(_11678_),
    .X(_11681_));
 sg13g2_nor2_1 _18505_ (.A(_11679_),
    .B(net86),
    .Y(_11682_));
 sg13g2_a221oi_1 _18506_ (.B2(_09392_),
    .C1(_11682_),
    .B1(_11681_),
    .A1(net535),
    .Y(_11683_),
    .A2(_11678_));
 sg13g2_nand2_1 _18507_ (.Y(_11684_),
    .A(\cpu.ex.r_mult[5] ),
    .B(_10271_));
 sg13g2_o21ai_1 _18508_ (.B1(_11684_),
    .Y(\cpu.ex.c_mult[5] ),
    .A1(net425),
    .A2(_11683_));
 sg13g2_buf_1 _18509_ (.A(_00151_),
    .X(_11685_));
 sg13g2_inv_1 _18510_ (.Y(_11686_),
    .A(_11685_));
 sg13g2_nand2_1 _18511_ (.Y(_11687_),
    .A(_11686_),
    .B(_11620_));
 sg13g2_inv_1 _18512_ (.Y(_11688_),
    .A(_11679_));
 sg13g2_nor2_1 _18513_ (.A(net794),
    .B(net264),
    .Y(_11689_));
 sg13g2_o21ai_1 _18514_ (.B1(_11689_),
    .Y(_11690_),
    .A1(_11688_),
    .A2(net225));
 sg13g2_o21ai_1 _18515_ (.B1(_11668_),
    .Y(_11691_),
    .A1(_11688_),
    .A2(_11125_));
 sg13g2_a21o_1 _18516_ (.A2(_11691_),
    .A1(_11690_),
    .B1(_11663_),
    .X(_11692_));
 sg13g2_buf_1 _18517_ (.A(_11692_),
    .X(_11693_));
 sg13g2_nor3_1 _18518_ (.A(_11679_),
    .B(net794),
    .C(_11261_),
    .Y(_11694_));
 sg13g2_nand2_1 _18519_ (.Y(_11695_),
    .A(net265),
    .B(_11668_));
 sg13g2_a21oi_1 _18520_ (.A1(_11679_),
    .A2(_11261_),
    .Y(_11696_),
    .B1(_11695_));
 sg13g2_nor2_2 _18521_ (.A(_11694_),
    .B(_11696_),
    .Y(_11697_));
 sg13g2_nand3_1 _18522_ (.B(_11693_),
    .C(_11697_),
    .A(net222),
    .Y(_11698_));
 sg13g2_a21o_1 _18523_ (.A2(_11697_),
    .A1(_11693_),
    .B1(net222),
    .X(_11699_));
 sg13g2_a21oi_1 _18524_ (.A1(_11698_),
    .A2(_11699_),
    .Y(_11700_),
    .B1(net77));
 sg13g2_mux2_1 _18525_ (.A0(_11687_),
    .A1(_11686_),
    .S(_11700_),
    .X(_11701_));
 sg13g2_a22oi_1 _18526_ (.Y(_11702_),
    .B1(_11700_),
    .B2(net535),
    .A2(_11629_),
    .A1(_11686_));
 sg13g2_o21ai_1 _18527_ (.B1(_11702_),
    .Y(_11703_),
    .A1(_10250_),
    .A2(_11701_));
 sg13g2_a22oi_1 _18528_ (.Y(_11704_),
    .B1(_11703_),
    .B2(net483),
    .A2(_10272_),
    .A1(\cpu.ex.r_mult[6] ));
 sg13g2_inv_1 _18529_ (.Y(\cpu.ex.c_mult[6] ),
    .A(_11704_));
 sg13g2_buf_1 _18530_ (.A(net77),
    .X(_11705_));
 sg13g2_nand2b_1 _18531_ (.Y(_11706_),
    .B(net483),
    .A_N(_11585_));
 sg13g2_buf_1 _18532_ (.A(_11706_),
    .X(_11707_));
 sg13g2_nor2_1 _18533_ (.A(_11685_),
    .B(net689),
    .Y(_11708_));
 sg13g2_nand3_1 _18534_ (.B(_11693_),
    .C(_11697_),
    .A(net337),
    .Y(_11709_));
 sg13g2_a21oi_1 _18535_ (.A1(_11693_),
    .A2(_11697_),
    .Y(_11710_),
    .B1(net337));
 sg13g2_a21o_1 _18536_ (.A2(_11709_),
    .A1(_11708_),
    .B1(_11710_),
    .X(_11711_));
 sg13g2_buf_1 _18537_ (.A(_11711_),
    .X(_11712_));
 sg13g2_xnor2_1 _18538_ (.Y(_11713_),
    .A(net224),
    .B(_11712_));
 sg13g2_buf_2 _18539_ (.A(_00163_),
    .X(_11714_));
 sg13g2_nor2_2 _18540_ (.A(_11714_),
    .B(net794),
    .Y(_11715_));
 sg13g2_or4_1 _18541_ (.A(net65),
    .B(_11707_),
    .C(_11713_),
    .D(_11715_),
    .X(_11716_));
 sg13g2_nor2_1 _18542_ (.A(_11585_),
    .B(_11592_),
    .Y(_11717_));
 sg13g2_buf_2 _18543_ (.A(_11717_),
    .X(_11718_));
 sg13g2_and2_1 _18544_ (.A(_11718_),
    .B(_11715_),
    .X(_11719_));
 sg13g2_o21ai_1 _18545_ (.B1(_11719_),
    .Y(_11720_),
    .A1(net65),
    .A2(_11713_));
 sg13g2_nor2_1 _18546_ (.A(_11592_),
    .B(_11583_),
    .Y(_11721_));
 sg13g2_inv_1 _18547_ (.Y(_11722_),
    .A(_11714_));
 sg13g2_a22oi_1 _18548_ (.Y(_11723_),
    .B1(_11721_),
    .B2(_11722_),
    .A2(_10271_),
    .A1(\cpu.ex.r_mult[7] ));
 sg13g2_nand3_1 _18549_ (.B(_11720_),
    .C(_11723_),
    .A(_11716_),
    .Y(\cpu.ex.c_mult[7] ));
 sg13g2_nand2_1 _18550_ (.Y(_11724_),
    .A(net224),
    .B(_11712_));
 sg13g2_o21ai_1 _18551_ (.B1(_11715_),
    .Y(_11725_),
    .A1(net224),
    .A2(_11712_));
 sg13g2_nand2_1 _18552_ (.Y(_11726_),
    .A(_11724_),
    .B(_11725_));
 sg13g2_xnor2_1 _18553_ (.Y(_11727_),
    .A(net208),
    .B(_11726_));
 sg13g2_buf_1 _18554_ (.A(_11721_),
    .X(_11728_));
 sg13g2_nor2_1 _18555_ (.A(net65),
    .B(net64),
    .Y(_11729_));
 sg13g2_nand2_1 _18556_ (.Y(_11730_),
    .A(net1141),
    .B(net536));
 sg13g2_buf_2 _18557_ (.A(_11730_),
    .X(_11731_));
 sg13g2_nor2_1 _18558_ (.A(_11592_),
    .B(_11731_),
    .Y(_11732_));
 sg13g2_buf_2 _18559_ (.A(_11732_),
    .X(_11733_));
 sg13g2_buf_1 _18560_ (.A(_00164_),
    .X(_11734_));
 sg13g2_inv_1 _18561_ (.Y(_11735_),
    .A(_11734_));
 sg13g2_o21ai_1 _18562_ (.B1(_11735_),
    .Y(_11736_),
    .A1(net64),
    .A2(_11733_));
 sg13g2_a21oi_1 _18563_ (.A1(_11727_),
    .A2(_11729_),
    .Y(_11737_),
    .B1(_11736_));
 sg13g2_nor2_1 _18564_ (.A(_11734_),
    .B(net794),
    .Y(_11738_));
 sg13g2_nor3_1 _18565_ (.A(net65),
    .B(_11707_),
    .C(_11738_),
    .Y(_11739_));
 sg13g2_a22oi_1 _18566_ (.Y(_11740_),
    .B1(_11727_),
    .B2(_11739_),
    .A2(net340),
    .A1(\cpu.ex.r_mult[8] ));
 sg13g2_nand2b_1 _18567_ (.Y(\cpu.ex.c_mult[8] ),
    .B(_11740_),
    .A_N(_11737_));
 sg13g2_buf_1 _18568_ (.A(_00165_),
    .X(_11741_));
 sg13g2_inv_1 _18569_ (.Y(_11742_),
    .A(_11741_));
 sg13g2_nand3_1 _18570_ (.B(_11742_),
    .C(net536),
    .A(net1141),
    .Y(_11743_));
 sg13g2_buf_1 _18571_ (.A(_11340_),
    .X(_11744_));
 sg13g2_buf_1 _18572_ (.A(_11567_),
    .X(_11745_));
 sg13g2_and2_1 _18573_ (.A(_11382_),
    .B(_11738_),
    .X(_11746_));
 sg13g2_a21o_1 _18574_ (.A2(_11567_),
    .A1(_11734_),
    .B1(_11746_),
    .X(_11747_));
 sg13g2_a22oi_1 _18575_ (.Y(_11748_),
    .B1(_11747_),
    .B2(_11714_),
    .A2(net205),
    .A1(net689));
 sg13g2_or2_1 _18576_ (.X(_11749_),
    .B(_11748_),
    .A(net263));
 sg13g2_nand2_1 _18577_ (.Y(_11750_),
    .A(_11735_),
    .B(net205));
 sg13g2_nand2_1 _18578_ (.Y(_11751_),
    .A(_11734_),
    .B(net208));
 sg13g2_nand4_1 _18579_ (.B(_11715_),
    .C(_11750_),
    .A(net263),
    .Y(_11752_),
    .D(_11751_));
 sg13g2_nand2_1 _18580_ (.Y(_11753_),
    .A(_11749_),
    .B(_11752_));
 sg13g2_nor2_1 _18581_ (.A(_11714_),
    .B(_11188_),
    .Y(_11754_));
 sg13g2_nor2_1 _18582_ (.A(_11734_),
    .B(net208),
    .Y(_11755_));
 sg13g2_a21oi_1 _18583_ (.A1(_11751_),
    .A2(_11754_),
    .Y(_11756_),
    .B1(_11755_));
 sg13g2_nor2_1 _18584_ (.A(_09394_),
    .B(_11756_),
    .Y(_11757_));
 sg13g2_a21oi_1 _18585_ (.A1(_11712_),
    .A2(_11753_),
    .Y(_11758_),
    .B1(_11757_));
 sg13g2_xnor2_1 _18586_ (.Y(_11759_),
    .A(net187),
    .B(_11758_));
 sg13g2_nor2_1 _18587_ (.A(net65),
    .B(_11759_),
    .Y(_11760_));
 sg13g2_mux2_1 _18588_ (.A0(_11743_),
    .A1(net536),
    .S(_11760_),
    .X(_11761_));
 sg13g2_buf_8 _18589_ (.A(_11629_),
    .X(_11762_));
 sg13g2_nor2_1 _18590_ (.A(_10250_),
    .B(_11742_),
    .Y(_11763_));
 sg13g2_a22oi_1 _18591_ (.Y(_11764_),
    .B1(_11760_),
    .B2(_11763_),
    .A2(net63),
    .A1(_11742_));
 sg13g2_a21o_1 _18592_ (.A2(_11764_),
    .A1(_11761_),
    .B1(net425),
    .X(_11765_));
 sg13g2_nand2_1 _18593_ (.Y(_11766_),
    .A(\cpu.ex.r_mult[9] ),
    .B(net340));
 sg13g2_nand2_1 _18594_ (.Y(\cpu.ex.c_mult[9] ),
    .A(_11765_),
    .B(_11766_));
 sg13g2_buf_2 _18595_ (.A(_00166_),
    .X(_11767_));
 sg13g2_inv_1 _18596_ (.Y(_11768_),
    .A(_11767_));
 sg13g2_nor2_1 _18597_ (.A(_11767_),
    .B(net794),
    .Y(_11769_));
 sg13g2_buf_1 _18598_ (.A(_11309_),
    .X(_11770_));
 sg13g2_a221oi_1 _18599_ (.B2(_11338_),
    .C1(_11741_),
    .B1(_11315_),
    .A1(_09373_),
    .Y(_11771_),
    .A2(_11223_));
 sg13g2_nor3_1 _18600_ (.A(_11742_),
    .B(_11344_),
    .C(_11346_),
    .Y(_11772_));
 sg13g2_o21ai_1 _18601_ (.B1(_11734_),
    .Y(_11773_),
    .A1(_11771_),
    .A2(_11772_));
 sg13g2_nand2_1 _18602_ (.Y(_11774_),
    .A(net794),
    .B(_11353_));
 sg13g2_a21o_1 _18603_ (.A2(_11774_),
    .A1(_11773_),
    .B1(net208),
    .X(_11775_));
 sg13g2_nor2_1 _18604_ (.A(_11741_),
    .B(_11353_),
    .Y(_11776_));
 sg13g2_o21ai_1 _18605_ (.B1(_11746_),
    .Y(_11777_),
    .A1(_11772_),
    .A2(_11776_));
 sg13g2_mux2_1 _18606_ (.A0(_11714_),
    .A1(_11715_),
    .S(_11188_),
    .X(_11778_));
 sg13g2_nor2_1 _18607_ (.A(_11620_),
    .B(net263),
    .Y(_11779_));
 sg13g2_a21o_1 _18608_ (.A2(_11778_),
    .A1(_11685_),
    .B1(_11779_),
    .X(_11780_));
 sg13g2_and2_1 _18609_ (.A(_11714_),
    .B(net263),
    .X(_11781_));
 sg13g2_nor4_1 _18610_ (.A(_11217_),
    .B(_11687_),
    .C(_11754_),
    .D(_11781_),
    .Y(_11782_));
 sg13g2_a21oi_1 _18611_ (.A1(_11217_),
    .A2(_11780_),
    .Y(_11783_),
    .B1(_11782_));
 sg13g2_a221oi_1 _18612_ (.B2(_11777_),
    .C1(_11783_),
    .B1(_11775_),
    .A1(_11693_),
    .Y(_11784_),
    .A2(_11697_));
 sg13g2_buf_1 _18613_ (.A(_11784_),
    .X(_11785_));
 sg13g2_nand2_1 _18614_ (.Y(_11786_),
    .A(_11714_),
    .B(_11188_));
 sg13g2_nor2_1 _18615_ (.A(_11685_),
    .B(net337),
    .Y(_11787_));
 sg13g2_a21o_1 _18616_ (.A2(_11787_),
    .A1(_11786_),
    .B1(_11754_),
    .X(_11788_));
 sg13g2_buf_1 _18617_ (.A(_11788_),
    .X(_11789_));
 sg13g2_a21oi_1 _18618_ (.A1(_11741_),
    .A2(_11340_),
    .Y(_11790_),
    .B1(_11734_));
 sg13g2_nand3_1 _18619_ (.B(_11789_),
    .C(_11790_),
    .A(_11620_),
    .Y(_11791_));
 sg13g2_nand4_1 _18620_ (.B(_11620_),
    .C(_11567_),
    .A(_11742_),
    .Y(_11792_),
    .D(_11789_));
 sg13g2_nor2_1 _18621_ (.A(_11741_),
    .B(net794),
    .Y(_11793_));
 sg13g2_nor2_1 _18622_ (.A(_09393_),
    .B(_11382_),
    .Y(_11794_));
 sg13g2_a22oi_1 _18623_ (.Y(_11795_),
    .B1(_11790_),
    .B2(_11794_),
    .A2(_11793_),
    .A1(_11353_));
 sg13g2_nand4_1 _18624_ (.B(_11567_),
    .C(_11353_),
    .A(_11620_),
    .Y(_11796_),
    .D(_11789_));
 sg13g2_nand4_1 _18625_ (.B(_11792_),
    .C(_11795_),
    .A(_11791_),
    .Y(_11797_),
    .D(_11796_));
 sg13g2_buf_1 _18626_ (.A(_11797_),
    .X(_11798_));
 sg13g2_or3_1 _18627_ (.A(net132),
    .B(_11785_),
    .C(_11798_),
    .X(_11799_));
 sg13g2_o21ai_1 _18628_ (.B1(net132),
    .Y(_11800_),
    .A1(_11785_),
    .A2(_11798_));
 sg13g2_nand3_1 _18629_ (.B(_11799_),
    .C(_11800_),
    .A(net78),
    .Y(_11801_));
 sg13g2_mux2_1 _18630_ (.A0(_11767_),
    .A1(_11769_),
    .S(_11801_),
    .X(_11802_));
 sg13g2_nor2_1 _18631_ (.A(_11622_),
    .B(_11801_),
    .Y(_11803_));
 sg13g2_a221oi_1 _18632_ (.B2(net1141),
    .C1(_11803_),
    .B1(_11802_),
    .A1(_11768_),
    .Y(_11804_),
    .A2(_11762_));
 sg13g2_nand2_1 _18633_ (.Y(_11805_),
    .A(\cpu.ex.r_mult[10] ),
    .B(_10272_));
 sg13g2_o21ai_1 _18634_ (.B1(_11805_),
    .Y(\cpu.ex.c_mult[10] ),
    .A1(_11593_),
    .A2(_11804_));
 sg13g2_buf_1 _18635_ (.A(_00167_),
    .X(_11806_));
 sg13g2_nor2_1 _18636_ (.A(_11806_),
    .B(_11731_),
    .Y(_11807_));
 sg13g2_inv_1 _18637_ (.Y(_11808_),
    .A(_11806_));
 sg13g2_nor2_1 _18638_ (.A(_10250_),
    .B(_11808_),
    .Y(_11809_));
 sg13g2_nor2_1 _18639_ (.A(net77),
    .B(net207),
    .Y(_11810_));
 sg13g2_nor2_1 _18640_ (.A(net77),
    .B(net190),
    .Y(_11811_));
 sg13g2_xnor2_1 _18641_ (.Y(_11812_),
    .A(_11767_),
    .B(_11309_));
 sg13g2_mux2_1 _18642_ (.A0(_11767_),
    .A1(_11769_),
    .S(net169),
    .X(_11813_));
 sg13g2_nor2_1 _18643_ (.A(net169),
    .B(_11774_),
    .Y(_11814_));
 sg13g2_a221oi_1 _18644_ (.B2(_11772_),
    .C1(_11814_),
    .B1(_11813_),
    .A1(_11771_),
    .Y(_11815_),
    .A2(_11812_));
 sg13g2_a21oi_1 _18645_ (.A1(_11749_),
    .A2(_11752_),
    .Y(_11816_),
    .B1(_11815_));
 sg13g2_o21ai_1 _18646_ (.B1(_11340_),
    .Y(_11817_),
    .A1(_09394_),
    .A2(_11756_));
 sg13g2_a21oi_1 _18647_ (.A1(_11767_),
    .A2(net169),
    .Y(_11818_),
    .B1(_11741_));
 sg13g2_nand2_1 _18648_ (.Y(_11819_),
    .A(_11621_),
    .B(net189));
 sg13g2_o21ai_1 _18649_ (.B1(net169),
    .Y(_11820_),
    .A1(_11756_),
    .A2(_11819_));
 sg13g2_a22oi_1 _18650_ (.Y(_11821_),
    .B1(_11820_),
    .B2(_11768_),
    .A2(_11818_),
    .A1(_11817_));
 sg13g2_nand3_1 _18651_ (.B(net189),
    .C(_11757_),
    .A(net132),
    .Y(_11822_));
 sg13g2_o21ai_1 _18652_ (.B1(_11822_),
    .Y(_11823_),
    .A1(net610),
    .A2(_11821_));
 sg13g2_a21o_1 _18653_ (.A2(_11816_),
    .A1(_11712_),
    .B1(_11823_),
    .X(_11824_));
 sg13g2_buf_1 _18654_ (.A(_11824_),
    .X(_11825_));
 sg13g2_mux2_1 _18655_ (.A0(_11810_),
    .A1(_11811_),
    .S(_11825_),
    .X(_11826_));
 sg13g2_mux2_1 _18656_ (.A0(_11807_),
    .A1(_11809_),
    .S(_11826_),
    .X(_11827_));
 sg13g2_nor2_1 _18657_ (.A(_11620_),
    .B(_11506_),
    .Y(_11828_));
 sg13g2_a22oi_1 _18658_ (.Y(_11829_),
    .B1(_11828_),
    .B2(_11588_),
    .A2(_11629_),
    .A1(_11808_));
 sg13g2_nor2_1 _18659_ (.A(_11593_),
    .B(_11829_),
    .Y(_11830_));
 sg13g2_a221oi_1 _18660_ (.B2(_10269_),
    .C1(_11830_),
    .B1(_11827_),
    .A1(\cpu.ex.r_mult[11] ),
    .Y(_11831_),
    .A2(net340));
 sg13g2_inv_1 _18661_ (.Y(\cpu.ex.c_mult[11] ),
    .A(_11831_));
 sg13g2_buf_8 _18662_ (.A(_11455_),
    .X(_11832_));
 sg13g2_nand3_1 _18663_ (.B(_11280_),
    .C(_11307_),
    .A(_11768_),
    .Y(_11833_));
 sg13g2_nand2_1 _18664_ (.Y(_11834_),
    .A(_11808_),
    .B(_11490_));
 sg13g2_nor2_1 _18665_ (.A(_11808_),
    .B(_11490_),
    .Y(_11835_));
 sg13g2_a21o_1 _18666_ (.A2(_11834_),
    .A1(_11833_),
    .B1(_11835_),
    .X(_11836_));
 sg13g2_buf_2 _18667_ (.A(_11836_),
    .X(_11837_));
 sg13g2_buf_1 _18668_ (.A(_00168_),
    .X(_11838_));
 sg13g2_nor2_1 _18669_ (.A(net1125),
    .B(net689),
    .Y(_11839_));
 sg13g2_and3_1 _18670_ (.X(_11840_),
    .A(net167),
    .B(_11837_),
    .C(_11839_));
 sg13g2_and4_1 _18671_ (.A(net1125),
    .B(net78),
    .C(net191),
    .D(_11837_),
    .X(_11841_));
 sg13g2_nand2_1 _18672_ (.Y(_11842_),
    .A(_11808_),
    .B(_11620_));
 sg13g2_a21o_1 _18673_ (.A2(_11488_),
    .A1(_11485_),
    .B1(_11842_),
    .X(_11843_));
 sg13g2_nand3_1 _18674_ (.B(_11485_),
    .C(_11488_),
    .A(_11806_),
    .Y(_11844_));
 sg13g2_a21oi_1 _18675_ (.A1(_11843_),
    .A2(_11844_),
    .Y(_11845_),
    .B1(_11768_));
 sg13g2_o21ai_1 _18676_ (.B1(_11309_),
    .Y(_11846_),
    .A1(_11828_),
    .A2(_11845_));
 sg13g2_nand2_1 _18677_ (.Y(_11847_),
    .A(_11806_),
    .B(_11506_));
 sg13g2_nand4_1 _18678_ (.B(_11769_),
    .C(_11834_),
    .A(_11355_),
    .Y(_11848_),
    .D(_11847_));
 sg13g2_a221oi_1 _18679_ (.B2(_11848_),
    .C1(_10931_),
    .B1(_11846_),
    .A1(_10610_),
    .Y(_11849_),
    .A2(_10744_));
 sg13g2_o21ai_1 _18680_ (.B1(_11849_),
    .Y(_11850_),
    .A1(_11785_),
    .A2(_11798_));
 sg13g2_buf_1 _18681_ (.A(_11850_),
    .X(_11851_));
 sg13g2_o21ai_1 _18682_ (.B1(_11851_),
    .Y(_11852_),
    .A1(_11840_),
    .A2(_11841_));
 sg13g2_nor2_1 _18683_ (.A(net597),
    .B(net167),
    .Y(_11853_));
 sg13g2_nand2_1 _18684_ (.Y(_11854_),
    .A(net78),
    .B(_11853_));
 sg13g2_nand2_1 _18685_ (.Y(_11855_),
    .A(net65),
    .B(_11839_));
 sg13g2_nand2_1 _18686_ (.Y(_11856_),
    .A(net1125),
    .B(net167));
 sg13g2_nor2_1 _18687_ (.A(_11851_),
    .B(_11856_),
    .Y(_11857_));
 sg13g2_nor4_1 _18688_ (.A(net1125),
    .B(net610),
    .C(net167),
    .D(_11851_),
    .Y(_11858_));
 sg13g2_nand3_1 _18689_ (.B(net536),
    .C(net167),
    .A(net1125),
    .Y(_11859_));
 sg13g2_nor3_1 _18690_ (.A(_11624_),
    .B(_11837_),
    .C(_11859_),
    .Y(_11860_));
 sg13g2_nor4_1 _18691_ (.A(net1125),
    .B(net535),
    .C(net167),
    .D(_11837_),
    .Y(_11861_));
 sg13g2_nor4_1 _18692_ (.A(_11857_),
    .B(_11858_),
    .C(_11860_),
    .D(_11861_),
    .Y(_11862_));
 sg13g2_and4_1 _18693_ (.A(_11852_),
    .B(_11854_),
    .C(_11855_),
    .D(_11862_),
    .X(_11863_));
 sg13g2_inv_1 _18694_ (.Y(_11864_),
    .A(_11838_));
 sg13g2_a22oi_1 _18695_ (.Y(_11865_),
    .B1(_11728_),
    .B2(_11864_),
    .A2(net340),
    .A1(\cpu.ex.r_mult[12] ));
 sg13g2_o21ai_1 _18696_ (.B1(_11865_),
    .Y(\cpu.ex.c_mult[12] ),
    .A1(_11707_),
    .A2(_11863_));
 sg13g2_mux2_1 _18697_ (.A0(net1125),
    .A1(_11839_),
    .S(_11455_),
    .X(_11866_));
 sg13g2_a21o_1 _18698_ (.A2(_11866_),
    .A1(_11806_),
    .B1(_11853_),
    .X(_11867_));
 sg13g2_nor2_1 _18699_ (.A(net190),
    .B(_11842_),
    .Y(_11868_));
 sg13g2_nand2_1 _18700_ (.Y(_11869_),
    .A(_11864_),
    .B(net191));
 sg13g2_and3_1 _18701_ (.X(_11870_),
    .A(_11868_),
    .B(_11856_),
    .C(_11869_));
 sg13g2_a21o_1 _18702_ (.A2(_11867_),
    .A1(net190),
    .B1(_11870_),
    .X(_11871_));
 sg13g2_a21o_1 _18703_ (.A2(net167),
    .A1(net1125),
    .B1(_11834_),
    .X(_11872_));
 sg13g2_a21oi_1 _18704_ (.A1(_11869_),
    .A2(_11872_),
    .Y(_11873_),
    .B1(_10247_));
 sg13g2_a21oi_1 _18705_ (.A1(_11825_),
    .A2(_11871_),
    .Y(_11874_),
    .B1(_11873_));
 sg13g2_nor2_1 _18706_ (.A(net65),
    .B(_11874_),
    .Y(_11875_));
 sg13g2_buf_2 _18707_ (.A(_00169_),
    .X(_11876_));
 sg13g2_nor2_2 _18708_ (.A(_11876_),
    .B(net689),
    .Y(_11877_));
 sg13g2_nand2_1 _18709_ (.Y(_11878_),
    .A(net78),
    .B(net133));
 sg13g2_xor2_1 _18710_ (.B(_11878_),
    .A(_11877_),
    .X(_11879_));
 sg13g2_xnor2_1 _18711_ (.Y(_11880_),
    .A(_11875_),
    .B(_11879_));
 sg13g2_nand2_1 _18712_ (.Y(_11881_),
    .A(_11718_),
    .B(_11880_));
 sg13g2_nand2_2 _18713_ (.Y(_11882_),
    .A(net483),
    .B(_11762_));
 sg13g2_nor2_1 _18714_ (.A(_11876_),
    .B(_11882_),
    .Y(_11883_));
 sg13g2_and2_1 _18715_ (.A(\cpu.ex.r_mult[13] ),
    .B(net340),
    .X(_11884_));
 sg13g2_nor2_1 _18716_ (.A(_11883_),
    .B(_11884_),
    .Y(_11885_));
 sg13g2_nand2_1 _18717_ (.Y(\cpu.ex.c_mult[13] ),
    .A(_11881_),
    .B(_11885_));
 sg13g2_nand2_1 _18718_ (.Y(_11886_),
    .A(_11423_),
    .B(_11449_));
 sg13g2_buf_2 _18719_ (.A(_11886_),
    .X(_11887_));
 sg13g2_mux2_1 _18720_ (.A0(_11876_),
    .A1(_11877_),
    .S(_11887_),
    .X(_11888_));
 sg13g2_a22oi_1 _18721_ (.Y(_11889_),
    .B1(_11888_),
    .B2(_11838_),
    .A2(_11453_),
    .A1(net689));
 sg13g2_xnor2_1 _18722_ (.Y(_11890_),
    .A(_11876_),
    .B(_11453_));
 sg13g2_nand3_1 _18723_ (.B(_11839_),
    .C(_11890_),
    .A(_11455_),
    .Y(_11891_));
 sg13g2_o21ai_1 _18724_ (.B1(_11891_),
    .Y(_11892_),
    .A1(net167),
    .A2(_11889_));
 sg13g2_nand2b_1 _18725_ (.Y(_11893_),
    .B(_11892_),
    .A_N(_11851_));
 sg13g2_a21oi_1 _18726_ (.A1(_11455_),
    .A2(_11837_),
    .Y(_11894_),
    .B1(_00168_));
 sg13g2_nor2_1 _18727_ (.A(_11455_),
    .B(_11837_),
    .Y(_11895_));
 sg13g2_nand2_1 _18728_ (.Y(_11896_),
    .A(_11876_),
    .B(_11887_));
 sg13g2_o21ai_1 _18729_ (.B1(_11896_),
    .Y(_11897_),
    .A1(_11894_),
    .A2(_11895_));
 sg13g2_nand2b_1 _18730_ (.Y(_11898_),
    .B(_11453_),
    .A_N(_11876_));
 sg13g2_nand2_1 _18731_ (.Y(_11899_),
    .A(net597),
    .B(_11587_));
 sg13g2_a21o_1 _18732_ (.A2(_11898_),
    .A1(_11897_),
    .B1(_11899_),
    .X(_11900_));
 sg13g2_buf_1 _18733_ (.A(_11900_),
    .X(_11901_));
 sg13g2_nor2_1 _18734_ (.A(_10841_),
    .B(_10880_),
    .Y(_11902_));
 sg13g2_nor2_1 _18735_ (.A(_10797_),
    .B(_10930_),
    .Y(_11903_));
 sg13g2_a221oi_1 _18736_ (.B2(_11903_),
    .C1(_11546_),
    .B1(_11902_),
    .A1(_10610_),
    .Y(_11904_),
    .A2(_10744_));
 sg13g2_inv_1 _18737_ (.Y(_11905_),
    .A(_00170_));
 sg13g2_nand2_1 _18738_ (.Y(_11906_),
    .A(_11905_),
    .B(net597));
 sg13g2_xnor2_1 _18739_ (.Y(_11907_),
    .A(_11904_),
    .B(_11906_));
 sg13g2_nand4_1 _18740_ (.B(_11893_),
    .C(_11901_),
    .A(_11718_),
    .Y(_11908_),
    .D(_11907_));
 sg13g2_or2_1 _18741_ (.X(_11909_),
    .B(_11907_),
    .A(_11707_));
 sg13g2_a21o_1 _18742_ (.A2(_11901_),
    .A1(_11893_),
    .B1(_11909_),
    .X(_11910_));
 sg13g2_a22oi_1 _18743_ (.Y(_11911_),
    .B1(_11721_),
    .B2(_11905_),
    .A2(_10271_),
    .A1(\cpu.ex.r_mult[14] ));
 sg13g2_nand3_1 _18744_ (.B(_11910_),
    .C(_11911_),
    .A(_11908_),
    .Y(\cpu.ex.c_mult[14] ));
 sg13g2_a221oi_1 _18745_ (.B2(_11903_),
    .C1(_10367_),
    .B1(_11902_),
    .A1(_10610_),
    .Y(_11912_),
    .A2(_10744_));
 sg13g2_buf_1 _18746_ (.A(_00171_),
    .X(_11913_));
 sg13g2_nor2_1 _18747_ (.A(_11913_),
    .B(net610),
    .Y(_11914_));
 sg13g2_xnor2_1 _18748_ (.Y(_11915_),
    .A(_11912_),
    .B(_11914_));
 sg13g2_nor2_1 _18749_ (.A(_11547_),
    .B(_11906_),
    .Y(_11916_));
 sg13g2_nor3_1 _18750_ (.A(_11707_),
    .B(_11915_),
    .C(_11916_),
    .Y(_11917_));
 sg13g2_and3_1 _18751_ (.X(_11918_),
    .A(net78),
    .B(_11718_),
    .C(_11915_));
 sg13g2_a21oi_1 _18752_ (.A1(net190),
    .A2(_11867_),
    .Y(_11919_),
    .B1(_11870_));
 sg13g2_nor4_1 _18753_ (.A(_11876_),
    .B(_11630_),
    .C(_11624_),
    .D(_11919_),
    .Y(_11920_));
 sg13g2_nor2_1 _18754_ (.A(_11919_),
    .B(_11878_),
    .Y(_11921_));
 sg13g2_o21ai_1 _18755_ (.B1(_11825_),
    .Y(_11922_),
    .A1(_11920_),
    .A2(_11921_));
 sg13g2_nand2_1 _18756_ (.Y(_11923_),
    .A(_11877_),
    .B(_11873_));
 sg13g2_nand2_1 _18757_ (.Y(_11924_),
    .A(net133),
    .B(_11873_));
 sg13g2_a21oi_1 _18758_ (.A1(_11923_),
    .A2(_11924_),
    .Y(_11925_),
    .B1(_11705_));
 sg13g2_a21oi_1 _18759_ (.A1(net133),
    .A2(_11877_),
    .Y(_11926_),
    .B1(_11925_));
 sg13g2_a22oi_1 _18760_ (.Y(_11927_),
    .B1(_11922_),
    .B2(_11926_),
    .A2(_11906_),
    .A1(_11547_));
 sg13g2_mux2_1 _18761_ (.A0(_11917_),
    .A1(_11918_),
    .S(_11927_),
    .X(_11928_));
 sg13g2_buf_1 _18762_ (.A(\cpu.ex.r_mult[15] ),
    .X(_11929_));
 sg13g2_inv_1 _18763_ (.Y(_11930_),
    .A(_11913_));
 sg13g2_a22oi_1 _18764_ (.Y(_11931_),
    .B1(_11728_),
    .B2(_11930_),
    .A2(net340),
    .A1(_11929_));
 sg13g2_nand3_1 _18765_ (.B(_11718_),
    .C(_11914_),
    .A(_11705_),
    .Y(_11932_));
 sg13g2_nand4_1 _18766_ (.B(_11718_),
    .C(_11915_),
    .A(_11588_),
    .Y(_11933_),
    .D(_11916_));
 sg13g2_nand3_1 _18767_ (.B(_11932_),
    .C(_11933_),
    .A(_11931_),
    .Y(_11934_));
 sg13g2_or2_1 _18768_ (.X(\cpu.ex.c_mult[15] ),
    .B(_11934_),
    .A(_11928_));
 sg13g2_inv_1 _18769_ (.Y(_00000_),
    .A(net2));
 sg13g2_buf_1 _18770_ (.A(\cpu.qspi.r_state[11] ),
    .X(_11935_));
 sg13g2_buf_1 _18771_ (.A(net916),
    .X(_11936_));
 sg13g2_and2_1 _18772_ (.A(_11935_),
    .B(net750),
    .X(_00004_));
 sg13g2_nor3_1 _18773_ (.A(net691),
    .B(_09881_),
    .C(_09882_),
    .Y(_00007_));
 sg13g2_buf_2 _18774_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11937_));
 sg13g2_and2_1 _18775_ (.A(_11937_),
    .B(net750),
    .X(_00003_));
 sg13g2_buf_2 _18776_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11938_));
 sg13g2_and2_1 _18777_ (.A(_11938_),
    .B(net750),
    .X(_00002_));
 sg13g2_inv_1 _18778_ (.Y(_11939_),
    .A(_09851_));
 sg13g2_nor3_1 _18779_ (.A(_11939_),
    .B(net682),
    .C(_09853_),
    .Y(_00001_));
 sg13g2_nand2_1 _18780_ (.Y(_11940_),
    .A(\cpu.dec.iready ),
    .B(_00199_));
 sg13g2_nor2_2 _18781_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11940_),
    .Y(_11941_));
 sg13g2_nand2_1 _18782_ (.Y(_11942_),
    .A(net1066),
    .B(_11941_));
 sg13g2_buf_2 _18783_ (.A(_11942_),
    .X(_11943_));
 sg13g2_inv_1 _18784_ (.Y(_11944_),
    .A(_00275_));
 sg13g2_buf_1 _18785_ (.A(_08402_),
    .X(_11945_));
 sg13g2_buf_1 _18786_ (.A(_08428_),
    .X(_11946_));
 sg13g2_nand2_1 _18787_ (.Y(_11947_),
    .A(_10481_),
    .B(_10857_));
 sg13g2_o21ai_1 _18788_ (.B1(_11947_),
    .Y(_11948_),
    .A1(net749),
    .A2(net539));
 sg13g2_nand2_1 _18789_ (.Y(_11949_),
    .A(_10770_),
    .B(_10793_));
 sg13g2_or2_1 _18790_ (.X(_11950_),
    .B(_10817_),
    .A(_10800_));
 sg13g2_buf_1 _18791_ (.A(_11950_),
    .X(_11951_));
 sg13g2_nand2b_1 _18792_ (.Y(_11952_),
    .B(net539),
    .A_N(_10877_));
 sg13g2_o21ai_1 _18793_ (.B1(_11952_),
    .Y(_11953_),
    .A1(net598),
    .A2(net539));
 sg13g2_nand3_1 _18794_ (.B(_11951_),
    .C(_11953_),
    .A(_11949_),
    .Y(_11954_));
 sg13g2_nor2b_1 _18795_ (.A(_10835_),
    .B_N(_10905_),
    .Y(_11955_));
 sg13g2_nand3b_1 _18796_ (.B(_10740_),
    .C(_11955_),
    .Y(_11956_),
    .A_N(_10592_));
 sg13g2_nor2_1 _18797_ (.A(_10669_),
    .B(_10705_),
    .Y(_11957_));
 sg13g2_nor3_1 _18798_ (.A(_10640_),
    .B(_10471_),
    .C(_10523_),
    .Y(_11958_));
 sg13g2_nand4_1 _18799_ (.B(_10927_),
    .C(_11957_),
    .A(_10563_),
    .Y(_11959_),
    .D(_11958_));
 sg13g2_nor4_1 _18800_ (.A(_11948_),
    .B(_11954_),
    .C(_11956_),
    .D(_11959_),
    .Y(_11960_));
 sg13g2_o21ai_1 _18801_ (.B1(_10768_),
    .Y(_11961_),
    .A1(\cpu.cond[1] ),
    .A2(_11960_));
 sg13g2_xnor2_1 _18802_ (.Y(_11962_),
    .A(_11945_),
    .B(_11961_));
 sg13g2_o21ai_1 _18803_ (.B1(net1039),
    .Y(_11963_),
    .A1(_11944_),
    .A2(_11962_));
 sg13g2_nor2b_1 _18804_ (.A(\cpu.dec.jmp ),
    .B_N(_11963_),
    .Y(_11964_));
 sg13g2_nor2_1 _18805_ (.A(_11943_),
    .B(_11964_),
    .Y(_00053_));
 sg13g2_and3_1 _18806_ (.X(_00005_),
    .A(net1137),
    .B(net797),
    .C(_09846_));
 sg13g2_buf_2 _18807_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11965_));
 sg13g2_and2_1 _18808_ (.A(_11965_),
    .B(net750),
    .X(_00006_));
 sg13g2_inv_1 _18809_ (.Y(_11966_),
    .A(_09856_));
 sg13g2_nor3_1 _18810_ (.A(_11966_),
    .B(_09889_),
    .C(net172),
    .Y(_00008_));
 sg13g2_buf_2 _18811_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11967_));
 sg13g2_and2_1 _18812_ (.A(_11967_),
    .B(_11936_),
    .X(_00009_));
 sg13g2_buf_2 _18813_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11968_));
 sg13g2_and2_1 _18814_ (.A(_11968_),
    .B(_11936_),
    .X(_00010_));
 sg13g2_and2_1 _18815_ (.A(net108),
    .B(net797),
    .X(_00052_));
 sg13g2_o21ai_1 _18816_ (.B1(_09216_),
    .Y(_11969_),
    .A1(net1064),
    .A2(net1143));
 sg13g2_or4_1 _18817_ (.A(net1144),
    .B(_09317_),
    .C(net1143),
    .D(_09357_),
    .X(_11970_));
 sg13g2_nand3_1 _18818_ (.B(_11969_),
    .C(_11970_),
    .A(_09305_),
    .Y(_11971_));
 sg13g2_buf_1 _18819_ (.A(_11971_),
    .X(_11972_));
 sg13g2_buf_1 _18820_ (.A(_00228_),
    .X(_11973_));
 sg13g2_nor2_1 _18821_ (.A(net1143),
    .B(_09357_),
    .Y(_11974_));
 sg13g2_buf_1 _18822_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11975_));
 sg13g2_inv_2 _18823_ (.Y(_11976_),
    .A(_11975_));
 sg13g2_buf_2 _18824_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11977_));
 sg13g2_buf_1 _18825_ (.A(_11977_),
    .X(_11978_));
 sg13g2_buf_1 _18826_ (.A(_11978_),
    .X(_11979_));
 sg13g2_buf_1 _18827_ (.A(_11977_),
    .X(_11980_));
 sg13g2_buf_1 _18828_ (.A(_00284_),
    .X(_11981_));
 sg13g2_nor2b_1 _18829_ (.A(_11980_),
    .B_N(_11981_),
    .Y(_11982_));
 sg13g2_a21oi_1 _18830_ (.A1(net874),
    .A2(_00285_),
    .Y(_11983_),
    .B1(_11982_));
 sg13g2_nand2b_1 _18831_ (.Y(_11984_),
    .B(_11980_),
    .A_N(_11981_));
 sg13g2_buf_1 _18832_ (.A(\cpu.spi.r_src[2] ),
    .X(_11985_));
 sg13g2_nand2b_1 _18833_ (.Y(_11986_),
    .B(_11985_),
    .A_N(net1028));
 sg13g2_a21oi_1 _18834_ (.A1(_11984_),
    .A2(_11986_),
    .Y(_11987_),
    .B1(_11976_));
 sg13g2_a21oi_2 _18835_ (.B1(_11987_),
    .Y(_11988_),
    .A2(_11983_),
    .A1(_11976_));
 sg13g2_a21oi_1 _18836_ (.A1(_11973_),
    .A2(_11974_),
    .Y(_11989_),
    .B1(_11988_));
 sg13g2_nor2_1 _18837_ (.A(net1064),
    .B(_09357_),
    .Y(_11990_));
 sg13g2_buf_1 _18838_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11991_));
 sg13g2_buf_1 _18839_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11992_));
 sg13g2_buf_1 _18840_ (.A(net1029),
    .X(_11993_));
 sg13g2_mux2_1 _18841_ (.A0(_11991_),
    .A1(_11992_),
    .S(_11993_),
    .X(_11994_));
 sg13g2_nor2_1 _18842_ (.A(_11976_),
    .B(_11977_),
    .Y(_11995_));
 sg13g2_buf_1 _18843_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11996_));
 sg13g2_a22oi_1 _18844_ (.Y(_11997_),
    .B1(_11995_),
    .B2(_11996_),
    .A2(_11994_),
    .A1(_11976_));
 sg13g2_xnor2_1 _18845_ (.Y(_11998_),
    .A(_11990_),
    .B(_11997_));
 sg13g2_nand2_1 _18846_ (.Y(_11999_),
    .A(_11973_),
    .B(_11974_));
 sg13g2_buf_1 _18847_ (.A(_10561_),
    .X(_12000_));
 sg13g2_buf_1 _18848_ (.A(_09524_),
    .X(_12001_));
 sg13g2_and2_1 _18849_ (.A(net748),
    .B(_00285_),
    .X(_12002_));
 sg13g2_a21oi_1 _18850_ (.A1(net774),
    .A2(_11981_),
    .Y(_12003_),
    .B1(_12002_));
 sg13g2_buf_1 _18851_ (.A(net748),
    .X(_12004_));
 sg13g2_nor2_1 _18852_ (.A(net872),
    .B(net663),
    .Y(_12005_));
 sg13g2_a22oi_1 _18853_ (.Y(_12006_),
    .B1(_12005_),
    .B2(_11985_),
    .A2(_12003_),
    .A1(net872));
 sg13g2_nor2_1 _18854_ (.A(_11999_),
    .B(_12006_),
    .Y(_12007_));
 sg13g2_buf_1 _18855_ (.A(net1058),
    .X(_12008_));
 sg13g2_buf_1 _18856_ (.A(net871),
    .X(_12009_));
 sg13g2_buf_2 _18857_ (.A(net747),
    .X(_12010_));
 sg13g2_buf_1 _18858_ (.A(net663),
    .X(_12011_));
 sg13g2_nand2b_1 _18859_ (.Y(_12012_),
    .B(net596),
    .A_N(_11991_));
 sg13g2_o21ai_1 _18860_ (.B1(_12012_),
    .Y(_12013_),
    .A1(net596),
    .A2(_11996_));
 sg13g2_buf_1 _18861_ (.A(net747),
    .X(_12014_));
 sg13g2_buf_1 _18862_ (.A(net748),
    .X(_12015_));
 sg13g2_mux2_1 _18863_ (.A0(_11991_),
    .A1(_11992_),
    .S(_12015_),
    .X(_12016_));
 sg13g2_nor2_1 _18864_ (.A(_12014_),
    .B(_12016_),
    .Y(_12017_));
 sg13g2_a21oi_1 _18865_ (.A1(net662),
    .A2(_12013_),
    .Y(_12018_),
    .B1(_12017_));
 sg13g2_a22oi_1 _18866_ (.Y(_12019_),
    .B1(_12007_),
    .B2(_12018_),
    .A2(_11998_),
    .A1(_11989_));
 sg13g2_nor2_1 _18867_ (.A(_11989_),
    .B(_12007_),
    .Y(_12020_));
 sg13g2_buf_1 _18868_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_12021_));
 sg13g2_o21ai_1 _18869_ (.B1(_12021_),
    .Y(_12022_),
    .A1(_11972_),
    .A2(_12020_));
 sg13g2_o21ai_1 _18870_ (.B1(_12022_),
    .Y(_00320_),
    .A1(_11972_),
    .A2(_12019_));
 sg13g2_nor2b_1 _18871_ (.A(_11972_),
    .B_N(_12020_),
    .Y(_12023_));
 sg13g2_buf_1 _18872_ (.A(_11999_),
    .X(_12024_));
 sg13g2_nor2b_1 _18873_ (.A(net746),
    .B_N(_12018_),
    .Y(_12025_));
 sg13g2_a21oi_1 _18874_ (.A1(net746),
    .A2(_11998_),
    .Y(_12026_),
    .B1(_12025_));
 sg13g2_buf_1 _18875_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_12027_));
 sg13g2_nor2_1 _18876_ (.A(_12027_),
    .B(_12023_),
    .Y(_12028_));
 sg13g2_a21oi_1 _18877_ (.A1(_12023_),
    .A2(_12026_),
    .Y(_00321_),
    .B1(_12028_));
 sg13g2_buf_1 _18878_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_12029_));
 sg13g2_buf_1 _18879_ (.A(net1065),
    .X(_12030_));
 sg13g2_mux2_1 _18880_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_10131_),
    .S(_12030_),
    .X(_12031_));
 sg13g2_nor2_1 _18881_ (.A(net917),
    .B(_09297_),
    .Y(_12032_));
 sg13g2_inv_1 _18882_ (.Y(_12033_),
    .A(_00226_));
 sg13g2_mux2_1 _18883_ (.A0(_12033_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_11977_),
    .X(_12034_));
 sg13g2_a22oi_1 _18884_ (.Y(_12035_),
    .B1(_12034_),
    .B2(_11976_),
    .A2(_11995_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18885_ (.A(_12035_),
    .X(_12036_));
 sg13g2_nand2_1 _18886_ (.Y(_12037_),
    .A(_09320_),
    .B(_12036_));
 sg13g2_a21o_1 _18887_ (.A2(_09324_),
    .A1(_00223_),
    .B1(net1143),
    .X(_12038_));
 sg13g2_o21ai_1 _18888_ (.B1(net1143),
    .Y(_12039_),
    .A1(_09216_),
    .A2(_12036_));
 sg13g2_nand2b_1 _18889_ (.Y(_12040_),
    .B(_12039_),
    .A_N(_09317_));
 sg13g2_o21ai_1 _18890_ (.B1(_12040_),
    .Y(_12041_),
    .A1(_12037_),
    .A2(_12038_));
 sg13g2_nand2_1 _18891_ (.Y(_12042_),
    .A(_12032_),
    .B(_12041_));
 sg13g2_nand2b_1 _18892_ (.Y(_12043_),
    .B(_11974_),
    .A_N(_09317_));
 sg13g2_buf_1 _18893_ (.A(_12036_),
    .X(_12044_));
 sg13g2_nand3b_1 _18894_ (.B(_09358_),
    .C(_09289_),
    .Y(_12045_),
    .A_N(net595));
 sg13g2_o21ai_1 _18895_ (.B1(_12045_),
    .Y(_12046_),
    .A1(net1145),
    .A2(_12043_));
 sg13g2_nor3_1 _18896_ (.A(_11988_),
    .B(_12042_),
    .C(_12046_),
    .Y(_12047_));
 sg13g2_mux2_1 _18897_ (.A0(_12029_),
    .A1(_12031_),
    .S(_12047_),
    .X(_00322_));
 sg13g2_buf_1 _18898_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_12048_));
 sg13g2_nor2_1 _18899_ (.A(_12042_),
    .B(_12046_),
    .Y(_12049_));
 sg13g2_nand2_1 _18900_ (.Y(_12050_),
    .A(_11988_),
    .B(_12049_));
 sg13g2_mux2_1 _18901_ (.A0(_12031_),
    .A1(_12048_),
    .S(_12050_),
    .X(_00323_));
 sg13g2_buf_1 _18902_ (.A(uio_in[0]),
    .X(_12051_));
 sg13g2_buf_2 _18903_ (.A(_12051_),
    .X(_12052_));
 sg13g2_nand2_1 _18904_ (.Y(_12053_),
    .A(net1061),
    .B(_09521_));
 sg13g2_buf_1 _18905_ (.A(_12053_),
    .X(_12054_));
 sg13g2_buf_1 _18906_ (.A(\cpu.d_wstrobe_d ),
    .X(_12055_));
 sg13g2_buf_1 _18907_ (.A(_00278_),
    .X(_12056_));
 sg13g2_buf_1 _18908_ (.A(_12056_),
    .X(_12057_));
 sg13g2_nand2_2 _18909_ (.Y(_12058_),
    .A(_12055_),
    .B(net1027));
 sg13g2_buf_2 _18910_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_12059_));
 sg13g2_inv_1 _18911_ (.Y(_12060_),
    .A(_12059_));
 sg13g2_buf_1 _18912_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12061_));
 sg13g2_buf_1 _18913_ (.A(_12061_),
    .X(_12062_));
 sg13g2_nand2_1 _18914_ (.Y(_12063_),
    .A(_12060_),
    .B(net1026));
 sg13g2_or2_1 _18915_ (.X(_12064_),
    .B(_12063_),
    .A(_12058_));
 sg13g2_buf_2 _18916_ (.A(_12064_),
    .X(_12065_));
 sg13g2_or2_1 _18917_ (.X(_12066_),
    .B(_12065_),
    .A(net659));
 sg13g2_buf_1 _18918_ (.A(_12066_),
    .X(_12067_));
 sg13g2_mux2_1 _18919_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][0] ),
    .S(_12067_),
    .X(_12068_));
 sg13g2_buf_1 _18920_ (.A(net1057),
    .X(_12069_));
 sg13g2_nand2_2 _18921_ (.Y(_12070_),
    .A(_12059_),
    .B(_12061_));
 sg13g2_buf_1 _18922_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_12071_));
 sg13g2_nand2_1 _18923_ (.Y(_12072_),
    .A(_12071_),
    .B(_12055_));
 sg13g2_buf_2 _18924_ (.A(_12072_),
    .X(_12073_));
 sg13g2_nor2_2 _18925_ (.A(_12070_),
    .B(_12073_),
    .Y(_12074_));
 sg13g2_and3_1 _18926_ (.X(_12075_),
    .A(_09399_),
    .B(_08355_),
    .C(_09286_));
 sg13g2_o21ai_1 _18927_ (.B1(_12075_),
    .Y(_12076_),
    .A1(_09831_),
    .A2(_12074_));
 sg13g2_buf_1 _18928_ (.A(_12076_),
    .X(_12077_));
 sg13g2_or2_1 _18929_ (.X(_12078_),
    .B(_12077_),
    .A(_12053_));
 sg13g2_buf_1 _18930_ (.A(_12078_),
    .X(_12079_));
 sg13g2_buf_1 _18931_ (.A(_08350_),
    .X(_12080_));
 sg13g2_nand2b_1 _18932_ (.Y(_12081_),
    .B(_08351_),
    .A_N(net1025));
 sg13g2_buf_1 _18933_ (.A(_00277_),
    .X(_12082_));
 sg13g2_o21ai_1 _18934_ (.B1(net1119),
    .Y(_12083_),
    .A1(net1154),
    .A2(_12081_));
 sg13g2_nor2_1 _18935_ (.A(_12079_),
    .B(_12083_),
    .Y(_12084_));
 sg13g2_buf_4 _18936_ (.X(_12085_),
    .A(_12084_));
 sg13g2_mux2_1 _18937_ (.A0(_12068_),
    .A1(_12069_),
    .S(_12085_),
    .X(_00324_));
 sg13g2_buf_1 _18938_ (.A(uio_in[2]),
    .X(_12086_));
 sg13g2_buf_2 _18939_ (.A(_12086_),
    .X(_12087_));
 sg13g2_or2_1 _18940_ (.X(_12088_),
    .B(_12058_),
    .A(_12070_));
 sg13g2_buf_2 _18941_ (.A(_12088_),
    .X(_12089_));
 sg13g2_or2_1 _18942_ (.X(_12090_),
    .B(_12089_),
    .A(net659));
 sg13g2_buf_1 _18943_ (.A(_12090_),
    .X(_12091_));
 sg13g2_mux2_1 _18944_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][10] ),
    .S(_12091_),
    .X(_12092_));
 sg13g2_nor2b_1 _18945_ (.A(net1025),
    .B_N(_08351_),
    .Y(_12093_));
 sg13g2_nand2_1 _18946_ (.Y(_12094_),
    .A(net1154),
    .B(_12093_));
 sg13g2_buf_4 _18947_ (.X(_12095_),
    .A(_12094_));
 sg13g2_mux2_1 _18948_ (.A0(_10215_),
    .A1(_10105_),
    .S(_12095_),
    .X(_12096_));
 sg13g2_buf_2 _18949_ (.A(_12096_),
    .X(_12097_));
 sg13g2_buf_1 _18950_ (.A(_12097_),
    .X(_12098_));
 sg13g2_mux2_1 _18951_ (.A0(net1119),
    .A1(_10091_),
    .S(net1154),
    .X(_12099_));
 sg13g2_nand2_1 _18952_ (.Y(_12100_),
    .A(_12093_),
    .B(_12099_));
 sg13g2_nor2_1 _18953_ (.A(_12079_),
    .B(_12100_),
    .Y(_12101_));
 sg13g2_buf_4 _18954_ (.X(_12102_),
    .A(_12101_));
 sg13g2_mux2_1 _18955_ (.A0(_12092_),
    .A1(net482),
    .S(_12102_),
    .X(_00325_));
 sg13g2_buf_1 _18956_ (.A(uio_in[3]),
    .X(_12103_));
 sg13g2_buf_1 _18957_ (.A(_12103_),
    .X(_12104_));
 sg13g2_mux2_1 _18958_ (.A0(_12104_),
    .A1(\cpu.dcache.r_data[0][11] ),
    .S(_12091_),
    .X(_12105_));
 sg13g2_mux2_1 _18959_ (.A0(_10222_),
    .A1(net1133),
    .S(_12095_),
    .X(_12106_));
 sg13g2_buf_2 _18960_ (.A(_12106_),
    .X(_12107_));
 sg13g2_buf_1 _18961_ (.A(_12107_),
    .X(_12108_));
 sg13g2_mux2_1 _18962_ (.A0(_12105_),
    .A1(net481),
    .S(_12102_),
    .X(_00326_));
 sg13g2_nand2b_1 _18963_ (.Y(_12109_),
    .B(_12059_),
    .A_N(net1026));
 sg13g2_or2_1 _18964_ (.X(_12110_),
    .B(_12109_),
    .A(_12058_));
 sg13g2_buf_2 _18965_ (.A(_12110_),
    .X(_12111_));
 sg13g2_or2_1 _18966_ (.X(_12112_),
    .B(_12111_),
    .A(_12054_));
 sg13g2_buf_1 _18967_ (.A(_12112_),
    .X(_12113_));
 sg13g2_mux2_1 _18968_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][12] ),
    .S(_12113_),
    .X(_12114_));
 sg13g2_mux2_1 _18969_ (.A0(_10227_),
    .A1(_10116_),
    .S(_12095_),
    .X(_12115_));
 sg13g2_buf_2 _18970_ (.A(_12115_),
    .X(_12116_));
 sg13g2_buf_1 _18971_ (.A(_12116_),
    .X(_12117_));
 sg13g2_mux2_1 _18972_ (.A0(_12114_),
    .A1(net480),
    .S(_12102_),
    .X(_00327_));
 sg13g2_buf_1 _18973_ (.A(uio_in[1]),
    .X(_12118_));
 sg13g2_buf_2 _18974_ (.A(_12118_),
    .X(_12119_));
 sg13g2_mux2_1 _18975_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][13] ),
    .S(_12113_),
    .X(_12120_));
 sg13g2_mux2_1 _18976_ (.A0(_10229_),
    .A1(_10122_),
    .S(_12095_),
    .X(_12121_));
 sg13g2_buf_2 _18977_ (.A(_12121_),
    .X(_12122_));
 sg13g2_buf_1 _18978_ (.A(_12122_),
    .X(_12123_));
 sg13g2_mux2_1 _18979_ (.A0(_12120_),
    .A1(net479),
    .S(_12102_),
    .X(_00328_));
 sg13g2_mux2_1 _18980_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][14] ),
    .S(_12113_),
    .X(_12124_));
 sg13g2_mux2_1 _18981_ (.A0(_10239_),
    .A1(_10128_),
    .S(_12095_),
    .X(_12125_));
 sg13g2_buf_2 _18982_ (.A(_12125_),
    .X(_12126_));
 sg13g2_buf_1 _18983_ (.A(_12126_),
    .X(_12127_));
 sg13g2_mux2_1 _18984_ (.A0(_12124_),
    .A1(net478),
    .S(_12102_),
    .X(_00329_));
 sg13g2_mux2_1 _18985_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][15] ),
    .S(_12113_),
    .X(_12128_));
 sg13g2_mux2_1 _18986_ (.A0(_10244_),
    .A1(_10131_),
    .S(_12095_),
    .X(_12129_));
 sg13g2_buf_2 _18987_ (.A(_12129_),
    .X(_12130_));
 sg13g2_buf_1 _18988_ (.A(_12130_),
    .X(_12131_));
 sg13g2_mux2_1 _18989_ (.A0(_12128_),
    .A1(net477),
    .S(_12102_),
    .X(_00330_));
 sg13g2_or2_1 _18990_ (.X(_12132_),
    .B(_12063_),
    .A(_12073_));
 sg13g2_buf_2 _18991_ (.A(_12132_),
    .X(_12133_));
 sg13g2_or2_1 _18992_ (.X(_12134_),
    .B(_12133_),
    .A(net659));
 sg13g2_buf_1 _18993_ (.A(_12134_),
    .X(_12135_));
 sg13g2_mux2_1 _18994_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][16] ),
    .S(_12135_),
    .X(_12136_));
 sg13g2_o21ai_1 _18995_ (.B1(_10020_),
    .Y(_12137_),
    .A1(net1154),
    .A2(_12081_));
 sg13g2_nor2_1 _18996_ (.A(_12079_),
    .B(_12137_),
    .Y(_12138_));
 sg13g2_buf_4 _18997_ (.X(_12139_),
    .A(_12138_));
 sg13g2_mux2_1 _18998_ (.A0(_12136_),
    .A1(_12069_),
    .S(_12139_),
    .X(_00331_));
 sg13g2_mux2_1 _18999_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][17] ),
    .S(_12135_),
    .X(_12140_));
 sg13g2_mux2_1 _19000_ (.A0(_12140_),
    .A1(net898),
    .S(_12139_),
    .X(_00332_));
 sg13g2_mux2_1 _19001_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][18] ),
    .S(_12135_),
    .X(_12141_));
 sg13g2_mux2_1 _19002_ (.A0(_12141_),
    .A1(_10165_),
    .S(_12139_),
    .X(_00333_));
 sg13g2_mux2_1 _19003_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][19] ),
    .S(_12135_),
    .X(_12142_));
 sg13g2_mux2_1 _19004_ (.A0(_12142_),
    .A1(net896),
    .S(_12139_),
    .X(_00334_));
 sg13g2_mux2_1 _19005_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][1] ),
    .S(_12067_),
    .X(_12143_));
 sg13g2_mux2_1 _19006_ (.A0(_12143_),
    .A1(_10145_),
    .S(_12085_),
    .X(_00335_));
 sg13g2_nor2_2 _19007_ (.A(_12059_),
    .B(_12061_),
    .Y(_12144_));
 sg13g2_nor2b_2 _19008_ (.A(_12073_),
    .B_N(_12144_),
    .Y(_12145_));
 sg13g2_nand2b_1 _19009_ (.Y(_12146_),
    .B(_12145_),
    .A_N(net659));
 sg13g2_buf_1 _19010_ (.A(_12146_),
    .X(_12147_));
 sg13g2_mux2_1 _19011_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][20] ),
    .S(_12147_),
    .X(_12148_));
 sg13g2_mux2_1 _19012_ (.A0(_12148_),
    .A1(net1047),
    .S(_12139_),
    .X(_00336_));
 sg13g2_mux2_1 _19013_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][21] ),
    .S(_12147_),
    .X(_12149_));
 sg13g2_mux2_1 _19014_ (.A0(_12149_),
    .A1(net895),
    .S(_12139_),
    .X(_00337_));
 sg13g2_mux2_1 _19015_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][22] ),
    .S(_12147_),
    .X(_12150_));
 sg13g2_mux2_1 _19016_ (.A0(_12150_),
    .A1(net894),
    .S(_12139_),
    .X(_00338_));
 sg13g2_mux2_1 _19017_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][23] ),
    .S(_12147_),
    .X(_12151_));
 sg13g2_mux2_1 _19018_ (.A0(_12151_),
    .A1(_10133_),
    .S(_12139_),
    .X(_00339_));
 sg13g2_nand2b_1 _19019_ (.Y(_12152_),
    .B(_12074_),
    .A_N(net659));
 sg13g2_buf_1 _19020_ (.A(_12152_),
    .X(_12153_));
 sg13g2_mux2_1 _19021_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net534),
    .X(_12154_));
 sg13g2_mux2_1 _19022_ (.A0(_10205_),
    .A1(_10080_),
    .S(_12095_),
    .X(_12155_));
 sg13g2_buf_2 _19023_ (.A(_12155_),
    .X(_12156_));
 sg13g2_buf_1 _19024_ (.A(_12156_),
    .X(_12157_));
 sg13g2_nor2_1 _19025_ (.A(net1154),
    .B(net772),
    .Y(_12158_));
 sg13g2_a21oi_1 _19026_ (.A1(net1154),
    .A2(_12082_),
    .Y(_12159_),
    .B1(_12158_));
 sg13g2_nand2_1 _19027_ (.Y(_12160_),
    .A(_12093_),
    .B(_12159_));
 sg13g2_nor2_1 _19028_ (.A(_12079_),
    .B(_12160_),
    .Y(_12161_));
 sg13g2_buf_4 _19029_ (.X(_12162_),
    .A(_12161_));
 sg13g2_mux2_1 _19030_ (.A0(_12154_),
    .A1(net476),
    .S(_12162_),
    .X(_00340_));
 sg13g2_mux2_1 _19031_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net534),
    .X(_12163_));
 sg13g2_mux2_1 _19032_ (.A0(_10210_),
    .A1(_10087_),
    .S(_12095_),
    .X(_12164_));
 sg13g2_buf_2 _19033_ (.A(_12164_),
    .X(_12165_));
 sg13g2_buf_1 _19034_ (.A(_12165_),
    .X(_12166_));
 sg13g2_mux2_1 _19035_ (.A0(_12163_),
    .A1(net475),
    .S(_12162_),
    .X(_00341_));
 sg13g2_mux2_1 _19036_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net534),
    .X(_12167_));
 sg13g2_mux2_1 _19037_ (.A0(_12167_),
    .A1(_12098_),
    .S(_12162_),
    .X(_00342_));
 sg13g2_mux2_1 _19038_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(net534),
    .X(_12168_));
 sg13g2_mux2_1 _19039_ (.A0(_12168_),
    .A1(_12108_),
    .S(_12162_),
    .X(_00343_));
 sg13g2_or2_1 _19040_ (.X(_12169_),
    .B(_12109_),
    .A(_12073_));
 sg13g2_buf_2 _19041_ (.A(_12169_),
    .X(_12170_));
 sg13g2_or2_1 _19042_ (.X(_12171_),
    .B(_12170_),
    .A(_12054_));
 sg13g2_buf_1 _19043_ (.A(_12171_),
    .X(_12172_));
 sg13g2_mux2_1 _19044_ (.A0(_12052_),
    .A1(\cpu.dcache.r_data[0][28] ),
    .S(_12172_),
    .X(_12173_));
 sg13g2_mux2_1 _19045_ (.A0(_12173_),
    .A1(net480),
    .S(_12162_),
    .X(_00344_));
 sg13g2_mux2_1 _19046_ (.A0(_12119_),
    .A1(\cpu.dcache.r_data[0][29] ),
    .S(_12172_),
    .X(_12174_));
 sg13g2_mux2_1 _19047_ (.A0(_12174_),
    .A1(net479),
    .S(_12162_),
    .X(_00345_));
 sg13g2_mux2_1 _19048_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][2] ),
    .S(_12067_),
    .X(_12175_));
 sg13g2_mux2_1 _19049_ (.A0(_12175_),
    .A1(net897),
    .S(_12085_),
    .X(_00346_));
 sg13g2_mux2_1 _19050_ (.A0(_12087_),
    .A1(\cpu.dcache.r_data[0][30] ),
    .S(_12172_),
    .X(_12176_));
 sg13g2_mux2_1 _19051_ (.A0(_12176_),
    .A1(_12127_),
    .S(_12162_),
    .X(_00347_));
 sg13g2_mux2_1 _19052_ (.A0(_12104_),
    .A1(\cpu.dcache.r_data[0][31] ),
    .S(_12172_),
    .X(_12177_));
 sg13g2_mux2_1 _19053_ (.A0(_12177_),
    .A1(_12131_),
    .S(_12162_),
    .X(_00348_));
 sg13g2_mux2_1 _19054_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][3] ),
    .S(_12067_),
    .X(_12178_));
 sg13g2_mux2_1 _19055_ (.A0(_12178_),
    .A1(_10170_),
    .S(_12085_),
    .X(_00349_));
 sg13g2_nor2b_2 _19056_ (.A(_12058_),
    .B_N(_12144_),
    .Y(_12179_));
 sg13g2_nand2b_1 _19057_ (.Y(_12180_),
    .B(_12179_),
    .A_N(net659));
 sg13g2_buf_1 _19058_ (.A(_12180_),
    .X(_12181_));
 sg13g2_mux2_1 _19059_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][4] ),
    .S(_12181_),
    .X(_12182_));
 sg13g2_mux2_1 _19060_ (.A0(_12182_),
    .A1(_10176_),
    .S(_12085_),
    .X(_00350_));
 sg13g2_mux2_1 _19061_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][5] ),
    .S(_12181_),
    .X(_12183_));
 sg13g2_mux2_1 _19062_ (.A0(_12183_),
    .A1(_10181_),
    .S(_12085_),
    .X(_00351_));
 sg13g2_mux2_1 _19063_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[0][6] ),
    .S(_12181_),
    .X(_12184_));
 sg13g2_mux2_1 _19064_ (.A0(_12184_),
    .A1(net894),
    .S(_12085_),
    .X(_00352_));
 sg13g2_mux2_1 _19065_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[0][7] ),
    .S(_12181_),
    .X(_12185_));
 sg13g2_mux2_1 _19066_ (.A0(_12185_),
    .A1(_10133_),
    .S(_12085_),
    .X(_00353_));
 sg13g2_mux2_1 _19067_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[0][8] ),
    .S(_12091_),
    .X(_12186_));
 sg13g2_mux2_1 _19068_ (.A0(_12186_),
    .A1(net476),
    .S(_12102_),
    .X(_00354_));
 sg13g2_mux2_1 _19069_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[0][9] ),
    .S(_12091_),
    .X(_12187_));
 sg13g2_mux2_1 _19070_ (.A0(_12187_),
    .A1(net475),
    .S(_12102_),
    .X(_00355_));
 sg13g2_buf_1 _19071_ (.A(_09788_),
    .X(_12188_));
 sg13g2_buf_1 _19072_ (.A(net745),
    .X(_12189_));
 sg13g2_or2_1 _19073_ (.X(_12190_),
    .B(_12083_),
    .A(_12077_));
 sg13g2_buf_2 _19074_ (.A(_12190_),
    .X(_12191_));
 sg13g2_nor2_1 _19075_ (.A(net658),
    .B(_12191_),
    .Y(_12192_));
 sg13g2_buf_2 _19076_ (.A(_12192_),
    .X(_12193_));
 sg13g2_buf_1 _19077_ (.A(_12193_),
    .X(_12194_));
 sg13g2_buf_1 _19078_ (.A(_12051_),
    .X(_12195_));
 sg13g2_buf_1 _19079_ (.A(net1115),
    .X(_12196_));
 sg13g2_nor2_1 _19080_ (.A(net658),
    .B(_12065_),
    .Y(_12197_));
 sg13g2_buf_2 _19081_ (.A(_12197_),
    .X(_12198_));
 sg13g2_nor2b_1 _19082_ (.A(_12198_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12199_));
 sg13g2_a21oi_1 _19083_ (.A1(net1024),
    .A2(_12198_),
    .Y(_12200_),
    .B1(_12199_));
 sg13g2_buf_1 _19084_ (.A(net1057),
    .X(_12201_));
 sg13g2_nand2_1 _19085_ (.Y(_12202_),
    .A(net868),
    .B(net57));
 sg13g2_o21ai_1 _19086_ (.B1(_12202_),
    .Y(_00356_),
    .A1(net57),
    .A2(_12200_));
 sg13g2_or2_1 _19087_ (.X(_12203_),
    .B(_12100_),
    .A(_12077_));
 sg13g2_buf_2 _19088_ (.A(_12203_),
    .X(_12204_));
 sg13g2_or2_1 _19089_ (.X(_12205_),
    .B(_12204_),
    .A(net745));
 sg13g2_buf_1 _19090_ (.A(_12205_),
    .X(_12206_));
 sg13g2_buf_1 _19091_ (.A(_12206_),
    .X(_12207_));
 sg13g2_buf_1 _19092_ (.A(_12086_),
    .X(_12208_));
 sg13g2_buf_2 _19093_ (.A(net1114),
    .X(_12209_));
 sg13g2_nor2_1 _19094_ (.A(net658),
    .B(_12089_),
    .Y(_12210_));
 sg13g2_buf_2 _19095_ (.A(_12210_),
    .X(_12211_));
 sg13g2_nor2b_1 _19096_ (.A(_12211_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12212_));
 sg13g2_a21oi_1 _19097_ (.A1(net1023),
    .A2(_12211_),
    .Y(_12213_),
    .B1(_12212_));
 sg13g2_nor2_1 _19098_ (.A(_12097_),
    .B(net56),
    .Y(_12214_));
 sg13g2_a21oi_1 _19099_ (.A1(net56),
    .A2(_12213_),
    .Y(_00357_),
    .B1(_12214_));
 sg13g2_buf_1 _19100_ (.A(_12103_),
    .X(_12215_));
 sg13g2_buf_2 _19101_ (.A(net1113),
    .X(_12216_));
 sg13g2_nor2b_1 _19102_ (.A(_12211_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12217_));
 sg13g2_a21oi_1 _19103_ (.A1(net1022),
    .A2(_12211_),
    .Y(_12218_),
    .B1(_12217_));
 sg13g2_nor2_1 _19104_ (.A(_12107_),
    .B(net56),
    .Y(_12219_));
 sg13g2_a21oi_1 _19105_ (.A1(net56),
    .A2(_12218_),
    .Y(_00358_),
    .B1(_12219_));
 sg13g2_buf_2 _19106_ (.A(net1115),
    .X(_12220_));
 sg13g2_nor2_1 _19107_ (.A(_12189_),
    .B(_12111_),
    .Y(_12221_));
 sg13g2_buf_2 _19108_ (.A(_12221_),
    .X(_12222_));
 sg13g2_nor2b_1 _19109_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[1][12] ),
    .Y(_12223_));
 sg13g2_a21oi_1 _19110_ (.A1(net1021),
    .A2(_12222_),
    .Y(_12224_),
    .B1(_12223_));
 sg13g2_nor2_1 _19111_ (.A(_12116_),
    .B(_12206_),
    .Y(_12225_));
 sg13g2_a21oi_1 _19112_ (.A1(_12207_),
    .A2(_12224_),
    .Y(_00359_),
    .B1(_12225_));
 sg13g2_buf_1 _19113_ (.A(_12118_),
    .X(_12226_));
 sg13g2_buf_2 _19114_ (.A(net1112),
    .X(_12227_));
 sg13g2_nor2b_1 _19115_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[1][13] ),
    .Y(_12228_));
 sg13g2_a21oi_1 _19116_ (.A1(net1020),
    .A2(_12222_),
    .Y(_12229_),
    .B1(_12228_));
 sg13g2_nor2_1 _19117_ (.A(_12122_),
    .B(_12206_),
    .Y(_12230_));
 sg13g2_a21oi_1 _19118_ (.A1(net56),
    .A2(_12229_),
    .Y(_00360_),
    .B1(_12230_));
 sg13g2_nor2b_1 _19119_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[1][14] ),
    .Y(_12231_));
 sg13g2_a21oi_1 _19120_ (.A1(net1023),
    .A2(_12222_),
    .Y(_12232_),
    .B1(_12231_));
 sg13g2_nor2_1 _19121_ (.A(_12126_),
    .B(_12206_),
    .Y(_12233_));
 sg13g2_a21oi_1 _19122_ (.A1(_12207_),
    .A2(_12232_),
    .Y(_00361_),
    .B1(_12233_));
 sg13g2_nor2b_1 _19123_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[1][15] ),
    .Y(_12234_));
 sg13g2_a21oi_1 _19124_ (.A1(net1022),
    .A2(_12222_),
    .Y(_12235_),
    .B1(_12234_));
 sg13g2_nor2_1 _19125_ (.A(_12130_),
    .B(_12206_),
    .Y(_12236_));
 sg13g2_a21oi_1 _19126_ (.A1(net56),
    .A2(_12235_),
    .Y(_00362_),
    .B1(_12236_));
 sg13g2_or2_1 _19127_ (.X(_12237_),
    .B(_12137_),
    .A(_12077_));
 sg13g2_buf_2 _19128_ (.A(_12237_),
    .X(_12238_));
 sg13g2_nor2_1 _19129_ (.A(net658),
    .B(_12238_),
    .Y(_12239_));
 sg13g2_buf_2 _19130_ (.A(_12239_),
    .X(_12240_));
 sg13g2_buf_1 _19131_ (.A(_12240_),
    .X(_12241_));
 sg13g2_nor2_1 _19132_ (.A(net658),
    .B(_12133_),
    .Y(_12242_));
 sg13g2_buf_2 _19133_ (.A(_12242_),
    .X(_12243_));
 sg13g2_nor2b_1 _19134_ (.A(_12243_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12244_));
 sg13g2_a21oi_1 _19135_ (.A1(net1024),
    .A2(_12243_),
    .Y(_12245_),
    .B1(_12244_));
 sg13g2_nand2_1 _19136_ (.Y(_12246_),
    .A(net868),
    .B(net55));
 sg13g2_o21ai_1 _19137_ (.B1(_12246_),
    .Y(_00363_),
    .A1(net55),
    .A2(_12245_));
 sg13g2_buf_1 _19138_ (.A(net1112),
    .X(_12247_));
 sg13g2_nor2b_1 _19139_ (.A(_12243_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_12248_));
 sg13g2_a21oi_1 _19140_ (.A1(net1019),
    .A2(_12243_),
    .Y(_12249_),
    .B1(_12248_));
 sg13g2_buf_1 _19141_ (.A(net1049),
    .X(_12250_));
 sg13g2_nand2_1 _19142_ (.Y(_12251_),
    .A(net867),
    .B(net55));
 sg13g2_o21ai_1 _19143_ (.B1(_12251_),
    .Y(_00364_),
    .A1(net55),
    .A2(_12249_));
 sg13g2_buf_1 _19144_ (.A(net1114),
    .X(_12252_));
 sg13g2_nor2b_1 _19145_ (.A(_12243_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_12253_));
 sg13g2_a21oi_1 _19146_ (.A1(net1018),
    .A2(_12243_),
    .Y(_12254_),
    .B1(_12253_));
 sg13g2_buf_1 _19147_ (.A(net1048),
    .X(_12255_));
 sg13g2_nand2_1 _19148_ (.Y(_12256_),
    .A(net866),
    .B(_12240_));
 sg13g2_o21ai_1 _19149_ (.B1(_12256_),
    .Y(_00365_),
    .A1(net55),
    .A2(_12254_));
 sg13g2_buf_1 _19150_ (.A(net1113),
    .X(_12257_));
 sg13g2_nor2b_1 _19151_ (.A(_12243_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_12258_));
 sg13g2_a21oi_1 _19152_ (.A1(net1017),
    .A2(_12243_),
    .Y(_12259_),
    .B1(_12258_));
 sg13g2_buf_1 _19153_ (.A(net1133),
    .X(_12260_));
 sg13g2_nand2_1 _19154_ (.Y(_12261_),
    .A(net1016),
    .B(_12240_));
 sg13g2_o21ai_1 _19155_ (.B1(_12261_),
    .Y(_00366_),
    .A1(_12241_),
    .A2(_12259_));
 sg13g2_nor2b_1 _19156_ (.A(_12198_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_12262_));
 sg13g2_a21oi_1 _19157_ (.A1(net1019),
    .A2(_12198_),
    .Y(_12263_),
    .B1(_12262_));
 sg13g2_nand2_1 _19158_ (.Y(_12264_),
    .A(net867),
    .B(net57));
 sg13g2_o21ai_1 _19159_ (.B1(_12264_),
    .Y(_00367_),
    .A1(net57),
    .A2(_12263_));
 sg13g2_nand2b_1 _19160_ (.Y(_12265_),
    .B(_12144_),
    .A_N(_12073_));
 sg13g2_buf_1 _19161_ (.A(_12265_),
    .X(_12266_));
 sg13g2_nor2_1 _19162_ (.A(net658),
    .B(_12266_),
    .Y(_12267_));
 sg13g2_buf_2 _19163_ (.A(_12267_),
    .X(_12268_));
 sg13g2_nor2b_1 _19164_ (.A(_12268_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_12269_));
 sg13g2_a21oi_1 _19165_ (.A1(net1024),
    .A2(_12268_),
    .Y(_12270_),
    .B1(_12269_));
 sg13g2_buf_1 _19166_ (.A(_10116_),
    .X(_12271_));
 sg13g2_nand2_1 _19167_ (.Y(_12272_),
    .A(net1015),
    .B(_12240_));
 sg13g2_o21ai_1 _19168_ (.B1(_12272_),
    .Y(_00368_),
    .A1(net55),
    .A2(_12270_));
 sg13g2_nor2b_1 _19169_ (.A(_12268_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_12273_));
 sg13g2_a21oi_1 _19170_ (.A1(net1019),
    .A2(_12268_),
    .Y(_12274_),
    .B1(_12273_));
 sg13g2_buf_1 _19171_ (.A(_10122_),
    .X(_12275_));
 sg13g2_nand2_1 _19172_ (.Y(_12276_),
    .A(_12275_),
    .B(_12240_));
 sg13g2_o21ai_1 _19173_ (.B1(_12276_),
    .Y(_00369_),
    .A1(net55),
    .A2(_12274_));
 sg13g2_nor2b_1 _19174_ (.A(_12268_),
    .B_N(\cpu.dcache.r_data[1][22] ),
    .Y(_12277_));
 sg13g2_a21oi_1 _19175_ (.A1(net1018),
    .A2(_12268_),
    .Y(_12278_),
    .B1(_12277_));
 sg13g2_buf_1 _19176_ (.A(_10128_),
    .X(_12279_));
 sg13g2_nand2_1 _19177_ (.Y(_12280_),
    .A(net1013),
    .B(_12240_));
 sg13g2_o21ai_1 _19178_ (.B1(_12280_),
    .Y(_00370_),
    .A1(net55),
    .A2(_12278_));
 sg13g2_nor2b_1 _19179_ (.A(_12268_),
    .B_N(\cpu.dcache.r_data[1][23] ),
    .Y(_12281_));
 sg13g2_a21oi_1 _19180_ (.A1(net1017),
    .A2(_12268_),
    .Y(_12282_),
    .B1(_12281_));
 sg13g2_buf_1 _19181_ (.A(_10131_),
    .X(_12283_));
 sg13g2_nand2_1 _19182_ (.Y(_12284_),
    .A(net1012),
    .B(_12240_));
 sg13g2_o21ai_1 _19183_ (.B1(_12284_),
    .Y(_00371_),
    .A1(_12241_),
    .A2(_12282_));
 sg13g2_or2_1 _19184_ (.X(_12285_),
    .B(_12160_),
    .A(_12077_));
 sg13g2_buf_2 _19185_ (.A(_12285_),
    .X(_12286_));
 sg13g2_or2_1 _19186_ (.X(_12287_),
    .B(_12286_),
    .A(net745));
 sg13g2_buf_1 _19187_ (.A(_12287_),
    .X(_12288_));
 sg13g2_buf_1 _19188_ (.A(_12288_),
    .X(_12289_));
 sg13g2_or2_1 _19189_ (.X(_12290_),
    .B(_12073_),
    .A(_12070_));
 sg13g2_buf_2 _19190_ (.A(_12290_),
    .X(_12291_));
 sg13g2_nor2_1 _19191_ (.A(_12188_),
    .B(_12291_),
    .Y(_12292_));
 sg13g2_buf_1 _19192_ (.A(_12292_),
    .X(_12293_));
 sg13g2_nor2b_1 _19193_ (.A(net533),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12294_));
 sg13g2_a21oi_1 _19194_ (.A1(net1021),
    .A2(net533),
    .Y(_12295_),
    .B1(_12294_));
 sg13g2_nor2_1 _19195_ (.A(_12156_),
    .B(net54),
    .Y(_12296_));
 sg13g2_a21oi_1 _19196_ (.A1(net54),
    .A2(_12295_),
    .Y(_00372_),
    .B1(_12296_));
 sg13g2_nor2b_1 _19197_ (.A(net533),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12297_));
 sg13g2_a21oi_1 _19198_ (.A1(net1020),
    .A2(net533),
    .Y(_12298_),
    .B1(_12297_));
 sg13g2_nor2_1 _19199_ (.A(_12165_),
    .B(_12289_),
    .Y(_12299_));
 sg13g2_a21oi_1 _19200_ (.A1(_12289_),
    .A2(_12298_),
    .Y(_00373_),
    .B1(_12299_));
 sg13g2_nor2b_1 _19201_ (.A(net533),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12300_));
 sg13g2_a21oi_1 _19202_ (.A1(net1023),
    .A2(net533),
    .Y(_12301_),
    .B1(_12300_));
 sg13g2_nor2_1 _19203_ (.A(_12097_),
    .B(_12288_),
    .Y(_12302_));
 sg13g2_a21oi_1 _19204_ (.A1(net54),
    .A2(_12301_),
    .Y(_00374_),
    .B1(_12302_));
 sg13g2_nor2b_1 _19205_ (.A(net533),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12303_));
 sg13g2_a21oi_1 _19206_ (.A1(net1022),
    .A2(_12293_),
    .Y(_12304_),
    .B1(_12303_));
 sg13g2_nor2_1 _19207_ (.A(_12107_),
    .B(_12288_),
    .Y(_12305_));
 sg13g2_a21oi_1 _19208_ (.A1(net54),
    .A2(_12304_),
    .Y(_00375_),
    .B1(_12305_));
 sg13g2_nor2_1 _19209_ (.A(_12189_),
    .B(_12170_),
    .Y(_12306_));
 sg13g2_buf_2 _19210_ (.A(_12306_),
    .X(_12307_));
 sg13g2_nor2b_1 _19211_ (.A(_12307_),
    .B_N(\cpu.dcache.r_data[1][28] ),
    .Y(_12308_));
 sg13g2_a21oi_1 _19212_ (.A1(net1021),
    .A2(_12307_),
    .Y(_12309_),
    .B1(_12308_));
 sg13g2_nor2_1 _19213_ (.A(_12116_),
    .B(_12288_),
    .Y(_12310_));
 sg13g2_a21oi_1 _19214_ (.A1(net54),
    .A2(_12309_),
    .Y(_00376_),
    .B1(_12310_));
 sg13g2_nor2b_1 _19215_ (.A(_12307_),
    .B_N(\cpu.dcache.r_data[1][29] ),
    .Y(_12311_));
 sg13g2_a21oi_1 _19216_ (.A1(net1020),
    .A2(_12307_),
    .Y(_12312_),
    .B1(_12311_));
 sg13g2_nor2_1 _19217_ (.A(_12122_),
    .B(_12288_),
    .Y(_12313_));
 sg13g2_a21oi_1 _19218_ (.A1(net54),
    .A2(_12312_),
    .Y(_00377_),
    .B1(_12313_));
 sg13g2_nor2b_1 _19219_ (.A(_12198_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12314_));
 sg13g2_a21oi_1 _19220_ (.A1(net1018),
    .A2(_12198_),
    .Y(_12315_),
    .B1(_12314_));
 sg13g2_nand2_1 _19221_ (.Y(_12316_),
    .A(net866),
    .B(_12193_));
 sg13g2_o21ai_1 _19222_ (.B1(_12316_),
    .Y(_00378_),
    .A1(net57),
    .A2(_12315_));
 sg13g2_nor2b_1 _19223_ (.A(_12307_),
    .B_N(\cpu.dcache.r_data[1][30] ),
    .Y(_12317_));
 sg13g2_a21oi_1 _19224_ (.A1(net1023),
    .A2(_12307_),
    .Y(_12318_),
    .B1(_12317_));
 sg13g2_nor2_1 _19225_ (.A(_12126_),
    .B(_12288_),
    .Y(_12319_));
 sg13g2_a21oi_1 _19226_ (.A1(net54),
    .A2(_12318_),
    .Y(_00379_),
    .B1(_12319_));
 sg13g2_nor2b_1 _19227_ (.A(_12307_),
    .B_N(\cpu.dcache.r_data[1][31] ),
    .Y(_12320_));
 sg13g2_a21oi_1 _19228_ (.A1(net1022),
    .A2(_12307_),
    .Y(_12321_),
    .B1(_12320_));
 sg13g2_nor2_1 _19229_ (.A(_12130_),
    .B(_12288_),
    .Y(_12322_));
 sg13g2_a21oi_1 _19230_ (.A1(net54),
    .A2(_12321_),
    .Y(_00380_),
    .B1(_12322_));
 sg13g2_nor2b_1 _19231_ (.A(_12198_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12323_));
 sg13g2_a21oi_1 _19232_ (.A1(net1017),
    .A2(_12198_),
    .Y(_12324_),
    .B1(_12323_));
 sg13g2_nand2_1 _19233_ (.Y(_12325_),
    .A(net1016),
    .B(_12193_));
 sg13g2_o21ai_1 _19234_ (.B1(_12325_),
    .Y(_00381_),
    .A1(_12194_),
    .A2(_12324_));
 sg13g2_nand2b_1 _19235_ (.Y(_12326_),
    .B(_12144_),
    .A_N(_12058_));
 sg13g2_buf_1 _19236_ (.A(_12326_),
    .X(_12327_));
 sg13g2_nor2_1 _19237_ (.A(net745),
    .B(_12327_),
    .Y(_12328_));
 sg13g2_buf_2 _19238_ (.A(_12328_),
    .X(_12329_));
 sg13g2_nor2b_1 _19239_ (.A(_12329_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12330_));
 sg13g2_a21oi_1 _19240_ (.A1(net1024),
    .A2(_12329_),
    .Y(_12331_),
    .B1(_12330_));
 sg13g2_nand2_1 _19241_ (.Y(_12332_),
    .A(net1015),
    .B(_12193_));
 sg13g2_o21ai_1 _19242_ (.B1(_12332_),
    .Y(_00382_),
    .A1(net57),
    .A2(_12331_));
 sg13g2_nor2b_1 _19243_ (.A(_12329_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12333_));
 sg13g2_a21oi_1 _19244_ (.A1(net1019),
    .A2(_12329_),
    .Y(_12334_),
    .B1(_12333_));
 sg13g2_buf_1 _19245_ (.A(_10122_),
    .X(_12335_));
 sg13g2_nand2_1 _19246_ (.Y(_12336_),
    .A(net1011),
    .B(_12193_));
 sg13g2_o21ai_1 _19247_ (.B1(_12336_),
    .Y(_00383_),
    .A1(_12194_),
    .A2(_12334_));
 sg13g2_nor2b_1 _19248_ (.A(_12329_),
    .B_N(\cpu.dcache.r_data[1][6] ),
    .Y(_12337_));
 sg13g2_a21oi_1 _19249_ (.A1(net1018),
    .A2(_12329_),
    .Y(_12338_),
    .B1(_12337_));
 sg13g2_buf_1 _19250_ (.A(_10128_),
    .X(_12339_));
 sg13g2_nand2_1 _19251_ (.Y(_12340_),
    .A(net1010),
    .B(_12193_));
 sg13g2_o21ai_1 _19252_ (.B1(_12340_),
    .Y(_00384_),
    .A1(net57),
    .A2(_12338_));
 sg13g2_nor2b_1 _19253_ (.A(_12329_),
    .B_N(\cpu.dcache.r_data[1][7] ),
    .Y(_12341_));
 sg13g2_a21oi_1 _19254_ (.A1(net1017),
    .A2(_12329_),
    .Y(_12342_),
    .B1(_12341_));
 sg13g2_nand2_1 _19255_ (.Y(_12343_),
    .A(net1012),
    .B(_12193_));
 sg13g2_o21ai_1 _19256_ (.B1(_12343_),
    .Y(_00385_),
    .A1(net57),
    .A2(_12342_));
 sg13g2_nor2b_1 _19257_ (.A(_12211_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12344_));
 sg13g2_a21oi_1 _19258_ (.A1(net1021),
    .A2(_12211_),
    .Y(_12345_),
    .B1(_12344_));
 sg13g2_nor2_1 _19259_ (.A(_12156_),
    .B(_12206_),
    .Y(_12346_));
 sg13g2_a21oi_1 _19260_ (.A1(net56),
    .A2(_12345_),
    .Y(_00386_),
    .B1(_12346_));
 sg13g2_nor2b_1 _19261_ (.A(_12211_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12347_));
 sg13g2_a21oi_1 _19262_ (.A1(net1020),
    .A2(_12211_),
    .Y(_12348_),
    .B1(_12347_));
 sg13g2_nor2_1 _19263_ (.A(_12165_),
    .B(_12206_),
    .Y(_12349_));
 sg13g2_a21oi_1 _19264_ (.A1(net56),
    .A2(_12348_),
    .Y(_00387_),
    .B1(_12349_));
 sg13g2_nand2_1 _19265_ (.Y(_12350_),
    .A(net1061),
    .B(_09728_));
 sg13g2_buf_1 _19266_ (.A(_12350_),
    .X(_12351_));
 sg13g2_buf_1 _19267_ (.A(_12351_),
    .X(_12352_));
 sg13g2_nor2_1 _19268_ (.A(net532),
    .B(_12191_),
    .Y(_12353_));
 sg13g2_buf_2 _19269_ (.A(_12353_),
    .X(_12354_));
 sg13g2_buf_1 _19270_ (.A(_12354_),
    .X(_12355_));
 sg13g2_nor2_1 _19271_ (.A(net532),
    .B(_12065_),
    .Y(_12356_));
 sg13g2_buf_2 _19272_ (.A(_12356_),
    .X(_12357_));
 sg13g2_nor2b_1 _19273_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12358_));
 sg13g2_a21oi_1 _19274_ (.A1(net1024),
    .A2(_12357_),
    .Y(_12359_),
    .B1(_12358_));
 sg13g2_nand2_1 _19275_ (.Y(_12360_),
    .A(net868),
    .B(net53));
 sg13g2_o21ai_1 _19276_ (.B1(_12360_),
    .Y(_00388_),
    .A1(net53),
    .A2(_12359_));
 sg13g2_nor2_1 _19277_ (.A(net532),
    .B(_12204_),
    .Y(_12361_));
 sg13g2_buf_2 _19278_ (.A(_12361_),
    .X(_12362_));
 sg13g2_buf_1 _19279_ (.A(_12362_),
    .X(_12363_));
 sg13g2_nor2_1 _19280_ (.A(net532),
    .B(_12089_),
    .Y(_12364_));
 sg13g2_buf_2 _19281_ (.A(_12364_),
    .X(_12365_));
 sg13g2_nor2b_1 _19282_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12366_));
 sg13g2_a21oi_1 _19283_ (.A1(net1018),
    .A2(_12365_),
    .Y(_12367_),
    .B1(_12366_));
 sg13g2_nand2_1 _19284_ (.Y(_12368_),
    .A(net482),
    .B(net52));
 sg13g2_o21ai_1 _19285_ (.B1(_12368_),
    .Y(_00389_),
    .A1(net52),
    .A2(_12367_));
 sg13g2_nor2b_1 _19286_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12369_));
 sg13g2_a21oi_1 _19287_ (.A1(net1017),
    .A2(_12365_),
    .Y(_12370_),
    .B1(_12369_));
 sg13g2_nand2_1 _19288_ (.Y(_12371_),
    .A(net481),
    .B(net52));
 sg13g2_o21ai_1 _19289_ (.B1(_12371_),
    .Y(_00390_),
    .A1(net52),
    .A2(_12370_));
 sg13g2_nor2_1 _19290_ (.A(_12352_),
    .B(_12111_),
    .Y(_12372_));
 sg13g2_buf_2 _19291_ (.A(_12372_),
    .X(_12373_));
 sg13g2_nor2b_1 _19292_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[2][12] ),
    .Y(_12374_));
 sg13g2_a21oi_1 _19293_ (.A1(net1024),
    .A2(_12373_),
    .Y(_12375_),
    .B1(_12374_));
 sg13g2_nand2_1 _19294_ (.Y(_12376_),
    .A(net480),
    .B(_12362_));
 sg13g2_o21ai_1 _19295_ (.B1(_12376_),
    .Y(_00391_),
    .A1(_12363_),
    .A2(_12375_));
 sg13g2_nor2b_1 _19296_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[2][13] ),
    .Y(_12377_));
 sg13g2_a21oi_1 _19297_ (.A1(net1019),
    .A2(_12373_),
    .Y(_12378_),
    .B1(_12377_));
 sg13g2_nand2_1 _19298_ (.Y(_12379_),
    .A(net479),
    .B(_12362_));
 sg13g2_o21ai_1 _19299_ (.B1(_12379_),
    .Y(_00392_),
    .A1(net52),
    .A2(_12378_));
 sg13g2_nor2b_1 _19300_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[2][14] ),
    .Y(_12380_));
 sg13g2_a21oi_1 _19301_ (.A1(net1018),
    .A2(_12373_),
    .Y(_12381_),
    .B1(_12380_));
 sg13g2_nand2_1 _19302_ (.Y(_12382_),
    .A(net478),
    .B(_12362_));
 sg13g2_o21ai_1 _19303_ (.B1(_12382_),
    .Y(_00393_),
    .A1(_12363_),
    .A2(_12381_));
 sg13g2_nor2b_1 _19304_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[2][15] ),
    .Y(_12383_));
 sg13g2_a21oi_1 _19305_ (.A1(net1017),
    .A2(_12373_),
    .Y(_12384_),
    .B1(_12383_));
 sg13g2_nand2_1 _19306_ (.Y(_12385_),
    .A(net477),
    .B(_12362_));
 sg13g2_o21ai_1 _19307_ (.B1(_12385_),
    .Y(_00394_),
    .A1(net52),
    .A2(_12384_));
 sg13g2_nor2_1 _19308_ (.A(net532),
    .B(_12238_),
    .Y(_12386_));
 sg13g2_buf_2 _19309_ (.A(_12386_),
    .X(_12387_));
 sg13g2_buf_1 _19310_ (.A(_12387_),
    .X(_12388_));
 sg13g2_nor2_1 _19311_ (.A(net532),
    .B(_12133_),
    .Y(_12389_));
 sg13g2_buf_2 _19312_ (.A(_12389_),
    .X(_12390_));
 sg13g2_nor2b_1 _19313_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12391_));
 sg13g2_a21oi_1 _19314_ (.A1(net1024),
    .A2(_12390_),
    .Y(_12392_),
    .B1(_12391_));
 sg13g2_nand2_1 _19315_ (.Y(_12393_),
    .A(net868),
    .B(net51));
 sg13g2_o21ai_1 _19316_ (.B1(_12393_),
    .Y(_00395_),
    .A1(net51),
    .A2(_12392_));
 sg13g2_nor2b_1 _19317_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12394_));
 sg13g2_a21oi_1 _19318_ (.A1(net1019),
    .A2(_12390_),
    .Y(_12395_),
    .B1(_12394_));
 sg13g2_nand2_1 _19319_ (.Y(_12396_),
    .A(net867),
    .B(_12388_));
 sg13g2_o21ai_1 _19320_ (.B1(_12396_),
    .Y(_00396_),
    .A1(_12388_),
    .A2(_12395_));
 sg13g2_nor2b_1 _19321_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12397_));
 sg13g2_a21oi_1 _19322_ (.A1(net1018),
    .A2(_12390_),
    .Y(_12398_),
    .B1(_12397_));
 sg13g2_nand2_1 _19323_ (.Y(_12399_),
    .A(net866),
    .B(_12387_));
 sg13g2_o21ai_1 _19324_ (.B1(_12399_),
    .Y(_00397_),
    .A1(net51),
    .A2(_12398_));
 sg13g2_nor2b_1 _19325_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12400_));
 sg13g2_a21oi_1 _19326_ (.A1(net1017),
    .A2(_12390_),
    .Y(_12401_),
    .B1(_12400_));
 sg13g2_nand2_1 _19327_ (.Y(_12402_),
    .A(net1016),
    .B(_12387_));
 sg13g2_o21ai_1 _19328_ (.B1(_12402_),
    .Y(_00398_),
    .A1(net51),
    .A2(_12401_));
 sg13g2_nor2b_1 _19329_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12403_));
 sg13g2_a21oi_1 _19330_ (.A1(net1019),
    .A2(_12357_),
    .Y(_12404_),
    .B1(_12403_));
 sg13g2_nand2_1 _19331_ (.Y(_12405_),
    .A(net867),
    .B(net53));
 sg13g2_o21ai_1 _19332_ (.B1(_12405_),
    .Y(_00399_),
    .A1(net53),
    .A2(_12404_));
 sg13g2_nor2_1 _19333_ (.A(_12351_),
    .B(_12266_),
    .Y(_12406_));
 sg13g2_buf_2 _19334_ (.A(_12406_),
    .X(_12407_));
 sg13g2_nor2b_1 _19335_ (.A(_12407_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12408_));
 sg13g2_a21oi_1 _19336_ (.A1(net1024),
    .A2(_12407_),
    .Y(_12409_),
    .B1(_12408_));
 sg13g2_nand2_1 _19337_ (.Y(_12410_),
    .A(net1015),
    .B(_12387_));
 sg13g2_o21ai_1 _19338_ (.B1(_12410_),
    .Y(_00400_),
    .A1(net51),
    .A2(_12409_));
 sg13g2_nor2b_1 _19339_ (.A(_12407_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12411_));
 sg13g2_a21oi_1 _19340_ (.A1(net1019),
    .A2(_12407_),
    .Y(_12412_),
    .B1(_12411_));
 sg13g2_nand2_1 _19341_ (.Y(_12413_),
    .A(net1011),
    .B(_12387_));
 sg13g2_o21ai_1 _19342_ (.B1(_12413_),
    .Y(_00401_),
    .A1(net51),
    .A2(_12412_));
 sg13g2_nor2b_1 _19343_ (.A(_12407_),
    .B_N(\cpu.dcache.r_data[2][22] ),
    .Y(_12414_));
 sg13g2_a21oi_1 _19344_ (.A1(net1018),
    .A2(_12407_),
    .Y(_12415_),
    .B1(_12414_));
 sg13g2_nand2_1 _19345_ (.Y(_12416_),
    .A(net1010),
    .B(_12387_));
 sg13g2_o21ai_1 _19346_ (.B1(_12416_),
    .Y(_00402_),
    .A1(net51),
    .A2(_12415_));
 sg13g2_nor2b_1 _19347_ (.A(_12407_),
    .B_N(\cpu.dcache.r_data[2][23] ),
    .Y(_12417_));
 sg13g2_a21oi_1 _19348_ (.A1(net1017),
    .A2(_12407_),
    .Y(_12418_),
    .B1(_12417_));
 sg13g2_nand2_1 _19349_ (.Y(_12419_),
    .A(net1012),
    .B(_12387_));
 sg13g2_o21ai_1 _19350_ (.B1(_12419_),
    .Y(_00403_),
    .A1(net51),
    .A2(_12418_));
 sg13g2_nor2_1 _19351_ (.A(_12352_),
    .B(_12286_),
    .Y(_12420_));
 sg13g2_buf_2 _19352_ (.A(_12420_),
    .X(_12421_));
 sg13g2_buf_1 _19353_ (.A(_12421_),
    .X(_12422_));
 sg13g2_nor2_1 _19354_ (.A(_12351_),
    .B(_12291_),
    .Y(_12423_));
 sg13g2_buf_1 _19355_ (.A(_12423_),
    .X(_12424_));
 sg13g2_nor2b_1 _19356_ (.A(net474),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12425_));
 sg13g2_a21oi_1 _19357_ (.A1(_12196_),
    .A2(net474),
    .Y(_12426_),
    .B1(_12425_));
 sg13g2_nand2_1 _19358_ (.Y(_12427_),
    .A(net476),
    .B(net50));
 sg13g2_o21ai_1 _19359_ (.B1(_12427_),
    .Y(_00404_),
    .A1(net50),
    .A2(_12426_));
 sg13g2_nor2b_1 _19360_ (.A(net474),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12428_));
 sg13g2_a21oi_1 _19361_ (.A1(_12247_),
    .A2(net474),
    .Y(_12429_),
    .B1(_12428_));
 sg13g2_nand2_1 _19362_ (.Y(_12430_),
    .A(_12166_),
    .B(net50));
 sg13g2_o21ai_1 _19363_ (.B1(_12430_),
    .Y(_00405_),
    .A1(net50),
    .A2(_12429_));
 sg13g2_nor2b_1 _19364_ (.A(net474),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12431_));
 sg13g2_a21oi_1 _19365_ (.A1(_12252_),
    .A2(net474),
    .Y(_12432_),
    .B1(_12431_));
 sg13g2_nand2_1 _19366_ (.Y(_12433_),
    .A(net482),
    .B(_12421_));
 sg13g2_o21ai_1 _19367_ (.B1(_12433_),
    .Y(_00406_),
    .A1(net50),
    .A2(_12432_));
 sg13g2_nor2b_1 _19368_ (.A(net474),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12434_));
 sg13g2_a21oi_1 _19369_ (.A1(_12257_),
    .A2(net474),
    .Y(_12435_),
    .B1(_12434_));
 sg13g2_nand2_1 _19370_ (.Y(_12436_),
    .A(net481),
    .B(_12421_));
 sg13g2_o21ai_1 _19371_ (.B1(_12436_),
    .Y(_00407_),
    .A1(net50),
    .A2(_12435_));
 sg13g2_buf_1 _19372_ (.A(net1115),
    .X(_12437_));
 sg13g2_nor2_1 _19373_ (.A(_12351_),
    .B(_12170_),
    .Y(_12438_));
 sg13g2_buf_2 _19374_ (.A(_12438_),
    .X(_12439_));
 sg13g2_nor2b_1 _19375_ (.A(_12439_),
    .B_N(\cpu.dcache.r_data[2][28] ),
    .Y(_12440_));
 sg13g2_a21oi_1 _19376_ (.A1(net1009),
    .A2(_12439_),
    .Y(_12441_),
    .B1(_12440_));
 sg13g2_nand2_1 _19377_ (.Y(_12442_),
    .A(net480),
    .B(_12421_));
 sg13g2_o21ai_1 _19378_ (.B1(_12442_),
    .Y(_00408_),
    .A1(net50),
    .A2(_12441_));
 sg13g2_buf_1 _19379_ (.A(net1112),
    .X(_12443_));
 sg13g2_nor2b_1 _19380_ (.A(_12439_),
    .B_N(\cpu.dcache.r_data[2][29] ),
    .Y(_12444_));
 sg13g2_a21oi_1 _19381_ (.A1(net1008),
    .A2(_12439_),
    .Y(_12445_),
    .B1(_12444_));
 sg13g2_nand2_1 _19382_ (.Y(_12446_),
    .A(_12123_),
    .B(_12421_));
 sg13g2_o21ai_1 _19383_ (.B1(_12446_),
    .Y(_00409_),
    .A1(net50),
    .A2(_12445_));
 sg13g2_buf_1 _19384_ (.A(net1114),
    .X(_12447_));
 sg13g2_nor2b_1 _19385_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12448_));
 sg13g2_a21oi_1 _19386_ (.A1(net1007),
    .A2(_12357_),
    .Y(_12449_),
    .B1(_12448_));
 sg13g2_nand2_1 _19387_ (.Y(_12450_),
    .A(net866),
    .B(_12354_));
 sg13g2_o21ai_1 _19388_ (.B1(_12450_),
    .Y(_00410_),
    .A1(net53),
    .A2(_12449_));
 sg13g2_nor2b_1 _19389_ (.A(_12439_),
    .B_N(\cpu.dcache.r_data[2][30] ),
    .Y(_12451_));
 sg13g2_a21oi_1 _19390_ (.A1(net1007),
    .A2(_12439_),
    .Y(_12452_),
    .B1(_12451_));
 sg13g2_nand2_1 _19391_ (.Y(_12453_),
    .A(net478),
    .B(_12421_));
 sg13g2_o21ai_1 _19392_ (.B1(_12453_),
    .Y(_00411_),
    .A1(_12422_),
    .A2(_12452_));
 sg13g2_buf_1 _19393_ (.A(net1113),
    .X(_12454_));
 sg13g2_nor2b_1 _19394_ (.A(_12439_),
    .B_N(\cpu.dcache.r_data[2][31] ),
    .Y(_12455_));
 sg13g2_a21oi_1 _19395_ (.A1(net1006),
    .A2(_12439_),
    .Y(_12456_),
    .B1(_12455_));
 sg13g2_nand2_1 _19396_ (.Y(_12457_),
    .A(_12131_),
    .B(_12421_));
 sg13g2_o21ai_1 _19397_ (.B1(_12457_),
    .Y(_00412_),
    .A1(_12422_),
    .A2(_12456_));
 sg13g2_nor2b_1 _19398_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12458_));
 sg13g2_a21oi_1 _19399_ (.A1(net1006),
    .A2(_12357_),
    .Y(_12459_),
    .B1(_12458_));
 sg13g2_nand2_1 _19400_ (.Y(_12460_),
    .A(net1016),
    .B(_12354_));
 sg13g2_o21ai_1 _19401_ (.B1(_12460_),
    .Y(_00413_),
    .A1(_12355_),
    .A2(_12459_));
 sg13g2_nor2_1 _19402_ (.A(_12351_),
    .B(_12327_),
    .Y(_12461_));
 sg13g2_buf_2 _19403_ (.A(_12461_),
    .X(_12462_));
 sg13g2_nor2b_1 _19404_ (.A(_12462_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12463_));
 sg13g2_a21oi_1 _19405_ (.A1(net1009),
    .A2(_12462_),
    .Y(_12464_),
    .B1(_12463_));
 sg13g2_nand2_1 _19406_ (.Y(_12465_),
    .A(net1015),
    .B(_12354_));
 sg13g2_o21ai_1 _19407_ (.B1(_12465_),
    .Y(_00414_),
    .A1(net53),
    .A2(_12464_));
 sg13g2_nor2b_1 _19408_ (.A(_12462_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12466_));
 sg13g2_a21oi_1 _19409_ (.A1(net1008),
    .A2(_12462_),
    .Y(_12467_),
    .B1(_12466_));
 sg13g2_nand2_1 _19410_ (.Y(_12468_),
    .A(net1011),
    .B(_12354_));
 sg13g2_o21ai_1 _19411_ (.B1(_12468_),
    .Y(_00415_),
    .A1(net53),
    .A2(_12467_));
 sg13g2_nor2b_1 _19412_ (.A(_12462_),
    .B_N(\cpu.dcache.r_data[2][6] ),
    .Y(_12469_));
 sg13g2_a21oi_1 _19413_ (.A1(net1007),
    .A2(_12462_),
    .Y(_12470_),
    .B1(_12469_));
 sg13g2_nand2_1 _19414_ (.Y(_12471_),
    .A(net1010),
    .B(_12354_));
 sg13g2_o21ai_1 _19415_ (.B1(_12471_),
    .Y(_00416_),
    .A1(net53),
    .A2(_12470_));
 sg13g2_nor2b_1 _19416_ (.A(_12462_),
    .B_N(\cpu.dcache.r_data[2][7] ),
    .Y(_12472_));
 sg13g2_a21oi_1 _19417_ (.A1(net1006),
    .A2(_12462_),
    .Y(_12473_),
    .B1(_12472_));
 sg13g2_nand2_1 _19418_ (.Y(_12474_),
    .A(net1012),
    .B(_12354_));
 sg13g2_o21ai_1 _19419_ (.B1(_12474_),
    .Y(_00417_),
    .A1(_12355_),
    .A2(_12473_));
 sg13g2_nor2b_1 _19420_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12475_));
 sg13g2_a21oi_1 _19421_ (.A1(net1009),
    .A2(_12365_),
    .Y(_12476_),
    .B1(_12475_));
 sg13g2_nand2_1 _19422_ (.Y(_12477_),
    .A(net476),
    .B(_12362_));
 sg13g2_o21ai_1 _19423_ (.B1(_12477_),
    .Y(_00418_),
    .A1(net52),
    .A2(_12476_));
 sg13g2_nor2b_1 _19424_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12478_));
 sg13g2_a21oi_1 _19425_ (.A1(_12443_),
    .A2(_12365_),
    .Y(_12479_),
    .B1(_12478_));
 sg13g2_nand2_1 _19426_ (.Y(_12480_),
    .A(net475),
    .B(_12362_));
 sg13g2_o21ai_1 _19427_ (.B1(_12480_),
    .Y(_00419_),
    .A1(net52),
    .A2(_12479_));
 sg13g2_nand2_1 _19428_ (.Y(_12481_),
    .A(net1061),
    .B(_10095_));
 sg13g2_buf_1 _19429_ (.A(_12481_),
    .X(_12482_));
 sg13g2_nor2_1 _19430_ (.A(net531),
    .B(_12191_),
    .Y(_12483_));
 sg13g2_buf_1 _19431_ (.A(_12483_),
    .X(_12484_));
 sg13g2_nor2_1 _19432_ (.A(net531),
    .B(_12065_),
    .Y(_12485_));
 sg13g2_buf_2 _19433_ (.A(_12485_),
    .X(_12486_));
 sg13g2_nor2b_1 _19434_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12487_));
 sg13g2_a21oi_1 _19435_ (.A1(net1009),
    .A2(_12486_),
    .Y(_12488_),
    .B1(_12487_));
 sg13g2_nand2_1 _19436_ (.Y(_12489_),
    .A(net868),
    .B(net62));
 sg13g2_o21ai_1 _19437_ (.B1(_12489_),
    .Y(_00420_),
    .A1(net62),
    .A2(_12488_));
 sg13g2_nor2_1 _19438_ (.A(net531),
    .B(_12204_),
    .Y(_12490_));
 sg13g2_buf_2 _19439_ (.A(_12490_),
    .X(_12491_));
 sg13g2_buf_1 _19440_ (.A(_12491_),
    .X(_12492_));
 sg13g2_nor2_1 _19441_ (.A(_12482_),
    .B(_12089_),
    .Y(_12493_));
 sg13g2_buf_2 _19442_ (.A(_12493_),
    .X(_12494_));
 sg13g2_nor2b_1 _19443_ (.A(_12494_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12495_));
 sg13g2_a21oi_1 _19444_ (.A1(net1007),
    .A2(_12494_),
    .Y(_12496_),
    .B1(_12495_));
 sg13g2_nand2_1 _19445_ (.Y(_12497_),
    .A(net482),
    .B(net49));
 sg13g2_o21ai_1 _19446_ (.B1(_12497_),
    .Y(_00421_),
    .A1(net49),
    .A2(_12496_));
 sg13g2_nor2b_1 _19447_ (.A(_12494_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12498_));
 sg13g2_a21oi_1 _19448_ (.A1(net1006),
    .A2(_12494_),
    .Y(_12499_),
    .B1(_12498_));
 sg13g2_nand2_1 _19449_ (.Y(_12500_),
    .A(net481),
    .B(net49));
 sg13g2_o21ai_1 _19450_ (.B1(_12500_),
    .Y(_00422_),
    .A1(net49),
    .A2(_12499_));
 sg13g2_nor2_1 _19451_ (.A(net531),
    .B(_12111_),
    .Y(_12501_));
 sg13g2_buf_2 _19452_ (.A(_12501_),
    .X(_12502_));
 sg13g2_nor2b_1 _19453_ (.A(_12502_),
    .B_N(\cpu.dcache.r_data[3][12] ),
    .Y(_12503_));
 sg13g2_a21oi_1 _19454_ (.A1(net1009),
    .A2(_12502_),
    .Y(_12504_),
    .B1(_12503_));
 sg13g2_nand2_1 _19455_ (.Y(_12505_),
    .A(net480),
    .B(_12491_));
 sg13g2_o21ai_1 _19456_ (.B1(_12505_),
    .Y(_00423_),
    .A1(net49),
    .A2(_12504_));
 sg13g2_nor2b_1 _19457_ (.A(_12502_),
    .B_N(\cpu.dcache.r_data[3][13] ),
    .Y(_12506_));
 sg13g2_a21oi_1 _19458_ (.A1(net1008),
    .A2(_12502_),
    .Y(_12507_),
    .B1(_12506_));
 sg13g2_nand2_1 _19459_ (.Y(_12508_),
    .A(net479),
    .B(_12491_));
 sg13g2_o21ai_1 _19460_ (.B1(_12508_),
    .Y(_00424_),
    .A1(net49),
    .A2(_12507_));
 sg13g2_nor2b_1 _19461_ (.A(_12502_),
    .B_N(\cpu.dcache.r_data[3][14] ),
    .Y(_12509_));
 sg13g2_a21oi_1 _19462_ (.A1(net1007),
    .A2(_12502_),
    .Y(_12510_),
    .B1(_12509_));
 sg13g2_nand2_1 _19463_ (.Y(_12511_),
    .A(net478),
    .B(_12491_));
 sg13g2_o21ai_1 _19464_ (.B1(_12511_),
    .Y(_00425_),
    .A1(net49),
    .A2(_12510_));
 sg13g2_nor2b_1 _19465_ (.A(_12502_),
    .B_N(\cpu.dcache.r_data[3][15] ),
    .Y(_12512_));
 sg13g2_a21oi_1 _19466_ (.A1(net1006),
    .A2(_12502_),
    .Y(_12513_),
    .B1(_12512_));
 sg13g2_nand2_1 _19467_ (.Y(_12514_),
    .A(net477),
    .B(_12491_));
 sg13g2_o21ai_1 _19468_ (.B1(_12514_),
    .Y(_00426_),
    .A1(net49),
    .A2(_12513_));
 sg13g2_nor2_1 _19469_ (.A(net531),
    .B(_12238_),
    .Y(_12515_));
 sg13g2_buf_1 _19470_ (.A(_12515_),
    .X(_12516_));
 sg13g2_nor2_1 _19471_ (.A(net531),
    .B(_12133_),
    .Y(_12517_));
 sg13g2_buf_2 _19472_ (.A(_12517_),
    .X(_12518_));
 sg13g2_nor2b_1 _19473_ (.A(_12518_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12519_));
 sg13g2_a21oi_1 _19474_ (.A1(net1009),
    .A2(_12518_),
    .Y(_12520_),
    .B1(_12519_));
 sg13g2_nand2_1 _19475_ (.Y(_12521_),
    .A(_12201_),
    .B(net61));
 sg13g2_o21ai_1 _19476_ (.B1(_12521_),
    .Y(_00427_),
    .A1(net61),
    .A2(_12520_));
 sg13g2_nor2b_1 _19477_ (.A(_12518_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12522_));
 sg13g2_a21oi_1 _19478_ (.A1(net1008),
    .A2(_12518_),
    .Y(_12523_),
    .B1(_12522_));
 sg13g2_nand2_1 _19479_ (.Y(_12524_),
    .A(net867),
    .B(net61));
 sg13g2_o21ai_1 _19480_ (.B1(_12524_),
    .Y(_00428_),
    .A1(net61),
    .A2(_12523_));
 sg13g2_nor2b_1 _19481_ (.A(_12518_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12525_));
 sg13g2_a21oi_1 _19482_ (.A1(net1007),
    .A2(_12518_),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nand2_1 _19483_ (.Y(_12527_),
    .A(net866),
    .B(_12515_));
 sg13g2_o21ai_1 _19484_ (.B1(_12527_),
    .Y(_00429_),
    .A1(_12516_),
    .A2(_12526_));
 sg13g2_nor2b_1 _19485_ (.A(_12518_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12528_));
 sg13g2_a21oi_1 _19486_ (.A1(net1006),
    .A2(_12518_),
    .Y(_12529_),
    .B1(_12528_));
 sg13g2_nand2_1 _19487_ (.Y(_12530_),
    .A(net1016),
    .B(_12515_));
 sg13g2_o21ai_1 _19488_ (.B1(_12530_),
    .Y(_00430_),
    .A1(_12516_),
    .A2(_12529_));
 sg13g2_nor2b_1 _19489_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12531_));
 sg13g2_a21oi_1 _19490_ (.A1(net1008),
    .A2(_12486_),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_nand2_1 _19491_ (.Y(_12533_),
    .A(net867),
    .B(_12484_));
 sg13g2_o21ai_1 _19492_ (.B1(_12533_),
    .Y(_00431_),
    .A1(_12484_),
    .A2(_12532_));
 sg13g2_buf_1 _19493_ (.A(net615),
    .X(_12534_));
 sg13g2_buf_1 _19494_ (.A(net530),
    .X(_12535_));
 sg13g2_nand2_2 _19495_ (.Y(_12536_),
    .A(net473),
    .B(_12145_));
 sg13g2_mux2_1 _19496_ (.A0(net1120),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12536_),
    .X(_12537_));
 sg13g2_mux2_1 _19497_ (.A0(_12537_),
    .A1(_10176_),
    .S(net61),
    .X(_00432_));
 sg13g2_mux2_1 _19498_ (.A0(net1116),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12536_),
    .X(_12538_));
 sg13g2_mux2_1 _19499_ (.A0(_12538_),
    .A1(net895),
    .S(net61),
    .X(_00433_));
 sg13g2_mux2_1 _19500_ (.A0(net1118),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12536_),
    .X(_12539_));
 sg13g2_mux2_1 _19501_ (.A0(_12539_),
    .A1(net894),
    .S(net61),
    .X(_00434_));
 sg13g2_mux2_1 _19502_ (.A0(net1117),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12536_),
    .X(_12540_));
 sg13g2_buf_1 _19503_ (.A(_10131_),
    .X(_12541_));
 sg13g2_mux2_1 _19504_ (.A0(_12540_),
    .A1(net1005),
    .S(net61),
    .X(_00435_));
 sg13g2_nor2_1 _19505_ (.A(_12482_),
    .B(_12286_),
    .Y(_12542_));
 sg13g2_buf_2 _19506_ (.A(_12542_),
    .X(_12543_));
 sg13g2_buf_1 _19507_ (.A(_12543_),
    .X(_12544_));
 sg13g2_nor2_1 _19508_ (.A(_12481_),
    .B(_12291_),
    .Y(_12545_));
 sg13g2_buf_1 _19509_ (.A(_12545_),
    .X(_12546_));
 sg13g2_nor2b_1 _19510_ (.A(net472),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12547_));
 sg13g2_a21oi_1 _19511_ (.A1(_12437_),
    .A2(net472),
    .Y(_12548_),
    .B1(_12547_));
 sg13g2_nand2_1 _19512_ (.Y(_12549_),
    .A(_12157_),
    .B(net48));
 sg13g2_o21ai_1 _19513_ (.B1(_12549_),
    .Y(_00436_),
    .A1(net48),
    .A2(_12548_));
 sg13g2_nor2b_1 _19514_ (.A(net472),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12550_));
 sg13g2_a21oi_1 _19515_ (.A1(net1008),
    .A2(net472),
    .Y(_12551_),
    .B1(_12550_));
 sg13g2_nand2_1 _19516_ (.Y(_12552_),
    .A(_12166_),
    .B(_12544_));
 sg13g2_o21ai_1 _19517_ (.B1(_12552_),
    .Y(_00437_),
    .A1(_12544_),
    .A2(_12551_));
 sg13g2_nor2b_1 _19518_ (.A(net472),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12553_));
 sg13g2_a21oi_1 _19519_ (.A1(_12447_),
    .A2(net472),
    .Y(_12554_),
    .B1(_12553_));
 sg13g2_nand2_1 _19520_ (.Y(_12555_),
    .A(_12098_),
    .B(_12543_));
 sg13g2_o21ai_1 _19521_ (.B1(_12555_),
    .Y(_00438_),
    .A1(net48),
    .A2(_12554_));
 sg13g2_nor2b_1 _19522_ (.A(net472),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12556_));
 sg13g2_a21oi_1 _19523_ (.A1(_12454_),
    .A2(net472),
    .Y(_12557_),
    .B1(_12556_));
 sg13g2_nand2_1 _19524_ (.Y(_12558_),
    .A(_12108_),
    .B(_12543_));
 sg13g2_o21ai_1 _19525_ (.B1(_12558_),
    .Y(_00439_),
    .A1(net48),
    .A2(_12557_));
 sg13g2_nor2_1 _19526_ (.A(_12481_),
    .B(_12170_),
    .Y(_12559_));
 sg13g2_buf_2 _19527_ (.A(_12559_),
    .X(_12560_));
 sg13g2_nor2b_1 _19528_ (.A(_12560_),
    .B_N(\cpu.dcache.r_data[3][28] ),
    .Y(_12561_));
 sg13g2_a21oi_1 _19529_ (.A1(net1009),
    .A2(_12560_),
    .Y(_12562_),
    .B1(_12561_));
 sg13g2_nand2_1 _19530_ (.Y(_12563_),
    .A(_12117_),
    .B(_12543_));
 sg13g2_o21ai_1 _19531_ (.B1(_12563_),
    .Y(_00440_),
    .A1(net48),
    .A2(_12562_));
 sg13g2_nor2b_1 _19532_ (.A(_12560_),
    .B_N(\cpu.dcache.r_data[3][29] ),
    .Y(_12564_));
 sg13g2_a21oi_1 _19533_ (.A1(net1008),
    .A2(_12560_),
    .Y(_12565_),
    .B1(_12564_));
 sg13g2_nand2_1 _19534_ (.Y(_12566_),
    .A(_12123_),
    .B(_12543_));
 sg13g2_o21ai_1 _19535_ (.B1(_12566_),
    .Y(_00441_),
    .A1(net48),
    .A2(_12565_));
 sg13g2_nor2b_1 _19536_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12567_));
 sg13g2_a21oi_1 _19537_ (.A1(net1007),
    .A2(_12486_),
    .Y(_12568_),
    .B1(_12567_));
 sg13g2_nand2_1 _19538_ (.Y(_12569_),
    .A(_12255_),
    .B(_12483_));
 sg13g2_o21ai_1 _19539_ (.B1(_12569_),
    .Y(_00442_),
    .A1(net62),
    .A2(_12568_));
 sg13g2_nor2b_1 _19540_ (.A(_12560_),
    .B_N(\cpu.dcache.r_data[3][30] ),
    .Y(_12570_));
 sg13g2_a21oi_1 _19541_ (.A1(_12447_),
    .A2(_12560_),
    .Y(_12571_),
    .B1(_12570_));
 sg13g2_nand2_1 _19542_ (.Y(_12572_),
    .A(net478),
    .B(_12543_));
 sg13g2_o21ai_1 _19543_ (.B1(_12572_),
    .Y(_00443_),
    .A1(net48),
    .A2(_12571_));
 sg13g2_nor2b_1 _19544_ (.A(_12560_),
    .B_N(\cpu.dcache.r_data[3][31] ),
    .Y(_12573_));
 sg13g2_a21oi_1 _19545_ (.A1(_12454_),
    .A2(_12560_),
    .Y(_12574_),
    .B1(_12573_));
 sg13g2_nand2_1 _19546_ (.Y(_12575_),
    .A(net477),
    .B(_12543_));
 sg13g2_o21ai_1 _19547_ (.B1(_12575_),
    .Y(_00444_),
    .A1(net48),
    .A2(_12574_));
 sg13g2_nor2b_1 _19548_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12576_));
 sg13g2_a21oi_1 _19549_ (.A1(net1006),
    .A2(_12486_),
    .Y(_12577_),
    .B1(_12576_));
 sg13g2_nand2_1 _19550_ (.Y(_12578_),
    .A(_12260_),
    .B(_12483_));
 sg13g2_o21ai_1 _19551_ (.B1(_12578_),
    .Y(_00445_),
    .A1(net62),
    .A2(_12577_));
 sg13g2_nand2_2 _19552_ (.Y(_12579_),
    .A(net473),
    .B(_12179_));
 sg13g2_mux2_1 _19553_ (.A0(net1115),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12579_),
    .X(_12580_));
 sg13g2_buf_1 _19554_ (.A(net1053),
    .X(_12581_));
 sg13g2_mux2_1 _19555_ (.A0(_12580_),
    .A1(net865),
    .S(net62),
    .X(_00446_));
 sg13g2_mux2_1 _19556_ (.A0(net1112),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12579_),
    .X(_12582_));
 sg13g2_mux2_1 _19557_ (.A0(_12582_),
    .A1(net895),
    .S(net62),
    .X(_00447_));
 sg13g2_mux2_1 _19558_ (.A0(net1114),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12579_),
    .X(_12583_));
 sg13g2_mux2_1 _19559_ (.A0(_12583_),
    .A1(net894),
    .S(net62),
    .X(_00448_));
 sg13g2_mux2_1 _19560_ (.A0(net1113),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12579_),
    .X(_12584_));
 sg13g2_mux2_1 _19561_ (.A0(_12584_),
    .A1(net1005),
    .S(net62),
    .X(_00449_));
 sg13g2_nor2b_1 _19562_ (.A(_12494_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12585_));
 sg13g2_a21oi_1 _19563_ (.A1(_12437_),
    .A2(_12494_),
    .Y(_12586_),
    .B1(_12585_));
 sg13g2_nand2_1 _19564_ (.Y(_12587_),
    .A(net476),
    .B(_12491_));
 sg13g2_o21ai_1 _19565_ (.B1(_12587_),
    .Y(_00450_),
    .A1(_12492_),
    .A2(_12586_));
 sg13g2_nor2b_1 _19566_ (.A(_12494_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12588_));
 sg13g2_a21oi_1 _19567_ (.A1(_12443_),
    .A2(_12494_),
    .Y(_12589_),
    .B1(_12588_));
 sg13g2_nand2_1 _19568_ (.Y(_12590_),
    .A(net475),
    .B(_12491_));
 sg13g2_o21ai_1 _19569_ (.B1(_12590_),
    .Y(_00451_),
    .A1(_12492_),
    .A2(_12589_));
 sg13g2_buf_1 _19570_ (.A(_10140_),
    .X(_12591_));
 sg13g2_nor2_1 _19571_ (.A(net594),
    .B(_12191_),
    .Y(_12592_));
 sg13g2_buf_2 _19572_ (.A(_12592_),
    .X(_12593_));
 sg13g2_buf_1 _19573_ (.A(_12593_),
    .X(_12594_));
 sg13g2_nor2_1 _19574_ (.A(net594),
    .B(_12065_),
    .Y(_12595_));
 sg13g2_buf_2 _19575_ (.A(_12595_),
    .X(_12596_));
 sg13g2_nor2b_1 _19576_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12597_));
 sg13g2_a21oi_1 _19577_ (.A1(net1009),
    .A2(_12596_),
    .Y(_12598_),
    .B1(_12597_));
 sg13g2_nand2_1 _19578_ (.Y(_12599_),
    .A(net868),
    .B(net47));
 sg13g2_o21ai_1 _19579_ (.B1(_12599_),
    .Y(_00452_),
    .A1(net47),
    .A2(_12598_));
 sg13g2_or2_1 _19580_ (.X(_12600_),
    .B(_12204_),
    .A(_10140_));
 sg13g2_buf_1 _19581_ (.A(_12600_),
    .X(_12601_));
 sg13g2_buf_1 _19582_ (.A(_12601_),
    .X(_12602_));
 sg13g2_nor2_1 _19583_ (.A(net594),
    .B(_12089_),
    .Y(_12603_));
 sg13g2_buf_2 _19584_ (.A(_12603_),
    .X(_12604_));
 sg13g2_nor2b_1 _19585_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12605_));
 sg13g2_a21oi_1 _19586_ (.A1(net1023),
    .A2(_12604_),
    .Y(_12606_),
    .B1(_12605_));
 sg13g2_nor2_1 _19587_ (.A(_12097_),
    .B(net46),
    .Y(_12607_));
 sg13g2_a21oi_1 _19588_ (.A1(net46),
    .A2(_12606_),
    .Y(_00453_),
    .B1(_12607_));
 sg13g2_nor2b_1 _19589_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12608_));
 sg13g2_a21oi_1 _19590_ (.A1(net1022),
    .A2(_12604_),
    .Y(_12609_),
    .B1(_12608_));
 sg13g2_nor2_1 _19591_ (.A(_12107_),
    .B(net46),
    .Y(_12610_));
 sg13g2_a21oi_1 _19592_ (.A1(net46),
    .A2(_12609_),
    .Y(_00454_),
    .B1(_12610_));
 sg13g2_nor2_1 _19593_ (.A(net594),
    .B(_12111_),
    .Y(_12611_));
 sg13g2_buf_2 _19594_ (.A(_12611_),
    .X(_12612_));
 sg13g2_nor2b_1 _19595_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][12] ),
    .Y(_12613_));
 sg13g2_a21oi_1 _19596_ (.A1(net1021),
    .A2(_12612_),
    .Y(_12614_),
    .B1(_12613_));
 sg13g2_nor2_1 _19597_ (.A(_12116_),
    .B(_12601_),
    .Y(_12615_));
 sg13g2_a21oi_1 _19598_ (.A1(net46),
    .A2(_12614_),
    .Y(_00455_),
    .B1(_12615_));
 sg13g2_nor2b_1 _19599_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][13] ),
    .Y(_12616_));
 sg13g2_a21oi_1 _19600_ (.A1(net1020),
    .A2(_12612_),
    .Y(_12617_),
    .B1(_12616_));
 sg13g2_nor2_1 _19601_ (.A(_12122_),
    .B(_12601_),
    .Y(_12618_));
 sg13g2_a21oi_1 _19602_ (.A1(_12602_),
    .A2(_12617_),
    .Y(_00456_),
    .B1(_12618_));
 sg13g2_nor2b_1 _19603_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][14] ),
    .Y(_12619_));
 sg13g2_a21oi_1 _19604_ (.A1(net1023),
    .A2(_12612_),
    .Y(_12620_),
    .B1(_12619_));
 sg13g2_nor2_1 _19605_ (.A(_12126_),
    .B(_12601_),
    .Y(_12621_));
 sg13g2_a21oi_1 _19606_ (.A1(net46),
    .A2(_12620_),
    .Y(_00457_),
    .B1(_12621_));
 sg13g2_nor2b_1 _19607_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][15] ),
    .Y(_12622_));
 sg13g2_a21oi_1 _19608_ (.A1(net1022),
    .A2(_12612_),
    .Y(_12623_),
    .B1(_12622_));
 sg13g2_nor2_1 _19609_ (.A(_12130_),
    .B(_12601_),
    .Y(_12624_));
 sg13g2_a21oi_1 _19610_ (.A1(_12602_),
    .A2(_12623_),
    .Y(_00458_),
    .B1(_12624_));
 sg13g2_nor2_1 _19611_ (.A(net594),
    .B(_12238_),
    .Y(_12625_));
 sg13g2_buf_2 _19612_ (.A(_12625_),
    .X(_12626_));
 sg13g2_buf_1 _19613_ (.A(_12626_),
    .X(_12627_));
 sg13g2_buf_1 _19614_ (.A(net1115),
    .X(_12628_));
 sg13g2_nor2_1 _19615_ (.A(net594),
    .B(_12133_),
    .Y(_12629_));
 sg13g2_buf_2 _19616_ (.A(_12629_),
    .X(_12630_));
 sg13g2_nor2b_1 _19617_ (.A(_12630_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12631_));
 sg13g2_a21oi_1 _19618_ (.A1(net1004),
    .A2(_12630_),
    .Y(_12632_),
    .B1(_12631_));
 sg13g2_nand2_1 _19619_ (.Y(_12633_),
    .A(_12201_),
    .B(_12627_));
 sg13g2_o21ai_1 _19620_ (.B1(_12633_),
    .Y(_00459_),
    .A1(net45),
    .A2(_12632_));
 sg13g2_nor2b_1 _19621_ (.A(_12630_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12634_));
 sg13g2_a21oi_1 _19622_ (.A1(net1008),
    .A2(_12630_),
    .Y(_12635_),
    .B1(_12634_));
 sg13g2_nand2_1 _19623_ (.Y(_12636_),
    .A(_12250_),
    .B(net45));
 sg13g2_o21ai_1 _19624_ (.B1(_12636_),
    .Y(_00460_),
    .A1(_12627_),
    .A2(_12635_));
 sg13g2_nor2b_1 _19625_ (.A(_12630_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12637_));
 sg13g2_a21oi_1 _19626_ (.A1(net1007),
    .A2(_12630_),
    .Y(_12638_),
    .B1(_12637_));
 sg13g2_nand2_1 _19627_ (.Y(_12639_),
    .A(_12255_),
    .B(_12626_));
 sg13g2_o21ai_1 _19628_ (.B1(_12639_),
    .Y(_00461_),
    .A1(net45),
    .A2(_12638_));
 sg13g2_nor2b_1 _19629_ (.A(_12630_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12640_));
 sg13g2_a21oi_1 _19630_ (.A1(net1006),
    .A2(_12630_),
    .Y(_12641_),
    .B1(_12640_));
 sg13g2_nand2_1 _19631_ (.Y(_12642_),
    .A(_12260_),
    .B(_12626_));
 sg13g2_o21ai_1 _19632_ (.B1(_12642_),
    .Y(_00462_),
    .A1(net45),
    .A2(_12641_));
 sg13g2_buf_1 _19633_ (.A(net1112),
    .X(_12643_));
 sg13g2_nor2b_1 _19634_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12644_));
 sg13g2_a21oi_1 _19635_ (.A1(net1003),
    .A2(_12596_),
    .Y(_12645_),
    .B1(_12644_));
 sg13g2_nand2_1 _19636_ (.Y(_12646_),
    .A(net867),
    .B(net47));
 sg13g2_o21ai_1 _19637_ (.B1(_12646_),
    .Y(_00463_),
    .A1(net47),
    .A2(_12645_));
 sg13g2_nor2_1 _19638_ (.A(net594),
    .B(_12266_),
    .Y(_12647_));
 sg13g2_buf_2 _19639_ (.A(_12647_),
    .X(_12648_));
 sg13g2_nor2b_1 _19640_ (.A(_12648_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12649_));
 sg13g2_a21oi_1 _19641_ (.A1(net1004),
    .A2(_12648_),
    .Y(_12650_),
    .B1(_12649_));
 sg13g2_nand2_1 _19642_ (.Y(_12651_),
    .A(net1015),
    .B(_12626_));
 sg13g2_o21ai_1 _19643_ (.B1(_12651_),
    .Y(_00464_),
    .A1(net45),
    .A2(_12650_));
 sg13g2_nor2b_1 _19644_ (.A(_12648_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12652_));
 sg13g2_a21oi_1 _19645_ (.A1(net1003),
    .A2(_12648_),
    .Y(_12653_),
    .B1(_12652_));
 sg13g2_nand2_1 _19646_ (.Y(_12654_),
    .A(_12335_),
    .B(_12626_));
 sg13g2_o21ai_1 _19647_ (.B1(_12654_),
    .Y(_00465_),
    .A1(net45),
    .A2(_12653_));
 sg13g2_buf_1 _19648_ (.A(net1114),
    .X(_12655_));
 sg13g2_nor2b_1 _19649_ (.A(_12648_),
    .B_N(\cpu.dcache.r_data[4][22] ),
    .Y(_12656_));
 sg13g2_a21oi_1 _19650_ (.A1(net1002),
    .A2(_12648_),
    .Y(_12657_),
    .B1(_12656_));
 sg13g2_nand2_1 _19651_ (.Y(_12658_),
    .A(_12339_),
    .B(_12626_));
 sg13g2_o21ai_1 _19652_ (.B1(_12658_),
    .Y(_00466_),
    .A1(net45),
    .A2(_12657_));
 sg13g2_buf_1 _19653_ (.A(net1113),
    .X(_12659_));
 sg13g2_nor2b_1 _19654_ (.A(_12648_),
    .B_N(\cpu.dcache.r_data[4][23] ),
    .Y(_12660_));
 sg13g2_a21oi_1 _19655_ (.A1(net1001),
    .A2(_12648_),
    .Y(_12661_),
    .B1(_12660_));
 sg13g2_nand2_1 _19656_ (.Y(_12662_),
    .A(net1012),
    .B(_12626_));
 sg13g2_o21ai_1 _19657_ (.B1(_12662_),
    .Y(_00467_),
    .A1(net45),
    .A2(_12661_));
 sg13g2_buf_1 _19658_ (.A(net617),
    .X(_12663_));
 sg13g2_buf_1 _19659_ (.A(net529),
    .X(_12664_));
 sg13g2_buf_1 _19660_ (.A(net471),
    .X(_12665_));
 sg13g2_nand2_1 _19661_ (.Y(_12666_),
    .A(net424),
    .B(_12074_));
 sg13g2_buf_1 _19662_ (.A(_12666_),
    .X(_12667_));
 sg13g2_mux2_1 _19663_ (.A0(net1115),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net335),
    .X(_12668_));
 sg13g2_or2_1 _19664_ (.X(_12669_),
    .B(_12286_),
    .A(_12591_));
 sg13g2_buf_1 _19665_ (.A(_12669_),
    .X(_12670_));
 sg13g2_buf_1 _19666_ (.A(_12670_),
    .X(_12671_));
 sg13g2_mux2_1 _19667_ (.A0(net476),
    .A1(_12668_),
    .S(net44),
    .X(_00468_));
 sg13g2_mux2_1 _19668_ (.A0(net1112),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net335),
    .X(_12672_));
 sg13g2_mux2_1 _19669_ (.A0(net475),
    .A1(_12672_),
    .S(net44),
    .X(_00469_));
 sg13g2_mux2_1 _19670_ (.A0(net1114),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net335),
    .X(_12673_));
 sg13g2_mux2_1 _19671_ (.A0(net482),
    .A1(_12673_),
    .S(net44),
    .X(_00470_));
 sg13g2_mux2_1 _19672_ (.A0(net1113),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(net335),
    .X(_12674_));
 sg13g2_mux2_1 _19673_ (.A0(net481),
    .A1(_12674_),
    .S(net44),
    .X(_00471_));
 sg13g2_nor2_1 _19674_ (.A(_12591_),
    .B(_12170_),
    .Y(_12675_));
 sg13g2_buf_2 _19675_ (.A(_12675_),
    .X(_12676_));
 sg13g2_nor2b_1 _19676_ (.A(_12676_),
    .B_N(\cpu.dcache.r_data[4][28] ),
    .Y(_12677_));
 sg13g2_a21oi_1 _19677_ (.A1(net1021),
    .A2(_12676_),
    .Y(_12678_),
    .B1(_12677_));
 sg13g2_nor2_1 _19678_ (.A(_12116_),
    .B(net44),
    .Y(_12679_));
 sg13g2_a21oi_1 _19679_ (.A1(net44),
    .A2(_12678_),
    .Y(_00472_),
    .B1(_12679_));
 sg13g2_nor2b_1 _19680_ (.A(_12676_),
    .B_N(\cpu.dcache.r_data[4][29] ),
    .Y(_12680_));
 sg13g2_a21oi_1 _19681_ (.A1(net1020),
    .A2(_12676_),
    .Y(_12681_),
    .B1(_12680_));
 sg13g2_nor2_1 _19682_ (.A(_12122_),
    .B(net44),
    .Y(_12682_));
 sg13g2_a21oi_1 _19683_ (.A1(net44),
    .A2(_12681_),
    .Y(_00473_),
    .B1(_12682_));
 sg13g2_nor2b_1 _19684_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12683_));
 sg13g2_a21oi_1 _19685_ (.A1(net1002),
    .A2(_12596_),
    .Y(_12684_),
    .B1(_12683_));
 sg13g2_nand2_1 _19686_ (.Y(_12685_),
    .A(net866),
    .B(_12593_));
 sg13g2_o21ai_1 _19687_ (.B1(_12685_),
    .Y(_00474_),
    .A1(_12594_),
    .A2(_12684_));
 sg13g2_nor2b_1 _19688_ (.A(_12676_),
    .B_N(\cpu.dcache.r_data[4][30] ),
    .Y(_12686_));
 sg13g2_a21oi_1 _19689_ (.A1(_12252_),
    .A2(_12676_),
    .Y(_12687_),
    .B1(_12686_));
 sg13g2_nor2_1 _19690_ (.A(_12126_),
    .B(_12670_),
    .Y(_12688_));
 sg13g2_a21oi_1 _19691_ (.A1(_12671_),
    .A2(_12687_),
    .Y(_00475_),
    .B1(_12688_));
 sg13g2_nor2b_1 _19692_ (.A(_12676_),
    .B_N(\cpu.dcache.r_data[4][31] ),
    .Y(_12689_));
 sg13g2_a21oi_1 _19693_ (.A1(_12257_),
    .A2(_12676_),
    .Y(_12690_),
    .B1(_12689_));
 sg13g2_nor2_1 _19694_ (.A(_12130_),
    .B(_12670_),
    .Y(_12691_));
 sg13g2_a21oi_1 _19695_ (.A1(_12671_),
    .A2(_12690_),
    .Y(_00476_),
    .B1(_12691_));
 sg13g2_nor2b_1 _19696_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12692_));
 sg13g2_a21oi_1 _19697_ (.A1(net1001),
    .A2(_12596_),
    .Y(_12693_),
    .B1(_12692_));
 sg13g2_buf_1 _19698_ (.A(_10110_),
    .X(_12694_));
 sg13g2_nand2_1 _19699_ (.Y(_12695_),
    .A(_12694_),
    .B(_12593_));
 sg13g2_o21ai_1 _19700_ (.B1(_12695_),
    .Y(_00477_),
    .A1(net47),
    .A2(_12693_));
 sg13g2_nor2_1 _19701_ (.A(_10140_),
    .B(_12327_),
    .Y(_12696_));
 sg13g2_buf_2 _19702_ (.A(_12696_),
    .X(_12697_));
 sg13g2_nor2b_1 _19703_ (.A(_12697_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12698_));
 sg13g2_a21oi_1 _19704_ (.A1(net1004),
    .A2(_12697_),
    .Y(_12699_),
    .B1(_12698_));
 sg13g2_nand2_1 _19705_ (.Y(_12700_),
    .A(net1015),
    .B(_12593_));
 sg13g2_o21ai_1 _19706_ (.B1(_12700_),
    .Y(_00478_),
    .A1(net47),
    .A2(_12699_));
 sg13g2_nor2b_1 _19707_ (.A(_12697_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12701_));
 sg13g2_a21oi_1 _19708_ (.A1(net1003),
    .A2(_12697_),
    .Y(_12702_),
    .B1(_12701_));
 sg13g2_nand2_1 _19709_ (.Y(_12703_),
    .A(net1011),
    .B(_12593_));
 sg13g2_o21ai_1 _19710_ (.B1(_12703_),
    .Y(_00479_),
    .A1(net47),
    .A2(_12702_));
 sg13g2_nor2b_1 _19711_ (.A(_12697_),
    .B_N(\cpu.dcache.r_data[4][6] ),
    .Y(_12704_));
 sg13g2_a21oi_1 _19712_ (.A1(net1002),
    .A2(_12697_),
    .Y(_12705_),
    .B1(_12704_));
 sg13g2_nand2_1 _19713_ (.Y(_12706_),
    .A(net1010),
    .B(_12593_));
 sg13g2_o21ai_1 _19714_ (.B1(_12706_),
    .Y(_00480_),
    .A1(net47),
    .A2(_12705_));
 sg13g2_nor2b_1 _19715_ (.A(_12697_),
    .B_N(\cpu.dcache.r_data[4][7] ),
    .Y(_12707_));
 sg13g2_a21oi_1 _19716_ (.A1(net1001),
    .A2(_12697_),
    .Y(_12708_),
    .B1(_12707_));
 sg13g2_nand2_1 _19717_ (.Y(_12709_),
    .A(net1012),
    .B(_12593_));
 sg13g2_o21ai_1 _19718_ (.B1(_12709_),
    .Y(_00481_),
    .A1(_12594_),
    .A2(_12708_));
 sg13g2_nor2b_1 _19719_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12710_));
 sg13g2_a21oi_1 _19720_ (.A1(_12196_),
    .A2(_12604_),
    .Y(_12711_),
    .B1(_12710_));
 sg13g2_nor2_1 _19721_ (.A(_12156_),
    .B(_12601_),
    .Y(_12712_));
 sg13g2_a21oi_1 _19722_ (.A1(net46),
    .A2(_12711_),
    .Y(_00482_),
    .B1(_12712_));
 sg13g2_nor2b_1 _19723_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12713_));
 sg13g2_a21oi_1 _19724_ (.A1(_12247_),
    .A2(_12604_),
    .Y(_12714_),
    .B1(_12713_));
 sg13g2_nor2_1 _19725_ (.A(_12165_),
    .B(_12601_),
    .Y(_12715_));
 sg13g2_a21oi_1 _19726_ (.A1(net46),
    .A2(_12714_),
    .Y(_00483_),
    .B1(_12715_));
 sg13g2_or2_1 _19727_ (.X(_12716_),
    .B(_09463_),
    .A(net785));
 sg13g2_buf_2 _19728_ (.A(_12716_),
    .X(_12717_));
 sg13g2_buf_1 _19729_ (.A(_12717_),
    .X(_12718_));
 sg13g2_nor2_1 _19730_ (.A(net528),
    .B(_12191_),
    .Y(_12719_));
 sg13g2_buf_2 _19731_ (.A(_12719_),
    .X(_12720_));
 sg13g2_buf_1 _19732_ (.A(_12720_),
    .X(_12721_));
 sg13g2_nor2_1 _19733_ (.A(net528),
    .B(_12065_),
    .Y(_12722_));
 sg13g2_buf_2 _19734_ (.A(_12722_),
    .X(_12723_));
 sg13g2_nor2b_1 _19735_ (.A(_12723_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12724_));
 sg13g2_a21oi_1 _19736_ (.A1(net1004),
    .A2(_12723_),
    .Y(_12725_),
    .B1(_12724_));
 sg13g2_nand2_1 _19737_ (.Y(_12726_),
    .A(net901),
    .B(net43));
 sg13g2_o21ai_1 _19738_ (.B1(_12726_),
    .Y(_00484_),
    .A1(net43),
    .A2(_12725_));
 sg13g2_nor2_1 _19739_ (.A(_12718_),
    .B(_12204_),
    .Y(_12727_));
 sg13g2_buf_2 _19740_ (.A(_12727_),
    .X(_12728_));
 sg13g2_buf_1 _19741_ (.A(_12728_),
    .X(_12729_));
 sg13g2_nor2_1 _19742_ (.A(net528),
    .B(_12089_),
    .Y(_12730_));
 sg13g2_buf_2 _19743_ (.A(_12730_),
    .X(_12731_));
 sg13g2_nor2b_1 _19744_ (.A(_12731_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12732_));
 sg13g2_a21oi_1 _19745_ (.A1(net1002),
    .A2(_12731_),
    .Y(_12733_),
    .B1(_12732_));
 sg13g2_nand2_1 _19746_ (.Y(_12734_),
    .A(net482),
    .B(net42));
 sg13g2_o21ai_1 _19747_ (.B1(_12734_),
    .Y(_00485_),
    .A1(net42),
    .A2(_12733_));
 sg13g2_nor2b_1 _19748_ (.A(_12731_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12735_));
 sg13g2_a21oi_1 _19749_ (.A1(net1001),
    .A2(_12731_),
    .Y(_12736_),
    .B1(_12735_));
 sg13g2_nand2_1 _19750_ (.Y(_12737_),
    .A(net481),
    .B(net42));
 sg13g2_o21ai_1 _19751_ (.B1(_12737_),
    .Y(_00486_),
    .A1(net42),
    .A2(_12736_));
 sg13g2_nor2_1 _19752_ (.A(net528),
    .B(_12111_),
    .Y(_12738_));
 sg13g2_buf_2 _19753_ (.A(_12738_),
    .X(_12739_));
 sg13g2_nor2b_1 _19754_ (.A(_12739_),
    .B_N(\cpu.dcache.r_data[5][12] ),
    .Y(_12740_));
 sg13g2_a21oi_1 _19755_ (.A1(net1004),
    .A2(_12739_),
    .Y(_12741_),
    .B1(_12740_));
 sg13g2_nand2_1 _19756_ (.Y(_12742_),
    .A(net480),
    .B(_12728_));
 sg13g2_o21ai_1 _19757_ (.B1(_12742_),
    .Y(_00487_),
    .A1(net42),
    .A2(_12741_));
 sg13g2_nor2b_1 _19758_ (.A(_12739_),
    .B_N(\cpu.dcache.r_data[5][13] ),
    .Y(_12743_));
 sg13g2_a21oi_1 _19759_ (.A1(net1003),
    .A2(_12739_),
    .Y(_12744_),
    .B1(_12743_));
 sg13g2_nand2_1 _19760_ (.Y(_12745_),
    .A(net479),
    .B(_12728_));
 sg13g2_o21ai_1 _19761_ (.B1(_12745_),
    .Y(_00488_),
    .A1(_12729_),
    .A2(_12744_));
 sg13g2_nor2b_1 _19762_ (.A(_12739_),
    .B_N(\cpu.dcache.r_data[5][14] ),
    .Y(_12746_));
 sg13g2_a21oi_1 _19763_ (.A1(_12655_),
    .A2(_12739_),
    .Y(_12747_),
    .B1(_12746_));
 sg13g2_nand2_1 _19764_ (.Y(_12748_),
    .A(net478),
    .B(_12728_));
 sg13g2_o21ai_1 _19765_ (.B1(_12748_),
    .Y(_00489_),
    .A1(_12729_),
    .A2(_12747_));
 sg13g2_nor2b_1 _19766_ (.A(_12739_),
    .B_N(\cpu.dcache.r_data[5][15] ),
    .Y(_12749_));
 sg13g2_a21oi_1 _19767_ (.A1(_12659_),
    .A2(_12739_),
    .Y(_12750_),
    .B1(_12749_));
 sg13g2_nand2_1 _19768_ (.Y(_12751_),
    .A(net477),
    .B(_12728_));
 sg13g2_o21ai_1 _19769_ (.B1(_12751_),
    .Y(_00490_),
    .A1(net42),
    .A2(_12750_));
 sg13g2_nor2_1 _19770_ (.A(net528),
    .B(_12238_),
    .Y(_12752_));
 sg13g2_buf_2 _19771_ (.A(_12752_),
    .X(_12753_));
 sg13g2_buf_1 _19772_ (.A(_12753_),
    .X(_12754_));
 sg13g2_nor2_1 _19773_ (.A(net528),
    .B(_12133_),
    .Y(_12755_));
 sg13g2_buf_2 _19774_ (.A(_12755_),
    .X(_12756_));
 sg13g2_nor2b_1 _19775_ (.A(_12756_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12757_));
 sg13g2_a21oi_1 _19776_ (.A1(net1004),
    .A2(_12756_),
    .Y(_12758_),
    .B1(_12757_));
 sg13g2_nand2_1 _19777_ (.Y(_12759_),
    .A(net901),
    .B(net41));
 sg13g2_o21ai_1 _19778_ (.B1(_12759_),
    .Y(_00491_),
    .A1(net41),
    .A2(_12758_));
 sg13g2_nor2b_1 _19779_ (.A(_12756_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12760_));
 sg13g2_a21oi_1 _19780_ (.A1(net1003),
    .A2(_12756_),
    .Y(_12761_),
    .B1(_12760_));
 sg13g2_buf_1 _19781_ (.A(_10087_),
    .X(_12762_));
 sg13g2_nand2_1 _19782_ (.Y(_12763_),
    .A(net999),
    .B(_12754_));
 sg13g2_o21ai_1 _19783_ (.B1(_12763_),
    .Y(_00492_),
    .A1(_12754_),
    .A2(_12761_));
 sg13g2_nor2b_1 _19784_ (.A(_12756_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12764_));
 sg13g2_a21oi_1 _19785_ (.A1(net1002),
    .A2(_12756_),
    .Y(_12765_),
    .B1(_12764_));
 sg13g2_buf_1 _19786_ (.A(net1048),
    .X(_12766_));
 sg13g2_nand2_1 _19787_ (.Y(_12767_),
    .A(net864),
    .B(_12753_));
 sg13g2_o21ai_1 _19788_ (.B1(_12767_),
    .Y(_00493_),
    .A1(net41),
    .A2(_12765_));
 sg13g2_nor2b_1 _19789_ (.A(_12756_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_12768_));
 sg13g2_a21oi_1 _19790_ (.A1(net1001),
    .A2(_12756_),
    .Y(_12769_),
    .B1(_12768_));
 sg13g2_nand2_1 _19791_ (.Y(_12770_),
    .A(net1000),
    .B(_12753_));
 sg13g2_o21ai_1 _19792_ (.B1(_12770_),
    .Y(_00494_),
    .A1(net41),
    .A2(_12769_));
 sg13g2_nor2b_1 _19793_ (.A(_12723_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12771_));
 sg13g2_a21oi_1 _19794_ (.A1(net1003),
    .A2(_12723_),
    .Y(_02686_),
    .B1(_12771_));
 sg13g2_nand2_1 _19795_ (.Y(_02687_),
    .A(net999),
    .B(net43));
 sg13g2_o21ai_1 _19796_ (.B1(_02687_),
    .Y(_00495_),
    .A1(net43),
    .A2(_02686_));
 sg13g2_nor2_1 _19797_ (.A(_12717_),
    .B(_12266_),
    .Y(_02688_));
 sg13g2_buf_2 _19798_ (.A(_02688_),
    .X(_02689_));
 sg13g2_nor2b_1 _19799_ (.A(_02689_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_02690_));
 sg13g2_a21oi_1 _19800_ (.A1(net1004),
    .A2(_02689_),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_nand2_1 _19801_ (.Y(_02692_),
    .A(_12271_),
    .B(_12753_));
 sg13g2_o21ai_1 _19802_ (.B1(_02692_),
    .Y(_00496_),
    .A1(net41),
    .A2(_02691_));
 sg13g2_nor2b_1 _19803_ (.A(_02689_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_02693_));
 sg13g2_a21oi_1 _19804_ (.A1(net1003),
    .A2(_02689_),
    .Y(_02694_),
    .B1(_02693_));
 sg13g2_nand2_1 _19805_ (.Y(_02695_),
    .A(_12335_),
    .B(_12753_));
 sg13g2_o21ai_1 _19806_ (.B1(_02695_),
    .Y(_00497_),
    .A1(net41),
    .A2(_02694_));
 sg13g2_nor2b_1 _19807_ (.A(_02689_),
    .B_N(\cpu.dcache.r_data[5][22] ),
    .Y(_02696_));
 sg13g2_a21oi_1 _19808_ (.A1(net1002),
    .A2(_02689_),
    .Y(_02697_),
    .B1(_02696_));
 sg13g2_nand2_1 _19809_ (.Y(_02698_),
    .A(_12339_),
    .B(_12753_));
 sg13g2_o21ai_1 _19810_ (.B1(_02698_),
    .Y(_00498_),
    .A1(net41),
    .A2(_02697_));
 sg13g2_nor2b_1 _19811_ (.A(_02689_),
    .B_N(\cpu.dcache.r_data[5][23] ),
    .Y(_02699_));
 sg13g2_a21oi_1 _19812_ (.A1(net1001),
    .A2(_02689_),
    .Y(_02700_),
    .B1(_02699_));
 sg13g2_nand2_1 _19813_ (.Y(_02701_),
    .A(_12283_),
    .B(_12753_));
 sg13g2_o21ai_1 _19814_ (.B1(_02701_),
    .Y(_00499_),
    .A1(net41),
    .A2(_02700_));
 sg13g2_nor2_1 _19815_ (.A(net528),
    .B(_12286_),
    .Y(_02702_));
 sg13g2_buf_2 _19816_ (.A(_02702_),
    .X(_02703_));
 sg13g2_buf_1 _19817_ (.A(_02703_),
    .X(_02704_));
 sg13g2_nor2_1 _19818_ (.A(_12717_),
    .B(_12291_),
    .Y(_02705_));
 sg13g2_buf_1 _19819_ (.A(_02705_),
    .X(_02706_));
 sg13g2_nor2b_1 _19820_ (.A(net470),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_02707_));
 sg13g2_a21oi_1 _19821_ (.A1(_12628_),
    .A2(net470),
    .Y(_02708_),
    .B1(_02707_));
 sg13g2_nand2_1 _19822_ (.Y(_02709_),
    .A(net476),
    .B(net40));
 sg13g2_o21ai_1 _19823_ (.B1(_02709_),
    .Y(_00500_),
    .A1(net40),
    .A2(_02708_));
 sg13g2_nor2b_1 _19824_ (.A(net470),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_02710_));
 sg13g2_a21oi_1 _19825_ (.A1(_12643_),
    .A2(net470),
    .Y(_02711_),
    .B1(_02710_));
 sg13g2_nand2_1 _19826_ (.Y(_02712_),
    .A(net475),
    .B(net40));
 sg13g2_o21ai_1 _19827_ (.B1(_02712_),
    .Y(_00501_),
    .A1(net40),
    .A2(_02711_));
 sg13g2_nor2b_1 _19828_ (.A(net470),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_02713_));
 sg13g2_a21oi_1 _19829_ (.A1(_12655_),
    .A2(net470),
    .Y(_02714_),
    .B1(_02713_));
 sg13g2_nand2_1 _19830_ (.Y(_02715_),
    .A(net482),
    .B(_02703_));
 sg13g2_o21ai_1 _19831_ (.B1(_02715_),
    .Y(_00502_),
    .A1(net40),
    .A2(_02714_));
 sg13g2_nor2b_1 _19832_ (.A(net470),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_02716_));
 sg13g2_a21oi_1 _19833_ (.A1(_12659_),
    .A2(net470),
    .Y(_02717_),
    .B1(_02716_));
 sg13g2_nand2_1 _19834_ (.Y(_02718_),
    .A(net481),
    .B(_02703_));
 sg13g2_o21ai_1 _19835_ (.B1(_02718_),
    .Y(_00503_),
    .A1(net40),
    .A2(_02717_));
 sg13g2_nor2_1 _19836_ (.A(_12717_),
    .B(_12170_),
    .Y(_02719_));
 sg13g2_buf_2 _19837_ (.A(_02719_),
    .X(_02720_));
 sg13g2_nor2b_1 _19838_ (.A(_02720_),
    .B_N(\cpu.dcache.r_data[5][28] ),
    .Y(_02721_));
 sg13g2_a21oi_1 _19839_ (.A1(_12628_),
    .A2(_02720_),
    .Y(_02722_),
    .B1(_02721_));
 sg13g2_nand2_1 _19840_ (.Y(_02723_),
    .A(net480),
    .B(_02703_));
 sg13g2_o21ai_1 _19841_ (.B1(_02723_),
    .Y(_00504_),
    .A1(net40),
    .A2(_02722_));
 sg13g2_nor2b_1 _19842_ (.A(_02720_),
    .B_N(\cpu.dcache.r_data[5][29] ),
    .Y(_02724_));
 sg13g2_a21oi_1 _19843_ (.A1(_12643_),
    .A2(_02720_),
    .Y(_02725_),
    .B1(_02724_));
 sg13g2_nand2_1 _19844_ (.Y(_02726_),
    .A(net479),
    .B(_02703_));
 sg13g2_o21ai_1 _19845_ (.B1(_02726_),
    .Y(_00505_),
    .A1(_02704_),
    .A2(_02725_));
 sg13g2_nor2b_1 _19846_ (.A(_12723_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_02727_));
 sg13g2_a21oi_1 _19847_ (.A1(net1002),
    .A2(_12723_),
    .Y(_02728_),
    .B1(_02727_));
 sg13g2_nand2_1 _19848_ (.Y(_02729_),
    .A(net864),
    .B(_12720_));
 sg13g2_o21ai_1 _19849_ (.B1(_02729_),
    .Y(_00506_),
    .A1(_12721_),
    .A2(_02728_));
 sg13g2_nor2b_1 _19850_ (.A(_02720_),
    .B_N(\cpu.dcache.r_data[5][30] ),
    .Y(_02730_));
 sg13g2_a21oi_1 _19851_ (.A1(net1002),
    .A2(_02720_),
    .Y(_02731_),
    .B1(_02730_));
 sg13g2_nand2_1 _19852_ (.Y(_02732_),
    .A(net478),
    .B(_02703_));
 sg13g2_o21ai_1 _19853_ (.B1(_02732_),
    .Y(_00507_),
    .A1(net40),
    .A2(_02731_));
 sg13g2_nor2b_1 _19854_ (.A(_02720_),
    .B_N(\cpu.dcache.r_data[5][31] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _19855_ (.A1(net1001),
    .A2(_02720_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2_1 _19856_ (.Y(_02735_),
    .A(net477),
    .B(_02703_));
 sg13g2_o21ai_1 _19857_ (.B1(_02735_),
    .Y(_00508_),
    .A1(_02704_),
    .A2(_02734_));
 sg13g2_nor2b_1 _19858_ (.A(_12723_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_02736_));
 sg13g2_a21oi_1 _19859_ (.A1(net1001),
    .A2(_12723_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_nand2_1 _19860_ (.Y(_02738_),
    .A(net1000),
    .B(_12720_));
 sg13g2_o21ai_1 _19861_ (.B1(_02738_),
    .Y(_00509_),
    .A1(net43),
    .A2(_02737_));
 sg13g2_nor2_1 _19862_ (.A(_12717_),
    .B(_12327_),
    .Y(_02739_));
 sg13g2_buf_2 _19863_ (.A(_02739_),
    .X(_02740_));
 sg13g2_nor2b_1 _19864_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_02741_));
 sg13g2_a21oi_1 _19865_ (.A1(net1004),
    .A2(_02740_),
    .Y(_02742_),
    .B1(_02741_));
 sg13g2_nand2_1 _19866_ (.Y(_02743_),
    .A(_12271_),
    .B(_12720_));
 sg13g2_o21ai_1 _19867_ (.B1(_02743_),
    .Y(_00510_),
    .A1(net43),
    .A2(_02742_));
 sg13g2_nor2b_1 _19868_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_02744_));
 sg13g2_a21oi_1 _19869_ (.A1(net1003),
    .A2(_02740_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_nand2_1 _19870_ (.Y(_02746_),
    .A(net1011),
    .B(_12720_));
 sg13g2_o21ai_1 _19871_ (.B1(_02746_),
    .Y(_00511_),
    .A1(net43),
    .A2(_02745_));
 sg13g2_buf_1 _19872_ (.A(_12208_),
    .X(_02747_));
 sg13g2_nor2b_1 _19873_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][6] ),
    .Y(_02748_));
 sg13g2_a21oi_1 _19874_ (.A1(net998),
    .A2(_02740_),
    .Y(_02749_),
    .B1(_02748_));
 sg13g2_nand2_1 _19875_ (.Y(_02750_),
    .A(net1010),
    .B(_12720_));
 sg13g2_o21ai_1 _19876_ (.B1(_02750_),
    .Y(_00512_),
    .A1(_12721_),
    .A2(_02749_));
 sg13g2_buf_1 _19877_ (.A(_12215_),
    .X(_02751_));
 sg13g2_nor2b_1 _19878_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][7] ),
    .Y(_02752_));
 sg13g2_a21oi_1 _19879_ (.A1(net997),
    .A2(_02740_),
    .Y(_02753_),
    .B1(_02752_));
 sg13g2_nand2_1 _19880_ (.Y(_02754_),
    .A(net1012),
    .B(_12720_));
 sg13g2_o21ai_1 _19881_ (.B1(_02754_),
    .Y(_00513_),
    .A1(net43),
    .A2(_02753_));
 sg13g2_buf_1 _19882_ (.A(_12195_),
    .X(_02755_));
 sg13g2_nor2b_1 _19883_ (.A(_12731_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_02756_));
 sg13g2_a21oi_1 _19884_ (.A1(net996),
    .A2(_12731_),
    .Y(_02757_),
    .B1(_02756_));
 sg13g2_nand2_1 _19885_ (.Y(_02758_),
    .A(net476),
    .B(_12728_));
 sg13g2_o21ai_1 _19886_ (.B1(_02758_),
    .Y(_00514_),
    .A1(net42),
    .A2(_02757_));
 sg13g2_buf_1 _19887_ (.A(_12226_),
    .X(_02759_));
 sg13g2_nor2b_1 _19888_ (.A(_12731_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_02760_));
 sg13g2_a21oi_1 _19889_ (.A1(net995),
    .A2(_12731_),
    .Y(_02761_),
    .B1(_02760_));
 sg13g2_nand2_1 _19890_ (.Y(_02762_),
    .A(net475),
    .B(_12728_));
 sg13g2_o21ai_1 _19891_ (.B1(_02762_),
    .Y(_00515_),
    .A1(net42),
    .A2(_02761_));
 sg13g2_nand2_1 _19892_ (.Y(_02763_),
    .A(net919),
    .B(_09451_));
 sg13g2_buf_2 _19893_ (.A(_02763_),
    .X(_02764_));
 sg13g2_buf_1 _19894_ (.A(_02764_),
    .X(_02765_));
 sg13g2_nor2_1 _19895_ (.A(net593),
    .B(_12191_),
    .Y(_02766_));
 sg13g2_buf_2 _19896_ (.A(_02766_),
    .X(_02767_));
 sg13g2_buf_1 _19897_ (.A(_02767_),
    .X(_02768_));
 sg13g2_nor2_1 _19898_ (.A(net593),
    .B(_12065_),
    .Y(_02769_));
 sg13g2_buf_2 _19899_ (.A(_02769_),
    .X(_02770_));
 sg13g2_nor2b_1 _19900_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_02771_));
 sg13g2_a21oi_1 _19901_ (.A1(net996),
    .A2(_02770_),
    .Y(_02772_),
    .B1(_02771_));
 sg13g2_nand2_1 _19902_ (.Y(_02773_),
    .A(_10082_),
    .B(net39));
 sg13g2_o21ai_1 _19903_ (.B1(_02773_),
    .Y(_00516_),
    .A1(net39),
    .A2(_02772_));
 sg13g2_nor2_1 _19904_ (.A(net593),
    .B(_12204_),
    .Y(_02774_));
 sg13g2_buf_2 _19905_ (.A(_02774_),
    .X(_02775_));
 sg13g2_buf_1 _19906_ (.A(_02775_),
    .X(_02776_));
 sg13g2_nor2_1 _19907_ (.A(net593),
    .B(_12089_),
    .Y(_02777_));
 sg13g2_buf_2 _19908_ (.A(_02777_),
    .X(_02778_));
 sg13g2_nor2b_1 _19909_ (.A(_02778_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_02779_));
 sg13g2_a21oi_1 _19910_ (.A1(net998),
    .A2(_02778_),
    .Y(_02780_),
    .B1(_02779_));
 sg13g2_nand2_1 _19911_ (.Y(_02781_),
    .A(net482),
    .B(net38));
 sg13g2_o21ai_1 _19912_ (.B1(_02781_),
    .Y(_00517_),
    .A1(net38),
    .A2(_02780_));
 sg13g2_nor2b_1 _19913_ (.A(_02778_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_02782_));
 sg13g2_a21oi_1 _19914_ (.A1(net997),
    .A2(_02778_),
    .Y(_02783_),
    .B1(_02782_));
 sg13g2_nand2_1 _19915_ (.Y(_02784_),
    .A(net481),
    .B(net38));
 sg13g2_o21ai_1 _19916_ (.B1(_02784_),
    .Y(_00518_),
    .A1(net38),
    .A2(_02783_));
 sg13g2_nor2_1 _19917_ (.A(_02765_),
    .B(_12111_),
    .Y(_02785_));
 sg13g2_buf_2 _19918_ (.A(_02785_),
    .X(_02786_));
 sg13g2_nor2b_1 _19919_ (.A(_02786_),
    .B_N(\cpu.dcache.r_data[6][12] ),
    .Y(_02787_));
 sg13g2_a21oi_1 _19920_ (.A1(net996),
    .A2(_02786_),
    .Y(_02788_),
    .B1(_02787_));
 sg13g2_nand2_1 _19921_ (.Y(_02789_),
    .A(net480),
    .B(_02775_));
 sg13g2_o21ai_1 _19922_ (.B1(_02789_),
    .Y(_00519_),
    .A1(net38),
    .A2(_02788_));
 sg13g2_nor2b_1 _19923_ (.A(_02786_),
    .B_N(\cpu.dcache.r_data[6][13] ),
    .Y(_02790_));
 sg13g2_a21oi_1 _19924_ (.A1(net995),
    .A2(_02786_),
    .Y(_02791_),
    .B1(_02790_));
 sg13g2_nand2_1 _19925_ (.Y(_02792_),
    .A(net479),
    .B(_02775_));
 sg13g2_o21ai_1 _19926_ (.B1(_02792_),
    .Y(_00520_),
    .A1(_02776_),
    .A2(_02791_));
 sg13g2_nor2b_1 _19927_ (.A(_02786_),
    .B_N(\cpu.dcache.r_data[6][14] ),
    .Y(_02793_));
 sg13g2_a21oi_1 _19928_ (.A1(net998),
    .A2(_02786_),
    .Y(_02794_),
    .B1(_02793_));
 sg13g2_nand2_1 _19929_ (.Y(_02795_),
    .A(net478),
    .B(_02775_));
 sg13g2_o21ai_1 _19930_ (.B1(_02795_),
    .Y(_00521_),
    .A1(_02776_),
    .A2(_02794_));
 sg13g2_nor2b_1 _19931_ (.A(_02786_),
    .B_N(\cpu.dcache.r_data[6][15] ),
    .Y(_02796_));
 sg13g2_a21oi_1 _19932_ (.A1(_02751_),
    .A2(_02786_),
    .Y(_02797_),
    .B1(_02796_));
 sg13g2_nand2_1 _19933_ (.Y(_02798_),
    .A(net477),
    .B(_02775_));
 sg13g2_o21ai_1 _19934_ (.B1(_02798_),
    .Y(_00522_),
    .A1(net38),
    .A2(_02797_));
 sg13g2_nor2_1 _19935_ (.A(net593),
    .B(_12238_),
    .Y(_02799_));
 sg13g2_buf_2 _19936_ (.A(_02799_),
    .X(_02800_));
 sg13g2_buf_1 _19937_ (.A(_02800_),
    .X(_02801_));
 sg13g2_nor2_1 _19938_ (.A(net593),
    .B(_12133_),
    .Y(_02802_));
 sg13g2_buf_2 _19939_ (.A(_02802_),
    .X(_02803_));
 sg13g2_nor2b_1 _19940_ (.A(_02803_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02804_));
 sg13g2_a21oi_1 _19941_ (.A1(net996),
    .A2(_02803_),
    .Y(_02805_),
    .B1(_02804_));
 sg13g2_nand2_1 _19942_ (.Y(_02806_),
    .A(net901),
    .B(net37));
 sg13g2_o21ai_1 _19943_ (.B1(_02806_),
    .Y(_00523_),
    .A1(net37),
    .A2(_02805_));
 sg13g2_nor2b_1 _19944_ (.A(_02803_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_02807_));
 sg13g2_a21oi_1 _19945_ (.A1(net995),
    .A2(_02803_),
    .Y(_02808_),
    .B1(_02807_));
 sg13g2_nand2_1 _19946_ (.Y(_02809_),
    .A(net999),
    .B(_02801_));
 sg13g2_o21ai_1 _19947_ (.B1(_02809_),
    .Y(_00524_),
    .A1(_02801_),
    .A2(_02808_));
 sg13g2_nor2b_1 _19948_ (.A(_02803_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_02810_));
 sg13g2_a21oi_1 _19949_ (.A1(net998),
    .A2(_02803_),
    .Y(_02811_),
    .B1(_02810_));
 sg13g2_nand2_1 _19950_ (.Y(_02812_),
    .A(net864),
    .B(_02800_));
 sg13g2_o21ai_1 _19951_ (.B1(_02812_),
    .Y(_00525_),
    .A1(net37),
    .A2(_02811_));
 sg13g2_nor2b_1 _19952_ (.A(_02803_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02813_));
 sg13g2_a21oi_1 _19953_ (.A1(net997),
    .A2(_02803_),
    .Y(_02814_),
    .B1(_02813_));
 sg13g2_nand2_1 _19954_ (.Y(_02815_),
    .A(net1000),
    .B(_02800_));
 sg13g2_o21ai_1 _19955_ (.B1(_02815_),
    .Y(_00526_),
    .A1(net37),
    .A2(_02814_));
 sg13g2_nor2b_1 _19956_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02816_));
 sg13g2_a21oi_1 _19957_ (.A1(net995),
    .A2(_02770_),
    .Y(_02817_),
    .B1(_02816_));
 sg13g2_nand2_1 _19958_ (.Y(_02818_),
    .A(net999),
    .B(net39));
 sg13g2_o21ai_1 _19959_ (.B1(_02818_),
    .Y(_00527_),
    .A1(net39),
    .A2(_02817_));
 sg13g2_nor2_1 _19960_ (.A(_02764_),
    .B(_12266_),
    .Y(_02819_));
 sg13g2_buf_2 _19961_ (.A(_02819_),
    .X(_02820_));
 sg13g2_nor2b_1 _19962_ (.A(_02820_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02821_));
 sg13g2_a21oi_1 _19963_ (.A1(net996),
    .A2(_02820_),
    .Y(_02822_),
    .B1(_02821_));
 sg13g2_nand2_1 _19964_ (.Y(_02823_),
    .A(net1015),
    .B(_02800_));
 sg13g2_o21ai_1 _19965_ (.B1(_02823_),
    .Y(_00528_),
    .A1(net37),
    .A2(_02822_));
 sg13g2_nor2b_1 _19966_ (.A(_02820_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02824_));
 sg13g2_a21oi_1 _19967_ (.A1(net995),
    .A2(_02820_),
    .Y(_02825_),
    .B1(_02824_));
 sg13g2_nand2_1 _19968_ (.Y(_02826_),
    .A(net1011),
    .B(_02800_));
 sg13g2_o21ai_1 _19969_ (.B1(_02826_),
    .Y(_00529_),
    .A1(net37),
    .A2(_02825_));
 sg13g2_nor2b_1 _19970_ (.A(_02820_),
    .B_N(\cpu.dcache.r_data[6][22] ),
    .Y(_02827_));
 sg13g2_a21oi_1 _19971_ (.A1(net998),
    .A2(_02820_),
    .Y(_02828_),
    .B1(_02827_));
 sg13g2_nand2_1 _19972_ (.Y(_02829_),
    .A(net1010),
    .B(_02800_));
 sg13g2_o21ai_1 _19973_ (.B1(_02829_),
    .Y(_00530_),
    .A1(net37),
    .A2(_02828_));
 sg13g2_nor2b_1 _19974_ (.A(_02820_),
    .B_N(\cpu.dcache.r_data[6][23] ),
    .Y(_02830_));
 sg13g2_a21oi_1 _19975_ (.A1(net997),
    .A2(_02820_),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_nand2_1 _19976_ (.Y(_02832_),
    .A(net1050),
    .B(_02800_));
 sg13g2_o21ai_1 _19977_ (.B1(_02832_),
    .Y(_00531_),
    .A1(net37),
    .A2(_02831_));
 sg13g2_nor2_1 _19978_ (.A(_02765_),
    .B(_12286_),
    .Y(_02833_));
 sg13g2_buf_2 _19979_ (.A(_02833_),
    .X(_02834_));
 sg13g2_buf_1 _19980_ (.A(_02834_),
    .X(_02835_));
 sg13g2_nor2_1 _19981_ (.A(_02764_),
    .B(_12291_),
    .Y(_02836_));
 sg13g2_buf_1 _19982_ (.A(_02836_),
    .X(_02837_));
 sg13g2_nor2b_1 _19983_ (.A(net527),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02838_));
 sg13g2_a21oi_1 _19984_ (.A1(net996),
    .A2(net527),
    .Y(_02839_),
    .B1(_02838_));
 sg13g2_nand2_1 _19985_ (.Y(_02840_),
    .A(_12157_),
    .B(net36));
 sg13g2_o21ai_1 _19986_ (.B1(_02840_),
    .Y(_00532_),
    .A1(net36),
    .A2(_02839_));
 sg13g2_nor2b_1 _19987_ (.A(net527),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02841_));
 sg13g2_a21oi_1 _19988_ (.A1(net995),
    .A2(net527),
    .Y(_02842_),
    .B1(_02841_));
 sg13g2_nand2_1 _19989_ (.Y(_02843_),
    .A(net475),
    .B(net36));
 sg13g2_o21ai_1 _19990_ (.B1(_02843_),
    .Y(_00533_),
    .A1(net36),
    .A2(_02842_));
 sg13g2_nor2b_1 _19991_ (.A(net527),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02844_));
 sg13g2_a21oi_1 _19992_ (.A1(_02747_),
    .A2(net527),
    .Y(_02845_),
    .B1(_02844_));
 sg13g2_nand2_1 _19993_ (.Y(_02846_),
    .A(_12097_),
    .B(_02834_));
 sg13g2_o21ai_1 _19994_ (.B1(_02846_),
    .Y(_00534_),
    .A1(net36),
    .A2(_02845_));
 sg13g2_nor2b_1 _19995_ (.A(net527),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02847_));
 sg13g2_a21oi_1 _19996_ (.A1(net997),
    .A2(net527),
    .Y(_02848_),
    .B1(_02847_));
 sg13g2_nand2_1 _19997_ (.Y(_02849_),
    .A(_12107_),
    .B(_02834_));
 sg13g2_o21ai_1 _19998_ (.B1(_02849_),
    .Y(_00535_),
    .A1(net36),
    .A2(_02848_));
 sg13g2_nor2_1 _19999_ (.A(_02764_),
    .B(_12170_),
    .Y(_02850_));
 sg13g2_buf_2 _20000_ (.A(_02850_),
    .X(_02851_));
 sg13g2_nor2b_1 _20001_ (.A(_02851_),
    .B_N(\cpu.dcache.r_data[6][28] ),
    .Y(_02852_));
 sg13g2_a21oi_1 _20002_ (.A1(_02755_),
    .A2(_02851_),
    .Y(_02853_),
    .B1(_02852_));
 sg13g2_nand2_1 _20003_ (.Y(_02854_),
    .A(_12117_),
    .B(_02834_));
 sg13g2_o21ai_1 _20004_ (.B1(_02854_),
    .Y(_00536_),
    .A1(_02835_),
    .A2(_02853_));
 sg13g2_nor2b_1 _20005_ (.A(_02851_),
    .B_N(\cpu.dcache.r_data[6][29] ),
    .Y(_02855_));
 sg13g2_a21oi_1 _20006_ (.A1(net995),
    .A2(_02851_),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_nand2_1 _20007_ (.Y(_02857_),
    .A(net479),
    .B(_02834_));
 sg13g2_o21ai_1 _20008_ (.B1(_02857_),
    .Y(_00537_),
    .A1(net36),
    .A2(_02856_));
 sg13g2_nor2b_1 _20009_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02858_));
 sg13g2_a21oi_1 _20010_ (.A1(net998),
    .A2(_02770_),
    .Y(_02859_),
    .B1(_02858_));
 sg13g2_nand2_1 _20011_ (.Y(_02860_),
    .A(net864),
    .B(_02767_));
 sg13g2_o21ai_1 _20012_ (.B1(_02860_),
    .Y(_00538_),
    .A1(_02768_),
    .A2(_02859_));
 sg13g2_nor2b_1 _20013_ (.A(_02851_),
    .B_N(\cpu.dcache.r_data[6][30] ),
    .Y(_02861_));
 sg13g2_a21oi_1 _20014_ (.A1(_02747_),
    .A2(_02851_),
    .Y(_02862_),
    .B1(_02861_));
 sg13g2_nand2_1 _20015_ (.Y(_02863_),
    .A(_12127_),
    .B(_02834_));
 sg13g2_o21ai_1 _20016_ (.B1(_02863_),
    .Y(_00539_),
    .A1(_02835_),
    .A2(_02862_));
 sg13g2_nor2b_1 _20017_ (.A(_02851_),
    .B_N(\cpu.dcache.r_data[6][31] ),
    .Y(_02864_));
 sg13g2_a21oi_1 _20018_ (.A1(_02751_),
    .A2(_02851_),
    .Y(_02865_),
    .B1(_02864_));
 sg13g2_nand2_1 _20019_ (.Y(_02866_),
    .A(net477),
    .B(_02834_));
 sg13g2_o21ai_1 _20020_ (.B1(_02866_),
    .Y(_00540_),
    .A1(net36),
    .A2(_02865_));
 sg13g2_nor2b_1 _20021_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02867_));
 sg13g2_a21oi_1 _20022_ (.A1(net997),
    .A2(_02770_),
    .Y(_02868_),
    .B1(_02867_));
 sg13g2_nand2_1 _20023_ (.Y(_02869_),
    .A(net1000),
    .B(_02767_));
 sg13g2_o21ai_1 _20024_ (.B1(_02869_),
    .Y(_00541_),
    .A1(_02768_),
    .A2(_02868_));
 sg13g2_nor2_1 _20025_ (.A(_02764_),
    .B(_12327_),
    .Y(_02870_));
 sg13g2_buf_2 _20026_ (.A(_02870_),
    .X(_02871_));
 sg13g2_nor2b_1 _20027_ (.A(_02871_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02872_));
 sg13g2_a21oi_1 _20028_ (.A1(net996),
    .A2(_02871_),
    .Y(_02873_),
    .B1(_02872_));
 sg13g2_nand2_1 _20029_ (.Y(_02874_),
    .A(_10117_),
    .B(_02767_));
 sg13g2_o21ai_1 _20030_ (.B1(_02874_),
    .Y(_00542_),
    .A1(net39),
    .A2(_02873_));
 sg13g2_nor2b_1 _20031_ (.A(_02871_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02875_));
 sg13g2_a21oi_1 _20032_ (.A1(net995),
    .A2(_02871_),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nand2_1 _20033_ (.Y(_02877_),
    .A(net1011),
    .B(_02767_));
 sg13g2_o21ai_1 _20034_ (.B1(_02877_),
    .Y(_00543_),
    .A1(net39),
    .A2(_02876_));
 sg13g2_nor2b_1 _20035_ (.A(_02871_),
    .B_N(\cpu.dcache.r_data[6][6] ),
    .Y(_02878_));
 sg13g2_a21oi_1 _20036_ (.A1(net998),
    .A2(_02871_),
    .Y(_02879_),
    .B1(_02878_));
 sg13g2_nand2_1 _20037_ (.Y(_02880_),
    .A(net1010),
    .B(_02767_));
 sg13g2_o21ai_1 _20038_ (.B1(_02880_),
    .Y(_00544_),
    .A1(net39),
    .A2(_02879_));
 sg13g2_nor2b_1 _20039_ (.A(_02871_),
    .B_N(\cpu.dcache.r_data[6][7] ),
    .Y(_02881_));
 sg13g2_a21oi_1 _20040_ (.A1(net997),
    .A2(_02871_),
    .Y(_02882_),
    .B1(_02881_));
 sg13g2_nand2_1 _20041_ (.Y(_02883_),
    .A(_10132_),
    .B(_02767_));
 sg13g2_o21ai_1 _20042_ (.B1(_02883_),
    .Y(_00545_),
    .A1(net39),
    .A2(_02882_));
 sg13g2_nor2b_1 _20043_ (.A(_02778_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02884_));
 sg13g2_a21oi_1 _20044_ (.A1(_02755_),
    .A2(_02778_),
    .Y(_02885_),
    .B1(_02884_));
 sg13g2_nand2_1 _20045_ (.Y(_02886_),
    .A(_12156_),
    .B(_02775_));
 sg13g2_o21ai_1 _20046_ (.B1(_02886_),
    .Y(_00546_),
    .A1(net38),
    .A2(_02885_));
 sg13g2_nor2b_1 _20047_ (.A(_02778_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02887_));
 sg13g2_a21oi_1 _20048_ (.A1(_02759_),
    .A2(_02778_),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_nand2_1 _20049_ (.Y(_02889_),
    .A(_12165_),
    .B(_02775_));
 sg13g2_o21ai_1 _20050_ (.B1(_02889_),
    .Y(_00547_),
    .A1(net38),
    .A2(_02888_));
 sg13g2_buf_1 _20051_ (.A(_10097_),
    .X(_02890_));
 sg13g2_nor2_1 _20052_ (.A(net469),
    .B(_12191_),
    .Y(_02891_));
 sg13g2_buf_1 _20053_ (.A(_02891_),
    .X(_02892_));
 sg13g2_nor2_1 _20054_ (.A(net469),
    .B(_12065_),
    .Y(_02893_));
 sg13g2_buf_2 _20055_ (.A(_02893_),
    .X(_02894_));
 sg13g2_nor2b_1 _20056_ (.A(_02894_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02895_));
 sg13g2_a21oi_1 _20057_ (.A1(net996),
    .A2(_02894_),
    .Y(_02896_),
    .B1(_02895_));
 sg13g2_nand2_1 _20058_ (.Y(_02897_),
    .A(_10082_),
    .B(net60));
 sg13g2_o21ai_1 _20059_ (.B1(_02897_),
    .Y(_00548_),
    .A1(net60),
    .A2(_02896_));
 sg13g2_nor2_1 _20060_ (.A(_02890_),
    .B(_12204_),
    .Y(_02898_));
 sg13g2_buf_2 _20061_ (.A(_02898_),
    .X(_02899_));
 sg13g2_buf_1 _20062_ (.A(_02899_),
    .X(_02900_));
 sg13g2_nor2_1 _20063_ (.A(net469),
    .B(_12089_),
    .Y(_02901_));
 sg13g2_buf_2 _20064_ (.A(_02901_),
    .X(_02902_));
 sg13g2_nor2b_1 _20065_ (.A(_02902_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02903_));
 sg13g2_a21oi_1 _20066_ (.A1(net998),
    .A2(_02902_),
    .Y(_02904_),
    .B1(_02903_));
 sg13g2_nand2_1 _20067_ (.Y(_02905_),
    .A(_12097_),
    .B(net35));
 sg13g2_o21ai_1 _20068_ (.B1(_02905_),
    .Y(_00549_),
    .A1(net35),
    .A2(_02904_));
 sg13g2_nor2b_1 _20069_ (.A(_02902_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02906_));
 sg13g2_a21oi_1 _20070_ (.A1(net997),
    .A2(_02902_),
    .Y(_02907_),
    .B1(_02906_));
 sg13g2_nand2_1 _20071_ (.Y(_02908_),
    .A(_12107_),
    .B(net35));
 sg13g2_o21ai_1 _20072_ (.B1(_02908_),
    .Y(_00550_),
    .A1(net35),
    .A2(_02907_));
 sg13g2_buf_2 _20073_ (.A(_12051_),
    .X(_02909_));
 sg13g2_nor2_1 _20074_ (.A(_02890_),
    .B(_12111_),
    .Y(_02910_));
 sg13g2_buf_2 _20075_ (.A(_02910_),
    .X(_02911_));
 sg13g2_nor2b_1 _20076_ (.A(_02911_),
    .B_N(\cpu.dcache.r_data[7][12] ),
    .Y(_02912_));
 sg13g2_a21oi_1 _20077_ (.A1(net1111),
    .A2(_02911_),
    .Y(_02913_),
    .B1(_02912_));
 sg13g2_nand2_1 _20078_ (.Y(_02914_),
    .A(_12116_),
    .B(_02899_));
 sg13g2_o21ai_1 _20079_ (.B1(_02914_),
    .Y(_00551_),
    .A1(net35),
    .A2(_02913_));
 sg13g2_nor2b_1 _20080_ (.A(_02911_),
    .B_N(\cpu.dcache.r_data[7][13] ),
    .Y(_02915_));
 sg13g2_a21oi_1 _20081_ (.A1(_02759_),
    .A2(_02911_),
    .Y(_02916_),
    .B1(_02915_));
 sg13g2_nand2_1 _20082_ (.Y(_02917_),
    .A(_12122_),
    .B(_02899_));
 sg13g2_o21ai_1 _20083_ (.B1(_02917_),
    .Y(_00552_),
    .A1(net35),
    .A2(_02916_));
 sg13g2_buf_2 _20084_ (.A(_12086_),
    .X(_02918_));
 sg13g2_nor2b_1 _20085_ (.A(_02911_),
    .B_N(\cpu.dcache.r_data[7][14] ),
    .Y(_02919_));
 sg13g2_a21oi_1 _20086_ (.A1(net1110),
    .A2(_02911_),
    .Y(_02920_),
    .B1(_02919_));
 sg13g2_nand2_1 _20087_ (.Y(_02921_),
    .A(_12126_),
    .B(_02899_));
 sg13g2_o21ai_1 _20088_ (.B1(_02921_),
    .Y(_00553_),
    .A1(net35),
    .A2(_02920_));
 sg13g2_buf_2 _20089_ (.A(_12103_),
    .X(_02922_));
 sg13g2_nor2b_1 _20090_ (.A(_02911_),
    .B_N(\cpu.dcache.r_data[7][15] ),
    .Y(_02923_));
 sg13g2_a21oi_1 _20091_ (.A1(net1109),
    .A2(_02911_),
    .Y(_02924_),
    .B1(_02923_));
 sg13g2_nand2_1 _20092_ (.Y(_02925_),
    .A(_12130_),
    .B(_02899_));
 sg13g2_o21ai_1 _20093_ (.B1(_02925_),
    .Y(_00554_),
    .A1(net35),
    .A2(_02924_));
 sg13g2_nor2_1 _20094_ (.A(net469),
    .B(_12238_),
    .Y(_02926_));
 sg13g2_buf_1 _20095_ (.A(_02926_),
    .X(_02927_));
 sg13g2_nor2_1 _20096_ (.A(net469),
    .B(_12133_),
    .Y(_02928_));
 sg13g2_buf_2 _20097_ (.A(_02928_),
    .X(_02929_));
 sg13g2_nor2b_1 _20098_ (.A(_02929_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02930_));
 sg13g2_a21oi_1 _20099_ (.A1(net1111),
    .A2(_02929_),
    .Y(_02931_),
    .B1(_02930_));
 sg13g2_nand2_1 _20100_ (.Y(_02932_),
    .A(net901),
    .B(net59));
 sg13g2_o21ai_1 _20101_ (.B1(_02932_),
    .Y(_00555_),
    .A1(net59),
    .A2(_02931_));
 sg13g2_buf_2 _20102_ (.A(_12118_),
    .X(_02933_));
 sg13g2_nor2b_1 _20103_ (.A(_02929_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02934_));
 sg13g2_a21oi_1 _20104_ (.A1(net1108),
    .A2(_02929_),
    .Y(_02935_),
    .B1(_02934_));
 sg13g2_nand2_1 _20105_ (.Y(_02936_),
    .A(_12762_),
    .B(net59));
 sg13g2_o21ai_1 _20106_ (.B1(_02936_),
    .Y(_00556_),
    .A1(net59),
    .A2(_02935_));
 sg13g2_nor2b_1 _20107_ (.A(_02929_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02937_));
 sg13g2_a21oi_1 _20108_ (.A1(net1110),
    .A2(_02929_),
    .Y(_02938_),
    .B1(_02937_));
 sg13g2_nand2_1 _20109_ (.Y(_02939_),
    .A(_12766_),
    .B(_02926_));
 sg13g2_o21ai_1 _20110_ (.B1(_02939_),
    .Y(_00557_),
    .A1(_02927_),
    .A2(_02938_));
 sg13g2_nor2b_1 _20111_ (.A(_02929_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02940_));
 sg13g2_a21oi_1 _20112_ (.A1(net1109),
    .A2(_02929_),
    .Y(_02941_),
    .B1(_02940_));
 sg13g2_nand2_1 _20113_ (.Y(_02942_),
    .A(net1000),
    .B(_02926_));
 sg13g2_o21ai_1 _20114_ (.B1(_02942_),
    .Y(_00558_),
    .A1(_02927_),
    .A2(_02941_));
 sg13g2_nor2b_1 _20115_ (.A(_02894_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02943_));
 sg13g2_a21oi_1 _20116_ (.A1(net1108),
    .A2(_02894_),
    .Y(_02944_),
    .B1(_02943_));
 sg13g2_nand2_1 _20117_ (.Y(_02945_),
    .A(_12762_),
    .B(_02892_));
 sg13g2_o21ai_1 _20118_ (.B1(_02945_),
    .Y(_00559_),
    .A1(_02892_),
    .A2(_02944_));
 sg13g2_nand2_2 _20119_ (.Y(_02946_),
    .A(net485),
    .B(_12145_));
 sg13g2_mux2_1 _20120_ (.A0(net1115),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02946_),
    .X(_02947_));
 sg13g2_mux2_1 _20121_ (.A0(_02947_),
    .A1(net865),
    .S(net59),
    .X(_00560_));
 sg13g2_mux2_1 _20122_ (.A0(net1112),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02946_),
    .X(_02948_));
 sg13g2_mux2_1 _20123_ (.A0(_02948_),
    .A1(net1014),
    .S(net59),
    .X(_00561_));
 sg13g2_mux2_1 _20124_ (.A0(net1114),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02946_),
    .X(_02949_));
 sg13g2_mux2_1 _20125_ (.A0(_02949_),
    .A1(net1013),
    .S(net59),
    .X(_00562_));
 sg13g2_mux2_1 _20126_ (.A0(net1113),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02946_),
    .X(_02950_));
 sg13g2_mux2_1 _20127_ (.A0(_02950_),
    .A1(net1005),
    .S(net59),
    .X(_00563_));
 sg13g2_nor2_1 _20128_ (.A(net469),
    .B(_12286_),
    .Y(_02951_));
 sg13g2_buf_2 _20129_ (.A(_02951_),
    .X(_02952_));
 sg13g2_buf_1 _20130_ (.A(_02952_),
    .X(_02953_));
 sg13g2_nor2_1 _20131_ (.A(_10097_),
    .B(_12291_),
    .Y(_02954_));
 sg13g2_buf_1 _20132_ (.A(_02954_),
    .X(_02955_));
 sg13g2_nor2b_1 _20133_ (.A(net423),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02956_));
 sg13g2_a21oi_1 _20134_ (.A1(net1111),
    .A2(net423),
    .Y(_02957_),
    .B1(_02956_));
 sg13g2_nand2_1 _20135_ (.Y(_02958_),
    .A(_12156_),
    .B(net34));
 sg13g2_o21ai_1 _20136_ (.B1(_02958_),
    .Y(_00564_),
    .A1(net34),
    .A2(_02957_));
 sg13g2_nor2b_1 _20137_ (.A(net423),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02959_));
 sg13g2_a21oi_1 _20138_ (.A1(net1108),
    .A2(net423),
    .Y(_02960_),
    .B1(_02959_));
 sg13g2_nand2_1 _20139_ (.Y(_02961_),
    .A(_12165_),
    .B(net34));
 sg13g2_o21ai_1 _20140_ (.B1(_02961_),
    .Y(_00565_),
    .A1(net34),
    .A2(_02960_));
 sg13g2_nor2b_1 _20141_ (.A(_02955_),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02962_));
 sg13g2_a21oi_1 _20142_ (.A1(net1110),
    .A2(_02955_),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_nand2_1 _20143_ (.Y(_02964_),
    .A(_12097_),
    .B(_02952_));
 sg13g2_o21ai_1 _20144_ (.B1(_02964_),
    .Y(_00566_),
    .A1(net34),
    .A2(_02963_));
 sg13g2_nor2b_1 _20145_ (.A(net423),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02965_));
 sg13g2_a21oi_1 _20146_ (.A1(net1109),
    .A2(net423),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_nand2_1 _20147_ (.Y(_02967_),
    .A(_12107_),
    .B(_02952_));
 sg13g2_o21ai_1 _20148_ (.B1(_02967_),
    .Y(_00567_),
    .A1(net34),
    .A2(_02966_));
 sg13g2_nor2_1 _20149_ (.A(_10097_),
    .B(_12170_),
    .Y(_02968_));
 sg13g2_buf_2 _20150_ (.A(_02968_),
    .X(_02969_));
 sg13g2_nor2b_1 _20151_ (.A(_02969_),
    .B_N(\cpu.dcache.r_data[7][28] ),
    .Y(_02970_));
 sg13g2_a21oi_1 _20152_ (.A1(net1111),
    .A2(_02969_),
    .Y(_02971_),
    .B1(_02970_));
 sg13g2_nand2_1 _20153_ (.Y(_02972_),
    .A(_12116_),
    .B(_02952_));
 sg13g2_o21ai_1 _20154_ (.B1(_02972_),
    .Y(_00568_),
    .A1(net34),
    .A2(_02971_));
 sg13g2_nor2b_1 _20155_ (.A(_02969_),
    .B_N(\cpu.dcache.r_data[7][29] ),
    .Y(_02973_));
 sg13g2_a21oi_1 _20156_ (.A1(net1108),
    .A2(_02969_),
    .Y(_02974_),
    .B1(_02973_));
 sg13g2_nand2_1 _20157_ (.Y(_02975_),
    .A(_12122_),
    .B(_02952_));
 sg13g2_o21ai_1 _20158_ (.B1(_02975_),
    .Y(_00569_),
    .A1(_02953_),
    .A2(_02974_));
 sg13g2_nor2b_1 _20159_ (.A(_02894_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02976_));
 sg13g2_a21oi_1 _20160_ (.A1(net1110),
    .A2(_02894_),
    .Y(_02977_),
    .B1(_02976_));
 sg13g2_nand2_1 _20161_ (.Y(_02978_),
    .A(_12766_),
    .B(_02891_));
 sg13g2_o21ai_1 _20162_ (.B1(_02978_),
    .Y(_00570_),
    .A1(net60),
    .A2(_02977_));
 sg13g2_nor2b_1 _20163_ (.A(_02969_),
    .B_N(\cpu.dcache.r_data[7][30] ),
    .Y(_02979_));
 sg13g2_a21oi_1 _20164_ (.A1(net1110),
    .A2(_02969_),
    .Y(_02980_),
    .B1(_02979_));
 sg13g2_nand2_1 _20165_ (.Y(_02981_),
    .A(_12126_),
    .B(_02952_));
 sg13g2_o21ai_1 _20166_ (.B1(_02981_),
    .Y(_00571_),
    .A1(_02953_),
    .A2(_02980_));
 sg13g2_nor2b_1 _20167_ (.A(_02969_),
    .B_N(\cpu.dcache.r_data[7][31] ),
    .Y(_02982_));
 sg13g2_a21oi_1 _20168_ (.A1(net1109),
    .A2(_02969_),
    .Y(_02983_),
    .B1(_02982_));
 sg13g2_nand2_1 _20169_ (.Y(_02984_),
    .A(_12130_),
    .B(_02952_));
 sg13g2_o21ai_1 _20170_ (.B1(_02984_),
    .Y(_00572_),
    .A1(net34),
    .A2(_02983_));
 sg13g2_nor2b_1 _20171_ (.A(_02894_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02985_));
 sg13g2_a21oi_1 _20172_ (.A1(net1109),
    .A2(_02894_),
    .Y(_02986_),
    .B1(_02985_));
 sg13g2_nand2_1 _20173_ (.Y(_02987_),
    .A(net1000),
    .B(_02891_));
 sg13g2_o21ai_1 _20174_ (.B1(_02987_),
    .Y(_00573_),
    .A1(net60),
    .A2(_02986_));
 sg13g2_nand2_2 _20175_ (.Y(_02988_),
    .A(_10025_),
    .B(_12179_));
 sg13g2_mux2_1 _20176_ (.A0(net1115),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02988_),
    .X(_02989_));
 sg13g2_mux2_1 _20177_ (.A0(_02989_),
    .A1(_12581_),
    .S(net60),
    .X(_00574_));
 sg13g2_mux2_1 _20178_ (.A0(net1112),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02988_),
    .X(_02990_));
 sg13g2_mux2_1 _20179_ (.A0(_02990_),
    .A1(_12275_),
    .S(net60),
    .X(_00575_));
 sg13g2_mux2_1 _20180_ (.A0(net1114),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02988_),
    .X(_02991_));
 sg13g2_mux2_1 _20181_ (.A0(_02991_),
    .A1(net1013),
    .S(net60),
    .X(_00576_));
 sg13g2_mux2_1 _20182_ (.A0(net1113),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02988_),
    .X(_02992_));
 sg13g2_mux2_1 _20183_ (.A0(_02992_),
    .A1(_12541_),
    .S(net60),
    .X(_00577_));
 sg13g2_nor2b_1 _20184_ (.A(_02902_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02993_));
 sg13g2_a21oi_1 _20185_ (.A1(net1111),
    .A2(_02902_),
    .Y(_02994_),
    .B1(_02993_));
 sg13g2_nand2_1 _20186_ (.Y(_02995_),
    .A(_12156_),
    .B(_02899_));
 sg13g2_o21ai_1 _20187_ (.B1(_02995_),
    .Y(_00578_),
    .A1(_02900_),
    .A2(_02994_));
 sg13g2_nor2b_1 _20188_ (.A(_02902_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02996_));
 sg13g2_a21oi_1 _20189_ (.A1(net1108),
    .A2(_02902_),
    .Y(_02997_),
    .B1(_02996_));
 sg13g2_nand2_1 _20190_ (.Y(_02998_),
    .A(_12165_),
    .B(_02899_));
 sg13g2_o21ai_1 _20191_ (.B1(_02998_),
    .Y(_00579_),
    .A1(_02900_),
    .A2(_02997_));
 sg13g2_and2_1 _20192_ (.A(_09831_),
    .B(_12075_),
    .X(_02999_));
 sg13g2_buf_1 _20193_ (.A(\cpu.d_rstrobe_d ),
    .X(_03000_));
 sg13g2_inv_1 _20194_ (.Y(_03001_),
    .A(_12055_));
 sg13g2_nor4_1 _20195_ (.A(_09398_),
    .B(_03000_),
    .C(_03001_),
    .D(_08409_),
    .Y(_03002_));
 sg13g2_or2_1 _20196_ (.X(_03003_),
    .B(_03002_),
    .A(_02999_));
 sg13g2_buf_2 _20197_ (.A(_03003_),
    .X(_03004_));
 sg13g2_buf_1 _20198_ (.A(_12071_),
    .X(_03005_));
 sg13g2_inv_1 _20199_ (.Y(_03006_),
    .A(net994));
 sg13g2_nor2_1 _20200_ (.A(_03006_),
    .B(_12070_),
    .Y(_03007_));
 sg13g2_xor2_1 _20201_ (.B(_12055_),
    .A(_03000_),
    .X(_03008_));
 sg13g2_a21oi_1 _20202_ (.A1(_03007_),
    .A2(_03008_),
    .Y(_03009_),
    .B1(_02999_));
 sg13g2_buf_2 _20203_ (.A(_03009_),
    .X(_03010_));
 sg13g2_nor2_1 _20204_ (.A(net659),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_mux2_1 _20205_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_03004_),
    .S(_03011_),
    .X(_00580_));
 sg13g2_nor2_1 _20206_ (.A(net658),
    .B(_03010_),
    .Y(_03012_));
 sg13g2_mux2_1 _20207_ (.A0(\cpu.dcache.r_dirty[1] ),
    .A1(_03004_),
    .S(_03012_),
    .X(_00581_));
 sg13g2_nor2_1 _20208_ (.A(net532),
    .B(_03010_),
    .Y(_03013_));
 sg13g2_mux2_1 _20209_ (.A0(\cpu.dcache.r_dirty[2] ),
    .A1(_03004_),
    .S(_03013_),
    .X(_00582_));
 sg13g2_nor2_1 _20210_ (.A(net531),
    .B(_03010_),
    .Y(_03014_));
 sg13g2_mux2_1 _20211_ (.A0(\cpu.dcache.r_dirty[3] ),
    .A1(_03004_),
    .S(_03014_),
    .X(_00583_));
 sg13g2_nor2_1 _20212_ (.A(net594),
    .B(_03010_),
    .Y(_03015_));
 sg13g2_mux2_1 _20213_ (.A0(\cpu.dcache.r_dirty[4] ),
    .A1(_03004_),
    .S(_03015_),
    .X(_00584_));
 sg13g2_nor2_1 _20214_ (.A(_12718_),
    .B(_03010_),
    .Y(_03016_));
 sg13g2_mux2_1 _20215_ (.A0(\cpu.dcache.r_dirty[5] ),
    .A1(_03004_),
    .S(_03016_),
    .X(_00585_));
 sg13g2_nor2_1 _20216_ (.A(net593),
    .B(_03010_),
    .Y(_03017_));
 sg13g2_mux2_1 _20217_ (.A0(\cpu.dcache.r_dirty[6] ),
    .A1(_03004_),
    .S(_03017_),
    .X(_00586_));
 sg13g2_nor2_1 _20218_ (.A(net469),
    .B(_03010_),
    .Y(_03018_));
 sg13g2_mux2_1 _20219_ (.A0(\cpu.dcache.r_dirty[7] ),
    .A1(_03004_),
    .S(_03018_),
    .X(_00587_));
 sg13g2_buf_1 _20220_ (.A(net872),
    .X(_03019_));
 sg13g2_buf_1 _20221_ (.A(net744),
    .X(_03020_));
 sg13g2_buf_1 _20222_ (.A(net534),
    .X(_03021_));
 sg13g2_buf_1 _20223_ (.A(net534),
    .X(_03022_));
 sg13g2_nand2_1 _20224_ (.Y(_03023_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net467));
 sg13g2_o21ai_1 _20225_ (.B1(_03023_),
    .Y(_00591_),
    .A1(_03020_),
    .A2(net468));
 sg13g2_mux2_1 _20226_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(_03021_),
    .X(_00592_));
 sg13g2_mux2_1 _20227_ (.A0(_09680_),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net468),
    .X(_00593_));
 sg13g2_mux2_1 _20228_ (.A0(net434),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net468),
    .X(_00594_));
 sg13g2_mux2_1 _20229_ (.A0(_09701_),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net468),
    .X(_00595_));
 sg13g2_mux2_1 _20230_ (.A0(net435),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net468),
    .X(_00596_));
 sg13g2_mux2_1 _20231_ (.A0(net433),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(_03021_),
    .X(_00597_));
 sg13g2_mux2_1 _20232_ (.A0(net427),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net468),
    .X(_00598_));
 sg13g2_mux2_1 _20233_ (.A0(net431),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net467),
    .X(_00599_));
 sg13g2_nand2_1 _20234_ (.Y(_03024_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(net534));
 sg13g2_o21ai_1 _20235_ (.B1(_03024_),
    .Y(_00600_),
    .A1(_09867_),
    .A2(net468));
 sg13g2_buf_1 _20236_ (.A(_10619_),
    .X(_03025_));
 sg13g2_buf_1 _20237_ (.A(_03025_),
    .X(_03026_));
 sg13g2_nand2_1 _20238_ (.Y(_03027_),
    .A(\cpu.dcache.r_tag[0][6] ),
    .B(_12153_));
 sg13g2_o21ai_1 _20239_ (.B1(_03027_),
    .Y(_00601_),
    .A1(_03026_),
    .A2(net468));
 sg13g2_buf_1 _20240_ (.A(net1069),
    .X(_03028_));
 sg13g2_buf_1 _20241_ (.A(net862),
    .X(_03029_));
 sg13g2_mux2_1 _20242_ (.A0(net742),
    .A1(\cpu.dcache.r_tag[0][7] ),
    .S(net467),
    .X(_00602_));
 sg13g2_buf_1 _20243_ (.A(net1070),
    .X(_03030_));
 sg13g2_buf_1 _20244_ (.A(net861),
    .X(_03031_));
 sg13g2_mux2_1 _20245_ (.A0(net741),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(net467),
    .X(_00603_));
 sg13g2_buf_1 _20246_ (.A(_10819_),
    .X(_03032_));
 sg13g2_buf_1 _20247_ (.A(net993),
    .X(_03033_));
 sg13g2_mux2_1 _20248_ (.A0(net860),
    .A1(\cpu.dcache.r_tag[0][9] ),
    .S(net467),
    .X(_00604_));
 sg13g2_buf_1 _20249_ (.A(_10903_),
    .X(_03034_));
 sg13g2_buf_1 _20250_ (.A(net992),
    .X(_03035_));
 sg13g2_mux2_1 _20251_ (.A0(_03035_),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net467),
    .X(_00605_));
 sg13g2_buf_1 _20252_ (.A(_10925_),
    .X(_03036_));
 sg13g2_buf_1 _20253_ (.A(net991),
    .X(_03037_));
 sg13g2_mux2_1 _20254_ (.A0(_03037_),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net467),
    .X(_00606_));
 sg13g2_mux2_1 _20255_ (.A0(_09657_),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net467),
    .X(_00607_));
 sg13g2_mux2_1 _20256_ (.A0(net386),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(_03022_),
    .X(_00608_));
 sg13g2_mux2_1 _20257_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(_03022_),
    .X(_00609_));
 sg13g2_buf_1 _20258_ (.A(net662),
    .X(_03038_));
 sg13g2_buf_1 _20259_ (.A(net592),
    .X(_03039_));
 sg13g2_buf_1 _20260_ (.A(net533),
    .X(_03040_));
 sg13g2_mux2_1 _20261_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net526),
    .S(net466),
    .X(_00610_));
 sg13g2_mux2_1 _20262_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net432),
    .S(net466),
    .X(_00611_));
 sg13g2_mux2_1 _20263_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net429),
    .S(net466),
    .X(_00612_));
 sg13g2_mux2_1 _20264_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net434),
    .S(net466),
    .X(_00613_));
 sg13g2_mux2_1 _20265_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net428),
    .S(net466),
    .X(_00614_));
 sg13g2_mux2_1 _20266_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net435),
    .S(_03040_),
    .X(_00615_));
 sg13g2_mux2_1 _20267_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net433),
    .S(net466),
    .X(_00616_));
 sg13g2_mux2_1 _20268_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net427),
    .S(_03040_),
    .X(_00617_));
 sg13g2_mux2_1 _20269_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net431),
    .S(net466),
    .X(_00618_));
 sg13g2_buf_1 _20270_ (.A(_12292_),
    .X(_03041_));
 sg13g2_mux2_1 _20271_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(_09426_),
    .S(net525),
    .X(_00619_));
 sg13g2_buf_1 _20272_ (.A(net1071),
    .X(_03042_));
 sg13g2_buf_1 _20273_ (.A(net857),
    .X(_03043_));
 sg13g2_mux2_1 _20274_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net740),
    .S(_03041_),
    .X(_00620_));
 sg13g2_buf_1 _20275_ (.A(net862),
    .X(_03044_));
 sg13g2_mux2_1 _20276_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net739),
    .S(net525),
    .X(_00621_));
 sg13g2_buf_1 _20277_ (.A(net861),
    .X(_03045_));
 sg13g2_mux2_1 _20278_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net738),
    .S(net525),
    .X(_00622_));
 sg13g2_buf_1 _20279_ (.A(net993),
    .X(_03046_));
 sg13g2_mux2_1 _20280_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net856),
    .S(net525),
    .X(_00623_));
 sg13g2_nand2_1 _20281_ (.Y(_03047_),
    .A(net992),
    .B(net525));
 sg13g2_o21ai_1 _20282_ (.B1(_03047_),
    .Y(_00624_),
    .A1(_09786_),
    .A2(net466));
 sg13g2_buf_1 _20283_ (.A(net991),
    .X(_03048_));
 sg13g2_mux2_1 _20284_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net855),
    .S(net525),
    .X(_00625_));
 sg13g2_mux2_1 _20285_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net385),
    .S(net525),
    .X(_00626_));
 sg13g2_mux2_1 _20286_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net386),
    .S(net525),
    .X(_00627_));
 sg13g2_mux2_1 _20287_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net430),
    .S(_03041_),
    .X(_00628_));
 sg13g2_buf_1 _20288_ (.A(_12424_),
    .X(_03049_));
 sg13g2_mux2_1 _20289_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net526),
    .S(net422),
    .X(_00629_));
 sg13g2_mux2_1 _20290_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net432),
    .S(_03049_),
    .X(_00630_));
 sg13g2_mux2_1 _20291_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net429),
    .S(net422),
    .X(_00631_));
 sg13g2_mux2_1 _20292_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net434),
    .S(net422),
    .X(_00632_));
 sg13g2_mux2_1 _20293_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net428),
    .S(net422),
    .X(_00633_));
 sg13g2_mux2_1 _20294_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net435),
    .S(net422),
    .X(_00634_));
 sg13g2_mux2_1 _20295_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net433),
    .S(_03049_),
    .X(_00635_));
 sg13g2_mux2_1 _20296_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net427),
    .S(net422),
    .X(_00636_));
 sg13g2_mux2_1 _20297_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net431),
    .S(net422),
    .X(_00637_));
 sg13g2_mux2_1 _20298_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(_09426_),
    .S(net422),
    .X(_00638_));
 sg13g2_buf_1 _20299_ (.A(_12424_),
    .X(_03050_));
 sg13g2_mux2_1 _20300_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net740),
    .S(_03050_),
    .X(_00639_));
 sg13g2_mux2_1 _20301_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net739),
    .S(net421),
    .X(_00640_));
 sg13g2_mux2_1 _20302_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(_03045_),
    .S(net421),
    .X(_00641_));
 sg13g2_mux2_1 _20303_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net856),
    .S(net421),
    .X(_00642_));
 sg13g2_buf_1 _20304_ (.A(net992),
    .X(_03051_));
 sg13g2_mux2_1 _20305_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net854),
    .S(net421),
    .X(_00643_));
 sg13g2_mux2_1 _20306_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net855),
    .S(net421),
    .X(_00644_));
 sg13g2_mux2_1 _20307_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net385),
    .S(net421),
    .X(_00645_));
 sg13g2_mux2_1 _20308_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net386),
    .S(net421),
    .X(_00646_));
 sg13g2_mux2_1 _20309_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net430),
    .S(_03050_),
    .X(_00647_));
 sg13g2_buf_1 _20310_ (.A(_12546_),
    .X(_03052_));
 sg13g2_mux2_1 _20311_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net526),
    .S(net420),
    .X(_00648_));
 sg13g2_mux2_1 _20312_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net432),
    .S(_03052_),
    .X(_00649_));
 sg13g2_mux2_1 _20313_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net429),
    .S(net420),
    .X(_00650_));
 sg13g2_mux2_1 _20314_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net434),
    .S(net420),
    .X(_00651_));
 sg13g2_mux2_1 _20315_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net428),
    .S(net420),
    .X(_00652_));
 sg13g2_mux2_1 _20316_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(_09485_),
    .S(net420),
    .X(_00653_));
 sg13g2_mux2_1 _20317_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net433),
    .S(_03052_),
    .X(_00654_));
 sg13g2_mux2_1 _20318_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net427),
    .S(net420),
    .X(_00655_));
 sg13g2_mux2_1 _20319_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net431),
    .S(net420),
    .X(_00656_));
 sg13g2_mux2_1 _20320_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(_09426_),
    .S(net420),
    .X(_00657_));
 sg13g2_buf_1 _20321_ (.A(_12546_),
    .X(_03053_));
 sg13g2_mux2_1 _20322_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net740),
    .S(net419),
    .X(_00658_));
 sg13g2_mux2_1 _20323_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(_03044_),
    .S(net419),
    .X(_00659_));
 sg13g2_mux2_1 _20324_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(_03045_),
    .S(net419),
    .X(_00660_));
 sg13g2_mux2_1 _20325_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(_03046_),
    .S(net419),
    .X(_00661_));
 sg13g2_mux2_1 _20326_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net854),
    .S(net419),
    .X(_00662_));
 sg13g2_mux2_1 _20327_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(_03048_),
    .S(net419),
    .X(_00663_));
 sg13g2_mux2_1 _20328_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(_09657_),
    .S(_03053_),
    .X(_00664_));
 sg13g2_mux2_1 _20329_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net386),
    .S(net419),
    .X(_00665_));
 sg13g2_mux2_1 _20330_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net430),
    .S(_03053_),
    .X(_00666_));
 sg13g2_buf_1 _20331_ (.A(net335),
    .X(_03054_));
 sg13g2_nand2_1 _20332_ (.Y(_03055_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net335));
 sg13g2_o21ai_1 _20333_ (.B1(_03055_),
    .Y(_00667_),
    .A1(_03020_),
    .A2(net259));
 sg13g2_mux2_1 _20334_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net259),
    .X(_00668_));
 sg13g2_mux2_1 _20335_ (.A0(net429),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net259),
    .X(_00669_));
 sg13g2_mux2_1 _20336_ (.A0(net434),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(_03054_),
    .X(_00670_));
 sg13g2_mux2_1 _20337_ (.A0(_09701_),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net259),
    .X(_00671_));
 sg13g2_mux2_1 _20338_ (.A0(net435),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net259),
    .X(_00672_));
 sg13g2_mux2_1 _20339_ (.A0(_09543_),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(_03054_),
    .X(_00673_));
 sg13g2_buf_1 _20340_ (.A(net335),
    .X(_03056_));
 sg13g2_mux2_1 _20341_ (.A0(_09724_),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net258),
    .X(_00674_));
 sg13g2_mux2_1 _20342_ (.A0(net431),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net258),
    .X(_00675_));
 sg13g2_nand2_1 _20343_ (.Y(_03057_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(net335));
 sg13g2_o21ai_1 _20344_ (.B1(_03057_),
    .Y(_00676_),
    .A1(_09867_),
    .A2(net259));
 sg13g2_nand2_1 _20345_ (.Y(_03058_),
    .A(\cpu.dcache.r_tag[4][6] ),
    .B(_12667_));
 sg13g2_o21ai_1 _20346_ (.B1(_03058_),
    .Y(_00677_),
    .A1(net743),
    .A2(net259));
 sg13g2_mux2_1 _20347_ (.A0(net742),
    .A1(\cpu.dcache.r_tag[4][7] ),
    .S(net258),
    .X(_00678_));
 sg13g2_mux2_1 _20348_ (.A0(net741),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(net258),
    .X(_00679_));
 sg13g2_mux2_1 _20349_ (.A0(net860),
    .A1(\cpu.dcache.r_tag[4][9] ),
    .S(net258),
    .X(_00680_));
 sg13g2_mux2_1 _20350_ (.A0(net859),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(net258),
    .X(_00681_));
 sg13g2_mux2_1 _20351_ (.A0(_03037_),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net258),
    .X(_00682_));
 sg13g2_mux2_1 _20352_ (.A0(net385),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net258),
    .X(_00683_));
 sg13g2_mux2_1 _20353_ (.A0(net386),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(_03056_),
    .X(_00684_));
 sg13g2_mux2_1 _20354_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(_03056_),
    .X(_00685_));
 sg13g2_buf_1 _20355_ (.A(_02706_),
    .X(_03059_));
 sg13g2_mux2_1 _20356_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net526),
    .S(net418),
    .X(_00686_));
 sg13g2_mux2_1 _20357_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net432),
    .S(_03059_),
    .X(_00687_));
 sg13g2_mux2_1 _20358_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(_09680_),
    .S(net418),
    .X(_00688_));
 sg13g2_mux2_1 _20359_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(_09513_),
    .S(net418),
    .X(_00689_));
 sg13g2_mux2_1 _20360_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net428),
    .S(net418),
    .X(_00690_));
 sg13g2_mux2_1 _20361_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net435),
    .S(net418),
    .X(_00691_));
 sg13g2_mux2_1 _20362_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net433),
    .S(_03059_),
    .X(_00692_));
 sg13g2_mux2_1 _20363_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net427),
    .S(net418),
    .X(_00693_));
 sg13g2_mux2_1 _20364_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net431),
    .S(net418),
    .X(_00694_));
 sg13g2_mux2_1 _20365_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(_09426_),
    .S(net418),
    .X(_00695_));
 sg13g2_buf_1 _20366_ (.A(_02706_),
    .X(_03060_));
 sg13g2_mux2_1 _20367_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(net740),
    .S(_03060_),
    .X(_00696_));
 sg13g2_mux2_1 _20368_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(_03044_),
    .S(net417),
    .X(_00697_));
 sg13g2_mux2_1 _20369_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net738),
    .S(net417),
    .X(_00698_));
 sg13g2_mux2_1 _20370_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(_03046_),
    .S(net417),
    .X(_00699_));
 sg13g2_mux2_1 _20371_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(_03051_),
    .S(net417),
    .X(_00700_));
 sg13g2_mux2_1 _20372_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(_03048_),
    .S(net417),
    .X(_00701_));
 sg13g2_mux2_1 _20373_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net385),
    .S(net417),
    .X(_00702_));
 sg13g2_mux2_1 _20374_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net386),
    .S(net417),
    .X(_00703_));
 sg13g2_mux2_1 _20375_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net430),
    .S(_03060_),
    .X(_00704_));
 sg13g2_buf_1 _20376_ (.A(_02837_),
    .X(_03061_));
 sg13g2_mux2_1 _20377_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net526),
    .S(net465),
    .X(_00705_));
 sg13g2_mux2_1 _20378_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net432),
    .S(net465),
    .X(_00706_));
 sg13g2_mux2_1 _20379_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(net429),
    .S(net465),
    .X(_00707_));
 sg13g2_mux2_1 _20380_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(_09513_),
    .S(net465),
    .X(_00708_));
 sg13g2_mux2_1 _20381_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net428),
    .S(net465),
    .X(_00709_));
 sg13g2_mux2_1 _20382_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(_09485_),
    .S(_03061_),
    .X(_00710_));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net433),
    .S(_03061_),
    .X(_00711_));
 sg13g2_mux2_1 _20384_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net427),
    .S(net465),
    .X(_00712_));
 sg13g2_mux2_1 _20385_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(_09589_),
    .S(net465),
    .X(_00713_));
 sg13g2_mux2_1 _20386_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(_09426_),
    .S(net465),
    .X(_00714_));
 sg13g2_buf_1 _20387_ (.A(_02837_),
    .X(_03062_));
 sg13g2_mux2_1 _20388_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net740),
    .S(_03062_),
    .X(_00715_));
 sg13g2_buf_1 _20389_ (.A(net862),
    .X(_03063_));
 sg13g2_mux2_1 _20390_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net737),
    .S(net464),
    .X(_00716_));
 sg13g2_buf_1 _20391_ (.A(net861),
    .X(_03064_));
 sg13g2_mux2_1 _20392_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net736),
    .S(net464),
    .X(_00717_));
 sg13g2_buf_1 _20393_ (.A(net993),
    .X(_03065_));
 sg13g2_mux2_1 _20394_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net853),
    .S(net464),
    .X(_00718_));
 sg13g2_mux2_1 _20395_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(_03051_),
    .S(net464),
    .X(_00719_));
 sg13g2_buf_1 _20396_ (.A(net991),
    .X(_03066_));
 sg13g2_mux2_1 _20397_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(_03066_),
    .S(net464),
    .X(_00720_));
 sg13g2_mux2_1 _20398_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net385),
    .S(net464),
    .X(_00721_));
 sg13g2_mux2_1 _20399_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(_09642_),
    .S(net464),
    .X(_00722_));
 sg13g2_mux2_1 _20400_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net430),
    .S(_03062_),
    .X(_00723_));
 sg13g2_buf_1 _20401_ (.A(net423),
    .X(_03067_));
 sg13g2_mux2_1 _20402_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net526),
    .S(net383),
    .X(_00724_));
 sg13g2_mux2_1 _20403_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net432),
    .S(net383),
    .X(_00725_));
 sg13g2_mux2_1 _20404_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net429),
    .S(net383),
    .X(_00726_));
 sg13g2_mux2_1 _20405_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net434),
    .S(net383),
    .X(_00727_));
 sg13g2_mux2_1 _20406_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(net428),
    .S(net383),
    .X(_00728_));
 sg13g2_mux2_1 _20407_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net435),
    .S(_03067_),
    .X(_00729_));
 sg13g2_mux2_1 _20408_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net433),
    .S(net383),
    .X(_00730_));
 sg13g2_mux2_1 _20409_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(net427),
    .S(net383),
    .X(_00731_));
 sg13g2_mux2_1 _20410_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net431),
    .S(net383),
    .X(_00732_));
 sg13g2_mux2_1 _20411_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09426_),
    .S(_03067_),
    .X(_00733_));
 sg13g2_buf_1 _20412_ (.A(net423),
    .X(_03068_));
 sg13g2_mux2_1 _20413_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net740),
    .S(_03068_),
    .X(_00734_));
 sg13g2_mux2_1 _20414_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net737),
    .S(net382),
    .X(_00735_));
 sg13g2_mux2_1 _20415_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net736),
    .S(net382),
    .X(_00736_));
 sg13g2_mux2_1 _20416_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net853),
    .S(net382),
    .X(_00737_));
 sg13g2_buf_1 _20417_ (.A(net992),
    .X(_03069_));
 sg13g2_mux2_1 _20418_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(_03069_),
    .S(net382),
    .X(_00738_));
 sg13g2_mux2_1 _20419_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(_03066_),
    .S(net382),
    .X(_00739_));
 sg13g2_mux2_1 _20420_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net385),
    .S(net382),
    .X(_00740_));
 sg13g2_mux2_1 _20421_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(_09642_),
    .S(net382),
    .X(_00741_));
 sg13g2_mux2_1 _20422_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(net430),
    .S(_03068_),
    .X(_00742_));
 sg13g2_buf_1 _20423_ (.A(_08941_),
    .X(_03070_));
 sg13g2_buf_1 _20424_ (.A(net220),
    .X(_03071_));
 sg13g2_buf_1 _20425_ (.A(_09898_),
    .X(_03072_));
 sg13g2_nand2_1 _20426_ (.Y(_03073_),
    .A(net219),
    .B(_09900_));
 sg13g2_buf_1 _20427_ (.A(_03073_),
    .X(_03074_));
 sg13g2_buf_1 _20428_ (.A(net347),
    .X(_03075_));
 sg13g2_buf_1 _20429_ (.A(net257),
    .X(_03076_));
 sg13g2_buf_1 _20430_ (.A(_09900_),
    .X(_03077_));
 sg13g2_buf_1 _20431_ (.A(net346),
    .X(_03078_));
 sg13g2_buf_1 _20432_ (.A(_08961_),
    .X(_03079_));
 sg13g2_nor2_1 _20433_ (.A(net270),
    .B(net216),
    .Y(_03080_));
 sg13g2_nor2_1 _20434_ (.A(net220),
    .B(net256),
    .Y(_03081_));
 sg13g2_a21oi_1 _20435_ (.A1(net256),
    .A2(_03080_),
    .Y(_03082_),
    .B1(_03081_));
 sg13g2_or3_1 _20436_ (.A(net218),
    .B(net217),
    .C(_03082_),
    .X(_03083_));
 sg13g2_o21ai_1 _20437_ (.B1(_03083_),
    .Y(_03084_),
    .A1(net204),
    .A2(net186));
 sg13g2_buf_1 _20438_ (.A(net174),
    .X(_03085_));
 sg13g2_mux2_1 _20439_ (.A0(_03084_),
    .A1(_10373_),
    .S(net131),
    .X(_00751_));
 sg13g2_buf_1 _20440_ (.A(net219),
    .X(_03086_));
 sg13g2_buf_1 _20441_ (.A(_08994_),
    .X(_03087_));
 sg13g2_o21ai_1 _20442_ (.B1(net202),
    .Y(_03088_),
    .A1(net204),
    .A2(_03086_));
 sg13g2_buf_1 _20443_ (.A(_08977_),
    .X(_03089_));
 sg13g2_buf_1 _20444_ (.A(net215),
    .X(_03090_));
 sg13g2_nand2_1 _20445_ (.Y(_03091_),
    .A(net257),
    .B(net201));
 sg13g2_buf_1 _20446_ (.A(_09901_),
    .X(_03092_));
 sg13g2_nand2_2 _20447_ (.Y(_03093_),
    .A(_09900_),
    .B(_03092_));
 sg13g2_o21ai_1 _20448_ (.B1(_03093_),
    .Y(_03094_),
    .A1(net343),
    .A2(_03091_));
 sg13g2_buf_1 _20449_ (.A(net216),
    .X(_03095_));
 sg13g2_nor2_1 _20450_ (.A(_03095_),
    .B(_03093_),
    .Y(_03096_));
 sg13g2_a221oi_1 _20451_ (.B2(net204),
    .C1(_03096_),
    .B1(_03094_),
    .A1(net231),
    .Y(_03097_),
    .A2(_03088_));
 sg13g2_buf_1 _20452_ (.A(_11945_),
    .X(_03098_));
 sg13g2_buf_1 _20453_ (.A(net850),
    .X(_03099_));
 sg13g2_nand2_1 _20454_ (.Y(_03100_),
    .A(_03099_),
    .B(net138));
 sg13g2_o21ai_1 _20455_ (.B1(_03100_),
    .Y(_00752_),
    .A1(net107),
    .A2(_03097_));
 sg13g2_nor2_1 _20456_ (.A(net216),
    .B(net215),
    .Y(_03101_));
 sg13g2_buf_2 _20457_ (.A(_03101_),
    .X(_03102_));
 sg13g2_nand2_1 _20458_ (.Y(_03103_),
    .A(_09113_),
    .B(_03102_));
 sg13g2_nand2_1 _20459_ (.Y(_03104_),
    .A(\cpu.cond[1] ),
    .B(_09941_));
 sg13g2_o21ai_1 _20460_ (.B1(_03104_),
    .Y(_00753_),
    .A1(_09121_),
    .A2(_03103_));
 sg13g2_a21oi_1 _20461_ (.A1(net204),
    .A2(net202),
    .Y(_03105_),
    .B1(net218));
 sg13g2_o21ai_1 _20462_ (.B1(_03105_),
    .Y(_03106_),
    .A1(net204),
    .A2(net186));
 sg13g2_nand2_1 _20463_ (.Y(_03107_),
    .A(\cpu.cond[2] ),
    .B(net138));
 sg13g2_o21ai_1 _20464_ (.B1(_03107_),
    .Y(_00754_),
    .A1(net107),
    .A2(_03106_));
 sg13g2_nand3_1 _20465_ (.B(_09118_),
    .C(_09134_),
    .A(net142),
    .Y(_03108_));
 sg13g2_o21ai_1 _20466_ (.B1(_03108_),
    .Y(_00755_),
    .A1(_09378_),
    .A2(net108));
 sg13g2_nand2_1 _20467_ (.Y(_03109_),
    .A(net194),
    .B(_09928_));
 sg13g2_nand2b_1 _20468_ (.Y(_03110_),
    .B(net547),
    .A_N(_00175_));
 sg13g2_mux2_1 _20469_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net802),
    .X(_03111_));
 sg13g2_a22oi_1 _20470_ (.Y(_03112_),
    .B1(_03111_),
    .B2(_08810_),
    .A2(net921),
    .A1(\cpu.icache.r_data[5][24] ));
 sg13g2_nand2b_1 _20471_ (.Y(_03113_),
    .B(_08534_),
    .A_N(_03112_));
 sg13g2_buf_1 _20472_ (.A(net634),
    .X(_03114_));
 sg13g2_buf_1 _20473_ (.A(net550),
    .X(_03115_));
 sg13g2_a22oi_1 _20474_ (.Y(_03116_),
    .B1(net463),
    .B2(\cpu.icache.r_data[2][24] ),
    .A2(net524),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_buf_1 _20475_ (.A(net628),
    .X(_03117_));
 sg13g2_buf_1 _20476_ (.A(_08511_),
    .X(_03118_));
 sg13g2_a22oi_1 _20477_ (.Y(_03119_),
    .B1(net522),
    .B2(\cpu.icache.r_data[4][24] ),
    .A2(net523),
    .A1(\cpu.icache.r_data[6][24] ));
 sg13g2_nand4_1 _20478_ (.B(_03113_),
    .C(_03116_),
    .A(_03110_),
    .Y(_03120_),
    .D(_03119_));
 sg13g2_nand2_1 _20479_ (.Y(_03121_),
    .A(_00174_),
    .B(net547));
 sg13g2_a22oi_1 _20480_ (.Y(_03122_),
    .B1(_08511_),
    .B2(\cpu.icache.r_data[4][8] ),
    .A2(_08506_),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_a22oi_1 _20481_ (.Y(_03123_),
    .B1(net546),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(_08516_),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_mux2_1 _20482_ (.A0(\cpu.icache.r_data[5][8] ),
    .A1(\cpu.icache.r_data[7][8] ),
    .S(net813),
    .X(_03124_));
 sg13g2_a22oi_1 _20483_ (.Y(_03125_),
    .B1(_03124_),
    .B2(_08534_),
    .A2(_08528_),
    .A1(\cpu.icache.r_data[6][8] ));
 sg13g2_or2_1 _20484_ (.X(_03126_),
    .B(_03125_),
    .A(_08525_));
 sg13g2_nand4_1 _20485_ (.B(_03122_),
    .C(_03123_),
    .A(_08500_),
    .Y(_03127_),
    .D(_03126_));
 sg13g2_a21o_1 _20486_ (.A2(_03127_),
    .A1(_03121_),
    .B1(net800),
    .X(_03128_));
 sg13g2_o21ai_1 _20487_ (.B1(_03128_),
    .Y(_03129_),
    .A1(net1077),
    .A2(_03120_));
 sg13g2_buf_1 _20488_ (.A(_03129_),
    .X(_03130_));
 sg13g2_buf_1 _20489_ (.A(_03130_),
    .X(_03131_));
 sg13g2_nand2b_1 _20490_ (.Y(_03132_),
    .B(net627),
    .A_N(_00177_));
 sg13g2_mux2_1 _20491_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(\cpu.icache.r_data[7][25] ),
    .S(net813),
    .X(_03133_));
 sg13g2_a22oi_1 _20492_ (.Y(_03134_),
    .B1(_03133_),
    .B2(net801),
    .A2(net814),
    .A1(\cpu.icache.r_data[6][25] ));
 sg13g2_or2_1 _20493_ (.X(_03135_),
    .B(_03134_),
    .A(net815));
 sg13g2_a22oi_1 _20494_ (.Y(_03136_),
    .B1(net635),
    .B2(\cpu.icache.r_data[4][25] ),
    .A2(net549),
    .A1(\cpu.icache.r_data[3][25] ));
 sg13g2_a22oi_1 _20495_ (.Y(_03137_),
    .B1(net550),
    .B2(\cpu.icache.r_data[2][25] ),
    .A2(net630),
    .A1(\cpu.icache.r_data[1][25] ));
 sg13g2_nand4_1 _20496_ (.B(_03135_),
    .C(_03136_),
    .A(_03132_),
    .Y(_03138_),
    .D(_03137_));
 sg13g2_nand2_1 _20497_ (.Y(_03139_),
    .A(_00176_),
    .B(net627));
 sg13g2_a22oi_1 _20498_ (.Y(_03140_),
    .B1(_08510_),
    .B2(\cpu.icache.r_data[4][9] ),
    .A2(_08505_),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_a22oi_1 _20499_ (.Y(_03141_),
    .B1(_08521_),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(_08515_),
    .A1(\cpu.icache.r_data[1][9] ));
 sg13g2_mux2_1 _20500_ (.A0(\cpu.icache.r_data[5][9] ),
    .A1(\cpu.icache.r_data[7][9] ),
    .S(net929),
    .X(_03142_));
 sg13g2_a22oi_1 _20501_ (.Y(_03143_),
    .B1(_03142_),
    .B2(net928),
    .A2(_08528_),
    .A1(\cpu.icache.r_data[6][9] ));
 sg13g2_or2_1 _20502_ (.X(_03144_),
    .B(_03143_),
    .A(_08719_));
 sg13g2_nand4_1 _20503_ (.B(_03140_),
    .C(_03141_),
    .A(_08499_),
    .Y(_03145_),
    .D(_03144_));
 sg13g2_a21o_1 _20504_ (.A2(_03145_),
    .A1(_03139_),
    .B1(_08899_),
    .X(_03146_));
 sg13g2_o21ai_1 _20505_ (.B1(_03146_),
    .Y(_03147_),
    .A1(_09006_),
    .A2(_03138_));
 sg13g2_buf_2 _20506_ (.A(_03147_),
    .X(_03148_));
 sg13g2_a22oi_1 _20507_ (.Y(_03149_),
    .B1(net699),
    .B2(\cpu.icache.r_data[6][7] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_a22oi_1 _20508_ (.Y(_03150_),
    .B1(_08509_),
    .B2(\cpu.icache.r_data[4][7] ),
    .A2(net709),
    .A1(\cpu.icache.r_data[1][7] ));
 sg13g2_mux2_1 _20509_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_08595_),
    .X(_03151_));
 sg13g2_a22oi_1 _20510_ (.Y(_03152_),
    .B1(_03151_),
    .B2(_08531_),
    .A2(_08875_),
    .A1(\cpu.icache.r_data[5][7] ));
 sg13g2_nand2b_1 _20511_ (.Y(_03153_),
    .B(net801),
    .A_N(_03152_));
 sg13g2_and4_1 _20512_ (.A(net551),
    .B(_03149_),
    .C(_03150_),
    .D(_03153_),
    .X(_03154_));
 sg13g2_a21oi_1 _20513_ (.A1(_00172_),
    .A2(net547),
    .Y(_03155_),
    .B1(_03154_));
 sg13g2_nand2b_1 _20514_ (.Y(_03156_),
    .B(net627),
    .A_N(_00173_));
 sg13g2_a22oi_1 _20515_ (.Y(_03157_),
    .B1(_08506_),
    .B2(\cpu.icache.r_data[2][23] ),
    .A2(_08516_),
    .A1(\cpu.icache.r_data[1][23] ));
 sg13g2_mux4_1 _20516_ (.S0(net928),
    .A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[5][23] ),
    .A2(\cpu.icache.r_data[6][23] ),
    .A3(\cpu.icache.r_data[7][23] ),
    .S1(_08617_),
    .X(_03158_));
 sg13g2_a22oi_1 _20517_ (.Y(_03159_),
    .B1(_03158_),
    .B2(_08619_),
    .A2(_08522_),
    .A1(\cpu.icache.r_data[3][23] ));
 sg13g2_nand4_1 _20518_ (.B(_03156_),
    .C(_03157_),
    .A(_08919_),
    .Y(_03160_),
    .D(_03159_));
 sg13g2_o21ai_1 _20519_ (.B1(_03160_),
    .Y(_03161_),
    .A1(net920),
    .A2(_03155_));
 sg13g2_buf_1 _20520_ (.A(_03161_),
    .X(_03162_));
 sg13g2_nand3_1 _20521_ (.B(_03148_),
    .C(_03162_),
    .A(net214),
    .Y(_03163_));
 sg13g2_buf_1 _20522_ (.A(_03163_),
    .X(_03164_));
 sg13g2_or3_1 _20523_ (.A(_09893_),
    .B(_03109_),
    .C(_03164_),
    .X(_03165_));
 sg13g2_buf_1 _20524_ (.A(_03165_),
    .X(_03166_));
 sg13g2_nand3b_1 _20525_ (.B(net272),
    .C(_09134_),
    .Y(_03167_),
    .A_N(_03166_));
 sg13g2_nand2_1 _20526_ (.Y(_03168_),
    .A(\cpu.dec.do_flush_all ),
    .B(_09941_));
 sg13g2_o21ai_1 _20527_ (.B1(_03168_),
    .Y(_00756_),
    .A1(net107),
    .A2(_03167_));
 sg13g2_nand2_1 _20528_ (.Y(_03169_),
    .A(_08918_),
    .B(_09930_));
 sg13g2_buf_1 _20529_ (.A(_03169_),
    .X(_03170_));
 sg13g2_nand2_1 _20530_ (.Y(_03171_),
    .A(net215),
    .B(net334));
 sg13g2_nor4_1 _20531_ (.A(_08896_),
    .B(net200),
    .C(_03170_),
    .D(_03171_),
    .Y(_03172_));
 sg13g2_a21o_1 _20532_ (.A2(net143),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03172_),
    .X(_00757_));
 sg13g2_nand2_1 _20533_ (.Y(_03173_),
    .A(_08918_),
    .B(_08941_));
 sg13g2_buf_1 _20534_ (.A(_03173_),
    .X(_03174_));
 sg13g2_nor2_1 _20535_ (.A(net217),
    .B(_03174_),
    .Y(_03175_));
 sg13g2_nand3_1 _20536_ (.B(_03078_),
    .C(net186),
    .A(_08943_),
    .Y(_03176_));
 sg13g2_nand2b_1 _20537_ (.Y(_03177_),
    .B(_03176_),
    .A_N(_03175_));
 sg13g2_nand2_1 _20538_ (.Y(_03178_),
    .A(_09901_),
    .B(_09157_));
 sg13g2_o21ai_1 _20539_ (.B1(net257),
    .Y(_03179_),
    .A1(_03090_),
    .A2(_03178_));
 sg13g2_nor2_1 _20540_ (.A(net219),
    .B(_09191_),
    .Y(_03180_));
 sg13g2_o21ai_1 _20541_ (.B1(net194),
    .Y(_03181_),
    .A1(net200),
    .A2(net341));
 sg13g2_nor3_1 _20542_ (.A(net202),
    .B(_03180_),
    .C(_03181_),
    .Y(_03182_));
 sg13g2_a221oi_1 _20543_ (.B2(_03071_),
    .C1(_03182_),
    .B1(_03179_),
    .A1(net341),
    .Y(_03183_),
    .A2(_03177_));
 sg13g2_nor2_1 _20544_ (.A(net347),
    .B(net270),
    .Y(_03184_));
 sg13g2_buf_1 _20545_ (.A(_03184_),
    .X(_03185_));
 sg13g2_o21ai_1 _20546_ (.B1(net199),
    .Y(_03186_),
    .A1(_09124_),
    .A2(_03093_));
 sg13g2_nand2b_1 _20547_ (.Y(_03187_),
    .B(_03186_),
    .A_N(_03183_));
 sg13g2_nand2_1 _20548_ (.Y(_03188_),
    .A(_11088_),
    .B(net138));
 sg13g2_o21ai_1 _20549_ (.B1(_03188_),
    .Y(_00758_),
    .A1(_08897_),
    .A2(_03187_));
 sg13g2_inv_1 _20550_ (.Y(_03189_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_buf_1 _20551_ (.A(_09120_),
    .X(_03190_));
 sg13g2_nor2_1 _20552_ (.A(_03072_),
    .B(net334),
    .Y(_03191_));
 sg13g2_buf_1 _20553_ (.A(_03191_),
    .X(_03192_));
 sg13g2_inv_1 _20554_ (.Y(_03193_),
    .A(_08943_));
 sg13g2_a21oi_1 _20555_ (.A1(net272),
    .A2(_03192_),
    .Y(_03194_),
    .B1(_03193_));
 sg13g2_buf_1 _20556_ (.A(_03194_),
    .X(_03195_));
 sg13g2_nand2_1 _20557_ (.Y(_03196_),
    .A(net216),
    .B(net346));
 sg13g2_o21ai_1 _20558_ (.B1(_03196_),
    .Y(_03197_),
    .A1(net214),
    .A2(_03171_));
 sg13g2_nor2_2 _20559_ (.A(_09898_),
    .B(_08977_),
    .Y(_03198_));
 sg13g2_nand2_1 _20560_ (.Y(_03199_),
    .A(net334),
    .B(_03198_));
 sg13g2_buf_1 _20561_ (.A(_03199_),
    .X(_03200_));
 sg13g2_nand2_1 _20562_ (.Y(_03201_),
    .A(net274),
    .B(_03102_));
 sg13g2_buf_2 _20563_ (.A(_03201_),
    .X(_03202_));
 sg13g2_o21ai_1 _20564_ (.B1(_03202_),
    .Y(_03203_),
    .A1(net272),
    .A2(net185));
 sg13g2_nor2_1 _20565_ (.A(_03170_),
    .B(_09928_),
    .Y(_03204_));
 sg13g2_buf_1 _20566_ (.A(_03204_),
    .X(_03205_));
 sg13g2_or2_1 _20567_ (.X(_03206_),
    .B(net129),
    .A(net130));
 sg13g2_a22oi_1 _20568_ (.Y(_03207_),
    .B1(_03203_),
    .B2(_03206_),
    .A2(_03197_),
    .A1(net130));
 sg13g2_nand2_1 _20569_ (.Y(_03208_),
    .A(net346),
    .B(_09157_));
 sg13g2_o21ai_1 _20570_ (.B1(_03208_),
    .Y(_03209_),
    .A1(_08993_),
    .A2(_09911_));
 sg13g2_nand2_1 _20571_ (.Y(_03210_),
    .A(_03089_),
    .B(_03178_));
 sg13g2_o21ai_1 _20572_ (.B1(_03210_),
    .Y(_03211_),
    .A1(net215),
    .A2(_03209_));
 sg13g2_nor3_1 _20573_ (.A(_03072_),
    .B(_03174_),
    .C(_03211_),
    .Y(_03212_));
 sg13g2_inv_1 _20574_ (.Y(_03213_),
    .A(_03148_));
 sg13g2_nor2_1 _20575_ (.A(_09900_),
    .B(net346),
    .Y(_03214_));
 sg13g2_nand2_1 _20576_ (.Y(_03215_),
    .A(_03213_),
    .B(_03214_));
 sg13g2_nand2_1 _20577_ (.Y(_03216_),
    .A(net346),
    .B(_09107_));
 sg13g2_o21ai_1 _20578_ (.B1(_03216_),
    .Y(_03217_),
    .A1(net346),
    .A2(_09069_));
 sg13g2_a22oi_1 _20579_ (.Y(_03218_),
    .B1(_03217_),
    .B2(net217),
    .A2(net273),
    .A1(_08996_));
 sg13g2_nand2_1 _20580_ (.Y(_03219_),
    .A(_08961_),
    .B(_09902_));
 sg13g2_nand2_1 _20581_ (.Y(_03220_),
    .A(_03219_),
    .B(_03184_));
 sg13g2_a21oi_1 _20582_ (.A1(_03215_),
    .A2(_03218_),
    .Y(_03221_),
    .B1(_03220_));
 sg13g2_nor3_1 _20583_ (.A(_08895_),
    .B(_03212_),
    .C(_03221_),
    .Y(_03222_));
 sg13g2_buf_2 _20584_ (.A(_03222_),
    .X(_03223_));
 sg13g2_a22oi_1 _20585_ (.Y(_00759_),
    .B1(_03207_),
    .B2(_03223_),
    .A2(net102),
    .A1(_03189_));
 sg13g2_inv_1 _20586_ (.Y(_03224_),
    .A(\cpu.dec.imm[11] ));
 sg13g2_inv_1 _20587_ (.Y(_03225_),
    .A(_03162_));
 sg13g2_or4_1 _20588_ (.A(_09034_),
    .B(_03130_),
    .C(_03213_),
    .D(_03225_),
    .X(_03226_));
 sg13g2_buf_1 _20589_ (.A(_03226_),
    .X(_03227_));
 sg13g2_nor3_2 _20590_ (.A(_09898_),
    .B(_08977_),
    .C(_08993_),
    .Y(_03228_));
 sg13g2_o21ai_1 _20591_ (.B1(_03228_),
    .Y(_03229_),
    .A1(_09158_),
    .A2(_03227_));
 sg13g2_buf_1 _20592_ (.A(_03229_),
    .X(_03230_));
 sg13g2_buf_1 _20593_ (.A(_03227_),
    .X(_03231_));
 sg13g2_and2_1 _20594_ (.A(net389),
    .B(net184),
    .X(_03232_));
 sg13g2_o21ai_1 _20595_ (.B1(net334),
    .Y(_03233_),
    .A1(net390),
    .A2(_03198_));
 sg13g2_o21ai_1 _20596_ (.B1(net219),
    .Y(_03234_),
    .A1(_09902_),
    .A2(net343));
 sg13g2_nand2_1 _20597_ (.Y(_03235_),
    .A(_03233_),
    .B(_03234_));
 sg13g2_o21ai_1 _20598_ (.B1(_03235_),
    .Y(_03236_),
    .A1(_03230_),
    .A2(_03232_));
 sg13g2_o21ai_1 _20599_ (.B1(_03202_),
    .Y(_03237_),
    .A1(net389),
    .A2(net185));
 sg13g2_a22oi_1 _20600_ (.Y(_03238_),
    .B1(_03237_),
    .B2(_03205_),
    .A2(_03236_),
    .A1(net130));
 sg13g2_a22oi_1 _20601_ (.Y(_00760_),
    .B1(_03223_),
    .B2(_03238_),
    .A2(net102),
    .A1(_03224_));
 sg13g2_and2_1 _20602_ (.A(_09137_),
    .B(net184),
    .X(_03239_));
 sg13g2_o21ai_1 _20603_ (.B1(_03235_),
    .Y(_03240_),
    .A1(_03230_),
    .A2(_03239_));
 sg13g2_o21ai_1 _20604_ (.B1(_03202_),
    .Y(_03241_),
    .A1(_09137_),
    .A2(net185));
 sg13g2_a22oi_1 _20605_ (.Y(_03242_),
    .B1(_03241_),
    .B2(net129),
    .A2(_03240_),
    .A1(net130));
 sg13g2_a22oi_1 _20606_ (.Y(_00761_),
    .B1(_03223_),
    .B2(_03242_),
    .A2(net102),
    .A1(_11416_));
 sg13g2_inv_1 _20607_ (.Y(_03243_),
    .A(\cpu.dec.imm[13] ));
 sg13g2_and2_1 _20608_ (.A(net343),
    .B(net184),
    .X(_03244_));
 sg13g2_o21ai_1 _20609_ (.B1(_03235_),
    .Y(_03245_),
    .A1(_03230_),
    .A2(_03244_));
 sg13g2_a21oi_1 _20610_ (.A1(net186),
    .A2(net185),
    .Y(_03246_),
    .B1(net343));
 sg13g2_a22oi_1 _20611_ (.Y(_03247_),
    .B1(_03246_),
    .B2(net129),
    .A2(_03245_),
    .A1(net130));
 sg13g2_a22oi_1 _20612_ (.Y(_00762_),
    .B1(_03223_),
    .B2(_03247_),
    .A2(_03190_),
    .A1(_03243_));
 sg13g2_inv_1 _20613_ (.Y(_03248_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_o21ai_1 _20614_ (.B1(_03202_),
    .Y(_03249_),
    .A1(_09892_),
    .A2(net185));
 sg13g2_nand2_1 _20615_ (.Y(_03250_),
    .A(net129),
    .B(_03249_));
 sg13g2_and2_1 _20616_ (.A(_09892_),
    .B(net184),
    .X(_03251_));
 sg13g2_o21ai_1 _20617_ (.B1(_03235_),
    .Y(_03252_),
    .A1(_03230_),
    .A2(_03251_));
 sg13g2_inv_1 _20618_ (.Y(_03253_),
    .A(_03223_));
 sg13g2_a21oi_1 _20619_ (.A1(net130),
    .A2(_03252_),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_a22oi_1 _20620_ (.Y(_00763_),
    .B1(_03250_),
    .B2(_03254_),
    .A2(net102),
    .A1(_03248_));
 sg13g2_inv_1 _20621_ (.Y(_03255_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_o21ai_1 _20622_ (.B1(_03202_),
    .Y(_03256_),
    .A1(net345),
    .A2(net185));
 sg13g2_nand2_1 _20623_ (.Y(_03257_),
    .A(net129),
    .B(_03256_));
 sg13g2_a22oi_1 _20624_ (.Y(_00764_),
    .B1(_03254_),
    .B2(_03257_),
    .A2(net102),
    .A1(_03255_));
 sg13g2_o21ai_1 _20625_ (.B1(net334),
    .Y(_03258_),
    .A1(net215),
    .A2(_03231_));
 sg13g2_buf_1 _20626_ (.A(_03214_),
    .X(_03259_));
 sg13g2_nor2_1 _20627_ (.A(net215),
    .B(net334),
    .Y(_03260_));
 sg13g2_a21o_1 _20628_ (.A2(net198),
    .A1(net347),
    .B1(_03260_),
    .X(_03261_));
 sg13g2_a21oi_1 _20629_ (.A1(net231),
    .A2(_03258_),
    .Y(_03262_),
    .B1(_03261_));
 sg13g2_nor2_1 _20630_ (.A(net220),
    .B(_08996_),
    .Y(_03263_));
 sg13g2_o21ai_1 _20631_ (.B1(_03263_),
    .Y(_03264_),
    .A1(net203),
    .A2(_03262_));
 sg13g2_nand2_1 _20632_ (.Y(_03265_),
    .A(_09089_),
    .B(_03264_));
 sg13g2_buf_1 _20633_ (.A(net270),
    .X(_03266_));
 sg13g2_nor2_1 _20634_ (.A(net347),
    .B(net346),
    .Y(_03267_));
 sg13g2_a21oi_1 _20635_ (.A1(net257),
    .A2(_03192_),
    .Y(_03268_),
    .B1(_03267_));
 sg13g2_o21ai_1 _20636_ (.B1(net186),
    .Y(_03269_),
    .A1(net217),
    .A2(_03268_));
 sg13g2_nand3_1 _20637_ (.B(net342),
    .C(_03269_),
    .A(net213),
    .Y(_03270_));
 sg13g2_a21oi_1 _20638_ (.A1(_03265_),
    .A2(_03270_),
    .Y(_03271_),
    .B1(net141));
 sg13g2_a21o_1 _20639_ (.A2(net131),
    .A1(_11051_),
    .B1(_03271_),
    .X(_00765_));
 sg13g2_nand2_1 _20640_ (.Y(_03272_),
    .A(_08943_),
    .B(_03196_));
 sg13g2_nand2b_1 _20641_ (.Y(_03273_),
    .B(_03272_),
    .A_N(net129));
 sg13g2_nand3_1 _20642_ (.B(net342),
    .C(_03273_),
    .A(net173),
    .Y(_03274_));
 sg13g2_inv_1 _20643_ (.Y(_03275_),
    .A(_03272_));
 sg13g2_nor2_1 _20644_ (.A(net185),
    .B(net184),
    .Y(_03276_));
 sg13g2_nand3_1 _20645_ (.B(_03275_),
    .C(_03276_),
    .A(net341),
    .Y(_03277_));
 sg13g2_nand3_1 _20646_ (.B(net273),
    .C(_03269_),
    .A(net213),
    .Y(_03278_));
 sg13g2_nand3_1 _20647_ (.B(net216),
    .C(_03261_),
    .A(net270),
    .Y(_03279_));
 sg13g2_o21ai_1 _20648_ (.B1(net231),
    .Y(_03280_),
    .A1(_08941_),
    .A2(_03192_));
 sg13g2_nand2_1 _20649_ (.Y(_03281_),
    .A(_03279_),
    .B(_03280_));
 sg13g2_nand2_1 _20650_ (.Y(_03282_),
    .A(net216),
    .B(_03092_));
 sg13g2_mux2_1 _20651_ (.A0(_09035_),
    .A1(_09911_),
    .S(_03282_),
    .X(_03283_));
 sg13g2_nand2_1 _20652_ (.Y(_03284_),
    .A(_03077_),
    .B(net341));
 sg13g2_o21ai_1 _20653_ (.B1(_03284_),
    .Y(_03285_),
    .A1(net217),
    .A2(_03283_));
 sg13g2_a22oi_1 _20654_ (.Y(_03286_),
    .B1(_03285_),
    .B2(_09931_),
    .A2(_03281_),
    .A1(net230));
 sg13g2_nand4_1 _20655_ (.B(_03277_),
    .C(_03278_),
    .A(_03274_),
    .Y(_03287_),
    .D(_03286_));
 sg13g2_mux2_1 _20656_ (.A0(_03287_),
    .A1(_11010_),
    .S(net131),
    .X(_00766_));
 sg13g2_buf_1 _20657_ (.A(net142),
    .X(_03288_));
 sg13g2_nand2_1 _20658_ (.Y(_03289_),
    .A(_03079_),
    .B(_03214_));
 sg13g2_nand2_1 _20659_ (.Y(_03290_),
    .A(_03089_),
    .B(_03289_));
 sg13g2_a221oi_1 _20660_ (.B2(_09931_),
    .C1(_03281_),
    .B1(_03290_),
    .A1(_03275_),
    .Y(_03291_),
    .A2(_03276_));
 sg13g2_a22oi_1 _20661_ (.Y(_03292_),
    .B1(_03102_),
    .B2(net230),
    .A2(net273),
    .A1(_08996_));
 sg13g2_inv_1 _20662_ (.Y(_03293_),
    .A(_03292_));
 sg13g2_o21ai_1 _20663_ (.B1(_03109_),
    .Y(_03294_),
    .A1(_03171_),
    .A2(_03272_));
 sg13g2_nor3_1 _20664_ (.A(_09907_),
    .B(_03174_),
    .C(_03290_),
    .Y(_03295_));
 sg13g2_a221oi_1 _20665_ (.B2(net341),
    .C1(_03295_),
    .B1(_03294_),
    .A1(_03273_),
    .Y(_03296_),
    .A2(_03293_));
 sg13g2_o21ai_1 _20666_ (.B1(_03296_),
    .Y(_03297_),
    .A1(_09892_),
    .A2(_03291_));
 sg13g2_nand2_1 _20667_ (.Y(_03298_),
    .A(_03288_),
    .B(_03297_));
 sg13g2_o21ai_1 _20668_ (.B1(_03298_),
    .Y(_00767_),
    .A1(_10973_),
    .A2(_09052_));
 sg13g2_nor2_1 _20669_ (.A(_03102_),
    .B(net198),
    .Y(_03299_));
 sg13g2_o21ai_1 _20670_ (.B1(_03103_),
    .Y(_03300_),
    .A1(_03272_),
    .A2(_03299_));
 sg13g2_nand3_1 _20671_ (.B(net200),
    .C(_03258_),
    .A(net231),
    .Y(_03301_));
 sg13g2_a21oi_1 _20672_ (.A1(_03263_),
    .A2(_03301_),
    .Y(_03302_),
    .B1(net343));
 sg13g2_a21oi_1 _20673_ (.A1(net345),
    .A2(_03300_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_nand2_1 _20674_ (.Y(_03304_),
    .A(\cpu.dec.imm[4] ),
    .B(net138));
 sg13g2_o21ai_1 _20675_ (.B1(_03304_),
    .Y(_00768_),
    .A1(net143),
    .A2(_03303_));
 sg13g2_nand2_1 _20676_ (.Y(_03305_),
    .A(net217),
    .B(_03217_));
 sg13g2_o21ai_1 _20677_ (.B1(net341),
    .Y(_03306_),
    .A1(_09928_),
    .A2(net198));
 sg13g2_nand2_1 _20678_ (.Y(_03307_),
    .A(net173),
    .B(net271));
 sg13g2_nand4_1 _20679_ (.B(_03305_),
    .C(_03306_),
    .A(net199),
    .Y(_03308_),
    .D(_03307_));
 sg13g2_nand2_1 _20680_ (.Y(_03309_),
    .A(_03228_),
    .B(net184));
 sg13g2_a21oi_1 _20681_ (.A1(net271),
    .A2(_03309_),
    .Y(_03310_),
    .B1(net204));
 sg13g2_nand2_1 _20682_ (.Y(_03311_),
    .A(net186),
    .B(_03263_));
 sg13g2_nand3_1 _20683_ (.B(net271),
    .C(_03311_),
    .A(net218),
    .Y(_03312_));
 sg13g2_o21ai_1 _20684_ (.B1(_03312_),
    .Y(_03313_),
    .A1(net218),
    .A2(_03310_));
 sg13g2_nand3_1 _20685_ (.B(_03308_),
    .C(_03313_),
    .A(net142),
    .Y(_03314_));
 sg13g2_o21ai_1 _20686_ (.B1(_03314_),
    .Y(_00769_),
    .A1(_11121_),
    .A2(_09052_));
 sg13g2_nand3_1 _20687_ (.B(net201),
    .C(net333),
    .A(net200),
    .Y(_03315_));
 sg13g2_nand3_1 _20688_ (.B(_09911_),
    .C(_03305_),
    .A(_03086_),
    .Y(_03316_));
 sg13g2_a21oi_1 _20689_ (.A1(_03315_),
    .A2(_03316_),
    .Y(_03317_),
    .B1(net334));
 sg13g2_o21ai_1 _20690_ (.B1(net201),
    .Y(_03318_),
    .A1(net256),
    .A2(_03225_));
 sg13g2_nand2_1 _20691_ (.Y(_03319_),
    .A(_03305_),
    .B(_03318_));
 sg13g2_nand3b_1 _20692_ (.B(net199),
    .C(_03319_),
    .Y(_03320_),
    .A_N(_03317_));
 sg13g2_a22oi_1 _20693_ (.Y(_03321_),
    .B1(_03225_),
    .B2(net198),
    .A2(_03102_),
    .A1(net341));
 sg13g2_o21ai_1 _20694_ (.B1(net342),
    .Y(_03322_),
    .A1(_03192_),
    .A2(_03276_));
 sg13g2_a21oi_1 _20695_ (.A1(_03321_),
    .A2(_03322_),
    .Y(_03323_),
    .B1(_03193_));
 sg13g2_nand3_1 _20696_ (.B(net342),
    .C(_03290_),
    .A(_03071_),
    .Y(_03324_));
 sg13g2_nor2_1 _20697_ (.A(_08941_),
    .B(net215),
    .Y(_03325_));
 sg13g2_nand3_1 _20698_ (.B(net341),
    .C(_03325_),
    .A(net203),
    .Y(_03326_));
 sg13g2_a21oi_1 _20699_ (.A1(_03324_),
    .A2(_03326_),
    .Y(_03327_),
    .B1(net231));
 sg13g2_nor3_1 _20700_ (.A(net141),
    .B(_03323_),
    .C(_03327_),
    .Y(_03328_));
 sg13g2_a22oi_1 _20701_ (.Y(_00770_),
    .B1(_03320_),
    .B2(_03328_),
    .A2(net102),
    .A1(_11213_));
 sg13g2_o21ai_1 _20702_ (.B1(net203),
    .Y(_03329_),
    .A1(_09902_),
    .A2(_09137_));
 sg13g2_nand2_1 _20703_ (.Y(_03330_),
    .A(_03195_),
    .B(_03329_));
 sg13g2_o21ai_1 _20704_ (.B1(_03198_),
    .Y(_03331_),
    .A1(net272),
    .A2(_03231_));
 sg13g2_nand2_1 _20705_ (.Y(_03332_),
    .A(net201),
    .B(_09137_));
 sg13g2_a21oi_1 _20706_ (.A1(_03331_),
    .A2(_03332_),
    .Y(_03333_),
    .B1(net256));
 sg13g2_nor2_1 _20707_ (.A(net231),
    .B(net186),
    .Y(_03334_));
 sg13g2_nand2_1 _20708_ (.Y(_03335_),
    .A(net270),
    .B(_09089_));
 sg13g2_o21ai_1 _20709_ (.B1(_03335_),
    .Y(_03336_),
    .A1(net270),
    .A2(_03208_));
 sg13g2_nor2_1 _20710_ (.A(_09928_),
    .B(net198),
    .Y(_03337_));
 sg13g2_o21ai_1 _20711_ (.B1(_03218_),
    .Y(_03338_),
    .A1(net214),
    .A2(_03337_));
 sg13g2_a221oi_1 _20712_ (.B2(net199),
    .C1(_03212_),
    .B1(_03338_),
    .A1(_03334_),
    .Y(_03339_),
    .A2(_03336_));
 sg13g2_o21ai_1 _20713_ (.B1(_03339_),
    .Y(_03340_),
    .A1(_03330_),
    .A2(_03333_));
 sg13g2_mux2_1 _20714_ (.A0(_03340_),
    .A1(\cpu.dec.imm[7] ),
    .S(net131),
    .X(_00771_));
 sg13g2_inv_1 _20715_ (.Y(_03341_),
    .A(\cpu.dec.imm[8] ));
 sg13g2_nand2b_1 _20716_ (.Y(_03342_),
    .B(net184),
    .A_N(net271));
 sg13g2_nand2b_1 _20717_ (.Y(_03343_),
    .B(_03342_),
    .A_N(_03230_));
 sg13g2_a21oi_1 _20718_ (.A1(net274),
    .A2(_03102_),
    .Y(_03344_),
    .B1(_03192_));
 sg13g2_nand3_1 _20719_ (.B(_03343_),
    .C(_03344_),
    .A(_03215_),
    .Y(_03345_));
 sg13g2_nor2b_1 _20720_ (.A(_03148_),
    .B_N(net199),
    .Y(_03346_));
 sg13g2_nand2_1 _20721_ (.Y(_03347_),
    .A(net271),
    .B(_03228_));
 sg13g2_a21oi_1 _20722_ (.A1(_03202_),
    .A2(_03347_),
    .Y(_03348_),
    .B1(_03170_));
 sg13g2_a221oi_1 _20723_ (.B2(_09928_),
    .C1(_03348_),
    .B1(_03346_),
    .A1(net130),
    .Y(_03349_),
    .A2(_03345_));
 sg13g2_a22oi_1 _20724_ (.Y(_00772_),
    .B1(_03223_),
    .B2(_03349_),
    .A2(_03190_),
    .A1(_03341_));
 sg13g2_inv_1 _20725_ (.Y(_03350_),
    .A(\cpu.dec.imm[9] ));
 sg13g2_a21o_1 _20726_ (.A2(net184),
    .A1(_09911_),
    .B1(_03230_),
    .X(_03351_));
 sg13g2_nand2_1 _20727_ (.Y(_03352_),
    .A(net230),
    .B(_03259_));
 sg13g2_nand3_1 _20728_ (.B(_03351_),
    .C(_03352_),
    .A(_03344_),
    .Y(_03353_));
 sg13g2_o21ai_1 _20729_ (.B1(_03202_),
    .Y(_03354_),
    .A1(_09911_),
    .A2(net185));
 sg13g2_a22oi_1 _20730_ (.Y(_03355_),
    .B1(_03354_),
    .B2(net129),
    .A2(_03353_),
    .A1(net130));
 sg13g2_a22oi_1 _20731_ (.Y(_00773_),
    .B1(_03223_),
    .B2(_03355_),
    .A2(net102),
    .A1(_03350_));
 sg13g2_buf_1 _20732_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03356_));
 sg13g2_nand2_1 _20733_ (.Y(_03357_),
    .A(_08484_),
    .B(net390));
 sg13g2_nor4_1 _20734_ (.A(_08896_),
    .B(_09137_),
    .C(_03166_),
    .D(_03357_),
    .Y(_03358_));
 sg13g2_a21o_1 _20735_ (.A2(net131),
    .A1(_03356_),
    .B1(_03358_),
    .X(_00774_));
 sg13g2_nor2_1 _20736_ (.A(net198),
    .B(_03260_),
    .Y(_03359_));
 sg13g2_nor4_1 _20737_ (.A(net174),
    .B(net203),
    .C(_03170_),
    .D(_03359_),
    .Y(_03360_));
 sg13g2_a21o_1 _20738_ (.A2(_03085_),
    .A1(\cpu.dec.io ),
    .B1(_03360_),
    .X(_00775_));
 sg13g2_nand3_1 _20739_ (.B(_09906_),
    .C(_09198_),
    .A(_09109_),
    .Y(_03361_));
 sg13g2_buf_1 _20740_ (.A(_03361_),
    .X(_03362_));
 sg13g2_nor3_1 _20741_ (.A(_09904_),
    .B(_03174_),
    .C(_03362_),
    .Y(_03363_));
 sg13g2_mux2_1 _20742_ (.A0(_03363_),
    .A1(\cpu.dec.jmp ),
    .S(_03085_),
    .X(_00776_));
 sg13g2_o21ai_1 _20743_ (.B1(net201),
    .Y(_03364_),
    .A1(net257),
    .A2(net256));
 sg13g2_a22oi_1 _20744_ (.Y(_03365_),
    .B1(_03364_),
    .B2(net204),
    .A2(_03260_),
    .A1(net218));
 sg13g2_nor3_1 _20745_ (.A(net141),
    .B(net203),
    .C(_03365_),
    .Y(_03366_));
 sg13g2_a21o_1 _20746_ (.A2(net131),
    .A1(_11595_),
    .B1(_03366_),
    .X(_00777_));
 sg13g2_nand4_1 _20747_ (.B(net343),
    .C(_09109_),
    .A(net142),
    .Y(_03367_),
    .D(_09118_));
 sg13g2_o21ai_1 _20748_ (.B1(_03367_),
    .Y(_00778_),
    .A1(_09374_),
    .A2(net108));
 sg13g2_nor2_1 _20749_ (.A(net345),
    .B(net274),
    .Y(_03368_));
 sg13g2_nor3_1 _20750_ (.A(net257),
    .B(_09904_),
    .C(_03368_),
    .Y(_03369_));
 sg13g2_nand2_1 _20751_ (.Y(_03370_),
    .A(_09918_),
    .B(_03369_));
 sg13g2_nand3_1 _20752_ (.B(net219),
    .C(_09116_),
    .A(net270),
    .Y(_03371_));
 sg13g2_nand3_1 _20753_ (.B(_03095_),
    .C(net343),
    .A(net220),
    .Y(_03372_));
 sg13g2_nand4_1 _20754_ (.B(_09902_),
    .C(_03371_),
    .A(net218),
    .Y(_03373_),
    .D(_03372_));
 sg13g2_a21oi_1 _20755_ (.A1(_03370_),
    .A2(_03373_),
    .Y(_03374_),
    .B1(_03185_));
 sg13g2_nand2_1 _20756_ (.Y(_03375_),
    .A(net101),
    .B(_03374_));
 sg13g2_o21ai_1 _20757_ (.B1(_03375_),
    .Y(_00779_),
    .A1(net877),
    .A2(net108));
 sg13g2_and3_1 _20758_ (.X(_03376_),
    .A(net256),
    .B(_09113_),
    .C(net271));
 sg13g2_a221oi_1 _20759_ (.B2(_03198_),
    .C1(net199),
    .B1(_03376_),
    .A1(net274),
    .Y(_03377_),
    .A2(_03363_));
 sg13g2_a21oi_1 _20760_ (.A1(net333),
    .A2(_03171_),
    .Y(_03378_),
    .B1(net347));
 sg13g2_nor2_1 _20761_ (.A(_03093_),
    .B(net333),
    .Y(_03379_));
 sg13g2_o21ai_1 _20762_ (.B1(net200),
    .Y(_03380_),
    .A1(_03378_),
    .A2(_03379_));
 sg13g2_o21ai_1 _20763_ (.B1(_03380_),
    .Y(_03381_),
    .A1(_09904_),
    .A2(net333));
 sg13g2_inv_1 _20764_ (.Y(_03382_),
    .A(_03362_));
 sg13g2_nor2_1 _20765_ (.A(net202),
    .B(_03382_),
    .Y(_03383_));
 sg13g2_o21ai_1 _20766_ (.B1(_09931_),
    .Y(_03384_),
    .A1(net216),
    .A2(_03383_));
 sg13g2_inv_1 _20767_ (.Y(_03385_),
    .A(_03384_));
 sg13g2_a22oi_1 _20768_ (.Y(_03386_),
    .B1(_03385_),
    .B2(_03225_),
    .A2(_03381_),
    .A1(net213));
 sg13g2_a21o_1 _20769_ (.A2(net202),
    .A1(net203),
    .B1(_03180_),
    .X(_03387_));
 sg13g2_a221oi_1 _20770_ (.B2(_03185_),
    .C1(net141),
    .B1(_03387_),
    .A1(_03377_),
    .Y(_03388_),
    .A2(_03386_));
 sg13g2_a21o_1 _20771_ (.A2(net131),
    .A1(\cpu.dec.r_rd[0] ),
    .B1(_03388_),
    .X(_00780_));
 sg13g2_nand4_1 _20772_ (.B(_09137_),
    .C(net389),
    .A(_09125_),
    .Y(_03389_),
    .D(net273));
 sg13g2_nor3_1 _20773_ (.A(_09937_),
    .B(_03166_),
    .C(_03389_),
    .Y(_03390_));
 sg13g2_a21oi_1 _20774_ (.A1(net194),
    .A2(_03260_),
    .Y(_03391_),
    .B1(_03184_));
 sg13g2_nor3_1 _20775_ (.A(net203),
    .B(_09911_),
    .C(_03391_),
    .Y(_03392_));
 sg13g2_a21oi_1 _20776_ (.A1(_08943_),
    .A2(_03299_),
    .Y(_03393_),
    .B1(_03385_));
 sg13g2_o21ai_1 _20777_ (.B1(net129),
    .Y(_03394_),
    .A1(net173),
    .A2(_03228_));
 sg13g2_a21oi_1 _20778_ (.A1(_03393_),
    .A2(_03394_),
    .Y(_03395_),
    .B1(net214));
 sg13g2_nor3_1 _20779_ (.A(_03390_),
    .B(_03392_),
    .C(_03395_),
    .Y(_03396_));
 sg13g2_nand2_1 _20780_ (.Y(_03397_),
    .A(\cpu.dec.r_rd[1] ),
    .B(net138));
 sg13g2_o21ai_1 _20781_ (.B1(_03397_),
    .Y(_00781_),
    .A1(net143),
    .A2(_03396_));
 sg13g2_nor3_1 _20782_ (.A(net213),
    .B(net203),
    .C(net272),
    .Y(_03398_));
 sg13g2_o21ai_1 _20783_ (.B1(_03208_),
    .Y(_03399_),
    .A1(net256),
    .A2(_03148_));
 sg13g2_nor3_1 _20784_ (.A(net200),
    .B(net202),
    .C(_03148_),
    .Y(_03400_));
 sg13g2_a21o_1 _20785_ (.A2(_03399_),
    .A1(_03198_),
    .B1(_03400_),
    .X(_03401_));
 sg13g2_a22oi_1 _20786_ (.Y(_03402_),
    .B1(_03401_),
    .B2(net194),
    .A2(_03398_),
    .A1(net231));
 sg13g2_o21ai_1 _20787_ (.B1(_03402_),
    .Y(_03403_),
    .A1(_03148_),
    .A2(_03393_));
 sg13g2_mux2_1 _20788_ (.A0(_03403_),
    .A1(\cpu.dec.r_rd[2] ),
    .S(net140),
    .X(_00782_));
 sg13g2_o21ai_1 _20789_ (.B1(net202),
    .Y(_03404_),
    .A1(net201),
    .A2(_09035_));
 sg13g2_a22oi_1 _20790_ (.Y(_03405_),
    .B1(_03404_),
    .B2(net200),
    .A2(_03383_),
    .A1(net230));
 sg13g2_o21ai_1 _20791_ (.B1(_03325_),
    .Y(_03406_),
    .A1(net256),
    .A2(net230));
 sg13g2_o21ai_1 _20792_ (.B1(_03406_),
    .Y(_03407_),
    .A1(net257),
    .A2(_03081_));
 sg13g2_a22oi_1 _20793_ (.Y(_03408_),
    .B1(_03407_),
    .B2(net200),
    .A2(net173),
    .A1(net213));
 sg13g2_o21ai_1 _20794_ (.B1(_03408_),
    .Y(_03409_),
    .A1(_03174_),
    .A2(_03405_));
 sg13g2_mux2_1 _20795_ (.A0(_03409_),
    .A1(\cpu.dec.r_rd[3] ),
    .S(net140),
    .X(_00783_));
 sg13g2_nand2_1 _20796_ (.Y(_03410_),
    .A(net202),
    .B(_03073_));
 sg13g2_nand4_1 _20797_ (.B(_09034_),
    .C(_09157_),
    .A(net345),
    .Y(_03411_),
    .D(_09199_));
 sg13g2_a21oi_1 _20798_ (.A1(net219),
    .A2(_03411_),
    .Y(_03412_),
    .B1(_03087_));
 sg13g2_nor3_1 _20799_ (.A(_03170_),
    .B(_03228_),
    .C(_03412_),
    .Y(_03413_));
 sg13g2_a21oi_1 _20800_ (.A1(_08943_),
    .A2(_03410_),
    .Y(_03414_),
    .B1(_03413_));
 sg13g2_nand2_1 _20801_ (.Y(_03415_),
    .A(net390),
    .B(_03362_));
 sg13g2_o21ai_1 _20802_ (.B1(_03175_),
    .Y(_03416_),
    .A1(_09904_),
    .A2(_03415_));
 sg13g2_and2_1 _20803_ (.A(_03414_),
    .B(_03416_),
    .X(_03417_));
 sg13g2_nor3_1 _20804_ (.A(net333),
    .B(net199),
    .C(_03417_),
    .Y(_03418_));
 sg13g2_a21oi_1 _20805_ (.A1(net217),
    .A2(net333),
    .Y(_03419_),
    .B1(_03220_));
 sg13g2_o21ai_1 _20806_ (.B1(_03288_),
    .Y(_03420_),
    .A1(_03418_),
    .A2(_03419_));
 sg13g2_o21ai_1 _20807_ (.B1(_03420_),
    .Y(_00784_),
    .A1(net759),
    .A2(net108));
 sg13g2_nand2b_1 _20808_ (.Y(_03421_),
    .B(_03413_),
    .A_N(net214));
 sg13g2_nor3_1 _20809_ (.A(_09904_),
    .B(_03413_),
    .C(_03415_),
    .Y(_03422_));
 sg13g2_a221oi_1 _20810_ (.B2(_03174_),
    .C1(_03422_),
    .B1(_03421_),
    .A1(net201),
    .Y(_03423_),
    .A2(net214));
 sg13g2_nand2_1 _20811_ (.Y(_03424_),
    .A(_03070_),
    .B(net215));
 sg13g2_a221oi_1 _20812_ (.B2(_03424_),
    .C1(net257),
    .B1(net214),
    .A1(_03070_),
    .Y(_03425_),
    .A2(_08996_));
 sg13g2_o21ai_1 _20813_ (.B1(_03425_),
    .Y(_03426_),
    .A1(net220),
    .A2(_03410_));
 sg13g2_nand2_1 _20814_ (.Y(_03427_),
    .A(_08943_),
    .B(_03276_));
 sg13g2_nand3_1 _20815_ (.B(_03426_),
    .C(_03427_),
    .A(_03109_),
    .Y(_03428_));
 sg13g2_o21ai_1 _20816_ (.B1(net142),
    .Y(_03429_),
    .A1(_03423_),
    .A2(_03428_));
 sg13g2_o21ai_1 _20817_ (.B1(_03429_),
    .Y(_00785_),
    .A1(net880),
    .A2(net108));
 sg13g2_nand2_1 _20818_ (.Y(_03430_),
    .A(net217),
    .B(_03184_));
 sg13g2_a21oi_1 _20819_ (.A1(_03417_),
    .A2(_03430_),
    .Y(_03431_),
    .B1(_03148_));
 sg13g2_a221oi_1 _20820_ (.B2(net199),
    .C1(_03431_),
    .B1(net198),
    .A1(net194),
    .Y(_03432_),
    .A2(_09928_));
 sg13g2_nand2_1 _20821_ (.Y(_03433_),
    .A(_10558_),
    .B(net138));
 sg13g2_o21ai_1 _20822_ (.B1(_03433_),
    .Y(_00786_),
    .A1(net143),
    .A2(_03432_));
 sg13g2_nand2_1 _20823_ (.Y(_03434_),
    .A(net347),
    .B(net219));
 sg13g2_a21oi_1 _20824_ (.A1(net230),
    .A2(_03415_),
    .Y(_03435_),
    .B1(_03434_));
 sg13g2_a21oi_1 _20825_ (.A1(_09111_),
    .A2(_03090_),
    .Y(_03436_),
    .B1(_03435_));
 sg13g2_a21oi_1 _20826_ (.A1(_03075_),
    .A2(_03290_),
    .Y(_03437_),
    .B1(net213));
 sg13g2_o21ai_1 _20827_ (.B1(_03437_),
    .Y(_03438_),
    .A1(net334),
    .A2(_03436_));
 sg13g2_and4_1 _20828_ (.A(_08458_),
    .B(_08894_),
    .C(_03414_),
    .D(_03438_),
    .X(_03439_));
 sg13g2_a21oi_1 _20829_ (.A1(_10421_),
    .A2(net102),
    .Y(_00787_),
    .B1(_03439_));
 sg13g2_nor2_1 _20830_ (.A(net342),
    .B(net333),
    .Y(_03440_));
 sg13g2_a21oi_1 _20831_ (.A1(_09908_),
    .A2(_03440_),
    .Y(_03441_),
    .B1(net271));
 sg13g2_nand2b_1 _20832_ (.Y(_03442_),
    .B(_09909_),
    .A_N(_09114_));
 sg13g2_o21ai_1 _20833_ (.B1(_03075_),
    .Y(_03443_),
    .A1(net220),
    .A2(_03289_));
 sg13g2_a22oi_1 _20834_ (.Y(_03444_),
    .B1(_03225_),
    .B2(_03334_),
    .A2(_03074_),
    .A1(_09912_));
 sg13g2_nor2_1 _20835_ (.A(_03266_),
    .B(_03444_),
    .Y(_03445_));
 sg13g2_a21oi_1 _20836_ (.A1(_09912_),
    .A2(_03443_),
    .Y(_03446_),
    .B1(_03445_));
 sg13g2_o21ai_1 _20837_ (.B1(_03446_),
    .Y(_03447_),
    .A1(_03441_),
    .A2(_03442_));
 sg13g2_nand2_1 _20838_ (.Y(_03448_),
    .A(net101),
    .B(_03447_));
 sg13g2_o21ai_1 _20839_ (.B1(_03448_),
    .Y(_00788_),
    .A1(_10337_),
    .A2(net101));
 sg13g2_inv_1 _20840_ (.Y(_03449_),
    .A(_03289_));
 sg13g2_a21oi_1 _20841_ (.A1(_09907_),
    .A2(_09908_),
    .Y(_03450_),
    .B1(_09904_));
 sg13g2_o21ai_1 _20842_ (.B1(_09175_),
    .Y(_03451_),
    .A1(_03449_),
    .A2(_03450_));
 sg13g2_nor2_1 _20843_ (.A(_09191_),
    .B(_03131_),
    .Y(_03452_));
 sg13g2_nand3_1 _20844_ (.B(_03452_),
    .C(_03450_),
    .A(_09908_),
    .Y(_03453_));
 sg13g2_nand2_1 _20845_ (.Y(_03454_),
    .A(_03451_),
    .B(_03453_));
 sg13g2_nand3_1 _20846_ (.B(_03102_),
    .C(net214),
    .A(net220),
    .Y(_03455_));
 sg13g2_o21ai_1 _20847_ (.B1(_03455_),
    .Y(_03456_),
    .A1(net220),
    .A2(_03454_));
 sg13g2_o21ai_1 _20848_ (.B1(net218),
    .Y(_03457_),
    .A1(net213),
    .A2(_03102_));
 sg13g2_a22oi_1 _20849_ (.Y(_03458_),
    .B1(_03457_),
    .B2(_09911_),
    .A2(_03456_),
    .A1(net218));
 sg13g2_nand2_1 _20850_ (.Y(_03459_),
    .A(net101),
    .B(_03458_));
 sg13g2_o21ai_1 _20851_ (.B1(_03459_),
    .Y(_00789_),
    .A1(_10334_),
    .A2(net101));
 sg13g2_nand4_1 _20852_ (.B(net230),
    .C(_09199_),
    .A(_09015_),
    .Y(_03460_),
    .D(_03148_));
 sg13g2_a21oi_1 _20853_ (.A1(net173),
    .A2(_03460_),
    .Y(_03461_),
    .B1(_03449_));
 sg13g2_o21ai_1 _20854_ (.B1(_03076_),
    .Y(_03462_),
    .A1(net204),
    .A2(_03461_));
 sg13g2_a22oi_1 _20855_ (.Y(_03463_),
    .B1(_03213_),
    .B2(_03334_),
    .A2(net186),
    .A1(net273));
 sg13g2_nor2_1 _20856_ (.A(net213),
    .B(_03463_),
    .Y(_03464_));
 sg13g2_a21oi_1 _20857_ (.A1(net273),
    .A2(_03462_),
    .Y(_03465_),
    .B1(_03464_));
 sg13g2_nand2_1 _20858_ (.Y(_03466_),
    .A(_10318_),
    .B(net138));
 sg13g2_o21ai_1 _20859_ (.B1(_03466_),
    .Y(_00790_),
    .A1(net143),
    .A2(_03465_));
 sg13g2_o21ai_1 _20860_ (.B1(_08997_),
    .Y(_03467_),
    .A1(_09198_),
    .A2(_09909_));
 sg13g2_nor2_1 _20861_ (.A(_03170_),
    .B(_03449_),
    .Y(_03468_));
 sg13g2_nand2_1 _20862_ (.Y(_03469_),
    .A(_08996_),
    .B(_09124_));
 sg13g2_o21ai_1 _20863_ (.B1(_03469_),
    .Y(_03470_),
    .A1(_09127_),
    .A2(_03074_));
 sg13g2_a22oi_1 _20864_ (.Y(_03471_),
    .B1(_03470_),
    .B2(_09931_),
    .A2(_03468_),
    .A1(_03467_));
 sg13g2_nand2_1 _20865_ (.Y(_03472_),
    .A(net101),
    .B(_03471_));
 sg13g2_o21ai_1 _20866_ (.B1(_03472_),
    .Y(_00791_),
    .A1(_10955_),
    .A2(net101));
 sg13g2_mux2_1 _20867_ (.A0(_09193_),
    .A1(_10274_),
    .S(_09132_),
    .X(_00792_));
 sg13g2_nand3_1 _20868_ (.B(_09198_),
    .C(_09939_),
    .A(net142),
    .Y(_03473_));
 sg13g2_o21ai_1 _20869_ (.B1(_03473_),
    .Y(_00793_),
    .A1(net1031),
    .A2(net101));
 sg13g2_nor4_1 _20870_ (.A(_08998_),
    .B(net343),
    .C(_09089_),
    .D(_09116_),
    .Y(_03474_));
 sg13g2_mux2_1 _20871_ (.A0(_03474_),
    .A1(\cpu.dec.r_set_cc ),
    .S(_09132_),
    .X(_00794_));
 sg13g2_a22oi_1 _20872_ (.Y(_03475_),
    .B1(_03364_),
    .B2(_03080_),
    .A2(net198),
    .A1(net194));
 sg13g2_buf_1 _20873_ (.A(\cpu.dec.r_store ),
    .X(_03476_));
 sg13g2_nand2_1 _20874_ (.Y(_03477_),
    .A(_03476_),
    .B(net141));
 sg13g2_o21ai_1 _20875_ (.B1(_03477_),
    .Y(_00795_),
    .A1(net143),
    .A2(_03475_));
 sg13g2_mux2_1 _20876_ (.A0(_03390_),
    .A1(\cpu.dec.r_swapsp ),
    .S(net140),
    .X(_00796_));
 sg13g2_nor3_1 _20877_ (.A(_09893_),
    .B(_03219_),
    .C(_03164_),
    .Y(_03478_));
 sg13g2_inv_1 _20878_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_nor4_1 _20879_ (.A(net174),
    .B(_09913_),
    .C(_03389_),
    .D(_03479_),
    .Y(_03480_));
 sg13g2_a21o_1 _20880_ (.A2(net131),
    .A1(\cpu.dec.r_sys_call ),
    .B1(_03480_),
    .X(_00797_));
 sg13g2_nand2b_1 _20881_ (.Y(_03481_),
    .B(net389),
    .A_N(_03164_));
 sg13g2_a22oi_1 _20882_ (.Y(_03482_),
    .B1(_03481_),
    .B2(_08997_),
    .A2(_03478_),
    .A1(_03382_));
 sg13g2_buf_1 _20883_ (.A(_08484_),
    .X(_03483_));
 sg13g2_nor2_1 _20884_ (.A(_03131_),
    .B(net333),
    .Y(_03484_));
 sg13g2_xnor2_1 _20885_ (.Y(_03485_),
    .A(_03213_),
    .B(_03484_));
 sg13g2_nor2_1 _20886_ (.A(_03483_),
    .B(_03485_),
    .Y(_03486_));
 sg13g2_nor2_1 _20887_ (.A(_09034_),
    .B(_03200_),
    .Y(_03487_));
 sg13g2_nor2_1 _20888_ (.A(net274),
    .B(_09191_),
    .Y(_03488_));
 sg13g2_a21oi_1 _20889_ (.A1(_09071_),
    .A2(_09109_),
    .Y(_03489_),
    .B1(_03488_));
 sg13g2_nand2_1 _20890_ (.Y(_03490_),
    .A(_09892_),
    .B(_03489_));
 sg13g2_nand3_1 _20891_ (.B(_09071_),
    .C(_09089_),
    .A(_09034_),
    .Y(_03491_));
 sg13g2_nand2_1 _20892_ (.Y(_03492_),
    .A(_03490_),
    .B(_03491_));
 sg13g2_a22oi_1 _20893_ (.Y(_03493_),
    .B1(_03492_),
    .B2(net173),
    .A2(_03487_),
    .A1(_03486_));
 sg13g2_a21oi_1 _20894_ (.A1(_08996_),
    .A2(_03415_),
    .Y(_03494_),
    .B1(_03077_));
 sg13g2_o21ai_1 _20895_ (.B1(_03289_),
    .Y(_03495_),
    .A1(_09127_),
    .A2(_03494_));
 sg13g2_nand2_1 _20896_ (.Y(_03496_),
    .A(_03192_),
    .B(_03489_));
 sg13g2_o21ai_1 _20897_ (.B1(_03496_),
    .Y(_03497_),
    .A1(_03079_),
    .A2(_03078_));
 sg13g2_nor2_1 _20898_ (.A(_03483_),
    .B(net390),
    .Y(_03498_));
 sg13g2_a21oi_1 _20899_ (.A1(_08308_),
    .A2(net390),
    .Y(_03499_),
    .B1(_03498_));
 sg13g2_xnor2_1 _20900_ (.Y(_03500_),
    .A(net272),
    .B(_09192_));
 sg13g2_nor3_1 _20901_ (.A(_03469_),
    .B(_03499_),
    .C(_03500_),
    .Y(_03501_));
 sg13g2_a221oi_1 _20902_ (.B2(net201),
    .C1(_03501_),
    .B1(_03497_),
    .A1(_03486_),
    .Y(_03502_),
    .A2(_03495_));
 sg13g2_nor3_1 _20903_ (.A(_09895_),
    .B(net272),
    .C(_09937_),
    .Y(_03503_));
 sg13g2_o21ai_1 _20904_ (.B1(_09137_),
    .Y(_03504_),
    .A1(net389),
    .A2(_09158_));
 sg13g2_o21ai_1 _20905_ (.B1(_03478_),
    .Y(_03505_),
    .A1(_03503_),
    .A2(_03504_));
 sg13g2_nand2_1 _20906_ (.Y(_03506_),
    .A(_03486_),
    .B(_03487_));
 sg13g2_or3_1 _20907_ (.A(_09893_),
    .B(_03357_),
    .C(_03362_),
    .X(_03507_));
 sg13g2_nand3_1 _20908_ (.B(_03259_),
    .C(_03507_),
    .A(net219),
    .Y(_03508_));
 sg13g2_o21ai_1 _20909_ (.B1(_03087_),
    .Y(_03509_),
    .A1(net734),
    .A2(_10721_));
 sg13g2_nand3_1 _20910_ (.B(_03093_),
    .C(_03509_),
    .A(net216),
    .Y(_03510_));
 sg13g2_nor4_1 _20911_ (.A(_09035_),
    .B(net390),
    .C(_09109_),
    .D(_09199_),
    .Y(_03511_));
 sg13g2_o21ai_1 _20912_ (.B1(_03450_),
    .Y(_03512_),
    .A1(_09892_),
    .A2(_03511_));
 sg13g2_nand4_1 _20913_ (.B(_03508_),
    .C(_03510_),
    .A(_03506_),
    .Y(_03513_),
    .D(_03512_));
 sg13g2_o21ai_1 _20914_ (.B1(_03513_),
    .Y(_03514_),
    .A1(_03357_),
    .A2(_03505_));
 sg13g2_mux4_1 _20915_ (.S0(_03266_),
    .A0(_03482_),
    .A1(_03493_),
    .A2(_03502_),
    .A3(_03514_),
    .S1(_03076_),
    .X(_03515_));
 sg13g2_nand2_1 _20916_ (.Y(_03516_),
    .A(_09241_),
    .B(net141));
 sg13g2_o21ai_1 _20917_ (.B1(_03516_),
    .Y(_00798_),
    .A1(net143),
    .A2(_03515_));
 sg13g2_buf_1 _20918_ (.A(net1151),
    .X(_03517_));
 sg13g2_buf_1 _20919_ (.A(_03517_),
    .X(_03518_));
 sg13g2_nand2b_1 _20920_ (.Y(_03519_),
    .B(net1131),
    .A_N(net1046));
 sg13g2_buf_1 _20921_ (.A(_03519_),
    .X(_03520_));
 sg13g2_nand3_1 _20922_ (.B(_10261_),
    .C(net1132),
    .A(net1130),
    .Y(_03521_));
 sg13g2_buf_1 _20923_ (.A(_03521_),
    .X(_03522_));
 sg13g2_nor2_1 _20924_ (.A(_03520_),
    .B(_03522_),
    .Y(_03523_));
 sg13g2_buf_2 _20925_ (.A(_03523_),
    .X(_03524_));
 sg13g2_buf_1 _20926_ (.A(_03524_),
    .X(_03525_));
 sg13g2_mux2_1 _20927_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net849),
    .S(net521),
    .X(_00803_));
 sg13g2_mux2_1 _20928_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net851),
    .S(net521),
    .X(_00804_));
 sg13g2_mux2_1 _20929_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net852),
    .S(net521),
    .X(_00805_));
 sg13g2_buf_1 _20930_ (.A(net664),
    .X(_03526_));
 sg13g2_mux2_1 _20931_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net591),
    .S(net521),
    .X(_00806_));
 sg13g2_buf_1 _20932_ (.A(_09710_),
    .X(_03527_));
 sg13g2_mux2_1 _20933_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net656),
    .S(net521),
    .X(_00807_));
 sg13g2_buf_8 _20934_ (.A(net598),
    .X(_03528_));
 sg13g2_buf_1 _20935_ (.A(net520),
    .X(_03529_));
 sg13g2_mux2_1 _20936_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net462),
    .S(_03525_),
    .X(_00808_));
 sg13g2_buf_1 _20937_ (.A(_09558_),
    .X(_03530_));
 sg13g2_mux2_1 _20938_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net733),
    .S(_03525_),
    .X(_00809_));
 sg13g2_buf_1 _20939_ (.A(net543),
    .X(_03531_));
 sg13g2_mux2_1 _20940_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net461),
    .S(net521),
    .X(_00810_));
 sg13g2_buf_1 _20941_ (.A(_09237_),
    .X(_03532_));
 sg13g2_buf_1 _20942_ (.A(net590),
    .X(_03533_));
 sg13g2_mux2_1 _20943_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net519),
    .S(net521),
    .X(_00811_));
 sg13g2_buf_1 _20944_ (.A(net624),
    .X(_03534_));
 sg13g2_mux2_1 _20945_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net518),
    .S(net521),
    .X(_00812_));
 sg13g2_buf_2 _20946_ (.A(net596),
    .X(_03535_));
 sg13g2_buf_1 _20947_ (.A(net517),
    .X(_03536_));
 sg13g2_mux2_1 _20948_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net460),
    .S(_03524_),
    .X(_00813_));
 sg13g2_mux2_1 _20949_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net526),
    .S(_03524_),
    .X(_00814_));
 sg13g2_mux2_1 _20950_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net740),
    .S(_03524_),
    .X(_00815_));
 sg13g2_mux2_1 _20951_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net737),
    .S(_03524_),
    .X(_00816_));
 sg13g2_mux2_1 _20952_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net736),
    .S(_03524_),
    .X(_00817_));
 sg13g2_mux2_1 _20953_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net853),
    .S(_03524_),
    .X(_00818_));
 sg13g2_nor2_1 _20954_ (.A(_10258_),
    .B(_03522_),
    .Y(_03537_));
 sg13g2_buf_2 _20955_ (.A(_03537_),
    .X(_03538_));
 sg13g2_buf_1 _20956_ (.A(_03538_),
    .X(_03539_));
 sg13g2_mux2_1 _20957_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net849),
    .S(net516),
    .X(_00819_));
 sg13g2_mux2_1 _20958_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net851),
    .S(net516),
    .X(_00820_));
 sg13g2_mux2_1 _20959_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net852),
    .S(net516),
    .X(_00821_));
 sg13g2_mux2_1 _20960_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net591),
    .S(net516),
    .X(_00822_));
 sg13g2_mux2_1 _20961_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net656),
    .S(net516),
    .X(_00823_));
 sg13g2_mux2_1 _20962_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net462),
    .S(_03539_),
    .X(_00824_));
 sg13g2_mux2_1 _20963_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net733),
    .S(_03539_),
    .X(_00825_));
 sg13g2_mux2_1 _20964_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net461),
    .S(net516),
    .X(_00826_));
 sg13g2_mux2_1 _20965_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net519),
    .S(net516),
    .X(_00827_));
 sg13g2_mux2_1 _20966_ (.A0(\cpu.ex.r_11[3] ),
    .A1(net518),
    .S(net516),
    .X(_00828_));
 sg13g2_mux2_1 _20967_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net460),
    .S(_03538_),
    .X(_00829_));
 sg13g2_mux2_1 _20968_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net526),
    .S(_03538_),
    .X(_00830_));
 sg13g2_mux2_1 _20969_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net740),
    .S(_03538_),
    .X(_00831_));
 sg13g2_mux2_1 _20970_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net737),
    .S(_03538_),
    .X(_00832_));
 sg13g2_mux2_1 _20971_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net736),
    .S(_03538_),
    .X(_00833_));
 sg13g2_mux2_1 _20972_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net853),
    .S(_03538_),
    .X(_00834_));
 sg13g2_nand3_1 _20973_ (.B(_10260_),
    .C(net1132),
    .A(net1130),
    .Y(_03540_));
 sg13g2_buf_1 _20974_ (.A(_03540_),
    .X(_03541_));
 sg13g2_nor3_1 _20975_ (.A(net1131),
    .B(net1046),
    .C(_03541_),
    .Y(_03542_));
 sg13g2_buf_2 _20976_ (.A(_03542_),
    .X(_03543_));
 sg13g2_buf_1 _20977_ (.A(_03543_),
    .X(_03544_));
 sg13g2_mux2_1 _20978_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net849),
    .S(net589),
    .X(_00835_));
 sg13g2_mux2_1 _20979_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net851),
    .S(net589),
    .X(_00836_));
 sg13g2_nand2_1 _20980_ (.Y(_03545_),
    .A(net991),
    .B(_03543_));
 sg13g2_o21ai_1 _20981_ (.B1(_03545_),
    .Y(_00837_),
    .A1(_11471_),
    .A2(net589));
 sg13g2_mux2_1 _20982_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net591),
    .S(net589),
    .X(_00838_));
 sg13g2_mux2_1 _20983_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net656),
    .S(net589),
    .X(_00839_));
 sg13g2_mux2_1 _20984_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net462),
    .S(_03544_),
    .X(_00840_));
 sg13g2_mux2_1 _20985_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net733),
    .S(_03544_),
    .X(_00841_));
 sg13g2_mux2_1 _20986_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net461),
    .S(net589),
    .X(_00842_));
 sg13g2_mux2_1 _20987_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net519),
    .S(net589),
    .X(_00843_));
 sg13g2_mux2_1 _20988_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net518),
    .S(net589),
    .X(_00844_));
 sg13g2_mux2_1 _20989_ (.A0(\cpu.ex.r_12[4] ),
    .A1(net460),
    .S(_03543_),
    .X(_00845_));
 sg13g2_mux2_1 _20990_ (.A0(\cpu.ex.r_12[5] ),
    .A1(_03039_),
    .S(_03543_),
    .X(_00846_));
 sg13g2_mux2_1 _20991_ (.A0(\cpu.ex.r_12[6] ),
    .A1(_03043_),
    .S(_03543_),
    .X(_00847_));
 sg13g2_mux2_1 _20992_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net737),
    .S(_03543_),
    .X(_00848_));
 sg13g2_mux2_1 _20993_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net736),
    .S(_03543_),
    .X(_00849_));
 sg13g2_mux2_1 _20994_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net853),
    .S(_03543_),
    .X(_00850_));
 sg13g2_inv_1 _20995_ (.Y(_03546_),
    .A(_10255_));
 sg13g2_nand2_1 _20996_ (.Y(_03547_),
    .A(_03546_),
    .B(_10257_));
 sg13g2_nor2_1 _20997_ (.A(_03541_),
    .B(_03547_),
    .Y(_03548_));
 sg13g2_buf_2 _20998_ (.A(_03548_),
    .X(_03549_));
 sg13g2_buf_1 _20999_ (.A(_03549_),
    .X(_03550_));
 sg13g2_mux2_1 _21000_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net849),
    .S(net588),
    .X(_00851_));
 sg13g2_mux2_1 _21001_ (.A0(\cpu.ex.r_13[10] ),
    .A1(net851),
    .S(net588),
    .X(_00852_));
 sg13g2_mux2_1 _21002_ (.A0(\cpu.ex.r_13[11] ),
    .A1(net852),
    .S(net588),
    .X(_00853_));
 sg13g2_mux2_1 _21003_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net591),
    .S(net588),
    .X(_00854_));
 sg13g2_mux2_1 _21004_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net656),
    .S(_03550_),
    .X(_00855_));
 sg13g2_mux2_1 _21005_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net462),
    .S(net588),
    .X(_00856_));
 sg13g2_mux2_1 _21006_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net733),
    .S(_03550_),
    .X(_00857_));
 sg13g2_mux2_1 _21007_ (.A0(\cpu.ex.r_13[1] ),
    .A1(_03531_),
    .S(net588),
    .X(_00858_));
 sg13g2_nand2_1 _21008_ (.Y(_03551_),
    .A(net590),
    .B(_03549_));
 sg13g2_o21ai_1 _21009_ (.B1(_03551_),
    .Y(_00859_),
    .A1(_10401_),
    .A2(net588));
 sg13g2_mux2_1 _21010_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net518),
    .S(net588),
    .X(_00860_));
 sg13g2_mux2_1 _21011_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net460),
    .S(_03549_),
    .X(_00861_));
 sg13g2_mux2_1 _21012_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_03039_),
    .S(_03549_),
    .X(_00862_));
 sg13g2_mux2_1 _21013_ (.A0(\cpu.ex.r_13[6] ),
    .A1(_03043_),
    .S(_03549_),
    .X(_00863_));
 sg13g2_mux2_1 _21014_ (.A0(\cpu.ex.r_13[7] ),
    .A1(net737),
    .S(_03549_),
    .X(_00864_));
 sg13g2_mux2_1 _21015_ (.A0(\cpu.ex.r_13[8] ),
    .A1(net736),
    .S(_03549_),
    .X(_00865_));
 sg13g2_mux2_1 _21016_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net853),
    .S(_03549_),
    .X(_00866_));
 sg13g2_nor2_1 _21017_ (.A(_03520_),
    .B(_03541_),
    .Y(_03552_));
 sg13g2_buf_2 _21018_ (.A(_03552_),
    .X(_03553_));
 sg13g2_buf_1 _21019_ (.A(_03553_),
    .X(_03554_));
 sg13g2_mux2_1 _21020_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net849),
    .S(net515),
    .X(_00867_));
 sg13g2_mux2_1 _21021_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net851),
    .S(net515),
    .X(_00868_));
 sg13g2_mux2_1 _21022_ (.A0(\cpu.ex.r_14[11] ),
    .A1(net852),
    .S(net515),
    .X(_00869_));
 sg13g2_mux2_1 _21023_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net591),
    .S(net515),
    .X(_00870_));
 sg13g2_mux2_1 _21024_ (.A0(\cpu.ex.r_14[13] ),
    .A1(_03527_),
    .S(net515),
    .X(_00871_));
 sg13g2_mux2_1 _21025_ (.A0(\cpu.ex.r_14[14] ),
    .A1(_03529_),
    .S(_03554_),
    .X(_00872_));
 sg13g2_mux2_1 _21026_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net733),
    .S(_03554_),
    .X(_00873_));
 sg13g2_mux2_1 _21027_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net461),
    .S(net515),
    .X(_00874_));
 sg13g2_mux2_1 _21028_ (.A0(\cpu.ex.r_14[2] ),
    .A1(net519),
    .S(net515),
    .X(_00875_));
 sg13g2_mux2_1 _21029_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net518),
    .S(net515),
    .X(_00876_));
 sg13g2_mux2_1 _21030_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net460),
    .S(_03553_),
    .X(_00877_));
 sg13g2_buf_1 _21031_ (.A(net592),
    .X(_03555_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_14[5] ),
    .A1(net514),
    .S(_03553_),
    .X(_00878_));
 sg13g2_buf_1 _21033_ (.A(net857),
    .X(_03556_));
 sg13g2_mux2_1 _21034_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net732),
    .S(_03553_),
    .X(_00879_));
 sg13g2_mux2_1 _21035_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net737),
    .S(_03553_),
    .X(_00880_));
 sg13g2_mux2_1 _21036_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net736),
    .S(_03553_),
    .X(_00881_));
 sg13g2_mux2_1 _21037_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net853),
    .S(_03553_),
    .X(_00882_));
 sg13g2_nor2_1 _21038_ (.A(_10258_),
    .B(_03541_),
    .Y(_03557_));
 sg13g2_buf_2 _21039_ (.A(_03557_),
    .X(_03558_));
 sg13g2_buf_1 _21040_ (.A(_03558_),
    .X(_03559_));
 sg13g2_mux2_1 _21041_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net849),
    .S(net587),
    .X(_00883_));
 sg13g2_mux2_1 _21042_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net851),
    .S(net587),
    .X(_00884_));
 sg13g2_mux2_1 _21043_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net852),
    .S(net587),
    .X(_00885_));
 sg13g2_mux2_1 _21044_ (.A0(\cpu.ex.r_15[12] ),
    .A1(_03526_),
    .S(net587),
    .X(_00886_));
 sg13g2_mux2_1 _21045_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net656),
    .S(_03559_),
    .X(_00887_));
 sg13g2_mux2_1 _21046_ (.A0(\cpu.ex.r_15[14] ),
    .A1(_03529_),
    .S(net587),
    .X(_00888_));
 sg13g2_mux2_1 _21047_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net733),
    .S(_03559_),
    .X(_00889_));
 sg13g2_mux2_1 _21048_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net461),
    .S(net587),
    .X(_00890_));
 sg13g2_mux2_1 _21049_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net519),
    .S(net587),
    .X(_00891_));
 sg13g2_mux2_1 _21050_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net518),
    .S(net587),
    .X(_00892_));
 sg13g2_mux2_1 _21051_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net460),
    .S(_03558_),
    .X(_00893_));
 sg13g2_mux2_1 _21052_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net514),
    .S(_03558_),
    .X(_00894_));
 sg13g2_mux2_1 _21053_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net732),
    .S(_03558_),
    .X(_00895_));
 sg13g2_mux2_1 _21054_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net737),
    .S(_03558_),
    .X(_00896_));
 sg13g2_mux2_1 _21055_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net736),
    .S(_03558_),
    .X(_00897_));
 sg13g2_mux2_1 _21056_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net853),
    .S(_03558_),
    .X(_00898_));
 sg13g2_nor3_1 _21057_ (.A(net1131),
    .B(net1046),
    .C(_03522_),
    .Y(_03560_));
 sg13g2_buf_2 _21058_ (.A(_03560_),
    .X(_03561_));
 sg13g2_buf_1 _21059_ (.A(_03561_),
    .X(_03562_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net849),
    .S(net513),
    .X(_00899_));
 sg13g2_mux2_1 _21061_ (.A0(\cpu.ex.r_8[10] ),
    .A1(_03069_),
    .S(net513),
    .X(_00900_));
 sg13g2_mux2_1 _21062_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net852),
    .S(net513),
    .X(_00901_));
 sg13g2_mux2_1 _21063_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net591),
    .S(net513),
    .X(_00902_));
 sg13g2_mux2_1 _21064_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net656),
    .S(net513),
    .X(_00903_));
 sg13g2_buf_1 _21065_ (.A(net598),
    .X(_03563_));
 sg13g2_mux2_1 _21066_ (.A0(\cpu.ex.r_8[14] ),
    .A1(net512),
    .S(_03562_),
    .X(_00904_));
 sg13g2_mux2_1 _21067_ (.A0(\cpu.ex.r_8[15] ),
    .A1(_03530_),
    .S(_03562_),
    .X(_00905_));
 sg13g2_mux2_1 _21068_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net461),
    .S(net513),
    .X(_00906_));
 sg13g2_mux2_1 _21069_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net519),
    .S(net513),
    .X(_00907_));
 sg13g2_mux2_1 _21070_ (.A0(\cpu.ex.r_8[3] ),
    .A1(_03534_),
    .S(net513),
    .X(_00908_));
 sg13g2_mux2_1 _21071_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net460),
    .S(_03561_),
    .X(_00909_));
 sg13g2_mux2_1 _21072_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net514),
    .S(_03561_),
    .X(_00910_));
 sg13g2_mux2_1 _21073_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net732),
    .S(_03561_),
    .X(_00911_));
 sg13g2_mux2_1 _21074_ (.A0(\cpu.ex.r_8[7] ),
    .A1(_03063_),
    .S(_03561_),
    .X(_00912_));
 sg13g2_mux2_1 _21075_ (.A0(\cpu.ex.r_8[8] ),
    .A1(_03064_),
    .S(_03561_),
    .X(_00913_));
 sg13g2_mux2_1 _21076_ (.A0(\cpu.ex.r_8[9] ),
    .A1(_03065_),
    .S(_03561_),
    .X(_00914_));
 sg13g2_nor2_1 _21077_ (.A(_03522_),
    .B(_03547_),
    .Y(_03564_));
 sg13g2_buf_2 _21078_ (.A(_03564_),
    .X(_03565_));
 sg13g2_buf_1 _21079_ (.A(_03565_),
    .X(_03566_));
 sg13g2_mux2_1 _21080_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net849),
    .S(net511),
    .X(_00915_));
 sg13g2_mux2_1 _21081_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net851),
    .S(_03566_),
    .X(_00916_));
 sg13g2_mux2_1 _21082_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net852),
    .S(net511),
    .X(_00917_));
 sg13g2_mux2_1 _21083_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net591),
    .S(net511),
    .X(_00918_));
 sg13g2_mux2_1 _21084_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net656),
    .S(net511),
    .X(_00919_));
 sg13g2_mux2_1 _21085_ (.A0(\cpu.ex.r_9[14] ),
    .A1(net512),
    .S(_03566_),
    .X(_00920_));
 sg13g2_mux2_1 _21086_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net733),
    .S(net511),
    .X(_00921_));
 sg13g2_mux2_1 _21087_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net461),
    .S(net511),
    .X(_00922_));
 sg13g2_mux2_1 _21088_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net519),
    .S(net511),
    .X(_00923_));
 sg13g2_mux2_1 _21089_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net518),
    .S(net511),
    .X(_00924_));
 sg13g2_mux2_1 _21090_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net460),
    .S(_03565_),
    .X(_00925_));
 sg13g2_mux2_1 _21091_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net514),
    .S(_03565_),
    .X(_00926_));
 sg13g2_mux2_1 _21092_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net732),
    .S(_03565_),
    .X(_00927_));
 sg13g2_mux2_1 _21093_ (.A0(\cpu.ex.r_9[7] ),
    .A1(_03063_),
    .S(_03565_),
    .X(_00928_));
 sg13g2_mux2_1 _21094_ (.A0(\cpu.ex.r_9[8] ),
    .A1(_03064_),
    .S(_03565_),
    .X(_00929_));
 sg13g2_mux2_1 _21095_ (.A0(\cpu.ex.r_9[9] ),
    .A1(_03065_),
    .S(_03565_),
    .X(_00930_));
 sg13g2_a21o_1 _21096_ (.A2(_11608_),
    .A1(_11596_),
    .B1(net917),
    .X(_03567_));
 sg13g2_buf_1 _21097_ (.A(_03567_),
    .X(_03568_));
 sg13g2_nand3b_1 _21098_ (.B(net1092),
    .C(_08406_),
    .Y(_03569_),
    .A_N(_11614_));
 sg13g2_buf_2 _21099_ (.A(_03569_),
    .X(_03570_));
 sg13g2_nand2_2 _21100_ (.Y(_03571_),
    .A(_03568_),
    .B(_03570_));
 sg13g2_or2_1 _21101_ (.X(_03572_),
    .B(_03571_),
    .A(\cpu.ex.r_cc ));
 sg13g2_buf_1 _21102_ (.A(net228),
    .X(_03573_));
 sg13g2_nor3_1 _21103_ (.A(net338),
    .B(net268),
    .C(_10768_),
    .Y(_03574_));
 sg13g2_a21oi_1 _21104_ (.A1(_10745_),
    .A2(_03573_),
    .Y(_03575_),
    .B1(_03574_));
 sg13g2_buf_1 _21105_ (.A(_03575_),
    .X(_03576_));
 sg13g2_inv_1 _21106_ (.Y(_03577_),
    .A(_00196_));
 sg13g2_nor3_1 _21107_ (.A(_10798_),
    .B(net268),
    .C(_11949_),
    .Y(_03578_));
 sg13g2_a21oi_2 _21108_ (.B1(_03578_),
    .Y(_03579_),
    .A2(net197),
    .A1(_03577_));
 sg13g2_a21oi_1 _21109_ (.A1(net339),
    .A2(net269),
    .Y(_03580_),
    .B1(_10612_));
 sg13g2_and3_1 _21110_ (.X(_03581_),
    .A(net339),
    .B(net269),
    .C(_10640_));
 sg13g2_buf_1 _21111_ (.A(_03581_),
    .X(_03582_));
 sg13g2_nor2_1 _21112_ (.A(_03580_),
    .B(_03582_),
    .Y(_03583_));
 sg13g2_buf_2 _21113_ (.A(_03583_),
    .X(_03584_));
 sg13g2_nor2_1 _21114_ (.A(net264),
    .B(_10679_),
    .Y(_03585_));
 sg13g2_nand2_1 _21115_ (.Y(_03586_),
    .A(_10392_),
    .B(_10473_));
 sg13g2_buf_2 _21116_ (.A(_03586_),
    .X(_03587_));
 sg13g2_nor2_1 _21117_ (.A(net264),
    .B(net267),
    .Y(_03588_));
 sg13g2_inv_1 _21118_ (.Y(_03589_),
    .A(_03588_));
 sg13g2_nor2_1 _21119_ (.A(net267),
    .B(_10679_),
    .Y(_03590_));
 sg13g2_inv_1 _21120_ (.Y(_03591_),
    .A(_03590_));
 sg13g2_and2_1 _21121_ (.A(_10392_),
    .B(_10473_),
    .X(_03592_));
 sg13g2_buf_1 _21122_ (.A(_03592_),
    .X(_03593_));
 sg13g2_inv_1 _21123_ (.Y(_03594_),
    .A(_10669_));
 sg13g2_nor3_1 _21124_ (.A(_08454_),
    .B(_10388_),
    .C(_03594_),
    .Y(_03595_));
 sg13g2_nor2b_1 _21125_ (.A(_10373_),
    .B_N(_10669_),
    .Y(_03596_));
 sg13g2_or3_1 _21126_ (.A(_10672_),
    .B(_10675_),
    .C(_03596_),
    .X(_03597_));
 sg13g2_nor3_1 _21127_ (.A(_03595_),
    .B(_03597_),
    .C(_11092_),
    .Y(_03598_));
 sg13g2_nand2_1 _21128_ (.Y(_03599_),
    .A(_11573_),
    .B(_10713_));
 sg13g2_nor2_1 _21129_ (.A(_11574_),
    .B(_10713_),
    .Y(_03600_));
 sg13g2_a221oi_1 _21130_ (.B2(_03599_),
    .C1(_03600_),
    .B1(_03598_),
    .A1(_11246_),
    .Y(_03601_),
    .A2(_03593_));
 sg13g2_buf_1 _21131_ (.A(_03601_),
    .X(_03602_));
 sg13g2_a221oi_1 _21132_ (.B2(_03591_),
    .C1(_03602_),
    .B1(_03589_),
    .A1(net223),
    .Y(_03603_),
    .A2(_03587_));
 sg13g2_a21oi_1 _21133_ (.A1(_10392_),
    .A2(_10473_),
    .Y(_03604_),
    .B1(net261));
 sg13g2_and2_1 _21134_ (.A(_10476_),
    .B(_10525_),
    .X(_03605_));
 sg13g2_buf_2 _21135_ (.A(_03605_),
    .X(_03606_));
 sg13g2_nand3b_1 _21136_ (.B(_03606_),
    .C(_11155_),
    .Y(_03607_),
    .A_N(_03604_));
 sg13g2_nand3b_1 _21137_ (.B(_10603_),
    .C(_03606_),
    .Y(_03608_),
    .A_N(_03604_));
 sg13g2_a21oi_1 _21138_ (.A1(_03607_),
    .A2(_03608_),
    .Y(_03609_),
    .B1(_03602_));
 sg13g2_nand2_1 _21139_ (.Y(_03610_),
    .A(_10476_),
    .B(_10525_));
 sg13g2_a21oi_1 _21140_ (.A1(_03589_),
    .A2(_03591_),
    .Y(_03611_),
    .B1(_03610_));
 sg13g2_or4_1 _21141_ (.A(_03585_),
    .B(_03603_),
    .C(_03609_),
    .D(_03611_),
    .X(_03612_));
 sg13g2_buf_1 _21142_ (.A(_03612_),
    .X(_03613_));
 sg13g2_nand2_1 _21143_ (.Y(_03614_),
    .A(net206),
    .B(_10566_));
 sg13g2_nor2_1 _21144_ (.A(net206),
    .B(_10566_),
    .Y(_03615_));
 sg13g2_a221oi_1 _21145_ (.B2(_03614_),
    .C1(_03615_),
    .B1(_03613_),
    .A1(_11255_),
    .Y(_03616_),
    .A2(_03584_));
 sg13g2_buf_2 _21146_ (.A(_03616_),
    .X(_03617_));
 sg13g2_inv_1 _21147_ (.Y(_03618_),
    .A(_00295_));
 sg13g2_o21ai_1 _21148_ (.B1(_03618_),
    .Y(_03619_),
    .A1(net338),
    .A2(net268));
 sg13g2_o21ai_1 _21149_ (.B1(_03619_),
    .Y(_03620_),
    .A1(_03573_),
    .A2(_11951_));
 sg13g2_buf_1 _21150_ (.A(_03620_),
    .X(_03621_));
 sg13g2_a21oi_2 _21151_ (.B1(_10714_),
    .Y(_03622_),
    .A2(net269),
    .A1(net339));
 sg13g2_nor3_2 _21152_ (.A(net338),
    .B(net268),
    .C(_10740_),
    .Y(_03623_));
 sg13g2_nor2_2 _21153_ (.A(_03622_),
    .B(_03623_),
    .Y(_03624_));
 sg13g2_nor2_1 _21154_ (.A(_11190_),
    .B(_03624_),
    .Y(_03625_));
 sg13g2_o21ai_1 _21155_ (.B1(_03625_),
    .Y(_03626_),
    .A1(net208),
    .A2(net165));
 sg13g2_nor2_1 _21156_ (.A(_11255_),
    .B(_03584_),
    .Y(_03627_));
 sg13g2_a21oi_1 _21157_ (.A1(net208),
    .A2(net165),
    .Y(_03628_),
    .B1(_03627_));
 sg13g2_nand2_1 _21158_ (.Y(_03629_),
    .A(_03626_),
    .B(_03628_));
 sg13g2_nor2_1 _21159_ (.A(net197),
    .B(_11951_),
    .Y(_03630_));
 sg13g2_a21oi_1 _21160_ (.A1(_03618_),
    .A2(net197),
    .Y(_03631_),
    .B1(_03630_));
 sg13g2_buf_2 _21161_ (.A(_03631_),
    .X(_03632_));
 sg13g2_or2_1 _21162_ (.X(_03633_),
    .B(_03623_),
    .A(_03622_));
 sg13g2_buf_1 _21163_ (.A(_03633_),
    .X(_03634_));
 sg13g2_nor2_1 _21164_ (.A(_11219_),
    .B(net183),
    .Y(_03635_));
 sg13g2_nor2_1 _21165_ (.A(_03632_),
    .B(_03635_),
    .Y(_03636_));
 sg13g2_a21oi_1 _21166_ (.A1(_03632_),
    .A2(_03635_),
    .Y(_03637_),
    .B1(net205));
 sg13g2_nor2_1 _21167_ (.A(_03636_),
    .B(_03637_),
    .Y(_03638_));
 sg13g2_nor3_1 _21168_ (.A(net338),
    .B(_10799_),
    .C(_10905_),
    .Y(_03639_));
 sg13g2_a21o_1 _21169_ (.A2(net228),
    .A1(_10881_),
    .B1(_03639_),
    .X(_03640_));
 sg13g2_buf_2 _21170_ (.A(_03640_),
    .X(_03641_));
 sg13g2_nand2_1 _21171_ (.Y(_03642_),
    .A(_11309_),
    .B(_03641_));
 sg13g2_buf_2 _21172_ (.A(_03642_),
    .X(_03643_));
 sg13g2_a21oi_1 _21173_ (.A1(_10881_),
    .A2(_10533_),
    .Y(_03644_),
    .B1(_03639_));
 sg13g2_buf_2 _21174_ (.A(_03644_),
    .X(_03645_));
 sg13g2_nand2_1 _21175_ (.Y(_03646_),
    .A(_11356_),
    .B(_03645_));
 sg13g2_and2_1 _21176_ (.A(_03643_),
    .B(_03646_),
    .X(_03647_));
 sg13g2_buf_1 _21177_ (.A(_03647_),
    .X(_03648_));
 sg13g2_and3_1 _21178_ (.X(_03649_),
    .A(net339),
    .B(net269),
    .C(_10835_));
 sg13g2_a21o_1 _21179_ (.A2(net228),
    .A1(_10838_),
    .B1(_03649_),
    .X(_03650_));
 sg13g2_buf_1 _21180_ (.A(_03650_),
    .X(_03651_));
 sg13g2_inv_1 _21181_ (.Y(_03652_),
    .A(_00292_));
 sg13g2_nor3_1 _21182_ (.A(net338),
    .B(net268),
    .C(_10927_),
    .Y(_03653_));
 sg13g2_a21oi_1 _21183_ (.A1(_03652_),
    .A2(_10533_),
    .Y(_03654_),
    .B1(_03653_));
 sg13g2_buf_2 _21184_ (.A(_03654_),
    .X(_03655_));
 sg13g2_nand2_2 _21185_ (.Y(_03656_),
    .A(net207),
    .B(_03655_));
 sg13g2_a21o_1 _21186_ (.A2(net228),
    .A1(_03652_),
    .B1(_03653_),
    .X(_03657_));
 sg13g2_buf_1 _21187_ (.A(_03657_),
    .X(_03658_));
 sg13g2_nand2_1 _21188_ (.Y(_03659_),
    .A(_11490_),
    .B(_03658_));
 sg13g2_nand2_1 _21189_ (.Y(_03660_),
    .A(_03656_),
    .B(_03659_));
 sg13g2_buf_2 _21190_ (.A(_03660_),
    .X(_03661_));
 sg13g2_o21ai_1 _21191_ (.B1(_03661_),
    .Y(_03662_),
    .A1(net187),
    .A2(_03651_));
 sg13g2_nor3_1 _21192_ (.A(_03638_),
    .B(_03648_),
    .C(_03662_),
    .Y(_03663_));
 sg13g2_o21ai_1 _21193_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_03617_),
    .A2(_03629_));
 sg13g2_nand2_1 _21194_ (.Y(_03665_),
    .A(_11340_),
    .B(_03651_));
 sg13g2_nand2_1 _21195_ (.Y(_03666_),
    .A(_03645_),
    .B(_03665_));
 sg13g2_o21ai_1 _21196_ (.B1(net132),
    .Y(_03667_),
    .A1(_03645_),
    .A2(_03665_));
 sg13g2_a22oi_1 _21197_ (.Y(_03668_),
    .B1(_03666_),
    .B2(_03667_),
    .A2(_03658_),
    .A1(net207));
 sg13g2_a21o_1 _21198_ (.A2(_03655_),
    .A1(_11491_),
    .B1(_03668_),
    .X(_03669_));
 sg13g2_nor3_1 _21199_ (.A(net338),
    .B(net268),
    .C(_11948_),
    .Y(_03670_));
 sg13g2_a21oi_1 _21200_ (.A1(_00291_),
    .A2(net197),
    .Y(_03671_),
    .B1(_03670_));
 sg13g2_buf_1 _21201_ (.A(_03671_),
    .X(_03672_));
 sg13g2_nand2_1 _21202_ (.Y(_03673_),
    .A(_11832_),
    .B(net164));
 sg13g2_and2_1 _21203_ (.A(_03669_),
    .B(_03673_),
    .X(_03674_));
 sg13g2_nor2_1 _21204_ (.A(_11832_),
    .B(net164),
    .Y(_03675_));
 sg13g2_a221oi_1 _21205_ (.B2(_03674_),
    .C1(_03675_),
    .B1(_03664_),
    .A1(_03579_),
    .Y(_03676_),
    .A2(net133));
 sg13g2_buf_1 _21206_ (.A(_03676_),
    .X(_03677_));
 sg13g2_inv_2 _21207_ (.Y(_03678_),
    .A(_11546_));
 sg13g2_o21ai_1 _21208_ (.B1(_10842_),
    .Y(_03679_),
    .A1(net338),
    .A2(net268));
 sg13g2_o21ai_1 _21209_ (.B1(_03679_),
    .Y(_03680_),
    .A1(net197),
    .A2(_11953_));
 sg13g2_buf_1 _21210_ (.A(_03680_),
    .X(_03681_));
 sg13g2_inv_1 _21211_ (.Y(_03682_),
    .A(net163));
 sg13g2_a21o_1 _21212_ (.A2(net197),
    .A1(_03577_),
    .B1(_03578_),
    .X(_03683_));
 sg13g2_buf_1 _21213_ (.A(_03683_),
    .X(_03684_));
 sg13g2_buf_1 _21214_ (.A(_03684_),
    .X(_03685_));
 sg13g2_nand2_1 _21215_ (.Y(_03686_),
    .A(net128),
    .B(_11887_));
 sg13g2_o21ai_1 _21216_ (.B1(_03686_),
    .Y(_03687_),
    .A1(_03678_),
    .A2(_03682_));
 sg13g2_nand2_1 _21217_ (.Y(_03688_),
    .A(_03678_),
    .B(_03682_));
 sg13g2_o21ai_1 _21218_ (.B1(_03688_),
    .Y(_03689_),
    .A1(_03677_),
    .A2(_03687_));
 sg13g2_o21ai_1 _21219_ (.B1(_03689_),
    .Y(_03690_),
    .A1(_11562_),
    .A2(net166));
 sg13g2_inv_1 _21220_ (.Y(_03691_),
    .A(_09202_));
 sg13g2_buf_1 _21221_ (.A(_03691_),
    .X(_03692_));
 sg13g2_a21oi_1 _21222_ (.A1(_11562_),
    .A2(net166),
    .Y(_03693_),
    .B1(net848));
 sg13g2_nand3_1 _21223_ (.B(_03690_),
    .C(_03693_),
    .A(_03571_),
    .Y(_03694_));
 sg13g2_nand2_2 _21224_ (.Y(_03695_),
    .A(_10367_),
    .B(net166));
 sg13g2_inv_1 _21225_ (.Y(_03696_),
    .A(_03695_));
 sg13g2_nand2_1 _21226_ (.Y(_03697_),
    .A(_03579_),
    .B(_11887_));
 sg13g2_nor2_1 _21227_ (.A(_11507_),
    .B(_03655_),
    .Y(_03698_));
 sg13g2_buf_1 _21228_ (.A(net164),
    .X(_03699_));
 sg13g2_a21oi_1 _21229_ (.A1(_03698_),
    .A2(net127),
    .Y(_03700_),
    .B1(net191));
 sg13g2_nor2_1 _21230_ (.A(_03698_),
    .B(net127),
    .Y(_03701_));
 sg13g2_nand2_1 _21231_ (.Y(_03702_),
    .A(_03684_),
    .B(_11458_));
 sg13g2_o21ai_1 _21232_ (.B1(_03702_),
    .Y(_03703_),
    .A1(_03700_),
    .A2(_03701_));
 sg13g2_nand2_1 _21233_ (.Y(_03704_),
    .A(_03697_),
    .B(_03703_));
 sg13g2_buf_1 _21234_ (.A(net165),
    .X(_03705_));
 sg13g2_buf_8 _21235_ (.A(_10713_),
    .X(_03706_));
 sg13g2_nor2_1 _21236_ (.A(_11248_),
    .B(net212),
    .Y(_03707_));
 sg13g2_o21ai_1 _21237_ (.B1(_11589_),
    .Y(_03708_),
    .A1(_03595_),
    .A2(_03597_));
 sg13g2_nor2_1 _21238_ (.A(_00299_),
    .B(net266),
    .Y(_03709_));
 sg13g2_and4_1 _21239_ (.A(net261),
    .B(net339),
    .C(net269),
    .D(_10471_),
    .X(_03710_));
 sg13g2_a221oi_1 _21240_ (.B2(net228),
    .C1(_03710_),
    .B1(_03709_),
    .A1(_11248_),
    .Y(_03711_),
    .A2(net212));
 sg13g2_o21ai_1 _21241_ (.B1(_03711_),
    .Y(_03712_),
    .A1(_03707_),
    .A2(_03708_));
 sg13g2_buf_1 _21242_ (.A(_03712_),
    .X(_03713_));
 sg13g2_nand2_1 _21243_ (.Y(_03714_),
    .A(_11161_),
    .B(_10603_));
 sg13g2_buf_2 _21244_ (.A(_03714_),
    .X(_03715_));
 sg13g2_nand3_1 _21245_ (.B(_10392_),
    .C(_10473_),
    .A(net266),
    .Y(_03716_));
 sg13g2_nand3_1 _21246_ (.B(_10476_),
    .C(_10525_),
    .A(_10980_),
    .Y(_03717_));
 sg13g2_buf_1 _21247_ (.A(_03717_),
    .X(_03718_));
 sg13g2_and3_1 _21248_ (.X(_03719_),
    .A(_03715_),
    .B(_03716_),
    .C(_03718_));
 sg13g2_buf_1 _21249_ (.A(_03719_),
    .X(_03720_));
 sg13g2_a21o_1 _21250_ (.A2(_10525_),
    .A1(_10476_),
    .B1(_10980_),
    .X(_03721_));
 sg13g2_buf_1 _21251_ (.A(_03721_),
    .X(_03722_));
 sg13g2_o21ai_1 _21252_ (.B1(_03722_),
    .Y(_03723_),
    .A1(_11161_),
    .A2(_10603_));
 sg13g2_a21oi_1 _21253_ (.A1(_10531_),
    .A2(net228),
    .Y(_03724_),
    .B1(_10564_));
 sg13g2_buf_1 _21254_ (.A(_03724_),
    .X(_03725_));
 sg13g2_o21ai_1 _21255_ (.B1(_11189_),
    .Y(_03726_),
    .A1(_03622_),
    .A2(_03623_));
 sg13g2_buf_1 _21256_ (.A(_03726_),
    .X(_03727_));
 sg13g2_o21ai_1 _21257_ (.B1(_11217_),
    .Y(_03728_),
    .A1(_03580_),
    .A2(_03582_));
 sg13g2_buf_2 _21258_ (.A(_03728_),
    .X(_03729_));
 sg13g2_nand3_1 _21259_ (.B(_03727_),
    .C(_03729_),
    .A(net182),
    .Y(_03730_));
 sg13g2_a221oi_1 _21260_ (.B2(_03715_),
    .C1(_03730_),
    .B1(_03723_),
    .A1(_03713_),
    .Y(_03731_),
    .A2(_03720_));
 sg13g2_nand2_1 _21261_ (.Y(_03732_),
    .A(_11222_),
    .B(_03584_));
 sg13g2_nor2b_1 _21262_ (.A(_03732_),
    .B_N(_03727_),
    .Y(_03733_));
 sg13g2_nand3_1 _21263_ (.B(_03727_),
    .C(_03729_),
    .A(net206),
    .Y(_03734_));
 sg13g2_a221oi_1 _21264_ (.B2(_03715_),
    .C1(_03734_),
    .B1(_03723_),
    .A1(_03713_),
    .Y(_03735_),
    .A2(_03720_));
 sg13g2_nand2_1 _21265_ (.Y(_03736_),
    .A(_11219_),
    .B(_03624_));
 sg13g2_o21ai_1 _21266_ (.B1(_03736_),
    .Y(_03737_),
    .A1(_10566_),
    .A2(_03734_));
 sg13g2_nor4_2 _21267_ (.A(_03731_),
    .B(_03733_),
    .C(_03735_),
    .Y(_03738_),
    .D(_03737_));
 sg13g2_nand2_1 _21268_ (.Y(_03739_),
    .A(net126),
    .B(_03738_));
 sg13g2_o21ai_1 _21269_ (.B1(net205),
    .Y(_03740_),
    .A1(net165),
    .A2(_03738_));
 sg13g2_buf_1 _21270_ (.A(_03740_),
    .X(_03741_));
 sg13g2_nand4_1 _21271_ (.B(net187),
    .C(_03739_),
    .A(_11356_),
    .Y(_03742_),
    .D(_03741_));
 sg13g2_buf_1 _21272_ (.A(_03651_),
    .X(_03743_));
 sg13g2_nor2_1 _21273_ (.A(net132),
    .B(net162),
    .Y(_03744_));
 sg13g2_nand3_1 _21274_ (.B(_03741_),
    .C(_03744_),
    .A(_03739_),
    .Y(_03745_));
 sg13g2_a21oi_1 _21275_ (.A1(net187),
    .A2(_03744_),
    .Y(_03746_),
    .B1(_03645_));
 sg13g2_nand2_1 _21276_ (.Y(_03747_),
    .A(_03697_),
    .B(_03702_));
 sg13g2_buf_1 _21277_ (.A(_03747_),
    .X(_03748_));
 sg13g2_nor2b_2 _21278_ (.A(_03675_),
    .B_N(_03673_),
    .Y(_03749_));
 sg13g2_nor2_1 _21279_ (.A(_03748_),
    .B(_03749_),
    .Y(_03750_));
 sg13g2_and2_1 _21280_ (.A(_03656_),
    .B(_03750_),
    .X(_03751_));
 sg13g2_nand4_1 _21281_ (.B(_03745_),
    .C(_03746_),
    .A(_03742_),
    .Y(_03752_),
    .D(_03751_));
 sg13g2_a21oi_1 _21282_ (.A1(_10838_),
    .A2(net197),
    .Y(_03753_),
    .B1(_03649_));
 sg13g2_buf_1 _21283_ (.A(_03753_),
    .X(_03754_));
 sg13g2_a22oi_1 _21284_ (.Y(_03755_),
    .B1(_03738_),
    .B2(net165),
    .A2(_03651_),
    .A1(net189));
 sg13g2_a22oi_1 _21285_ (.Y(_03756_),
    .B1(_03741_),
    .B2(_03755_),
    .A2(net161),
    .A1(net187));
 sg13g2_buf_1 _21286_ (.A(_03756_),
    .X(_03757_));
 sg13g2_nand4_1 _21287_ (.B(_03656_),
    .C(_03750_),
    .A(_11770_),
    .Y(_03758_),
    .D(_03757_));
 sg13g2_nand3_1 _21288_ (.B(_03752_),
    .C(_03758_),
    .A(_03704_),
    .Y(_03759_));
 sg13g2_buf_1 _21289_ (.A(_03759_),
    .X(_03760_));
 sg13g2_nand2_1 _21290_ (.Y(_03761_),
    .A(net168),
    .B(_03682_));
 sg13g2_nand2_2 _21291_ (.Y(_03762_),
    .A(_03678_),
    .B(net163));
 sg13g2_inv_1 _21292_ (.Y(_03763_),
    .A(_03762_));
 sg13g2_a21oi_1 _21293_ (.A1(_03760_),
    .A2(_03761_),
    .Y(_03764_),
    .B1(_03763_));
 sg13g2_a21o_1 _21294_ (.A2(net197),
    .A1(_10745_),
    .B1(_03574_),
    .X(_03765_));
 sg13g2_buf_2 _21295_ (.A(_03765_),
    .X(_03766_));
 sg13g2_buf_1 _21296_ (.A(_03766_),
    .X(_03767_));
 sg13g2_nand2_2 _21297_ (.Y(_03768_),
    .A(_11562_),
    .B(net125));
 sg13g2_and3_1 _21298_ (.X(_03769_),
    .A(net848),
    .B(_03571_),
    .C(_03768_));
 sg13g2_o21ai_1 _21299_ (.B1(_03769_),
    .Y(_03770_),
    .A1(_03696_),
    .A2(_03764_));
 sg13g2_and3_1 _21300_ (.X(_00931_),
    .A(_03572_),
    .B(_03694_),
    .C(_03770_));
 sg13g2_nor2_1 _21301_ (.A(_10259_),
    .B(_10260_),
    .Y(_03771_));
 sg13g2_nand4_1 _21302_ (.B(net1046),
    .C(net1132),
    .A(_10255_),
    .Y(_03772_),
    .D(_03771_));
 sg13g2_nand2b_1 _21303_ (.Y(_03773_),
    .B(_08309_),
    .A_N(_03772_));
 sg13g2_buf_1 _21304_ (.A(_03773_),
    .X(_03774_));
 sg13g2_buf_1 _21305_ (.A(_03774_),
    .X(_03775_));
 sg13g2_buf_1 _21306_ (.A(_03774_),
    .X(_03776_));
 sg13g2_nand2_1 _21307_ (.Y(_03777_),
    .A(\cpu.ex.r_epc[1] ),
    .B(_03776_));
 sg13g2_o21ai_1 _21308_ (.B1(_03777_),
    .Y(_00933_),
    .A1(net484),
    .A2(net586));
 sg13g2_mux2_1 _21309_ (.A0(net858),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net586),
    .X(_00934_));
 sg13g2_buf_1 _21310_ (.A(net749),
    .X(_03778_));
 sg13g2_nand2_1 _21311_ (.Y(_03779_),
    .A(\cpu.ex.r_epc[12] ),
    .B(net585));
 sg13g2_o21ai_1 _21312_ (.B1(_03779_),
    .Y(_00935_),
    .A1(_03778_),
    .A2(net586));
 sg13g2_buf_1 _21313_ (.A(net875),
    .X(_03780_));
 sg13g2_nand2_1 _21314_ (.Y(_03781_),
    .A(\cpu.ex.r_epc[13] ),
    .B(net585));
 sg13g2_o21ai_1 _21315_ (.B1(_03781_),
    .Y(_00936_),
    .A1(net731),
    .A2(net586));
 sg13g2_buf_1 _21316_ (.A(net520),
    .X(_03782_));
 sg13g2_mux2_1 _21317_ (.A0(net459),
    .A1(\cpu.ex.r_epc[14] ),
    .S(net585),
    .X(_00937_));
 sg13g2_buf_1 _21318_ (.A(net666),
    .X(_03783_));
 sg13g2_nand2_1 _21319_ (.Y(_03784_),
    .A(\cpu.ex.r_epc[15] ),
    .B(net585));
 sg13g2_o21ai_1 _21320_ (.B1(_03784_),
    .Y(_00938_),
    .A1(_03783_),
    .A2(net586));
 sg13g2_buf_1 _21321_ (.A(_09460_),
    .X(_03785_));
 sg13g2_nand2_1 _21322_ (.Y(_03786_),
    .A(\cpu.ex.r_epc[2] ),
    .B(net585));
 sg13g2_o21ai_1 _21323_ (.B1(_03786_),
    .Y(_00939_),
    .A1(net654),
    .A2(net586));
 sg13g2_nand2_1 _21324_ (.Y(_03787_),
    .A(\cpu.ex.r_epc[3] ),
    .B(_03774_));
 sg13g2_o21ai_1 _21325_ (.B1(_03787_),
    .Y(_00940_),
    .A1(net796),
    .A2(net586));
 sg13g2_buf_1 _21326_ (.A(net774),
    .X(_03788_));
 sg13g2_buf_1 _21327_ (.A(net653),
    .X(_03789_));
 sg13g2_nand2_1 _21328_ (.Y(_03790_),
    .A(\cpu.ex.r_epc[4] ),
    .B(_03774_));
 sg13g2_o21ai_1 _21329_ (.B1(_03790_),
    .Y(_00941_),
    .A1(_03789_),
    .A2(_03775_));
 sg13g2_nand2_1 _21330_ (.Y(_03791_),
    .A(\cpu.ex.r_epc[5] ),
    .B(_03774_));
 sg13g2_o21ai_1 _21331_ (.B1(_03791_),
    .Y(_00942_),
    .A1(net657),
    .A2(net586));
 sg13g2_nand2_1 _21332_ (.Y(_03792_),
    .A(\cpu.ex.r_epc[6] ),
    .B(_03774_));
 sg13g2_o21ai_1 _21333_ (.B1(_03792_),
    .Y(_00943_),
    .A1(_03026_),
    .A2(_03775_));
 sg13g2_mux2_1 _21334_ (.A0(_03029_),
    .A1(\cpu.ex.r_epc[7] ),
    .S(net585),
    .X(_00944_));
 sg13g2_mux2_1 _21335_ (.A0(_03031_),
    .A1(\cpu.ex.r_epc[8] ),
    .S(_03776_),
    .X(_00945_));
 sg13g2_mux2_1 _21336_ (.A0(_03033_),
    .A1(\cpu.ex.r_epc[9] ),
    .S(net585),
    .X(_00946_));
 sg13g2_mux2_1 _21337_ (.A0(net859),
    .A1(\cpu.ex.r_epc[10] ),
    .S(net585),
    .X(_00947_));
 sg13g2_nand4_1 _21338_ (.B(_10257_),
    .C(net1132),
    .A(_03546_),
    .Y(_03793_),
    .D(_03771_));
 sg13g2_buf_1 _21339_ (.A(_03793_),
    .X(_03794_));
 sg13g2_buf_1 _21340_ (.A(_03794_),
    .X(_03795_));
 sg13g2_buf_1 _21341_ (.A(_03794_),
    .X(_03796_));
 sg13g2_nand2_1 _21342_ (.Y(_03797_),
    .A(\cpu.ex.r_lr[1] ),
    .B(_03796_));
 sg13g2_o21ai_1 _21343_ (.B1(_03797_),
    .Y(_00953_),
    .A1(_10204_),
    .A2(net652));
 sg13g2_mux2_1 _21344_ (.A0(net858),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net652),
    .X(_00954_));
 sg13g2_nand2_1 _21345_ (.Y(_03798_),
    .A(\cpu.ex.r_lr[12] ),
    .B(net651));
 sg13g2_o21ai_1 _21346_ (.B1(_03798_),
    .Y(_00955_),
    .A1(_03778_),
    .A2(net652));
 sg13g2_nand2_1 _21347_ (.Y(_03799_),
    .A(\cpu.ex.r_lr[13] ),
    .B(net651));
 sg13g2_o21ai_1 _21348_ (.B1(_03799_),
    .Y(_00956_),
    .A1(net731),
    .A2(net652));
 sg13g2_mux2_1 _21349_ (.A0(net459),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net651),
    .X(_00957_));
 sg13g2_nand2_1 _21350_ (.Y(_03800_),
    .A(\cpu.ex.r_lr[15] ),
    .B(net651));
 sg13g2_o21ai_1 _21351_ (.B1(_03800_),
    .Y(_00958_),
    .A1(_03783_),
    .A2(net652));
 sg13g2_nand2_1 _21352_ (.Y(_03801_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net651));
 sg13g2_o21ai_1 _21353_ (.B1(_03801_),
    .Y(_00959_),
    .A1(net654),
    .A2(net652));
 sg13g2_nand2_1 _21354_ (.Y(_03802_),
    .A(\cpu.ex.r_lr[3] ),
    .B(_03794_));
 sg13g2_o21ai_1 _21355_ (.B1(_03802_),
    .Y(_00960_),
    .A1(net796),
    .A2(net652));
 sg13g2_nand2_1 _21356_ (.Y(_03803_),
    .A(\cpu.ex.r_lr[4] ),
    .B(_03794_));
 sg13g2_o21ai_1 _21357_ (.B1(_03803_),
    .Y(_00961_),
    .A1(_03789_),
    .A2(net652));
 sg13g2_nand2_1 _21358_ (.Y(_03804_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03794_));
 sg13g2_o21ai_1 _21359_ (.B1(_03804_),
    .Y(_00962_),
    .A1(net657),
    .A2(_03795_));
 sg13g2_nand2_1 _21360_ (.Y(_03805_),
    .A(\cpu.ex.r_lr[6] ),
    .B(_03794_));
 sg13g2_o21ai_1 _21361_ (.B1(_03805_),
    .Y(_00963_),
    .A1(net743),
    .A2(_03795_));
 sg13g2_mux2_1 _21362_ (.A0(_03029_),
    .A1(\cpu.ex.r_lr[7] ),
    .S(net651),
    .X(_00964_));
 sg13g2_mux2_1 _21363_ (.A0(_03031_),
    .A1(\cpu.ex.r_lr[8] ),
    .S(_03796_),
    .X(_00965_));
 sg13g2_mux2_1 _21364_ (.A0(_03033_),
    .A1(\cpu.ex.r_lr[9] ),
    .S(net651),
    .X(_00966_));
 sg13g2_mux2_1 _21365_ (.A0(_03035_),
    .A1(\cpu.ex.r_lr[10] ),
    .S(net651),
    .X(_00967_));
 sg13g2_and2_1 _21366_ (.A(_11549_),
    .B(_11565_),
    .X(_03806_));
 sg13g2_buf_2 _21367_ (.A(_03806_),
    .X(_03807_));
 sg13g2_nor2_1 _21368_ (.A(net226),
    .B(_03807_),
    .Y(_03808_));
 sg13g2_xnor2_1 _21369_ (.Y(_03809_),
    .A(net78),
    .B(_03808_));
 sg13g2_buf_1 _21370_ (.A(_10265_),
    .X(_03810_));
 sg13g2_buf_1 _21371_ (.A(net510),
    .X(_03811_));
 sg13g2_a22oi_1 _21372_ (.Y(_03812_),
    .B1(_03678_),
    .B2(_11905_),
    .A2(_11562_),
    .A1(_11930_));
 sg13g2_a21oi_1 _21373_ (.A1(_11913_),
    .A2(_10367_),
    .Y(_03813_),
    .B1(_03812_));
 sg13g2_nand2b_1 _21374_ (.Y(_03814_),
    .B(_03813_),
    .A_N(_11899_));
 sg13g2_nand3_1 _21375_ (.B(_11901_),
    .C(_03814_),
    .A(_11893_),
    .Y(_03815_));
 sg13g2_buf_2 _21376_ (.A(_03815_),
    .X(_03816_));
 sg13g2_o21ai_1 _21377_ (.B1(_11905_),
    .Y(_03817_),
    .A1(_11930_),
    .A2(_11912_));
 sg13g2_a21o_1 _21378_ (.A2(_11546_),
    .A1(_10367_),
    .B1(_11913_),
    .X(_03818_));
 sg13g2_a221oi_1 _21379_ (.B2(_11903_),
    .C1(_03818_),
    .B1(_11902_),
    .A1(_10610_),
    .Y(_03819_),
    .A2(_10744_));
 sg13g2_a22oi_1 _21380_ (.Y(_03820_),
    .B1(_03819_),
    .B2(net597),
    .A2(_11904_),
    .A1(_11562_));
 sg13g2_o21ai_1 _21381_ (.B1(_03820_),
    .Y(_03821_),
    .A1(net610),
    .A2(_03817_));
 sg13g2_and2_1 _21382_ (.A(_03816_),
    .B(_03821_),
    .X(_03822_));
 sg13g2_nand2_1 _21383_ (.Y(_03823_),
    .A(_11929_),
    .B(net536));
 sg13g2_xnor2_1 _21384_ (.Y(_03824_),
    .A(_03822_),
    .B(_03823_));
 sg13g2_nand3_1 _21385_ (.B(_10266_),
    .C(\cpu.ex.r_cc ),
    .A(net1132),
    .Y(_03825_));
 sg13g2_nand3_1 _21386_ (.B(_10267_),
    .C(_10252_),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_03826_));
 sg13g2_a21oi_1 _21387_ (.A1(_03825_),
    .A2(_03826_),
    .Y(_03827_),
    .B1(net510));
 sg13g2_a221oi_1 _21388_ (.B2(_03824_),
    .C1(_03827_),
    .B1(_11718_),
    .A1(net990),
    .Y(_03828_),
    .A2(net458));
 sg13g2_o21ai_1 _21389_ (.B1(_03828_),
    .Y(_00968_),
    .A1(_11882_),
    .A2(_03809_));
 sg13g2_inv_1 _21390_ (.Y(_03829_),
    .A(\cpu.ex.r_mult[17] ));
 sg13g2_and2_1 _21391_ (.A(net483),
    .B(_10252_),
    .X(_03830_));
 sg13g2_buf_1 _21392_ (.A(_03830_),
    .X(_03831_));
 sg13g2_buf_1 _21393_ (.A(_03831_),
    .X(_03832_));
 sg13g2_inv_1 _21394_ (.Y(_03833_),
    .A(_11058_));
 sg13g2_a21o_1 _21395_ (.A2(_03822_),
    .A1(_11929_),
    .B1(_03833_),
    .X(_03834_));
 sg13g2_and4_1 _21396_ (.A(_03833_),
    .B(_11929_),
    .C(net536),
    .D(_03821_),
    .X(_03835_));
 sg13g2_buf_8 _21397_ (.A(_03835_),
    .X(_03836_));
 sg13g2_a21oi_1 _21398_ (.A1(_03816_),
    .A2(_03836_),
    .Y(_03837_),
    .B1(_11731_));
 sg13g2_buf_8 _21399_ (.A(_11549_),
    .X(_03838_));
 sg13g2_buf_8 _21400_ (.A(_11565_),
    .X(_03839_));
 sg13g2_o21ai_1 _21401_ (.B1(net260),
    .Y(_03840_),
    .A1(net78),
    .A2(net226));
 sg13g2_nor2_1 _21402_ (.A(_11587_),
    .B(net226),
    .Y(_03841_));
 sg13g2_nand2_1 _21403_ (.Y(_03842_),
    .A(net336),
    .B(_03841_));
 sg13g2_nor2_1 _21404_ (.A(_11058_),
    .B(_09380_),
    .Y(_03843_));
 sg13g2_or2_1 _21405_ (.X(_03844_),
    .B(_03843_),
    .A(net86));
 sg13g2_a221oi_1 _21406_ (.B2(_03842_),
    .C1(_03844_),
    .B1(_03840_),
    .A1(net28),
    .Y(_03845_),
    .A2(net27));
 sg13g2_a21o_1 _21407_ (.A2(_03837_),
    .A1(_03834_),
    .B1(_03845_),
    .X(_03846_));
 sg13g2_nand2_1 _21408_ (.Y(_03847_),
    .A(_11549_),
    .B(_11565_));
 sg13g2_nand2_1 _21409_ (.Y(_03848_),
    .A(_03840_),
    .B(_03842_));
 sg13g2_nand2_1 _21410_ (.Y(_03849_),
    .A(net63),
    .B(_03843_));
 sg13g2_a21oi_1 _21411_ (.A1(_03847_),
    .A2(_03848_),
    .Y(_03850_),
    .B1(_03849_));
 sg13g2_o21ai_1 _21412_ (.B1(net483),
    .Y(_03851_),
    .A1(_03846_),
    .A2(_03850_));
 sg13g2_nand2_2 _21413_ (.Y(_03852_),
    .A(_10267_),
    .B(_10252_));
 sg13g2_nand4_1 _21414_ (.B(_10253_),
    .C(_10266_),
    .A(_09202_),
    .Y(_03853_),
    .D(\cpu.ex.r_cc ));
 sg13g2_a21oi_1 _21415_ (.A1(_03852_),
    .A2(_03853_),
    .Y(_03854_),
    .B1(_10265_));
 sg13g2_buf_8 _21416_ (.A(_03854_),
    .X(_03855_));
 sg13g2_buf_1 _21417_ (.A(_03855_),
    .X(_03856_));
 sg13g2_a21oi_1 _21418_ (.A1(_03531_),
    .A2(net458),
    .Y(_03857_),
    .B1(net331));
 sg13g2_a22oi_1 _21419_ (.Y(_00969_),
    .B1(_03851_),
    .B2(_03857_),
    .A2(net332),
    .A1(_03829_));
 sg13g2_inv_1 _21420_ (.Y(_03858_),
    .A(\cpu.ex.r_mult[18] ));
 sg13g2_nand2_1 _21421_ (.Y(_03859_),
    .A(net260),
    .B(_03841_));
 sg13g2_o21ai_1 _21422_ (.B1(net336),
    .Y(_03860_),
    .A1(_11587_),
    .A2(net226));
 sg13g2_nand2b_1 _21423_ (.Y(_03861_),
    .B(_03860_),
    .A_N(_03843_));
 sg13g2_nand2_1 _21424_ (.Y(_03862_),
    .A(_03859_),
    .B(_03861_));
 sg13g2_xnor2_1 _21425_ (.Y(_03863_),
    .A(net221),
    .B(_03862_));
 sg13g2_a21oi_1 _21426_ (.A1(net28),
    .A2(net27),
    .Y(_03864_),
    .B1(_03863_));
 sg13g2_nand2_2 _21427_ (.Y(_03865_),
    .A(_03816_),
    .B(_03836_));
 sg13g2_o21ai_1 _21428_ (.B1(_11234_),
    .Y(_03866_),
    .A1(_11731_),
    .A2(_03865_));
 sg13g2_a21o_1 _21429_ (.A2(_03864_),
    .A1(net63),
    .B1(_03866_),
    .X(_03867_));
 sg13g2_nand2_1 _21430_ (.Y(_03868_),
    .A(net537),
    .B(net63));
 sg13g2_nor2_1 _21431_ (.A(_11234_),
    .B(_03837_),
    .Y(_03869_));
 sg13g2_o21ai_1 _21432_ (.B1(_03869_),
    .Y(_03870_),
    .A1(_03864_),
    .A2(_03868_));
 sg13g2_nand3_1 _21433_ (.B(_03867_),
    .C(_03870_),
    .A(net483),
    .Y(_03871_));
 sg13g2_a21oi_1 _21434_ (.A1(net590),
    .A2(net458),
    .Y(_03872_),
    .B1(net331));
 sg13g2_a22oi_1 _21435_ (.Y(_00970_),
    .B1(_03871_),
    .B2(_03872_),
    .A2(net332),
    .A1(_03858_));
 sg13g2_inv_1 _21436_ (.Y(_03873_),
    .A(\cpu.ex.r_mult[19] ));
 sg13g2_nor2_1 _21437_ (.A(_11061_),
    .B(_11234_),
    .Y(_03874_));
 sg13g2_nor2b_1 _21438_ (.A(_03865_),
    .B_N(_03874_),
    .Y(_03875_));
 sg13g2_o21ai_1 _21439_ (.B1(_11061_),
    .Y(_03876_),
    .A1(_11234_),
    .A2(_03865_));
 sg13g2_nor2b_1 _21440_ (.A(_03875_),
    .B_N(_03876_),
    .Y(_03877_));
 sg13g2_a221oi_1 _21441_ (.B2(_03877_),
    .C1(net331),
    .B1(_11733_),
    .A1(net624),
    .Y(_03878_),
    .A2(net510));
 sg13g2_a221oi_1 _21442_ (.B2(_03841_),
    .C1(_11058_),
    .B1(net260),
    .A1(_11234_),
    .Y(_03879_),
    .A2(net221));
 sg13g2_a21oi_1 _21443_ (.A1(net221),
    .A2(_03860_),
    .Y(_03880_),
    .B1(_11234_));
 sg13g2_o21ai_1 _21444_ (.B1(net537),
    .Y(_03881_),
    .A1(_03879_),
    .A2(_03880_));
 sg13g2_o21ai_1 _21445_ (.B1(_03881_),
    .Y(_03882_),
    .A1(net221),
    .A2(_03860_));
 sg13g2_xnor2_1 _21446_ (.Y(_03883_),
    .A(net227),
    .B(_03882_));
 sg13g2_nor2_1 _21447_ (.A(_11061_),
    .B(_09380_),
    .Y(_03884_));
 sg13g2_o21ai_1 _21448_ (.B1(_03884_),
    .Y(_03885_),
    .A1(_03807_),
    .A2(_03883_));
 sg13g2_or3_1 _21449_ (.A(_03807_),
    .B(_03883_),
    .C(_03884_),
    .X(_03886_));
 sg13g2_a21o_1 _21450_ (.A2(_03886_),
    .A1(_03885_),
    .B1(_11882_),
    .X(_03887_));
 sg13g2_a22oi_1 _21451_ (.Y(_00971_),
    .B1(_03878_),
    .B2(_03887_),
    .A2(net332),
    .A1(_03873_));
 sg13g2_inv_1 _21452_ (.Y(_03888_),
    .A(\cpu.ex.r_mult[20] ));
 sg13g2_nor2_1 _21453_ (.A(_11158_),
    .B(_09380_),
    .Y(_03889_));
 sg13g2_nand2_1 _21454_ (.Y(_03890_),
    .A(net65),
    .B(_11094_));
 sg13g2_a21oi_1 _21455_ (.A1(_03890_),
    .A2(_11252_),
    .Y(_03891_),
    .B1(_11276_));
 sg13g2_xnor2_1 _21456_ (.Y(_03892_),
    .A(net265),
    .B(_03891_));
 sg13g2_a21oi_1 _21457_ (.A1(net28),
    .A2(net27),
    .Y(_03893_),
    .B1(_03892_));
 sg13g2_xor2_1 _21458_ (.B(_03893_),
    .A(_03889_),
    .X(_03894_));
 sg13g2_nand2_1 _21459_ (.Y(_03895_),
    .A(net64),
    .B(_03894_));
 sg13g2_nand2_1 _21460_ (.Y(_03896_),
    .A(_11159_),
    .B(net536));
 sg13g2_xnor2_1 _21461_ (.Y(_03897_),
    .A(_03875_),
    .B(_03896_));
 sg13g2_a221oi_1 _21462_ (.B2(_03897_),
    .C1(net331),
    .B1(_11718_),
    .A1(net517),
    .Y(_03898_),
    .A2(net458));
 sg13g2_a22oi_1 _21463_ (.Y(_00972_),
    .B1(_03895_),
    .B2(_03898_),
    .A2(net332),
    .A1(_03888_));
 sg13g2_inv_1 _21464_ (.Y(_03899_),
    .A(\cpu.ex.r_mult[21] ));
 sg13g2_buf_8 _21465_ (.A(_11157_),
    .X(_03900_));
 sg13g2_inv_1 _21466_ (.Y(_03901_),
    .A(_03900_));
 sg13g2_nand4_1 _21467_ (.B(_03816_),
    .C(_03836_),
    .A(_11159_),
    .Y(_03902_),
    .D(_03874_));
 sg13g2_buf_2 _21468_ (.A(_03902_),
    .X(_03903_));
 sg13g2_xnor2_1 _21469_ (.Y(_03904_),
    .A(_03901_),
    .B(_03903_));
 sg13g2_a22oi_1 _21470_ (.Y(_03905_),
    .B1(_11733_),
    .B2(_03904_),
    .A2(net458),
    .A1(net592));
 sg13g2_nand3_1 _21471_ (.B(_11057_),
    .C(_03843_),
    .A(_11055_),
    .Y(_03906_));
 sg13g2_a21o_1 _21472_ (.A2(_11057_),
    .A1(_11055_),
    .B1(_03833_),
    .X(_03907_));
 sg13g2_a21oi_1 _21473_ (.A1(_03906_),
    .A2(_03907_),
    .Y(_03908_),
    .B1(_11235_));
 sg13g2_nor2_1 _21474_ (.A(_11225_),
    .B(net260),
    .Y(_03909_));
 sg13g2_o21ai_1 _21475_ (.B1(net223),
    .Y(_03910_),
    .A1(_03908_),
    .A2(_03909_));
 sg13g2_xnor2_1 _21476_ (.Y(_03911_),
    .A(_03833_),
    .B(net260));
 sg13g2_nand4_1 _21477_ (.B(_11225_),
    .C(net261),
    .A(_11235_),
    .Y(_03912_),
    .D(_03911_));
 sg13g2_o21ai_1 _21478_ (.B1(_09380_),
    .Y(_03913_),
    .A1(_11237_),
    .A2(_11240_));
 sg13g2_nand4_1 _21479_ (.B(_10934_),
    .C(_10978_),
    .A(_11158_),
    .Y(_03914_),
    .D(_03884_));
 sg13g2_nor2_1 _21480_ (.A(_11159_),
    .B(_11062_),
    .Y(_03915_));
 sg13g2_o21ai_1 _21481_ (.B1(_03915_),
    .Y(_03916_),
    .A1(_11237_),
    .A2(_11240_));
 sg13g2_nand3_1 _21482_ (.B(_03914_),
    .C(_03916_),
    .A(_03913_),
    .Y(_03917_));
 sg13g2_xnor2_1 _21483_ (.Y(_03918_),
    .A(_11062_),
    .B(_11241_));
 sg13g2_and2_1 _21484_ (.A(net265),
    .B(_03889_),
    .X(_03919_));
 sg13g2_a22oi_1 _21485_ (.Y(_03920_),
    .B1(_03918_),
    .B2(_03919_),
    .A2(_03917_),
    .A1(net264));
 sg13g2_a21o_1 _21486_ (.A2(_03912_),
    .A1(_03910_),
    .B1(_03920_),
    .X(_03921_));
 sg13g2_a221oi_1 _21487_ (.B2(_11903_),
    .C1(_03921_),
    .B1(_11902_),
    .A1(_10610_),
    .Y(_03922_),
    .A2(_10744_));
 sg13g2_buf_2 _21488_ (.A(_03922_),
    .X(_03923_));
 sg13g2_a221oi_1 _21489_ (.B2(_11059_),
    .C1(_11235_),
    .B1(net266),
    .A1(_11062_),
    .Y(_03924_),
    .A2(net267));
 sg13g2_a221oi_1 _21490_ (.B2(_03833_),
    .C1(net266),
    .B1(net336),
    .A1(_11062_),
    .Y(_03925_),
    .A2(net267));
 sg13g2_nor4_1 _21491_ (.A(_11162_),
    .B(_11275_),
    .C(_03924_),
    .D(_03925_),
    .Y(_03926_));
 sg13g2_o21ai_1 _21492_ (.B1(net599),
    .Y(_03927_),
    .A1(_11262_),
    .A2(_03926_));
 sg13g2_o21ai_1 _21493_ (.B1(_03927_),
    .Y(_03928_),
    .A1(_11589_),
    .A2(_03921_));
 sg13g2_buf_2 _21494_ (.A(_03928_),
    .X(_03929_));
 sg13g2_nor2_1 _21495_ (.A(_03923_),
    .B(_03929_),
    .Y(_03930_));
 sg13g2_xnor2_1 _21496_ (.Y(_03931_),
    .A(net225),
    .B(_03930_));
 sg13g2_a21oi_1 _21497_ (.A1(net28),
    .A2(net27),
    .Y(_03932_),
    .B1(_03931_));
 sg13g2_xor2_1 _21498_ (.B(_03932_),
    .A(_11264_),
    .X(_03933_));
 sg13g2_a21oi_1 _21499_ (.A1(net64),
    .A2(_03933_),
    .Y(_03934_),
    .B1(net331));
 sg13g2_a22oi_1 _21500_ (.Y(_00973_),
    .B1(_03905_),
    .B2(_03934_),
    .A2(net332),
    .A1(_03899_));
 sg13g2_nor2_1 _21501_ (.A(net989),
    .B(_03903_),
    .Y(_03935_));
 sg13g2_xnor2_1 _21502_ (.Y(_03936_),
    .A(net1127),
    .B(_03935_));
 sg13g2_a221oi_1 _21503_ (.B2(_03936_),
    .C1(net331),
    .B1(_11733_),
    .A1(_09225_),
    .Y(_03937_),
    .A2(_03810_));
 sg13g2_nand2_1 _21504_ (.Y(_03938_),
    .A(_11156_),
    .B(_11163_));
 sg13g2_and2_1 _21505_ (.A(_11263_),
    .B(_11265_),
    .X(_03939_));
 sg13g2_o21ai_1 _21506_ (.B1(_03939_),
    .Y(_03940_),
    .A1(_03938_),
    .A2(_03891_));
 sg13g2_xnor2_1 _21507_ (.Y(_03941_),
    .A(net337),
    .B(_03940_));
 sg13g2_a21oi_1 _21508_ (.A1(net28),
    .A2(net27),
    .Y(_03942_),
    .B1(_03941_));
 sg13g2_xor2_1 _21509_ (.B(_03942_),
    .A(_11268_),
    .X(_03943_));
 sg13g2_nand2_1 _21510_ (.Y(_03944_),
    .A(net64),
    .B(_03943_));
 sg13g2_a22oi_1 _21511_ (.Y(_00974_),
    .B1(_03937_),
    .B2(_03944_),
    .A2(net332),
    .A1(_11164_));
 sg13g2_inv_1 _21512_ (.Y(_03945_),
    .A(\cpu.ex.r_mult[23] ));
 sg13g2_a21oi_1 _21513_ (.A1(_09229_),
    .A2(_10265_),
    .Y(_03946_),
    .B1(_03855_));
 sg13g2_nand2_1 _21514_ (.Y(_03947_),
    .A(net222),
    .B(net225));
 sg13g2_nor3_1 _21515_ (.A(_03947_),
    .B(_03923_),
    .C(_03929_),
    .Y(_03948_));
 sg13g2_nor4_1 _21516_ (.A(_03901_),
    .B(net337),
    .C(_03923_),
    .D(_03929_),
    .Y(_03949_));
 sg13g2_inv_1 _21517_ (.Y(_03950_),
    .A(_11218_));
 sg13g2_nor4_1 _21518_ (.A(_03950_),
    .B(net206),
    .C(_03923_),
    .D(_03929_),
    .Y(_03951_));
 sg13g2_o21ai_1 _21519_ (.B1(_11218_),
    .Y(_03952_),
    .A1(net989),
    .A2(net222));
 sg13g2_o21ai_1 _21520_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_03901_),
    .A2(_03947_));
 sg13g2_nor4_1 _21521_ (.A(_03948_),
    .B(_03949_),
    .C(_03951_),
    .D(_03953_),
    .Y(_03954_));
 sg13g2_o21ai_1 _21522_ (.B1(net206),
    .Y(_03955_),
    .A1(_03923_),
    .A2(_03929_));
 sg13g2_nor2_1 _21523_ (.A(net222),
    .B(_03955_),
    .Y(_03956_));
 sg13g2_a21oi_1 _21524_ (.A1(_11516_),
    .A2(_03954_),
    .Y(_03957_),
    .B1(_03956_));
 sg13g2_xnor2_1 _21525_ (.Y(_03958_),
    .A(net224),
    .B(_03957_));
 sg13g2_a21oi_1 _21526_ (.A1(_11549_),
    .A2(_11565_),
    .Y(_03959_),
    .B1(_03958_));
 sg13g2_xnor2_1 _21527_ (.Y(_03960_),
    .A(_11258_),
    .B(_03959_));
 sg13g2_nor3_1 _21528_ (.A(net1127),
    .B(net989),
    .C(_03903_),
    .Y(_03961_));
 sg13g2_xnor2_1 _21529_ (.Y(_03962_),
    .A(_11164_),
    .B(_03961_));
 sg13g2_a22oi_1 _21530_ (.Y(_03963_),
    .B1(_03962_),
    .B2(_11634_),
    .A2(_03960_),
    .A1(net63));
 sg13g2_and2_1 _21531_ (.A(net425),
    .B(_03946_),
    .X(_03964_));
 sg13g2_a221oi_1 _21532_ (.B2(_03963_),
    .C1(_03964_),
    .B1(_03946_),
    .A1(_03945_),
    .Y(_00975_),
    .A2(_03831_));
 sg13g2_inv_1 _21533_ (.Y(_03965_),
    .A(\cpu.ex.r_mult[24] ));
 sg13g2_xnor2_1 _21534_ (.Y(_03966_),
    .A(net205),
    .B(_11551_));
 sg13g2_a21oi_1 _21535_ (.A1(net28),
    .A2(net27),
    .Y(_03967_),
    .B1(_03966_));
 sg13g2_xor2_1 _21536_ (.B(_03967_),
    .A(_11385_),
    .X(_03968_));
 sg13g2_a221oi_1 _21537_ (.B2(_03968_),
    .C1(_03856_),
    .B1(net64),
    .A1(net1070),
    .Y(_03969_),
    .A2(net510));
 sg13g2_nor4_1 _21538_ (.A(_11164_),
    .B(net1127),
    .C(net989),
    .D(_03903_),
    .Y(_03970_));
 sg13g2_xnor2_1 _21539_ (.Y(_03971_),
    .A(_11384_),
    .B(_03970_));
 sg13g2_nand2_1 _21540_ (.Y(_03972_),
    .A(_11733_),
    .B(_03971_));
 sg13g2_a22oi_1 _21541_ (.Y(_00976_),
    .B1(_03969_),
    .B2(_03972_),
    .A2(net332),
    .A1(_03965_));
 sg13g2_or2_1 _21542_ (.X(_03973_),
    .B(_03855_),
    .A(_10267_));
 sg13g2_nor2b_1 _21543_ (.A(net510),
    .B_N(_03973_),
    .Y(_03974_));
 sg13g2_o21ai_1 _21544_ (.B1(_03974_),
    .Y(_03975_),
    .A1(\cpu.ex.r_mult[25] ),
    .A2(_03852_));
 sg13g2_nor2_1 _21545_ (.A(_11312_),
    .B(_11731_),
    .Y(_03976_));
 sg13g2_nor2_1 _21546_ (.A(_11498_),
    .B(_11731_),
    .Y(_03977_));
 sg13g2_nand2_1 _21547_ (.Y(_03978_),
    .A(_10620_),
    .B(_11495_));
 sg13g2_nor4_1 _21548_ (.A(net1127),
    .B(net989),
    .C(_03903_),
    .D(_03978_),
    .Y(_03979_));
 sg13g2_mux2_1 _21549_ (.A0(_03976_),
    .A1(_03977_),
    .S(_03979_),
    .X(_03980_));
 sg13g2_nor3_1 _21550_ (.A(net206),
    .B(_03923_),
    .C(_03929_),
    .Y(_03981_));
 sg13g2_nand2_1 _21551_ (.Y(_03982_),
    .A(_03950_),
    .B(net337));
 sg13g2_o21ai_1 _21552_ (.B1(_03982_),
    .Y(_03983_),
    .A1(_03900_),
    .A2(_03981_));
 sg13g2_nand3_1 _21553_ (.B(_11257_),
    .C(net263),
    .A(_10620_),
    .Y(_03984_));
 sg13g2_nand3b_1 _21554_ (.B(_03984_),
    .C(_11227_),
    .Y(_03985_),
    .A_N(_11386_));
 sg13g2_nor2_1 _21555_ (.A(net609),
    .B(_03985_),
    .Y(_03986_));
 sg13g2_nor3_1 _21556_ (.A(_11495_),
    .B(_11377_),
    .C(_11380_),
    .Y(_03987_));
 sg13g2_nand3b_1 _21557_ (.B(net263),
    .C(_10620_),
    .Y(_03988_),
    .A_N(_03987_));
 sg13g2_a21o_1 _21558_ (.A2(_03988_),
    .A1(_11496_),
    .B1(_10248_),
    .X(_03989_));
 sg13g2_buf_1 _21559_ (.A(_03989_),
    .X(_03990_));
 sg13g2_o21ai_1 _21560_ (.B1(_03990_),
    .Y(_03991_),
    .A1(_03955_),
    .A2(_03985_));
 sg13g2_a21oi_1 _21561_ (.A1(_03983_),
    .A2(_03986_),
    .Y(_03992_),
    .B1(_03991_));
 sg13g2_xnor2_1 _21562_ (.Y(_03993_),
    .A(net187),
    .B(_03992_));
 sg13g2_and4_1 _21563_ (.A(_11312_),
    .B(_03847_),
    .C(net63),
    .D(_03993_),
    .X(_03994_));
 sg13g2_nand3_1 _21564_ (.B(net537),
    .C(net63),
    .A(_11498_),
    .Y(_03995_));
 sg13g2_a21oi_1 _21565_ (.A1(_03847_),
    .A2(_03993_),
    .Y(_03996_),
    .B1(_03995_));
 sg13g2_nor4_1 _21566_ (.A(_03855_),
    .B(_03980_),
    .C(_03994_),
    .D(_03996_),
    .Y(_03997_));
 sg13g2_nand2_1 _21567_ (.Y(_03998_),
    .A(net993),
    .B(net458));
 sg13g2_o21ai_1 _21568_ (.B1(_03998_),
    .Y(_00977_),
    .A1(_03975_),
    .A2(_03997_));
 sg13g2_nor3_1 _21569_ (.A(_11312_),
    .B(net1127),
    .C(_03978_),
    .Y(_03999_));
 sg13g2_nand3b_1 _21570_ (.B(_03999_),
    .C(_03901_),
    .Y(_04000_),
    .A_N(_03903_));
 sg13g2_xnor2_1 _21571_ (.Y(_04001_),
    .A(_11350_),
    .B(_04000_));
 sg13g2_a21oi_1 _21572_ (.A1(net205),
    .A2(_11551_),
    .Y(_04002_),
    .B1(_11384_));
 sg13g2_o21ai_1 _21573_ (.B1(net189),
    .Y(_04003_),
    .A1(net205),
    .A2(_11551_));
 sg13g2_o21ai_1 _21574_ (.B1(_11348_),
    .Y(_04004_),
    .A1(_04002_),
    .A2(_04003_));
 sg13g2_nand2b_1 _21575_ (.Y(_04005_),
    .B(net187),
    .A_N(_03992_));
 sg13g2_a21oi_1 _21576_ (.A1(_04004_),
    .A2(_04005_),
    .Y(_04006_),
    .B1(net169));
 sg13g2_and3_1 _21577_ (.X(_04007_),
    .A(net169),
    .B(_04004_),
    .C(_04005_));
 sg13g2_o21ai_1 _21578_ (.B1(_03847_),
    .Y(_04008_),
    .A1(_04006_),
    .A2(_04007_));
 sg13g2_and2_1 _21579_ (.A(_11311_),
    .B(net64),
    .X(_04009_));
 sg13g2_a21o_1 _21580_ (.A2(_03810_),
    .A1(_10903_),
    .B1(_03855_),
    .X(_04010_));
 sg13g2_a221oi_1 _21581_ (.B2(_04009_),
    .C1(_04010_),
    .B1(_04008_),
    .A1(_11733_),
    .Y(_04011_),
    .A2(_04001_));
 sg13g2_or3_1 _21582_ (.A(_11311_),
    .B(_11882_),
    .C(_04008_),
    .X(_04012_));
 sg13g2_a22oi_1 _21583_ (.Y(_00978_),
    .B1(_04011_),
    .B2(_04012_),
    .A2(net332),
    .A1(_10888_));
 sg13g2_inv_1 _21584_ (.Y(_04013_),
    .A(\cpu.ex.r_mult[27] ));
 sg13g2_nor2_1 _21585_ (.A(_11310_),
    .B(net989),
    .Y(_04014_));
 sg13g2_nand4_1 _21586_ (.B(_03874_),
    .C(_03999_),
    .A(_11159_),
    .Y(_04015_),
    .D(_04014_));
 sg13g2_nor2_1 _21587_ (.A(_03865_),
    .B(_04015_),
    .Y(_04016_));
 sg13g2_xnor2_1 _21588_ (.Y(_04017_),
    .A(_10888_),
    .B(_04016_));
 sg13g2_a221oi_1 _21589_ (.B2(_04017_),
    .C1(net331),
    .B1(_11733_),
    .A1(_10925_),
    .Y(_04018_),
    .A2(net510));
 sg13g2_nand2_1 _21590_ (.Y(_04019_),
    .A(net224),
    .B(_11258_));
 sg13g2_and3_1 _21591_ (.X(_04020_),
    .A(_11387_),
    .B(_03984_),
    .C(_04019_));
 sg13g2_and2_1 _21592_ (.A(_11516_),
    .B(_04020_),
    .X(_04021_));
 sg13g2_o21ai_1 _21593_ (.B1(net132),
    .Y(_04022_),
    .A1(net189),
    .A2(_03990_));
 sg13g2_a221oi_1 _21594_ (.B2(_03990_),
    .C1(_11312_),
    .B1(net189),
    .A1(_11310_),
    .Y(_04023_),
    .A2(_11309_));
 sg13g2_a21oi_1 _21595_ (.A1(_11350_),
    .A2(_04022_),
    .Y(_04024_),
    .B1(_04023_));
 sg13g2_or2_1 _21596_ (.X(_04025_),
    .B(_04024_),
    .A(_10248_));
 sg13g2_o21ai_1 _21597_ (.B1(_04025_),
    .Y(_04026_),
    .A1(_11571_),
    .A2(_03990_));
 sg13g2_a221oi_1 _21598_ (.B2(_03954_),
    .C1(_04026_),
    .B1(_04021_),
    .A1(_03956_),
    .Y(_04027_),
    .A2(_04020_));
 sg13g2_buf_1 _21599_ (.A(_04027_),
    .X(_04028_));
 sg13g2_xnor2_1 _21600_ (.Y(_04029_),
    .A(net190),
    .B(_04028_));
 sg13g2_a21oi_1 _21601_ (.A1(_03838_),
    .A2(_03839_),
    .Y(_04030_),
    .B1(_04029_));
 sg13g2_xnor2_1 _21602_ (.Y(_04031_),
    .A(_11492_),
    .B(_04030_));
 sg13g2_nand2_1 _21603_ (.Y(_04032_),
    .A(net64),
    .B(_04031_));
 sg13g2_a22oi_1 _21604_ (.Y(_00979_),
    .B1(_04018_),
    .B2(_04032_),
    .A2(_03832_),
    .A1(_04013_));
 sg13g2_nand2_1 _21605_ (.Y(_04033_),
    .A(net664),
    .B(net458));
 sg13g2_o21ai_1 _21606_ (.B1(_03974_),
    .Y(_04034_),
    .A1(_10852_),
    .A2(_03852_));
 sg13g2_and2_1 _21607_ (.A(net207),
    .B(_11492_),
    .X(_04035_));
 sg13g2_nor2_1 _21608_ (.A(_10888_),
    .B(net207),
    .Y(_04036_));
 sg13g2_nand2_1 _21609_ (.Y(_04037_),
    .A(_11505_),
    .B(_11509_));
 sg13g2_a21o_1 _21610_ (.A2(_04036_),
    .A1(_11389_),
    .B1(_04037_),
    .X(_04038_));
 sg13g2_a22oi_1 _21611_ (.Y(_04039_),
    .B1(_04038_),
    .B2(net537),
    .A2(_04035_),
    .A1(_11389_));
 sg13g2_xnor2_1 _21612_ (.Y(_04040_),
    .A(net191),
    .B(_04039_));
 sg13g2_o21ai_1 _21613_ (.B1(_11513_),
    .Y(_04041_),
    .A1(_03807_),
    .A2(_04040_));
 sg13g2_or3_1 _21614_ (.A(_11513_),
    .B(_03807_),
    .C(_04040_),
    .X(_04042_));
 sg13g2_a21o_1 _21615_ (.A2(_04042_),
    .A1(_04041_),
    .B1(net86),
    .X(_04043_));
 sg13g2_nor4_1 _21616_ (.A(_10888_),
    .B(_11630_),
    .C(_03865_),
    .D(_04015_),
    .Y(_04044_));
 sg13g2_xnor2_1 _21617_ (.Y(_04045_),
    .A(_11419_),
    .B(_04044_));
 sg13g2_a221oi_1 _21618_ (.B2(_04045_),
    .C1(net331),
    .B1(_11634_),
    .A1(net664),
    .Y(_04046_),
    .A2(net458));
 sg13g2_a22oi_1 _21619_ (.Y(_00980_),
    .B1(_04043_),
    .B2(_04046_),
    .A2(_04034_),
    .A1(_04033_));
 sg13g2_inv_1 _21620_ (.Y(_04047_),
    .A(_10789_));
 sg13g2_nor3_1 _21621_ (.A(_10888_),
    .B(_11419_),
    .C(_11310_),
    .Y(_04048_));
 sg13g2_nand3_1 _21622_ (.B(_03999_),
    .C(_04048_),
    .A(net536),
    .Y(_04049_));
 sg13g2_nor3_1 _21623_ (.A(net989),
    .B(_03903_),
    .C(_04049_),
    .Y(_04050_));
 sg13g2_xnor2_1 _21624_ (.Y(_04051_),
    .A(_11461_),
    .B(_04050_));
 sg13g2_a21oi_1 _21625_ (.A1(net28),
    .A2(net27),
    .Y(_04052_),
    .B1(_11887_));
 sg13g2_a21oi_1 _21626_ (.A1(net28),
    .A2(net27),
    .Y(_04053_),
    .B1(net133));
 sg13g2_nand2_1 _21627_ (.Y(_04054_),
    .A(_11419_),
    .B(net191));
 sg13g2_nand3_1 _21628_ (.B(net537),
    .C(_04054_),
    .A(_10887_),
    .Y(_04055_));
 sg13g2_nand2_1 _21629_ (.Y(_04056_),
    .A(net207),
    .B(_11513_));
 sg13g2_a21oi_1 _21630_ (.A1(_04055_),
    .A2(_04056_),
    .Y(_04057_),
    .B1(_04028_));
 sg13g2_nor3_1 _21631_ (.A(net191),
    .B(net190),
    .C(_04028_),
    .Y(_04058_));
 sg13g2_and4_1 _21632_ (.A(_10887_),
    .B(net537),
    .C(net207),
    .D(_04054_),
    .X(_04059_));
 sg13g2_nor4_2 _21633_ (.A(_11518_),
    .B(_04057_),
    .C(_04058_),
    .Y(_04060_),
    .D(_04059_));
 sg13g2_mux2_1 _21634_ (.A0(_04052_),
    .A1(_04053_),
    .S(_04060_),
    .X(_04061_));
 sg13g2_o21ai_1 _21635_ (.B1(net483),
    .Y(_04062_),
    .A1(_11461_),
    .A2(net609));
 sg13g2_nor2_1 _21636_ (.A(net86),
    .B(_04062_),
    .Y(_04063_));
 sg13g2_a22oi_1 _21637_ (.Y(_04064_),
    .B1(_04061_),
    .B2(_04063_),
    .A2(_04051_),
    .A1(_11733_));
 sg13g2_a21o_1 _21638_ (.A2(_03839_),
    .A1(_03838_),
    .B1(_11887_),
    .X(_04065_));
 sg13g2_a21o_1 _21639_ (.A2(_11565_),
    .A1(_11549_),
    .B1(net133),
    .X(_04066_));
 sg13g2_mux2_1 _21640_ (.A0(_04065_),
    .A1(_04066_),
    .S(_04060_),
    .X(_04067_));
 sg13g2_nor4_1 _21641_ (.A(_11461_),
    .B(net609),
    .C(net425),
    .D(net86),
    .Y(_04068_));
 sg13g2_a221oi_1 _21642_ (.B2(_04068_),
    .C1(_03856_),
    .B1(_04067_),
    .A1(net776),
    .Y(_04069_),
    .A2(_03811_));
 sg13g2_a22oi_1 _21643_ (.Y(_00981_),
    .B1(_04064_),
    .B2(_04069_),
    .A2(_03832_),
    .A1(_04047_));
 sg13g2_o21ai_1 _21644_ (.B1(_03974_),
    .Y(_04070_),
    .A1(\cpu.ex.r_mult[30] ),
    .A2(_03852_));
 sg13g2_nor4_2 _21645_ (.A(_11461_),
    .B(net989),
    .C(_03903_),
    .Y(_04071_),
    .D(_04049_));
 sg13g2_xnor2_1 _21646_ (.Y(_04072_),
    .A(_04047_),
    .B(_04071_));
 sg13g2_nand2_1 _21647_ (.Y(_04073_),
    .A(_10789_),
    .B(net537));
 sg13g2_xnor2_1 _21648_ (.Y(_04074_),
    .A(_11522_),
    .B(net168));
 sg13g2_a21oi_1 _21649_ (.A1(_11549_),
    .A2(_11565_),
    .Y(_04075_),
    .B1(_04074_));
 sg13g2_xnor2_1 _21650_ (.Y(_04076_),
    .A(_04073_),
    .B(_04075_));
 sg13g2_a221oi_1 _21651_ (.B2(net63),
    .C1(_03855_),
    .B1(_04076_),
    .A1(_11634_),
    .Y(_04077_),
    .A2(_04072_));
 sg13g2_nand2_1 _21652_ (.Y(_04078_),
    .A(net520),
    .B(_03811_));
 sg13g2_o21ai_1 _21653_ (.B1(_04078_),
    .Y(_00982_),
    .A1(_04070_),
    .A2(_04077_));
 sg13g2_and2_1 _21654_ (.A(net907),
    .B(net510),
    .X(_04079_));
 sg13g2_o21ai_1 _21655_ (.B1(_03973_),
    .Y(_04080_),
    .A1(\cpu.ex.r_mult[31] ),
    .A2(_03852_));
 sg13g2_a21oi_1 _21656_ (.A1(_11522_),
    .A2(net168),
    .Y(_04081_),
    .B1(_11559_));
 sg13g2_xnor2_1 _21657_ (.Y(_04082_),
    .A(_11562_),
    .B(_04081_));
 sg13g2_nor2_1 _21658_ (.A(_11555_),
    .B(_03868_),
    .Y(_04083_));
 sg13g2_a21oi_1 _21659_ (.A1(_04082_),
    .A2(_04083_),
    .Y(_04084_),
    .B1(_03855_));
 sg13g2_nor3_1 _21660_ (.A(net510),
    .B(_04080_),
    .C(_04084_),
    .Y(_04085_));
 sg13g2_nand2_1 _21661_ (.Y(_04086_),
    .A(_10789_),
    .B(_04071_));
 sg13g2_nor4_1 _21662_ (.A(_11555_),
    .B(_10265_),
    .C(_11731_),
    .D(_04080_),
    .Y(_04087_));
 sg13g2_and2_1 _21663_ (.A(_04086_),
    .B(_04087_),
    .X(_04088_));
 sg13g2_nand2b_1 _21664_ (.Y(_04089_),
    .B(_11555_),
    .A_N(_10265_));
 sg13g2_nor4_1 _21665_ (.A(_11731_),
    .B(_04080_),
    .C(_04086_),
    .D(_04089_),
    .Y(_04090_));
 sg13g2_or4_1 _21666_ (.A(_04079_),
    .B(_04085_),
    .C(_04088_),
    .D(_04090_),
    .X(_00983_));
 sg13g2_inv_1 _21667_ (.Y(_04091_),
    .A(_00260_));
 sg13g2_nand2_1 _21668_ (.Y(_04092_),
    .A(net1152),
    .B(_04091_));
 sg13g2_mux2_1 _21669_ (.A0(_08362_),
    .A1(_04092_),
    .S(_11963_),
    .X(_04093_));
 sg13g2_and2_1 _21670_ (.A(net275),
    .B(_10674_),
    .X(_04094_));
 sg13g2_buf_1 _21671_ (.A(_04094_),
    .X(_04095_));
 sg13g2_nand3b_1 _21672_ (.B(net196),
    .C(net751),
    .Y(_04096_),
    .A_N(_04093_));
 sg13g2_buf_1 _21673_ (.A(_04096_),
    .X(_04097_));
 sg13g2_buf_1 _21674_ (.A(_04097_),
    .X(_04098_));
 sg13g2_buf_1 _21675_ (.A(net188),
    .X(_04099_));
 sg13g2_nand2_1 _21676_ (.Y(_04100_),
    .A(_10670_),
    .B(_10676_));
 sg13g2_buf_1 _21677_ (.A(_04100_),
    .X(_04101_));
 sg13g2_buf_1 _21678_ (.A(net181),
    .X(_04102_));
 sg13g2_inv_1 _21679_ (.Y(_04103_),
    .A(net159));
 sg13g2_nand2b_1 _21680_ (.Y(_04104_),
    .B(net336),
    .A_N(net212));
 sg13g2_nand2_1 _21681_ (.Y(_04105_),
    .A(net260),
    .B(net212));
 sg13g2_nand2_1 _21682_ (.Y(_04106_),
    .A(_04104_),
    .B(_04105_));
 sg13g2_nor2_1 _21683_ (.A(_09916_),
    .B(\cpu.dec.r_op[7] ),
    .Y(_04107_));
 sg13g2_nor2_1 _21684_ (.A(_08295_),
    .B(net1135),
    .Y(_04108_));
 sg13g2_buf_1 _21685_ (.A(_04108_),
    .X(_04109_));
 sg13g2_nor4_1 _21686_ (.A(net1148),
    .B(net1147),
    .C(net1134),
    .D(_09924_),
    .Y(_04110_));
 sg13g2_and2_1 _21687_ (.A(net847),
    .B(_04110_),
    .X(_04111_));
 sg13g2_buf_1 _21688_ (.A(_04111_),
    .X(_04112_));
 sg13g2_nor4_2 _21689_ (.A(_09195_),
    .B(_09202_),
    .C(_09916_),
    .Y(_04113_),
    .D(\cpu.dec.r_op[7] ));
 sg13g2_nand2_1 _21690_ (.Y(_04114_),
    .A(_04112_),
    .B(_04113_));
 sg13g2_buf_1 _21691_ (.A(_04114_),
    .X(_04115_));
 sg13g2_a22oi_1 _21692_ (.Y(_04116_),
    .B1(_04107_),
    .B2(net509),
    .A2(_04106_),
    .A1(_04103_));
 sg13g2_nand2_1 _21693_ (.Y(_04117_),
    .A(_04107_),
    .B(net509));
 sg13g2_buf_2 _21694_ (.A(_04117_),
    .X(_04118_));
 sg13g2_o21ai_1 _21695_ (.B1(_11589_),
    .Y(_04119_),
    .A1(_04103_),
    .A2(_04118_));
 sg13g2_nor2_1 _21696_ (.A(net181),
    .B(_04118_),
    .Y(_04120_));
 sg13g2_a21oi_1 _21697_ (.A1(net848),
    .A2(net159),
    .Y(_04121_),
    .B1(_04120_));
 sg13g2_nor2_1 _21698_ (.A(_04106_),
    .B(_04121_),
    .Y(_04122_));
 sg13g2_a22oi_1 _21699_ (.Y(_04123_),
    .B1(_04122_),
    .B2(_11589_),
    .A2(_04119_),
    .A1(_04106_));
 sg13g2_o21ai_1 _21700_ (.B1(_04123_),
    .Y(_04124_),
    .A1(net1073),
    .A2(_04116_));
 sg13g2_a21oi_1 _21701_ (.A1(net1076),
    .A2(net189),
    .Y(_04125_),
    .B1(net188));
 sg13g2_nor2_1 _21702_ (.A(net262),
    .B(net261),
    .Y(_04126_));
 sg13g2_buf_2 _21703_ (.A(_04126_),
    .X(_04127_));
 sg13g2_nor2_2 _21704_ (.A(_11249_),
    .B(_11092_),
    .Y(_04128_));
 sg13g2_and2_1 _21705_ (.A(_04127_),
    .B(_04128_),
    .X(_04129_));
 sg13g2_buf_1 _21706_ (.A(_04129_),
    .X(_04130_));
 sg13g2_buf_1 _21707_ (.A(net158),
    .X(_04131_));
 sg13g2_buf_1 _21708_ (.A(net124),
    .X(_04132_));
 sg13g2_nand3_1 _21709_ (.B(net159),
    .C(net100),
    .A(_09924_),
    .Y(_04133_));
 sg13g2_mux2_1 _21710_ (.A0(net1147),
    .A1(net1074),
    .S(_04105_),
    .X(_04134_));
 sg13g2_o21ai_1 _21711_ (.B1(_04104_),
    .Y(_04135_),
    .A1(net1134),
    .A2(_04134_));
 sg13g2_nand3_1 _21712_ (.B(_04133_),
    .C(_04135_),
    .A(_04125_),
    .Y(_04136_));
 sg13g2_nor4_1 _21713_ (.A(net262),
    .B(net223),
    .C(net336),
    .D(net226),
    .Y(_04137_));
 sg13g2_buf_1 _21714_ (.A(_04137_),
    .X(_04138_));
 sg13g2_buf_1 _21715_ (.A(net180),
    .X(_04139_));
 sg13g2_nor2_1 _21716_ (.A(net227),
    .B(net261),
    .Y(_04140_));
 sg13g2_nor2b_1 _21717_ (.A(_11576_),
    .B_N(_04140_),
    .Y(_04141_));
 sg13g2_buf_2 _21718_ (.A(_04141_),
    .X(_04142_));
 sg13g2_a22oi_1 _21719_ (.Y(_04143_),
    .B1(_04142_),
    .B2(net162),
    .A2(net157),
    .A1(net126));
 sg13g2_nand2_1 _21720_ (.Y(_04144_),
    .A(_11242_),
    .B(net221));
 sg13g2_nor2_1 _21721_ (.A(_11576_),
    .B(_04144_),
    .Y(_04145_));
 sg13g2_buf_2 _21722_ (.A(_04145_),
    .X(_04146_));
 sg13g2_nor4_1 _21723_ (.A(net262),
    .B(net223),
    .C(net260),
    .D(net226),
    .Y(_04147_));
 sg13g2_buf_1 _21724_ (.A(_04147_),
    .X(_04148_));
 sg13g2_buf_1 _21725_ (.A(net179),
    .X(_04149_));
 sg13g2_or2_1 _21726_ (.X(_04150_),
    .B(_03582_),
    .A(_03580_));
 sg13g2_buf_1 _21727_ (.A(_04150_),
    .X(_04151_));
 sg13g2_a22oi_1 _21728_ (.Y(_04152_),
    .B1(net156),
    .B2(net155),
    .A2(_04146_),
    .A1(net128));
 sg13g2_buf_1 _21729_ (.A(_03658_),
    .X(_04153_));
 sg13g2_nand3_1 _21730_ (.B(_11038_),
    .C(_11049_),
    .A(_11026_),
    .Y(_04154_));
 sg13g2_nor2b_1 _21731_ (.A(net1041),
    .B_N(_11051_),
    .Y(_04155_));
 sg13g2_a221oi_1 _21732_ (.B2(net541),
    .C1(_04155_),
    .B1(_11052_),
    .A1(_11149_),
    .Y(_04156_),
    .A2(_04154_));
 sg13g2_o21ai_1 _21733_ (.B1(net1031),
    .Y(_04157_),
    .A1(_10274_),
    .A2(_04156_));
 sg13g2_and3_1 _21734_ (.X(_04158_),
    .A(_11057_),
    .B(_11092_),
    .C(_04157_));
 sg13g2_buf_1 _21735_ (.A(_04158_),
    .X(_04159_));
 sg13g2_and2_1 _21736_ (.A(_04140_),
    .B(_04159_),
    .X(_04160_));
 sg13g2_buf_1 _21737_ (.A(_04160_),
    .X(_04161_));
 sg13g2_buf_1 _21738_ (.A(_04161_),
    .X(_04162_));
 sg13g2_and2_1 _21739_ (.A(_04128_),
    .B(_04140_),
    .X(_04163_));
 sg13g2_buf_1 _21740_ (.A(_04163_),
    .X(_04164_));
 sg13g2_buf_1 _21741_ (.A(_04164_),
    .X(_04165_));
 sg13g2_buf_1 _21742_ (.A(_03641_),
    .X(_04166_));
 sg13g2_a22oi_1 _21743_ (.Y(_04167_),
    .B1(net122),
    .B2(net153),
    .A2(net123),
    .A1(net154));
 sg13g2_nor2_1 _21744_ (.A(net227),
    .B(net223),
    .Y(_04168_));
 sg13g2_and2_1 _21745_ (.A(_04168_),
    .B(_04159_),
    .X(_04169_));
 sg13g2_buf_1 _21746_ (.A(_04169_),
    .X(_04170_));
 sg13g2_nor2_2 _21747_ (.A(net336),
    .B(_11092_),
    .Y(_04171_));
 sg13g2_and2_1 _21748_ (.A(_04171_),
    .B(_04140_),
    .X(_04172_));
 sg13g2_buf_2 _21749_ (.A(_04172_),
    .X(_04173_));
 sg13g2_a22oi_1 _21750_ (.Y(_04174_),
    .B1(_04173_),
    .B2(net164),
    .A2(_04170_),
    .A1(net125));
 sg13g2_nand4_1 _21751_ (.B(_04152_),
    .C(_04167_),
    .A(_04143_),
    .Y(_04175_),
    .D(_04174_));
 sg13g2_buf_1 _21752_ (.A(_10566_),
    .X(_04176_));
 sg13g2_nor3_1 _21753_ (.A(net262),
    .B(_11229_),
    .C(_11576_),
    .Y(_04177_));
 sg13g2_buf_1 _21754_ (.A(_04177_),
    .X(_04178_));
 sg13g2_nand2_1 _21755_ (.Y(_04179_),
    .A(net152),
    .B(net151));
 sg13g2_buf_1 _21756_ (.A(_03610_),
    .X(_04180_));
 sg13g2_and2_1 _21757_ (.A(_04127_),
    .B(_04159_),
    .X(_04181_));
 sg13g2_buf_1 _21758_ (.A(_04181_),
    .X(_04182_));
 sg13g2_buf_1 _21759_ (.A(_04182_),
    .X(_04183_));
 sg13g2_nand2_1 _21760_ (.Y(_04184_),
    .A(net150),
    .B(net121));
 sg13g2_and3_1 _21761_ (.X(_04185_),
    .A(net227),
    .B(net261),
    .C(_04159_));
 sg13g2_buf_1 _21762_ (.A(_04185_),
    .X(_04186_));
 sg13g2_a21oi_1 _21763_ (.A1(net183),
    .A2(net149),
    .Y(_04187_),
    .B1(net158));
 sg13g2_nand3_1 _21764_ (.B(_04184_),
    .C(_04187_),
    .A(_04179_),
    .Y(_04188_));
 sg13g2_nor2_1 _21765_ (.A(_11572_),
    .B(_11576_),
    .Y(_04189_));
 sg13g2_nand2_1 _21766_ (.Y(_04190_),
    .A(_04171_),
    .B(_04168_));
 sg13g2_inv_1 _21767_ (.Y(_04191_),
    .A(_04190_));
 sg13g2_and2_1 _21768_ (.A(_08295_),
    .B(_03766_),
    .X(_04192_));
 sg13g2_buf_1 _21769_ (.A(_04192_),
    .X(_04193_));
 sg13g2_o21ai_1 _21770_ (.B1(_04193_),
    .Y(_04194_),
    .A1(_04189_),
    .A2(_04191_));
 sg13g2_buf_1 _21771_ (.A(net163),
    .X(_04195_));
 sg13g2_and2_1 _21772_ (.A(_04128_),
    .B(_04168_),
    .X(_04196_));
 sg13g2_buf_1 _21773_ (.A(_04196_),
    .X(_04197_));
 sg13g2_and2_1 _21774_ (.A(_04127_),
    .B(_04171_),
    .X(_04198_));
 sg13g2_buf_2 _21775_ (.A(_04198_),
    .X(_04199_));
 sg13g2_buf_1 _21776_ (.A(_04199_),
    .X(_04200_));
 sg13g2_buf_1 _21777_ (.A(_10679_),
    .X(_04201_));
 sg13g2_a22oi_1 _21778_ (.Y(_04202_),
    .B1(net119),
    .B2(net211),
    .A2(_04197_),
    .A1(net120));
 sg13g2_nand2_1 _21779_ (.Y(_04203_),
    .A(_04194_),
    .B(_04202_));
 sg13g2_nor3_1 _21780_ (.A(_04175_),
    .B(_04188_),
    .C(_04203_),
    .Y(_04204_));
 sg13g2_buf_1 _21781_ (.A(_03587_),
    .X(_04205_));
 sg13g2_nand2_1 _21782_ (.Y(_04206_),
    .A(_04127_),
    .B(_04128_));
 sg13g2_buf_1 _21783_ (.A(_04206_),
    .X(_04207_));
 sg13g2_nor2_1 _21784_ (.A(net148),
    .B(net147),
    .Y(_04208_));
 sg13g2_nor3_1 _21785_ (.A(net847),
    .B(_04204_),
    .C(_04208_),
    .Y(_04209_));
 sg13g2_nor2_1 _21786_ (.A(_04136_),
    .B(_04209_),
    .Y(_04210_));
 sg13g2_a22oi_1 _21787_ (.Y(_04211_),
    .B1(_04124_),
    .B2(_04210_),
    .A2(_11633_),
    .A1(net160));
 sg13g2_inv_1 _21788_ (.Y(_04212_),
    .A(_04211_));
 sg13g2_and4_1 _21789_ (.A(net1152),
    .B(_11580_),
    .C(_11964_),
    .D(net196),
    .X(_04213_));
 sg13g2_buf_1 _21790_ (.A(_04213_),
    .X(_04214_));
 sg13g2_nand2_1 _21791_ (.Y(_04215_),
    .A(net275),
    .B(_10674_));
 sg13g2_buf_2 _21792_ (.A(_04215_),
    .X(_04216_));
 sg13g2_nor3_1 _21793_ (.A(_11943_),
    .B(_04093_),
    .C(_04216_),
    .Y(_04217_));
 sg13g2_nand2_1 _21794_ (.Y(_04218_),
    .A(_09241_),
    .B(_08456_));
 sg13g2_nor2_1 _21795_ (.A(_09376_),
    .B(_04218_),
    .Y(_04219_));
 sg13g2_a21oi_1 _21796_ (.A1(_08457_),
    .A2(_09376_),
    .Y(_04220_),
    .B1(_04219_));
 sg13g2_nand3_1 _21797_ (.B(_09284_),
    .C(net751),
    .A(net1152),
    .Y(_04221_));
 sg13g2_nor3_1 _21798_ (.A(_09241_),
    .B(_08457_),
    .C(_04221_),
    .Y(_04222_));
 sg13g2_nor2_1 _21799_ (.A(net917),
    .B(_04222_),
    .Y(_04223_));
 sg13g2_o21ai_1 _21800_ (.B1(_04223_),
    .Y(_04224_),
    .A1(net1092),
    .A2(_04220_));
 sg13g2_nor3_1 _21801_ (.A(_04217_),
    .B(net84),
    .C(_04224_),
    .Y(_04225_));
 sg13g2_buf_1 _21802_ (.A(_04225_),
    .X(_04226_));
 sg13g2_buf_1 _21803_ (.A(_04226_),
    .X(_04227_));
 sg13g2_a22oi_1 _21804_ (.Y(_04228_),
    .B1(net33),
    .B2(net696),
    .A2(net84),
    .A1(_00200_));
 sg13g2_o21ai_1 _21805_ (.B1(_04228_),
    .Y(_00984_),
    .A1(net76),
    .A2(_04212_));
 sg13g2_buf_1 _21806_ (.A(_08872_),
    .X(_04229_));
 sg13g2_nand2_1 _21807_ (.Y(_04230_),
    .A(_08898_),
    .B(net810));
 sg13g2_nor2_1 _21808_ (.A(_08839_),
    .B(_04230_),
    .Y(_04231_));
 sg13g2_nand3_1 _21809_ (.B(_08863_),
    .C(_04231_),
    .A(_08815_),
    .Y(_04232_));
 sg13g2_or2_1 _21810_ (.X(_04233_),
    .B(_04232_),
    .A(net988));
 sg13g2_buf_1 _21811_ (.A(_04233_),
    .X(_04234_));
 sg13g2_nor2_1 _21812_ (.A(_08852_),
    .B(_04234_),
    .Y(_04235_));
 sg13g2_nand3_1 _21813_ (.B(_08841_),
    .C(_04235_),
    .A(_08824_),
    .Y(_04236_));
 sg13g2_xnor2_1 _21814_ (.Y(_04237_),
    .A(_03652_),
    .B(_04236_));
 sg13g2_buf_1 _21815_ (.A(net84),
    .X(_04238_));
 sg13g2_a22oi_1 _21816_ (.Y(_04239_),
    .B1(_04237_),
    .B2(_04238_),
    .A2(net33),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_nor2_1 _21817_ (.A(_03638_),
    .B(net161),
    .Y(_04240_));
 sg13g2_o21ai_1 _21818_ (.B1(_04240_),
    .Y(_04241_),
    .A1(_03617_),
    .A2(_03629_));
 sg13g2_nor2_1 _21819_ (.A(_11570_),
    .B(_03638_),
    .Y(_04242_));
 sg13g2_o21ai_1 _21820_ (.B1(_04242_),
    .Y(_04243_),
    .A1(_03617_),
    .A2(_03629_));
 sg13g2_nand3_1 _21821_ (.B(_04241_),
    .C(_04243_),
    .A(_03665_),
    .Y(_04244_));
 sg13g2_nand2_1 _21822_ (.Y(_04245_),
    .A(_11770_),
    .B(_03645_));
 sg13g2_o21ai_1 _21823_ (.B1(_09202_),
    .Y(_04246_),
    .A1(_03661_),
    .A2(_04245_));
 sg13g2_a21oi_1 _21824_ (.A1(_03661_),
    .A2(_04245_),
    .Y(_04247_),
    .B1(_04246_));
 sg13g2_a22oi_1 _21825_ (.Y(_04248_),
    .B1(_03723_),
    .B2(_03715_),
    .A2(_03720_),
    .A1(_03713_));
 sg13g2_buf_8 _21826_ (.A(_04248_),
    .X(_04249_));
 sg13g2_nand2_1 _21827_ (.Y(_04250_),
    .A(_10566_),
    .B(_03732_));
 sg13g2_o21ai_1 _21828_ (.B1(_03729_),
    .Y(_04251_),
    .A1(_04249_),
    .A2(_04250_));
 sg13g2_a221oi_1 _21829_ (.B2(net182),
    .C1(net206),
    .B1(_04249_),
    .A1(_11222_),
    .Y(_04252_),
    .A2(_03584_));
 sg13g2_buf_1 _21830_ (.A(_04252_),
    .X(_04253_));
 sg13g2_nand2_1 _21831_ (.Y(_04254_),
    .A(_03727_),
    .B(_03736_));
 sg13g2_inv_1 _21832_ (.Y(_04255_),
    .A(_04254_));
 sg13g2_nor3_1 _21833_ (.A(_04251_),
    .B(_04253_),
    .C(_04255_),
    .Y(_04256_));
 sg13g2_o21ai_1 _21834_ (.B1(_04255_),
    .Y(_04257_),
    .A1(_04251_),
    .A2(_04253_));
 sg13g2_nand3b_1 _21835_ (.B(_09916_),
    .C(_04257_),
    .Y(_04258_),
    .A_N(_04256_));
 sg13g2_buf_1 _21836_ (.A(_04258_),
    .X(_04259_));
 sg13g2_nor2_1 _21837_ (.A(net127),
    .B(net147),
    .Y(_04260_));
 sg13g2_inv_1 _21838_ (.Y(_04261_),
    .A(net151));
 sg13g2_a221oi_1 _21839_ (.B2(net163),
    .C1(net158),
    .B1(_04199_),
    .A1(_03684_),
    .Y(_04262_),
    .A2(_04183_));
 sg13g2_o21ai_1 _21840_ (.B1(_04262_),
    .Y(_04263_),
    .A1(net166),
    .A2(_04261_));
 sg13g2_a21oi_1 _21841_ (.A1(_04127_),
    .A2(_11576_),
    .Y(_04264_),
    .B1(net166));
 sg13g2_nand2b_1 _21842_ (.Y(_04265_),
    .B(_04262_),
    .A_N(_04264_));
 sg13g2_a22oi_1 _21843_ (.Y(_04266_),
    .B1(_04265_),
    .B2(net1097),
    .A2(_04263_),
    .A1(net1135));
 sg13g2_or2_1 _21844_ (.X(_04267_),
    .B(_04266_),
    .A(_04260_));
 sg13g2_mux2_1 _21845_ (.A0(_09130_),
    .A1(_09195_),
    .S(_03659_),
    .X(_04268_));
 sg13g2_or2_1 _21846_ (.X(_04269_),
    .B(_04268_),
    .A(_09921_));
 sg13g2_a22oi_1 _21847_ (.Y(_04270_),
    .B1(_04161_),
    .B2(net212),
    .A2(net151),
    .A1(net183));
 sg13g2_a22oi_1 _21848_ (.Y(_04271_),
    .B1(_04164_),
    .B2(_03587_),
    .A2(net179),
    .A1(net155));
 sg13g2_nand2_1 _21849_ (.Y(_04272_),
    .A(_10679_),
    .B(net180));
 sg13g2_a22oi_1 _21850_ (.Y(_04273_),
    .B1(net149),
    .B2(net152),
    .A2(_04173_),
    .A1(net181));
 sg13g2_and4_1 _21851_ (.A(_04270_),
    .B(_04271_),
    .C(_04272_),
    .D(_04273_),
    .X(_04274_));
 sg13g2_a21oi_1 _21852_ (.A1(net165),
    .A2(_04199_),
    .Y(_04275_),
    .B1(net124));
 sg13g2_buf_1 _21853_ (.A(_04142_),
    .X(_04276_));
 sg13g2_nand2_1 _21854_ (.Y(_04277_),
    .A(_04180_),
    .B(_04276_));
 sg13g2_nand2_1 _21855_ (.Y(_04278_),
    .A(net162),
    .B(net121));
 sg13g2_nand4_1 _21856_ (.B(_04275_),
    .C(_04277_),
    .A(_04274_),
    .Y(_04279_),
    .D(_04278_));
 sg13g2_a21oi_1 _21857_ (.A1(_03645_),
    .A2(_04131_),
    .Y(_04280_),
    .B1(_09926_));
 sg13g2_nand2_1 _21858_ (.Y(_04281_),
    .A(net169),
    .B(_03641_));
 sg13g2_nor3_1 _21859_ (.A(net848),
    .B(_03661_),
    .C(_04281_),
    .Y(_04282_));
 sg13g2_a21o_1 _21860_ (.A2(net262),
    .A1(net1148),
    .B1(_04282_),
    .X(_04283_));
 sg13g2_a221oi_1 _21861_ (.B2(_04280_),
    .C1(_04283_),
    .B1(_04279_),
    .A1(_03656_),
    .Y(_04284_),
    .A2(_04269_));
 sg13g2_nand4_1 _21862_ (.B(_04259_),
    .C(_04267_),
    .A(net509),
    .Y(_04285_),
    .D(_04284_));
 sg13g2_a21oi_1 _21863_ (.A1(_04244_),
    .A2(_04247_),
    .Y(_04286_),
    .B1(_04285_));
 sg13g2_and3_1 _21864_ (.X(_04287_),
    .A(_03665_),
    .B(_04241_),
    .C(_04243_));
 sg13g2_nand4_1 _21865_ (.B(_03661_),
    .C(_04281_),
    .A(net1073),
    .Y(_04288_),
    .D(_04287_));
 sg13g2_inv_1 _21866_ (.Y(_04289_),
    .A(_03643_));
 sg13g2_a21oi_1 _21867_ (.A1(_03646_),
    .A2(_03757_),
    .Y(_04290_),
    .B1(_04289_));
 sg13g2_xnor2_1 _21868_ (.Y(_04291_),
    .A(_03661_),
    .B(_04290_));
 sg13g2_and2_1 _21869_ (.A(_04112_),
    .B(_04113_),
    .X(_04292_));
 sg13g2_buf_2 _21870_ (.A(_04292_),
    .X(_04293_));
 sg13g2_a221oi_1 _21871_ (.B2(_04293_),
    .C1(net160),
    .B1(_04291_),
    .A1(_04286_),
    .Y(_04294_),
    .A2(_04288_));
 sg13g2_o21ai_1 _21872_ (.B1(_10251_),
    .Y(_04295_),
    .A1(_09303_),
    .A2(_09389_));
 sg13g2_buf_1 _21873_ (.A(_04295_),
    .X(_04296_));
 sg13g2_buf_1 _21874_ (.A(_04296_),
    .X(_04297_));
 sg13g2_nor2_1 _21875_ (.A(_04297_),
    .B(_11831_),
    .Y(_04298_));
 sg13g2_o21ai_1 _21876_ (.B1(_04217_),
    .Y(_04299_),
    .A1(_04294_),
    .A2(_04298_));
 sg13g2_nand2_1 _21877_ (.Y(_00985_),
    .A(_04239_),
    .B(_04299_));
 sg13g2_nor2_1 _21878_ (.A(net178),
    .B(\cpu.ex.c_mult[12] ),
    .Y(_04300_));
 sg13g2_nand2_1 _21879_ (.Y(_04301_),
    .A(_03664_),
    .B(_03669_));
 sg13g2_xor2_1 _21880_ (.B(_03749_),
    .A(_04301_),
    .X(_04302_));
 sg13g2_o21ai_1 _21881_ (.B1(_11507_),
    .Y(_04303_),
    .A1(_03643_),
    .A2(_03655_));
 sg13g2_nand2_1 _21882_ (.Y(_04304_),
    .A(_03643_),
    .B(_03655_));
 sg13g2_o21ai_1 _21883_ (.B1(_03656_),
    .Y(_04305_),
    .A1(net132),
    .A2(net153));
 sg13g2_inv_1 _21884_ (.Y(_04306_),
    .A(_04305_));
 sg13g2_a22oi_1 _21885_ (.Y(_04307_),
    .B1(_04306_),
    .B2(_03757_),
    .A2(_04304_),
    .A1(_04303_));
 sg13g2_xor2_1 _21886_ (.B(_04307_),
    .A(_03749_),
    .X(_04308_));
 sg13g2_and2_1 _21887_ (.A(_04296_),
    .B(_04259_),
    .X(_04309_));
 sg13g2_buf_1 _21888_ (.A(_04309_),
    .X(_04310_));
 sg13g2_and2_1 _21889_ (.A(net181),
    .B(_04146_),
    .X(_04311_));
 sg13g2_a221oi_1 _21890_ (.B2(net148),
    .C1(_04311_),
    .B1(net123),
    .A1(net211),
    .Y(_04312_),
    .A2(net118));
 sg13g2_buf_1 _21891_ (.A(net121),
    .X(_04313_));
 sg13g2_nand2_2 _21892_ (.Y(_04314_),
    .A(_04127_),
    .B(_04171_));
 sg13g2_nor2_1 _21893_ (.A(net161),
    .B(_04314_),
    .Y(_04315_));
 sg13g2_a221oi_1 _21894_ (.B2(net153),
    .C1(_04315_),
    .B1(net99),
    .A1(net152),
    .Y(_04316_),
    .A2(net157));
 sg13g2_a21oi_1 _21895_ (.A1(net155),
    .A2(net149),
    .Y(_04317_),
    .B1(net158));
 sg13g2_buf_1 _21896_ (.A(_04178_),
    .X(_04318_));
 sg13g2_a22oi_1 _21897_ (.Y(_04319_),
    .B1(net122),
    .B2(net150),
    .A2(net117),
    .A1(net126));
 sg13g2_buf_1 _21898_ (.A(net212),
    .X(_04320_));
 sg13g2_a22oi_1 _21899_ (.Y(_04321_),
    .B1(_04173_),
    .B2(net195),
    .A2(net156),
    .A1(net183));
 sg13g2_and2_1 _21900_ (.A(_04319_),
    .B(_04321_),
    .X(_04322_));
 sg13g2_nand4_1 _21901_ (.B(_04316_),
    .C(_04317_),
    .A(_04312_),
    .Y(_04323_),
    .D(_04322_));
 sg13g2_nor2_1 _21902_ (.A(net154),
    .B(net147),
    .Y(_04324_));
 sg13g2_nor2_1 _21903_ (.A(net903),
    .B(_04324_),
    .Y(_04325_));
 sg13g2_o21ai_1 _21904_ (.B1(net147),
    .Y(_04326_),
    .A1(net166),
    .A2(_04314_));
 sg13g2_a221oi_1 _21905_ (.B2(net1097),
    .C1(_04326_),
    .B1(_04264_),
    .A1(net120),
    .Y(_04327_),
    .A2(net99));
 sg13g2_buf_1 _21906_ (.A(net124),
    .X(_04328_));
 sg13g2_a21o_1 _21907_ (.A2(_04328_),
    .A1(_03579_),
    .B1(net847),
    .X(_04329_));
 sg13g2_nand2_1 _21908_ (.Y(_04330_),
    .A(net191),
    .B(net164));
 sg13g2_mux2_1 _21909_ (.A0(net1075),
    .A1(net1074),
    .S(_04330_),
    .X(_04331_));
 sg13g2_or2_1 _21910_ (.X(_04332_),
    .B(net164),
    .A(_11460_));
 sg13g2_buf_1 _21911_ (.A(_04332_),
    .X(_04333_));
 sg13g2_o21ai_1 _21912_ (.B1(_04333_),
    .Y(_04334_),
    .A1(net1059),
    .A2(_04331_));
 sg13g2_o21ai_1 _21913_ (.B1(_04334_),
    .Y(_04335_),
    .A1(_04327_),
    .A2(_04329_));
 sg13g2_a221oi_1 _21914_ (.B2(_04325_),
    .C1(_04335_),
    .B1(_04323_),
    .A1(net1076),
    .Y(_04336_),
    .A2(_11155_));
 sg13g2_nand2_1 _21915_ (.Y(_04337_),
    .A(_04310_),
    .B(_04336_));
 sg13g2_a221oi_1 _21916_ (.B2(_04293_),
    .C1(_04337_),
    .B1(_04308_),
    .A1(net1073),
    .Y(_04338_),
    .A2(_04302_));
 sg13g2_or2_1 _21917_ (.X(_04339_),
    .B(_04338_),
    .A(_04300_));
 sg13g2_nor2_2 _21918_ (.A(_08883_),
    .B(_04236_),
    .Y(_04340_));
 sg13g2_xnor2_1 _21919_ (.Y(_04341_),
    .A(_00291_),
    .B(_04340_));
 sg13g2_a22oi_1 _21920_ (.Y(_04342_),
    .B1(_04341_),
    .B2(net75),
    .A2(net33),
    .A1(net821));
 sg13g2_o21ai_1 _21921_ (.B1(_04342_),
    .Y(_00986_),
    .A1(net76),
    .A2(_04339_));
 sg13g2_nor3_1 _21922_ (.A(net178),
    .B(_11883_),
    .C(_11884_),
    .Y(_04343_));
 sg13g2_and2_1 _21923_ (.A(_03748_),
    .B(_04333_),
    .X(_04344_));
 sg13g2_nor2b_1 _21924_ (.A(_03748_),
    .B_N(_04330_),
    .Y(_04345_));
 sg13g2_mux2_1 _21925_ (.A0(_04344_),
    .A1(_04345_),
    .S(_04307_),
    .X(_04346_));
 sg13g2_a21oi_1 _21926_ (.A1(_03664_),
    .A2(_03674_),
    .Y(_04347_),
    .B1(_03675_));
 sg13g2_xor2_1 _21927_ (.B(_03748_),
    .A(_04347_),
    .X(_04348_));
 sg13g2_nand2b_1 _21928_ (.Y(_04349_),
    .B(_03748_),
    .A_N(_04330_));
 sg13g2_o21ai_1 _21929_ (.B1(_04349_),
    .Y(_04350_),
    .A1(_03748_),
    .A2(_04333_));
 sg13g2_nor2_1 _21930_ (.A(net161),
    .B(_04261_),
    .Y(_04351_));
 sg13g2_nand2_1 _21931_ (.Y(_04352_),
    .A(_04127_),
    .B(_04159_));
 sg13g2_nor2_1 _21932_ (.A(_03655_),
    .B(_04352_),
    .Y(_04353_));
 sg13g2_nand3_1 _21933_ (.B(net221),
    .C(_04128_),
    .A(_11064_),
    .Y(_04354_));
 sg13g2_buf_1 _21934_ (.A(_04354_),
    .X(_04355_));
 sg13g2_nand2_1 _21935_ (.Y(_04356_),
    .A(_04180_),
    .B(net123));
 sg13g2_o21ai_1 _21936_ (.B1(_04356_),
    .Y(_04357_),
    .A1(_03632_),
    .A2(_04355_));
 sg13g2_nand2_1 _21937_ (.Y(_04358_),
    .A(_04171_),
    .B(_04140_));
 sg13g2_a22oi_1 _21938_ (.Y(_04359_),
    .B1(net122),
    .B2(net211),
    .A2(_04197_),
    .A1(_04101_));
 sg13g2_o21ai_1 _21939_ (.B1(_04359_),
    .Y(_04360_),
    .A1(_03593_),
    .A2(_04358_));
 sg13g2_nor4_1 _21940_ (.A(_04351_),
    .B(_04353_),
    .C(_04357_),
    .D(_04360_),
    .Y(_04361_));
 sg13g2_a22oi_1 _21941_ (.Y(_04362_),
    .B1(_04146_),
    .B2(net195),
    .A2(net157),
    .A1(net155));
 sg13g2_a22oi_1 _21942_ (.Y(_04363_),
    .B1(net119),
    .B2(_04166_),
    .A2(net118),
    .A1(net152));
 sg13g2_nand4_1 _21943_ (.B(_04361_),
    .C(_04362_),
    .A(_04187_),
    .Y(_04364_),
    .D(_04363_));
 sg13g2_nor2_1 _21944_ (.A(net903),
    .B(_04260_),
    .Y(_04365_));
 sg13g2_a22oi_1 _21945_ (.Y(_04366_),
    .B1(net99),
    .B2(net125),
    .A2(_04328_),
    .A1(net120));
 sg13g2_nand2b_1 _21946_ (.Y(_04367_),
    .B(net1135),
    .A_N(_04366_));
 sg13g2_nand2_1 _21947_ (.Y(_04368_),
    .A(_03576_),
    .B(_04207_));
 sg13g2_nand2_1 _21948_ (.Y(_04369_),
    .A(_03682_),
    .B(net124));
 sg13g2_nand3_1 _21949_ (.B(_04368_),
    .C(_04369_),
    .A(net1097),
    .Y(_04370_));
 sg13g2_nand2_1 _21950_ (.Y(_04371_),
    .A(net1076),
    .B(net225));
 sg13g2_mux2_1 _21951_ (.A0(net1075),
    .A1(net1074),
    .S(_03702_),
    .X(_04372_));
 sg13g2_o21ai_1 _21952_ (.B1(_03697_),
    .Y(_04373_),
    .A1(net1059),
    .A2(_04372_));
 sg13g2_nand4_1 _21953_ (.B(_04370_),
    .C(_04371_),
    .A(_04367_),
    .Y(_04374_),
    .D(_04373_));
 sg13g2_a221oi_1 _21954_ (.B2(_04365_),
    .C1(_04374_),
    .B1(_04364_),
    .A1(_04293_),
    .Y(_04375_),
    .A2(_04350_));
 sg13g2_nand2_1 _21955_ (.Y(_04376_),
    .A(_04310_),
    .B(_04375_));
 sg13g2_a221oi_1 _21956_ (.B2(_09203_),
    .C1(_04376_),
    .B1(_04348_),
    .A1(_04293_),
    .Y(_04377_),
    .A2(_04346_));
 sg13g2_a21o_1 _21957_ (.A2(_04343_),
    .A1(_11881_),
    .B1(_04377_),
    .X(_04378_));
 sg13g2_nand2_1 _21958_ (.Y(_04379_),
    .A(net821),
    .B(_04340_));
 sg13g2_xnor2_1 _21959_ (.Y(_04380_),
    .A(_03577_),
    .B(_04379_));
 sg13g2_a22oi_1 _21960_ (.Y(_04381_),
    .B1(_04380_),
    .B2(net75),
    .A2(net33),
    .A1(net714));
 sg13g2_o21ai_1 _21961_ (.B1(_04381_),
    .Y(_00987_),
    .A1(_04098_),
    .A2(_04378_));
 sg13g2_or2_1 _21962_ (.X(_04382_),
    .B(\cpu.ex.c_mult[14] ),
    .A(net178));
 sg13g2_inv_1 _21963_ (.Y(_04383_),
    .A(_03686_));
 sg13g2_and2_1 _21964_ (.A(_03762_),
    .B(_03761_),
    .X(_04384_));
 sg13g2_buf_1 _21965_ (.A(_04384_),
    .X(_04385_));
 sg13g2_or4_1 _21966_ (.A(_03692_),
    .B(_03677_),
    .C(_04383_),
    .D(_04385_),
    .X(_04386_));
 sg13g2_inv_1 _21967_ (.Y(_04387_),
    .A(_04385_));
 sg13g2_nor2_1 _21968_ (.A(_03692_),
    .B(_04387_),
    .Y(_04388_));
 sg13g2_o21ai_1 _21969_ (.B1(_04388_),
    .Y(_04389_),
    .A1(_03677_),
    .A2(_04383_));
 sg13g2_buf_1 _21970_ (.A(net149),
    .X(_04390_));
 sg13g2_a22oi_1 _21971_ (.Y(_04391_),
    .B1(net116),
    .B2(net126),
    .A2(net117),
    .A1(net153));
 sg13g2_a22oi_1 _21972_ (.Y(_04392_),
    .B1(_04146_),
    .B2(net148),
    .A2(_04197_),
    .A1(net195));
 sg13g2_nand2_1 _21973_ (.Y(_04393_),
    .A(net183),
    .B(net180));
 sg13g2_a22oi_1 _21974_ (.Y(_04394_),
    .B1(net122),
    .B2(net152),
    .A2(net118),
    .A1(net155));
 sg13g2_and4_1 _21975_ (.A(_04391_),
    .B(_04392_),
    .C(_04393_),
    .D(_04394_),
    .X(_04395_));
 sg13g2_nor2_1 _21976_ (.A(_03606_),
    .B(_04358_),
    .Y(_04396_));
 sg13g2_a221oi_1 _21977_ (.B2(_04102_),
    .C1(_04396_),
    .B1(_04170_),
    .A1(_04201_),
    .Y(_04397_),
    .A2(net123));
 sg13g2_a21oi_1 _21978_ (.A1(_04153_),
    .A2(_04200_),
    .Y(_04398_),
    .B1(net98));
 sg13g2_a22oi_1 _21979_ (.Y(_04399_),
    .B1(net99),
    .B2(net127),
    .A2(_04149_),
    .A1(net162));
 sg13g2_nand4_1 _21980_ (.B(_04397_),
    .C(_04398_),
    .A(_04395_),
    .Y(_04400_),
    .D(_04399_));
 sg13g2_a21oi_1 _21981_ (.A1(_03579_),
    .A2(net100),
    .Y(_04401_),
    .B1(_09926_));
 sg13g2_nand2_1 _21982_ (.Y(_04402_),
    .A(_09038_),
    .B(net222));
 sg13g2_nand3_1 _21983_ (.B(net125),
    .C(net100),
    .A(net1135),
    .Y(_04403_));
 sg13g2_mux2_1 _21984_ (.A0(_09131_),
    .A1(_09196_),
    .S(_03762_),
    .X(_04404_));
 sg13g2_o21ai_1 _21985_ (.B1(_03761_),
    .Y(_04405_),
    .A1(_09922_),
    .A2(_04404_));
 sg13g2_nand3_1 _21986_ (.B(_04403_),
    .C(_04405_),
    .A(_04402_),
    .Y(_04406_));
 sg13g2_a21oi_1 _21987_ (.A1(_04400_),
    .A2(_04401_),
    .Y(_04407_),
    .B1(_04406_));
 sg13g2_nor2_1 _21988_ (.A(_04251_),
    .B(_04253_),
    .Y(_04408_));
 sg13g2_xnor2_1 _21989_ (.Y(_04409_),
    .A(_04408_),
    .B(_04255_));
 sg13g2_a221oi_1 _21990_ (.B2(_09916_),
    .C1(net160),
    .B1(_04409_),
    .A1(_08296_),
    .Y(_04410_),
    .A2(net125));
 sg13g2_nand4_1 _21991_ (.B(_04389_),
    .C(_04407_),
    .A(_04386_),
    .Y(_04411_),
    .D(_04410_));
 sg13g2_and4_1 _21992_ (.A(_11607_),
    .B(_11908_),
    .C(_11910_),
    .D(_11911_),
    .X(_04412_));
 sg13g2_nor3_1 _21993_ (.A(net509),
    .B(_04412_),
    .C(_04387_),
    .Y(_04413_));
 sg13g2_nor3_1 _21994_ (.A(net509),
    .B(_04412_),
    .C(_04385_),
    .Y(_04414_));
 sg13g2_mux2_1 _21995_ (.A0(_04413_),
    .A1(_04414_),
    .S(_03760_),
    .X(_04415_));
 sg13g2_a21oi_1 _21996_ (.A1(_04382_),
    .A2(_04411_),
    .Y(_04416_),
    .B1(_04415_));
 sg13g2_nand3_1 _21997_ (.B(net714),
    .C(_04340_),
    .A(_08463_),
    .Y(_04417_));
 sg13g2_xnor2_1 _21998_ (.Y(_04418_),
    .A(_10842_),
    .B(_04417_));
 sg13g2_a22oi_1 _21999_ (.Y(_04419_),
    .B1(_04418_),
    .B2(net75),
    .A2(_04227_),
    .A1(net817));
 sg13g2_o21ai_1 _22000_ (.B1(_04419_),
    .Y(_00988_),
    .A1(net76),
    .A2(_04416_));
 sg13g2_nand2_1 _22001_ (.Y(_04420_),
    .A(_03695_),
    .B(_03768_));
 sg13g2_nand3_1 _22002_ (.B(_03689_),
    .C(_04420_),
    .A(net1073),
    .Y(_04421_));
 sg13g2_nand2b_1 _22003_ (.Y(_04422_),
    .B(_03686_),
    .A_N(_03677_));
 sg13g2_and4_1 _22004_ (.A(_09203_),
    .B(_03688_),
    .C(_03695_),
    .D(_03768_),
    .X(_04423_));
 sg13g2_nand2_1 _22005_ (.Y(_04424_),
    .A(_09202_),
    .B(net120));
 sg13g2_o21ai_1 _22006_ (.B1(_04424_),
    .Y(_04425_),
    .A1(net120),
    .A2(net509));
 sg13g2_a21o_1 _22007_ (.A2(_04425_),
    .A1(net168),
    .B1(_04420_),
    .X(_04426_));
 sg13g2_o21ai_1 _22008_ (.B1(_04420_),
    .Y(_04427_),
    .A1(_03762_),
    .A2(_04115_));
 sg13g2_a22oi_1 _22009_ (.Y(_04428_),
    .B1(_04426_),
    .B2(_04427_),
    .A2(_11190_),
    .A1(_09038_));
 sg13g2_mux2_1 _22010_ (.A0(_09131_),
    .A1(_09196_),
    .S(_03768_),
    .X(_04429_));
 sg13g2_o21ai_1 _22011_ (.B1(_03695_),
    .Y(_04430_),
    .A1(_09922_),
    .A2(_04429_));
 sg13g2_a21oi_1 _22012_ (.A1(net128),
    .A2(_04313_),
    .Y(_04431_),
    .B1(net100));
 sg13g2_a22oi_1 _22013_ (.Y(_04432_),
    .B1(_04170_),
    .B2(net195),
    .A2(net117),
    .A1(_04153_));
 sg13g2_a22oi_1 _22014_ (.Y(_04433_),
    .B1(net119),
    .B2(net127),
    .A2(net118),
    .A1(net183));
 sg13g2_a22oi_1 _22015_ (.Y(_04434_),
    .B1(net122),
    .B2(_04151_),
    .A2(net123),
    .A1(net152));
 sg13g2_a22oi_1 _22016_ (.Y(_04435_),
    .B1(net116),
    .B2(net162),
    .A2(_04197_),
    .A1(net148));
 sg13g2_and4_1 _22017_ (.A(_04432_),
    .B(_04433_),
    .C(_04434_),
    .D(_04435_),
    .X(_04436_));
 sg13g2_nor2_1 _22018_ (.A(_10603_),
    .B(_04358_),
    .Y(_04437_));
 sg13g2_a221oi_1 _22019_ (.B2(_04102_),
    .C1(_04437_),
    .B1(_04191_),
    .A1(net150),
    .Y(_04438_),
    .A2(_04146_));
 sg13g2_nor2_1 _22020_ (.A(_03645_),
    .B(_04355_),
    .Y(_04439_));
 sg13g2_a21oi_1 _22021_ (.A1(net126),
    .A2(net157),
    .Y(_04440_),
    .B1(_04439_));
 sg13g2_nand4_1 _22022_ (.B(_04436_),
    .C(_04438_),
    .A(_04431_),
    .Y(_04441_),
    .D(_04440_));
 sg13g2_nand3_1 _22023_ (.B(_04369_),
    .C(_04441_),
    .A(_09924_),
    .Y(_04442_));
 sg13g2_nand4_1 _22024_ (.B(_04428_),
    .C(_04430_),
    .A(_04410_),
    .Y(_04443_),
    .D(_04442_));
 sg13g2_a21oi_1 _22025_ (.A1(_04422_),
    .A2(_04423_),
    .Y(_04444_),
    .B1(_04443_));
 sg13g2_nand4_1 _22026_ (.B(_03762_),
    .C(_03768_),
    .A(_03695_),
    .Y(_04445_),
    .D(_04293_));
 sg13g2_nand3_1 _22027_ (.B(_04293_),
    .C(_04420_),
    .A(_03761_),
    .Y(_04446_));
 sg13g2_mux2_1 _22028_ (.A0(_04445_),
    .A1(_04446_),
    .S(_03760_),
    .X(_04447_));
 sg13g2_nand3_1 _22029_ (.B(_04444_),
    .C(_04447_),
    .A(_04421_),
    .Y(_04448_));
 sg13g2_nor3_1 _22030_ (.A(net178),
    .B(_11928_),
    .C(_11934_),
    .Y(_04449_));
 sg13g2_nor2_1 _22031_ (.A(_04097_),
    .B(_04449_),
    .Y(_04450_));
 sg13g2_nand4_1 _22032_ (.B(net714),
    .C(net817),
    .A(_08463_),
    .Y(_04451_),
    .D(_04340_));
 sg13g2_xnor2_1 _22033_ (.Y(_04452_),
    .A(_10745_),
    .B(_04451_));
 sg13g2_a22oi_1 _22034_ (.Y(_04453_),
    .B1(_04452_),
    .B2(net84),
    .A2(_04226_),
    .A1(_08375_));
 sg13g2_inv_1 _22035_ (.Y(_04454_),
    .A(_04453_));
 sg13g2_a21o_1 _22036_ (.A2(_04450_),
    .A1(_04448_),
    .B1(_04454_),
    .X(_00989_));
 sg13g2_o21ai_1 _22037_ (.B1(_11578_),
    .Y(_04455_),
    .A1(_11574_),
    .A2(_04144_));
 sg13g2_o21ai_1 _22038_ (.B1(net147),
    .Y(_04456_),
    .A1(net182),
    .A2(_04314_));
 sg13g2_a21oi_1 _22039_ (.A1(_04193_),
    .A2(_04455_),
    .Y(_04457_),
    .B1(_04456_));
 sg13g2_a22oi_1 _22040_ (.Y(_04458_),
    .B1(net116),
    .B2(net126),
    .A2(net156),
    .A1(net183));
 sg13g2_a22oi_1 _22041_ (.Y(_04459_),
    .B1(net99),
    .B2(_04201_),
    .A2(net118),
    .A1(net153));
 sg13g2_nand3_1 _22042_ (.B(_04458_),
    .C(_04459_),
    .A(_04457_),
    .Y(_04460_));
 sg13g2_nand2_1 _22043_ (.Y(_04461_),
    .A(net128),
    .B(_04173_));
 sg13g2_a22oi_1 _22044_ (.Y(_04462_),
    .B1(_04146_),
    .B2(net120),
    .A2(_04197_),
    .A1(net125));
 sg13g2_a22oi_1 _22045_ (.Y(_04463_),
    .B1(_04165_),
    .B2(net154),
    .A2(_04162_),
    .A1(net127));
 sg13g2_a22oi_1 _22046_ (.Y(_04464_),
    .B1(net117),
    .B2(net155),
    .A2(net157),
    .A1(net162));
 sg13g2_nand4_1 _22047_ (.B(_04462_),
    .C(_04463_),
    .A(_04461_),
    .Y(_04465_),
    .D(_04464_));
 sg13g2_a21oi_1 _22048_ (.A1(_03606_),
    .A2(_04132_),
    .Y(_04466_),
    .B1(_04109_));
 sg13g2_o21ai_1 _22049_ (.B1(_04466_),
    .Y(_04467_),
    .A1(_04460_),
    .A2(_04465_));
 sg13g2_a22oi_1 _22050_ (.Y(_04468_),
    .B1(net99),
    .B2(net159),
    .A2(net98),
    .A1(net195));
 sg13g2_inv_1 _22051_ (.Y(_04469_),
    .A(_04468_));
 sg13g2_nor2_1 _22052_ (.A(net221),
    .B(_03587_),
    .Y(_04470_));
 sg13g2_nand2_1 _22053_ (.Y(_04471_),
    .A(_11638_),
    .B(net148));
 sg13g2_a21oi_1 _22054_ (.A1(net1074),
    .A2(_04471_),
    .Y(_04472_),
    .B1(net1134));
 sg13g2_nor2_1 _22055_ (.A(_11229_),
    .B(_03593_),
    .Y(_04473_));
 sg13g2_a221oi_1 _22056_ (.B2(net1075),
    .C1(net188),
    .B1(_04473_),
    .A1(net1148),
    .Y(_04474_),
    .A2(net132));
 sg13g2_o21ai_1 _22057_ (.B1(_04474_),
    .Y(_04475_),
    .A1(_04470_),
    .A2(_04472_));
 sg13g2_a21oi_1 _22058_ (.A1(_09924_),
    .A2(_04469_),
    .Y(_04476_),
    .B1(_04475_));
 sg13g2_a21oi_1 _22059_ (.A1(_03598_),
    .A2(_03599_),
    .Y(_04477_),
    .B1(_03600_));
 sg13g2_nor2_1 _22060_ (.A(_04473_),
    .B(_04470_),
    .Y(_04478_));
 sg13g2_xnor2_1 _22061_ (.Y(_04479_),
    .A(_04477_),
    .B(_04478_));
 sg13g2_o21ai_1 _22062_ (.B1(_04105_),
    .Y(_04480_),
    .A1(_03707_),
    .A2(_03708_));
 sg13g2_xor2_1 _22063_ (.B(_04478_),
    .A(_04480_),
    .X(_04481_));
 sg13g2_a22oi_1 _22064_ (.Y(_04482_),
    .B1(_04481_),
    .B2(_04118_),
    .A2(_04479_),
    .A1(_09202_));
 sg13g2_nand3_1 _22065_ (.B(_04476_),
    .C(_04482_),
    .A(_04467_),
    .Y(_04483_));
 sg13g2_o21ai_1 _22066_ (.B1(_04483_),
    .Y(_04484_),
    .A1(net178),
    .A2(\cpu.ex.c_mult[2] ));
 sg13g2_a21o_1 _22067_ (.A2(net84),
    .A1(net1077),
    .B1(_04226_),
    .X(_04485_));
 sg13g2_nor2_1 _22068_ (.A(net812),
    .B(net1077),
    .Y(_04486_));
 sg13g2_nor3_1 _22069_ (.A(_08362_),
    .B(_11943_),
    .C(_04218_),
    .Y(_04487_));
 sg13g2_a221oi_1 _22070_ (.B2(net84),
    .C1(_04487_),
    .B1(_04486_),
    .A1(net812),
    .Y(_04488_),
    .A2(_04485_));
 sg13g2_o21ai_1 _22071_ (.B1(_04488_),
    .Y(_00990_),
    .A1(net76),
    .A2(_04484_));
 sg13g2_a22oi_1 _22072_ (.Y(_04489_),
    .B1(net119),
    .B2(net159),
    .A2(net121),
    .A1(net195));
 sg13g2_nand2_1 _22073_ (.Y(_04490_),
    .A(net147),
    .B(_04489_));
 sg13g2_nor2_1 _22074_ (.A(net903),
    .B(_04208_),
    .Y(_04491_));
 sg13g2_a221oi_1 _22075_ (.B2(_04491_),
    .C1(_04099_),
    .B1(_04490_),
    .A1(net1076),
    .Y(_04492_),
    .A2(_11491_));
 sg13g2_mux2_1 _22076_ (.A0(net1075),
    .A1(net1074),
    .S(_03722_),
    .X(_04493_));
 sg13g2_o21ai_1 _22077_ (.B1(_03718_),
    .Y(_04494_),
    .A1(net1059),
    .A2(_04493_));
 sg13g2_a22oi_1 _22078_ (.Y(_04495_),
    .B1(net116),
    .B2(net162),
    .A2(net156),
    .A1(_03705_));
 sg13g2_a22oi_1 _22079_ (.Y(_04496_),
    .B1(_04146_),
    .B2(net125),
    .A2(net157),
    .A1(net153));
 sg13g2_a22oi_1 _22080_ (.Y(_04497_),
    .B1(net123),
    .B2(net128),
    .A2(net118),
    .A1(net154));
 sg13g2_a22oi_1 _22081_ (.Y(_04498_),
    .B1(_04173_),
    .B2(net120),
    .A2(net122),
    .A1(net127));
 sg13g2_nand4_1 _22082_ (.B(_04496_),
    .C(_04497_),
    .A(_04495_),
    .Y(_04499_),
    .D(_04498_));
 sg13g2_nand2_1 _22083_ (.Y(_04500_),
    .A(net183),
    .B(net117));
 sg13g2_nand2_1 _22084_ (.Y(_04501_),
    .A(_04176_),
    .B(net121));
 sg13g2_a21oi_1 _22085_ (.A1(_11576_),
    .A2(_04168_),
    .Y(_04502_),
    .B1(_04189_));
 sg13g2_nand2b_1 _22086_ (.Y(_04503_),
    .B(_04193_),
    .A_N(_04502_));
 sg13g2_a21oi_1 _22087_ (.A1(net155),
    .A2(net119),
    .Y(_04504_),
    .B1(net124));
 sg13g2_nand4_1 _22088_ (.B(_04501_),
    .C(_04503_),
    .A(_04500_),
    .Y(_04505_),
    .D(_04504_));
 sg13g2_a21oi_1 _22089_ (.A1(_10603_),
    .A2(net98),
    .Y(_04506_),
    .B1(net847));
 sg13g2_o21ai_1 _22090_ (.B1(_04506_),
    .Y(_04507_),
    .A1(_04499_),
    .A2(_04505_));
 sg13g2_nor2_1 _22091_ (.A(_03602_),
    .B(_03604_),
    .Y(_04508_));
 sg13g2_and2_1 _22092_ (.A(_03718_),
    .B(_03722_),
    .X(_04509_));
 sg13g2_xor2_1 _22093_ (.B(_04509_),
    .A(_04508_),
    .X(_04510_));
 sg13g2_and2_1 _22094_ (.A(_03713_),
    .B(_03716_),
    .X(_04511_));
 sg13g2_xor2_1 _22095_ (.B(_04511_),
    .A(_04509_),
    .X(_04512_));
 sg13g2_a22oi_1 _22096_ (.Y(_04513_),
    .B1(_04512_),
    .B2(_04118_),
    .A2(_04510_),
    .A1(_09202_));
 sg13g2_nand4_1 _22097_ (.B(_04494_),
    .C(_04507_),
    .A(_04492_),
    .Y(_04514_),
    .D(_04513_));
 sg13g2_o21ai_1 _22098_ (.B1(_04514_),
    .Y(_04515_),
    .A1(_04296_),
    .A2(\cpu.ex.c_mult[3] ));
 sg13g2_nand2_1 _22099_ (.Y(_04516_),
    .A(net812),
    .B(net696));
 sg13g2_a21o_1 _22100_ (.A2(_04516_),
    .A1(_04214_),
    .B1(_04226_),
    .X(_04517_));
 sg13g2_nor2_1 _22101_ (.A(net698),
    .B(_04516_),
    .Y(_04518_));
 sg13g2_inv_1 _22102_ (.Y(_04519_),
    .A(_00276_));
 sg13g2_a21o_1 _22103_ (.A2(_04487_),
    .A1(_04519_),
    .B1(_04222_),
    .X(_04520_));
 sg13g2_a221oi_1 _22104_ (.B2(_04214_),
    .C1(_04520_),
    .B1(_04518_),
    .A1(net698),
    .Y(_04521_),
    .A2(_04517_));
 sg13g2_o21ai_1 _22105_ (.B1(_04521_),
    .Y(_00991_),
    .A1(net76),
    .A2(_04515_));
 sg13g2_a21oi_1 _22106_ (.A1(_11578_),
    .A2(_04144_),
    .Y(_04522_),
    .B1(net166));
 sg13g2_o21ai_1 _22107_ (.B1(net147),
    .Y(_04523_),
    .A1(_03624_),
    .A2(_04314_));
 sg13g2_a221oi_1 _22108_ (.B2(net164),
    .C1(_04523_),
    .B1(_04142_),
    .A1(net154),
    .Y(_04524_),
    .A2(_04138_));
 sg13g2_nor2_1 _22109_ (.A(_03575_),
    .B(_04358_),
    .Y(_04525_));
 sg13g2_a21oi_1 _22110_ (.A1(_03641_),
    .A2(net149),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_a22oi_1 _22111_ (.Y(_04527_),
    .B1(_04164_),
    .B2(net128),
    .A2(net123),
    .A1(net163));
 sg13g2_nor2_1 _22112_ (.A(_03584_),
    .B(_04352_),
    .Y(_04528_));
 sg13g2_a221oi_1 _22113_ (.B2(_03743_),
    .C1(_04528_),
    .B1(net179),
    .A1(net165),
    .Y(_04529_),
    .A2(net151));
 sg13g2_nand4_1 _22114_ (.B(_04526_),
    .C(_04527_),
    .A(_04524_),
    .Y(_04530_),
    .D(_04529_));
 sg13g2_o21ai_1 _22115_ (.B1(net1097),
    .Y(_04531_),
    .A1(_04522_),
    .A2(_04530_));
 sg13g2_nand2_1 _22116_ (.Y(_04532_),
    .A(net1135),
    .B(_04530_));
 sg13g2_a22oi_1 _22117_ (.Y(_04533_),
    .B1(_04531_),
    .B2(_04532_),
    .A2(_04132_),
    .A1(_03725_));
 sg13g2_nand2_1 _22118_ (.Y(_04534_),
    .A(net265),
    .B(net211));
 sg13g2_mux2_1 _22119_ (.A0(net1147),
    .A1(_09195_),
    .S(_04534_),
    .X(_04535_));
 sg13g2_o21ai_1 _22120_ (.B1(_03715_),
    .Y(_04536_),
    .A1(net1134),
    .A2(_04535_));
 sg13g2_a21oi_1 _22121_ (.A1(net1148),
    .A2(_11460_),
    .Y(_04537_),
    .B1(net188));
 sg13g2_nand2_1 _22122_ (.Y(_04538_),
    .A(_04536_),
    .B(_04537_));
 sg13g2_a22oi_1 _22123_ (.Y(_04539_),
    .B1(net99),
    .B2(net148),
    .A2(net117),
    .A1(net159));
 sg13g2_a21oi_1 _22124_ (.A1(net195),
    .A2(net119),
    .Y(_04540_),
    .B1(net98));
 sg13g2_a221oi_1 _22125_ (.B2(_04540_),
    .C1(net903),
    .B1(_04539_),
    .A1(_03606_),
    .Y(_04541_),
    .A2(net100));
 sg13g2_nor3_1 _22126_ (.A(_04533_),
    .B(_04538_),
    .C(_04541_),
    .Y(_04542_));
 sg13g2_a21o_1 _22127_ (.A2(_04508_),
    .A1(_03606_),
    .B1(net262),
    .X(_04543_));
 sg13g2_o21ai_1 _22128_ (.B1(_04543_),
    .Y(_04544_),
    .A1(_03606_),
    .A2(_04508_));
 sg13g2_and2_1 _22129_ (.A(_03715_),
    .B(_04534_),
    .X(_04545_));
 sg13g2_xnor2_1 _22130_ (.Y(_04546_),
    .A(_04544_),
    .B(_04545_));
 sg13g2_nor2_1 _22131_ (.A(_11064_),
    .B(_03606_),
    .Y(_04547_));
 sg13g2_o21ai_1 _22132_ (.B1(_03718_),
    .Y(_04548_),
    .A1(_04547_),
    .A2(_04511_));
 sg13g2_xnor2_1 _22133_ (.Y(_04549_),
    .A(_04545_),
    .B(_04548_));
 sg13g2_a22oi_1 _22134_ (.Y(_04550_),
    .B1(_04549_),
    .B2(_04118_),
    .A2(_04546_),
    .A1(net1073));
 sg13g2_nor2_1 _22135_ (.A(_04296_),
    .B(\cpu.ex.c_mult[4] ),
    .Y(_04551_));
 sg13g2_a21o_1 _22136_ (.A2(_04550_),
    .A1(_04542_),
    .B1(_04551_),
    .X(_04552_));
 sg13g2_a21o_1 _22137_ (.A2(_04230_),
    .A1(net84),
    .B1(_04226_),
    .X(_04553_));
 sg13g2_nor2_1 _22138_ (.A(net1150),
    .B(_04230_),
    .Y(_04554_));
 sg13g2_nor4_1 _22139_ (.A(net1092),
    .B(_08456_),
    .C(net795),
    .D(_11941_),
    .Y(_04555_));
 sg13g2_a221oi_1 _22140_ (.B2(net84),
    .C1(_04555_),
    .B1(_04554_),
    .A1(net1150),
    .Y(_04556_),
    .A2(_04553_));
 sg13g2_o21ai_1 _22141_ (.B1(_04556_),
    .Y(_00992_),
    .A1(net76),
    .A2(_04552_));
 sg13g2_xnor2_1 _22142_ (.Y(_04557_),
    .A(net225),
    .B(net182));
 sg13g2_xnor2_1 _22143_ (.Y(_04558_),
    .A(_03613_),
    .B(_04557_));
 sg13g2_a22oi_1 _22144_ (.Y(_04559_),
    .B1(_04162_),
    .B2(net125),
    .A2(net118),
    .A1(_03685_));
 sg13g2_a21oi_1 _22145_ (.A1(_03634_),
    .A2(net99),
    .Y(_04560_),
    .B1(_04351_));
 sg13g2_a22oi_1 _22146_ (.Y(_04561_),
    .B1(net116),
    .B2(net154),
    .A2(_04139_),
    .A1(_03699_));
 sg13g2_a21oi_1 _22147_ (.A1(_04195_),
    .A2(_04165_),
    .Y(_04562_),
    .B1(_04439_));
 sg13g2_o21ai_1 _22148_ (.B1(_08295_),
    .Y(_04563_),
    .A1(_04522_),
    .A2(_04525_));
 sg13g2_and3_1 _22149_ (.X(_04564_),
    .A(_04561_),
    .B(_04562_),
    .C(_04563_));
 sg13g2_nand4_1 _22150_ (.B(_04559_),
    .C(_04560_),
    .A(_04275_),
    .Y(_04565_),
    .D(_04564_));
 sg13g2_a21oi_1 _22151_ (.A1(_03584_),
    .A2(net100),
    .Y(_04566_),
    .B1(net847));
 sg13g2_xnor2_1 _22152_ (.Y(_04567_),
    .A(_04249_),
    .B(_04557_));
 sg13g2_nand2_1 _22153_ (.Y(_04568_),
    .A(net212),
    .B(net117));
 sg13g2_a221oi_1 _22154_ (.B2(_03587_),
    .C1(net124),
    .B1(net119),
    .A1(net181),
    .Y(_04569_),
    .A2(net179));
 sg13g2_nand3_1 _22155_ (.B(_04568_),
    .C(_04569_),
    .A(_04184_),
    .Y(_04570_));
 sg13g2_a21oi_1 _22156_ (.A1(_10603_),
    .A2(_04131_),
    .Y(_04571_),
    .B1(net903));
 sg13g2_a221oi_1 _22157_ (.B2(_04571_),
    .C1(net188),
    .B1(_04570_),
    .A1(net1148),
    .Y(_04572_),
    .A2(_11458_));
 sg13g2_nand3_1 _22158_ (.B(_11126_),
    .C(net152),
    .A(net1147),
    .Y(_04573_));
 sg13g2_o21ai_1 _22159_ (.B1(_09195_),
    .Y(_04574_),
    .A1(_11673_),
    .A2(net182));
 sg13g2_nand3b_1 _22160_ (.B(_04573_),
    .C(_04574_),
    .Y(_04575_),
    .A_N(net1134));
 sg13g2_o21ai_1 _22161_ (.B1(_04575_),
    .Y(_04576_),
    .A1(_11126_),
    .A2(net152));
 sg13g2_nand2_1 _22162_ (.Y(_04577_),
    .A(_04572_),
    .B(_04576_));
 sg13g2_a221oi_1 _22163_ (.B2(_04118_),
    .C1(_04577_),
    .B1(_04567_),
    .A1(_04565_),
    .Y(_04578_),
    .A2(_04566_));
 sg13g2_o21ai_1 _22164_ (.B1(_04578_),
    .Y(_04579_),
    .A1(net848),
    .A2(_04558_));
 sg13g2_o21ai_1 _22165_ (.B1(_04579_),
    .Y(_04580_),
    .A1(net178),
    .A2(\cpu.ex.c_mult[5] ));
 sg13g2_buf_1 _22166_ (.A(_08815_),
    .X(_04581_));
 sg13g2_xnor2_1 _22167_ (.Y(_04582_),
    .A(_00298_),
    .B(_04231_));
 sg13g2_a22oi_1 _22168_ (.Y(_04583_),
    .B1(_04582_),
    .B2(net75),
    .A2(net33),
    .A1(net987));
 sg13g2_o21ai_1 _22169_ (.B1(_04583_),
    .Y(_00993_),
    .A1(net76),
    .A2(_04580_));
 sg13g2_nor2_1 _22170_ (.A(net182),
    .B(_04249_),
    .Y(_04584_));
 sg13g2_a21oi_1 _22171_ (.A1(net182),
    .A2(_04249_),
    .Y(_04585_),
    .B1(_11673_));
 sg13g2_nor2_1 _22172_ (.A(_04584_),
    .B(_04585_),
    .Y(_04586_));
 sg13g2_nand2_1 _22173_ (.Y(_04587_),
    .A(_03729_),
    .B(_03732_));
 sg13g2_xor2_1 _22174_ (.B(_04587_),
    .A(_04586_),
    .X(_04588_));
 sg13g2_a21oi_1 _22175_ (.A1(_03613_),
    .A2(_03614_),
    .Y(_04589_),
    .B1(_03615_));
 sg13g2_xor2_1 _22176_ (.B(_04587_),
    .A(_04589_),
    .X(_04590_));
 sg13g2_a22oi_1 _22177_ (.Y(_04591_),
    .B1(_04164_),
    .B2(_03766_),
    .A2(net180),
    .A1(_03684_));
 sg13g2_a22oi_1 _22178_ (.Y(_04592_),
    .B1(_04186_),
    .B2(net164),
    .A2(_04183_),
    .A1(net165));
 sg13g2_a21oi_1 _22179_ (.A1(_03658_),
    .A2(_04148_),
    .Y(_04593_),
    .B1(net158));
 sg13g2_and3_1 _22180_ (.X(_04594_),
    .A(_04591_),
    .B(_04592_),
    .C(_04593_));
 sg13g2_a221oi_1 _22181_ (.B2(net163),
    .C1(_04315_),
    .B1(_04142_),
    .A1(net153),
    .Y(_04595_),
    .A2(net151));
 sg13g2_a21oi_1 _22182_ (.A1(_04594_),
    .A2(_04595_),
    .Y(_04596_),
    .B1(net847));
 sg13g2_o21ai_1 _22183_ (.B1(_03766_),
    .Y(_04597_),
    .A1(_04161_),
    .A2(_04173_));
 sg13g2_nand2b_1 _22184_ (.Y(_04598_),
    .B(_04597_),
    .A_N(_04522_));
 sg13g2_and2_1 _22185_ (.A(net1097),
    .B(_04598_),
    .X(_04599_));
 sg13g2_nand2_1 _22186_ (.Y(_04600_),
    .A(_03624_),
    .B(net98));
 sg13g2_o21ai_1 _22187_ (.B1(_04600_),
    .Y(_04601_),
    .A1(_04596_),
    .A2(_04599_));
 sg13g2_nand2_1 _22188_ (.Y(_04602_),
    .A(_04320_),
    .B(net156));
 sg13g2_a22oi_1 _22189_ (.Y(_04603_),
    .B1(net119),
    .B2(net150),
    .A2(net117),
    .A1(net148));
 sg13g2_a221oi_1 _22190_ (.B2(net181),
    .C1(net124),
    .B1(net116),
    .A1(net211),
    .Y(_04604_),
    .A2(net121));
 sg13g2_nand3_1 _22191_ (.B(_04603_),
    .C(_04604_),
    .A(_04602_),
    .Y(_04605_));
 sg13g2_a21oi_1 _22192_ (.A1(net182),
    .A2(net98),
    .Y(_04606_),
    .B1(net903));
 sg13g2_nand2_1 _22193_ (.Y(_04607_),
    .A(_04605_),
    .B(_04606_));
 sg13g2_a21oi_1 _22194_ (.A1(_09037_),
    .A2(_03678_),
    .Y(_04608_),
    .B1(net188));
 sg13g2_mux2_1 _22195_ (.A0(net1147),
    .A1(_09195_),
    .S(_03729_),
    .X(_04609_));
 sg13g2_o21ai_1 _22196_ (.B1(_03732_),
    .Y(_04610_),
    .A1(net1134),
    .A2(_04609_));
 sg13g2_nand4_1 _22197_ (.B(_04607_),
    .C(_04608_),
    .A(_04601_),
    .Y(_04611_),
    .D(_04610_));
 sg13g2_a221oi_1 _22198_ (.B2(net1073),
    .C1(_04611_),
    .B1(_04590_),
    .A1(_04118_),
    .Y(_04612_),
    .A2(_04588_));
 sg13g2_a21o_1 _22199_ (.A2(_11704_),
    .A1(net160),
    .B1(_04612_),
    .X(_04613_));
 sg13g2_buf_1 _22200_ (.A(_08863_),
    .X(_04614_));
 sg13g2_nand2_1 _22201_ (.Y(_04615_),
    .A(_08815_),
    .B(_04231_));
 sg13g2_xor2_1 _22202_ (.B(_04615_),
    .A(_10612_),
    .X(_04616_));
 sg13g2_a22oi_1 _22203_ (.Y(_04617_),
    .B1(_04616_),
    .B2(net75),
    .A2(net33),
    .A1(net986));
 sg13g2_o21ai_1 _22204_ (.B1(_04617_),
    .Y(_00994_),
    .A1(net76),
    .A2(_04613_));
 sg13g2_or2_1 _22205_ (.X(_04618_),
    .B(\cpu.ex.c_mult[7] ),
    .A(_04297_));
 sg13g2_nor2_1 _22206_ (.A(_03617_),
    .B(_03627_),
    .Y(_04619_));
 sg13g2_xnor2_1 _22207_ (.Y(_04620_),
    .A(_04619_),
    .B(_04255_));
 sg13g2_nand2_1 _22208_ (.Y(_04621_),
    .A(_03632_),
    .B(net98));
 sg13g2_a21oi_1 _22209_ (.A1(net163),
    .A2(net180),
    .Y(_04622_),
    .B1(net158));
 sg13g2_a22oi_1 _22210_ (.Y(_04623_),
    .B1(_04186_),
    .B2(_03685_),
    .A2(net179),
    .A1(_03672_));
 sg13g2_a22oi_1 _22211_ (.Y(_04624_),
    .B1(_04199_),
    .B2(_03641_),
    .A2(_04178_),
    .A1(net154));
 sg13g2_nand4_1 _22212_ (.B(_04622_),
    .C(_04623_),
    .A(_04278_),
    .Y(_04625_),
    .D(_04624_));
 sg13g2_a21oi_1 _22213_ (.A1(_03767_),
    .A2(_04276_),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_a21oi_1 _22214_ (.A1(net1097),
    .A2(_04625_),
    .Y(_04627_),
    .B1(net1135));
 sg13g2_o21ai_1 _22215_ (.B1(_04193_),
    .Y(_04628_),
    .A1(net262),
    .A2(_04189_));
 sg13g2_o21ai_1 _22216_ (.B1(_04628_),
    .Y(_04629_),
    .A1(_04626_),
    .A2(_04627_));
 sg13g2_mux2_1 _22217_ (.A0(net1075),
    .A1(net1074),
    .S(_03727_),
    .X(_04630_));
 sg13g2_o21ai_1 _22218_ (.B1(_03736_),
    .Y(_04631_),
    .A1(net1059),
    .A2(_04630_));
 sg13g2_nand2_1 _22219_ (.Y(_04632_),
    .A(net150),
    .B(net151));
 sg13g2_a22oi_1 _22220_ (.Y(_04633_),
    .B1(net116),
    .B2(net212),
    .A2(net156),
    .A1(_03587_));
 sg13g2_a221oi_1 _22221_ (.B2(net211),
    .C1(net158),
    .B1(_04199_),
    .A1(net181),
    .Y(_04634_),
    .A2(net180));
 sg13g2_nand4_1 _22222_ (.B(_04632_),
    .C(_04633_),
    .A(_04501_),
    .Y(_04635_),
    .D(_04634_));
 sg13g2_a21oi_1 _22223_ (.A1(_03584_),
    .A2(net124),
    .Y(_04636_),
    .B1(net903));
 sg13g2_a221oi_1 _22224_ (.B2(_04636_),
    .C1(net188),
    .B1(_04635_),
    .A1(net1148),
    .Y(_04637_),
    .A2(_11562_));
 sg13g2_nand2_1 _22225_ (.Y(_04638_),
    .A(_04631_),
    .B(_04637_));
 sg13g2_a221oi_1 _22226_ (.B2(_04629_),
    .C1(_04638_),
    .B1(_04621_),
    .A1(_04118_),
    .Y(_04639_),
    .A2(_04409_));
 sg13g2_o21ai_1 _22227_ (.B1(_04639_),
    .Y(_04640_),
    .A1(net848),
    .A2(_04620_));
 sg13g2_nand2_1 _22228_ (.Y(_04641_),
    .A(_04618_),
    .B(_04640_));
 sg13g2_xor2_1 _22229_ (.B(_04232_),
    .A(_10714_),
    .X(_04642_));
 sg13g2_a22oi_1 _22230_ (.Y(_04643_),
    .B1(_04642_),
    .B2(_04238_),
    .A2(_04227_),
    .A1(\cpu.ex.pc[7] ));
 sg13g2_o21ai_1 _22231_ (.B1(_04643_),
    .Y(_00995_),
    .A1(_04098_),
    .A2(_04641_));
 sg13g2_xnor2_1 _22232_ (.Y(_04644_),
    .A(_11383_),
    .B(_03632_));
 sg13g2_inv_1 _22233_ (.Y(_04645_),
    .A(_03625_));
 sg13g2_a21oi_1 _22234_ (.A1(_04645_),
    .A2(_04619_),
    .Y(_04646_),
    .B1(_03635_));
 sg13g2_xnor2_1 _22235_ (.Y(_04647_),
    .A(_04644_),
    .B(_04646_));
 sg13g2_nor2_1 _22236_ (.A(_03579_),
    .B(_04355_),
    .Y(_04648_));
 sg13g2_a221oi_1 _22237_ (.B2(_03699_),
    .C1(_04648_),
    .B1(_04318_),
    .A1(_03767_),
    .Y(_04649_),
    .A2(_04139_));
 sg13g2_a22oi_1 _22238_ (.Y(_04650_),
    .B1(_04390_),
    .B2(net120),
    .A2(_04313_),
    .A1(net153));
 sg13g2_nand4_1 _22239_ (.B(_04628_),
    .C(_04649_),
    .A(_04398_),
    .Y(_04651_),
    .D(_04650_));
 sg13g2_a21oi_1 _22240_ (.A1(net161),
    .A2(net100),
    .Y(_04652_),
    .B1(net847));
 sg13g2_nand2_1 _22241_ (.Y(_04653_),
    .A(net211),
    .B(net151));
 sg13g2_a221oi_1 _22242_ (.B2(net148),
    .C1(_04456_),
    .B1(net149),
    .A1(_04101_),
    .Y(_04654_),
    .A2(_04142_));
 sg13g2_nand2_1 _22243_ (.Y(_04655_),
    .A(_03706_),
    .B(net157));
 sg13g2_a21oi_1 _22244_ (.A1(net150),
    .A2(net156),
    .Y(_04656_),
    .B1(_04528_));
 sg13g2_nand4_1 _22245_ (.B(_04654_),
    .C(_04655_),
    .A(_04653_),
    .Y(_04657_),
    .D(_04656_));
 sg13g2_nand3_1 _22246_ (.B(_04600_),
    .C(_04657_),
    .A(_09924_),
    .Y(_04658_));
 sg13g2_nand3_1 _22247_ (.B(net205),
    .C(net126),
    .A(net1147),
    .Y(_04659_));
 sg13g2_o21ai_1 _22248_ (.B1(_09195_),
    .Y(_04660_),
    .A1(_11383_),
    .A2(_03632_));
 sg13g2_nand3b_1 _22249_ (.B(_04659_),
    .C(_04660_),
    .Y(_04661_),
    .A_N(net1134));
 sg13g2_o21ai_1 _22250_ (.B1(_04661_),
    .Y(_04662_),
    .A1(_11745_),
    .A2(net126));
 sg13g2_nand2_1 _22251_ (.Y(_04663_),
    .A(_04658_),
    .B(_04662_));
 sg13g2_a221oi_1 _22252_ (.B2(_04652_),
    .C1(_04663_),
    .B1(_04651_),
    .A1(net1076),
    .Y(_04664_),
    .A2(_11589_));
 sg13g2_and3_1 _22253_ (.X(_04665_),
    .A(_04115_),
    .B(_04259_),
    .C(_04664_));
 sg13g2_o21ai_1 _22254_ (.B1(_04665_),
    .Y(_04666_),
    .A1(net848),
    .A2(_04647_));
 sg13g2_xor2_1 _22255_ (.B(_04644_),
    .A(_03738_),
    .X(_04667_));
 sg13g2_a21oi_1 _22256_ (.A1(_04293_),
    .A2(_04667_),
    .Y(_04668_),
    .B1(net160));
 sg13g2_a22oi_1 _22257_ (.Y(_04669_),
    .B1(_04666_),
    .B2(_04668_),
    .A2(\cpu.ex.c_mult[8] ),
    .A1(net160));
 sg13g2_xnor2_1 _22258_ (.Y(_04670_),
    .A(_03618_),
    .B(_04234_));
 sg13g2_a22oi_1 _22259_ (.Y(_04671_),
    .B1(_04670_),
    .B2(net75),
    .A2(net33),
    .A1(_08850_));
 sg13g2_o21ai_1 _22260_ (.B1(_04671_),
    .Y(_00996_),
    .A1(_04097_),
    .A2(_04669_));
 sg13g2_and3_1 _22261_ (.X(_04672_),
    .A(net160),
    .B(_11765_),
    .C(_11766_));
 sg13g2_nor2_1 _22262_ (.A(_03617_),
    .B(_03629_),
    .Y(_04673_));
 sg13g2_nor2_1 _22263_ (.A(_04673_),
    .B(_03638_),
    .Y(_04674_));
 sg13g2_xnor2_1 _22264_ (.Y(_04675_),
    .A(net187),
    .B(net161));
 sg13g2_xor2_1 _22265_ (.B(_04675_),
    .A(_04674_),
    .X(_04676_));
 sg13g2_nand2_1 _22266_ (.Y(_04677_),
    .A(_03739_),
    .B(_03741_));
 sg13g2_xnor2_1 _22267_ (.Y(_04678_),
    .A(_04677_),
    .B(_04675_));
 sg13g2_a21oi_1 _22268_ (.A1(net128),
    .A2(_04318_),
    .Y(_04679_),
    .B1(net98));
 sg13g2_a221oi_1 _22269_ (.B2(net127),
    .C1(_04353_),
    .B1(_04200_),
    .A1(_04195_),
    .Y(_04680_),
    .A2(_04149_));
 sg13g2_nand2_1 _22270_ (.Y(_04681_),
    .A(_04679_),
    .B(_04680_));
 sg13g2_or3_1 _22271_ (.A(net262),
    .B(_04189_),
    .C(net180),
    .X(_04682_));
 sg13g2_a21oi_1 _22272_ (.A1(_08296_),
    .A2(_04682_),
    .Y(_04683_),
    .B1(_04390_));
 sg13g2_nor2_1 _22273_ (.A(_03576_),
    .B(_04683_),
    .Y(_04684_));
 sg13g2_a21oi_1 _22274_ (.A1(_03645_),
    .A2(net100),
    .Y(_04685_),
    .B1(net847));
 sg13g2_o21ai_1 _22275_ (.B1(_04685_),
    .Y(_04686_),
    .A1(_04681_),
    .A2(_04684_));
 sg13g2_o21ai_1 _22276_ (.B1(_04179_),
    .Y(_04687_),
    .A1(_03624_),
    .A2(_04352_));
 sg13g2_a221oi_1 _22277_ (.B2(_04320_),
    .C1(_04687_),
    .B1(net118),
    .A1(_04205_),
    .Y(_04688_),
    .A2(net157));
 sg13g2_nand2_1 _22278_ (.Y(_04689_),
    .A(net150),
    .B(net116));
 sg13g2_a22oi_1 _22279_ (.Y(_04690_),
    .B1(net122),
    .B2(net159),
    .A2(net156),
    .A1(net211));
 sg13g2_nand4_1 _22280_ (.B(_04688_),
    .C(_04689_),
    .A(_04504_),
    .Y(_04691_),
    .D(_04690_));
 sg13g2_nand3_1 _22281_ (.B(_04621_),
    .C(_04691_),
    .A(_09924_),
    .Y(_04692_));
 sg13g2_nand2_1 _22282_ (.Y(_04693_),
    .A(_11744_),
    .B(net161));
 sg13g2_nand3_1 _22283_ (.B(_11570_),
    .C(net162),
    .A(net1075),
    .Y(_04694_));
 sg13g2_o21ai_1 _22284_ (.B1(net1074),
    .Y(_04695_),
    .A1(_11744_),
    .A2(net161));
 sg13g2_nand3b_1 _22285_ (.B(_04694_),
    .C(_04695_),
    .Y(_04696_),
    .A_N(net1059));
 sg13g2_a22oi_1 _22286_ (.Y(_04697_),
    .B1(_04693_),
    .B2(_04696_),
    .A2(_11249_),
    .A1(net1076));
 sg13g2_nand4_1 _22287_ (.B(_04686_),
    .C(_04692_),
    .A(_04310_),
    .Y(_04698_),
    .D(_04697_));
 sg13g2_a221oi_1 _22288_ (.B2(_04293_),
    .C1(_04698_),
    .B1(_04678_),
    .A1(net1073),
    .Y(_04699_),
    .A2(_04676_));
 sg13g2_nand2b_1 _22289_ (.Y(_04700_),
    .B(_04217_),
    .A_N(_04699_));
 sg13g2_xnor2_1 _22290_ (.Y(_04701_),
    .A(_00294_),
    .B(_04235_));
 sg13g2_a22oi_1 _22291_ (.Y(_04702_),
    .B1(_04701_),
    .B2(net75),
    .A2(_04226_),
    .A1(_08824_));
 sg13g2_o21ai_1 _22292_ (.B1(_04702_),
    .Y(_00997_),
    .A1(_04672_),
    .A2(_04700_));
 sg13g2_nand2_1 _22293_ (.Y(_04703_),
    .A(net160),
    .B(\cpu.ex.c_mult[10] ));
 sg13g2_a22oi_1 _22294_ (.Y(_04704_),
    .B1(_04182_),
    .B2(_03671_),
    .A2(net179),
    .A1(_03766_));
 sg13g2_nand2_1 _22295_ (.Y(_04705_),
    .A(_03684_),
    .B(_04199_));
 sg13g2_a21oi_1 _22296_ (.A1(net163),
    .A2(_04177_),
    .Y(_04706_),
    .B1(_04130_));
 sg13g2_nand3_1 _22297_ (.B(_04705_),
    .C(_04706_),
    .A(_04704_),
    .Y(_04707_));
 sg13g2_o21ai_1 _22298_ (.B1(_03766_),
    .Y(_04708_),
    .A1(net149),
    .A2(_04682_));
 sg13g2_nand2b_1 _22299_ (.Y(_04709_),
    .B(_04708_),
    .A_N(_04707_));
 sg13g2_a22oi_1 _22300_ (.Y(_04710_),
    .B1(_04709_),
    .B2(_08295_),
    .A2(_04707_),
    .A1(_09890_));
 sg13g2_nand2_1 _22301_ (.Y(_04711_),
    .A(net155),
    .B(net151));
 sg13g2_and2_1 _22302_ (.A(_03587_),
    .B(_04142_),
    .X(_04712_));
 sg13g2_a221oi_1 _22303_ (.B2(_10679_),
    .C1(_04712_),
    .B1(net149),
    .A1(net181),
    .Y(_04713_),
    .A2(_04161_));
 sg13g2_a221oi_1 _22304_ (.B2(_10566_),
    .C1(_04523_),
    .B1(net179),
    .A1(_03610_),
    .Y(_04714_),
    .A2(net180));
 sg13g2_a22oi_1 _22305_ (.Y(_04715_),
    .B1(net121),
    .B2(_03621_),
    .A2(_04164_),
    .A1(_03706_));
 sg13g2_nand4_1 _22306_ (.B(_04713_),
    .C(_04714_),
    .A(_04711_),
    .Y(_04716_),
    .D(_04715_));
 sg13g2_a21oi_1 _22307_ (.A1(_03754_),
    .A2(net158),
    .Y(_04717_),
    .B1(_09925_));
 sg13g2_mux2_1 _22308_ (.A0(net1147),
    .A1(_09195_),
    .S(_03643_),
    .X(_04718_));
 sg13g2_or2_1 _22309_ (.X(_04719_),
    .B(_04718_),
    .A(_09921_));
 sg13g2_and2_1 _22310_ (.A(net1148),
    .B(_11638_),
    .X(_04720_));
 sg13g2_a221oi_1 _22311_ (.B2(_03646_),
    .C1(_04720_),
    .B1(_04719_),
    .A1(_04716_),
    .Y(_04721_),
    .A2(_04717_));
 sg13g2_o21ai_1 _22312_ (.B1(_04721_),
    .Y(_04722_),
    .A1(_04324_),
    .A2(_04710_));
 sg13g2_a221oi_1 _22313_ (.B2(_09916_),
    .C1(_04722_),
    .B1(_04409_),
    .A1(_04112_),
    .Y(_04723_),
    .A2(_04113_));
 sg13g2_buf_1 _22314_ (.A(_04723_),
    .X(_04724_));
 sg13g2_nand3_1 _22315_ (.B(_04287_),
    .C(_04724_),
    .A(_03648_),
    .Y(_04725_));
 sg13g2_nand2_1 _22316_ (.Y(_04726_),
    .A(_03643_),
    .B(_03646_));
 sg13g2_nand3_1 _22317_ (.B(_04244_),
    .C(_04724_),
    .A(_04726_),
    .Y(_04727_));
 sg13g2_nor2_1 _22318_ (.A(_04726_),
    .B(net509),
    .Y(_04728_));
 sg13g2_nor3_1 _22319_ (.A(_03648_),
    .B(_03757_),
    .C(net509),
    .Y(_04729_));
 sg13g2_a221oi_1 _22320_ (.B2(_03757_),
    .C1(_04729_),
    .B1(_04728_),
    .A1(net848),
    .Y(_04730_),
    .A2(_04724_));
 sg13g2_nand4_1 _22321_ (.B(_04725_),
    .C(_04727_),
    .A(net178),
    .Y(_04731_),
    .D(_04730_));
 sg13g2_a21oi_1 _22322_ (.A1(_04703_),
    .A2(_04731_),
    .Y(_04732_),
    .B1(_04097_));
 sg13g2_buf_1 _22323_ (.A(_08841_),
    .X(_04733_));
 sg13g2_nand2_1 _22324_ (.Y(_04734_),
    .A(_08824_),
    .B(_04235_));
 sg13g2_xnor2_1 _22325_ (.Y(_04735_),
    .A(_10881_),
    .B(_04734_));
 sg13g2_a22oi_1 _22326_ (.Y(_04736_),
    .B1(_04735_),
    .B2(net75),
    .A2(net33),
    .A1(net985));
 sg13g2_nand2b_1 _22327_ (.Y(_00998_),
    .B(_04736_),
    .A_N(_04732_));
 sg13g2_mux2_1 _22328_ (.A0(_10266_),
    .A1(\cpu.dec.r_set_cc ),
    .S(_03571_),
    .X(_01001_));
 sg13g2_buf_1 _22329_ (.A(_00258_),
    .X(_04737_));
 sg13g2_nor4_1 _22330_ (.A(net1130),
    .B(_10260_),
    .C(_04737_),
    .D(_03520_),
    .Y(_04738_));
 sg13g2_buf_2 _22331_ (.A(_04738_),
    .X(_04739_));
 sg13g2_buf_1 _22332_ (.A(_04739_),
    .X(_04740_));
 sg13g2_mux2_1 _22333_ (.A0(_10698_),
    .A1(net461),
    .S(net508),
    .X(_01002_));
 sg13g2_mux2_1 _22334_ (.A0(_10907_),
    .A1(net852),
    .S(net508),
    .X(_01003_));
 sg13g2_mux2_1 _22335_ (.A0(_10854_),
    .A1(net591),
    .S(net508),
    .X(_01004_));
 sg13g2_mux2_1 _22336_ (.A0(_10783_),
    .A1(net656),
    .S(net508),
    .X(_01005_));
 sg13g2_mux2_1 _22337_ (.A0(_10861_),
    .A1(net512),
    .S(net508),
    .X(_01006_));
 sg13g2_mux2_1 _22338_ (.A0(_10322_),
    .A1(net733),
    .S(_04740_),
    .X(_01007_));
 sg13g2_mux2_1 _22339_ (.A0(_10443_),
    .A1(net519),
    .S(net508),
    .X(_01008_));
 sg13g2_mux2_1 _22340_ (.A0(_10515_),
    .A1(net518),
    .S(net508),
    .X(_01009_));
 sg13g2_mux2_1 _22341_ (.A0(_10582_),
    .A1(_03536_),
    .S(_04739_),
    .X(_01010_));
 sg13g2_mux2_1 _22342_ (.A0(_10547_),
    .A1(net514),
    .S(_04739_),
    .X(_01011_));
 sg13g2_nand2_1 _22343_ (.Y(_04741_),
    .A(net857),
    .B(_04739_));
 sg13g2_o21ai_1 _22344_ (.B1(_04741_),
    .Y(_01012_),
    .A1(_11198_),
    .A2(net508));
 sg13g2_buf_1 _22345_ (.A(net862),
    .X(_04742_));
 sg13g2_mux2_1 _22346_ (.A0(_10725_),
    .A1(_04742_),
    .S(_04739_),
    .X(_01013_));
 sg13g2_buf_1 _22347_ (.A(net861),
    .X(_04743_));
 sg13g2_mux2_1 _22348_ (.A0(_10802_),
    .A1(_04743_),
    .S(_04739_),
    .X(_01014_));
 sg13g2_nand2_1 _22349_ (.Y(_04744_),
    .A(net993),
    .B(_04739_));
 sg13g2_o21ai_1 _22350_ (.B1(_04744_),
    .Y(_01015_),
    .A1(_10822_),
    .A2(_04740_));
 sg13g2_mux2_1 _22351_ (.A0(_10891_),
    .A1(net851),
    .S(_04739_),
    .X(_01016_));
 sg13g2_or2_1 _22352_ (.X(_04745_),
    .B(_03520_),
    .A(_10263_));
 sg13g2_buf_2 _22353_ (.A(_04745_),
    .X(_04746_));
 sg13g2_buf_1 _22354_ (.A(_04746_),
    .X(_04747_));
 sg13g2_nor2b_1 _22355_ (.A(_04737_),
    .B_N(net932),
    .Y(_04748_));
 sg13g2_nand2_1 _22356_ (.Y(_04749_),
    .A(_03518_),
    .B(_04748_));
 sg13g2_and2_1 _22357_ (.A(net932),
    .B(_10260_),
    .X(_04750_));
 sg13g2_a21oi_1 _22358_ (.A1(_10261_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04751_),
    .B1(_04750_));
 sg13g2_or4_1 _22359_ (.A(net1130),
    .B(_04737_),
    .C(_03520_),
    .D(_04751_),
    .X(_04752_));
 sg13g2_buf_2 _22360_ (.A(_04752_),
    .X(_04753_));
 sg13g2_buf_1 _22361_ (.A(_04753_),
    .X(_04754_));
 sg13g2_nand2_1 _22362_ (.Y(_04755_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net457));
 sg13g2_o21ai_1 _22363_ (.B1(_04755_),
    .Y(_01017_),
    .A1(net507),
    .A2(_04749_));
 sg13g2_buf_1 _22364_ (.A(_04746_),
    .X(_04756_));
 sg13g2_mux2_1 _22365_ (.A0(_10903_),
    .A1(_10891_),
    .S(_04756_),
    .X(_04757_));
 sg13g2_mux2_1 _22366_ (.A0(_04757_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net457),
    .X(_01018_));
 sg13g2_buf_1 _22367_ (.A(_04753_),
    .X(_04758_));
 sg13g2_mux2_1 _22368_ (.A0(_10925_),
    .A1(_10907_),
    .S(_04746_),
    .X(_04759_));
 sg13g2_nor2_1 _22369_ (.A(_04753_),
    .B(_04759_),
    .Y(_04760_));
 sg13g2_a21oi_1 _22370_ (.A1(_10917_),
    .A2(net456),
    .Y(_01019_),
    .B1(_04760_));
 sg13g2_nor2_1 _22371_ (.A(_11946_),
    .B(net506),
    .Y(_04761_));
 sg13g2_a21oi_1 _22372_ (.A1(_10854_),
    .A2(_04747_),
    .Y(_04762_),
    .B1(_04761_));
 sg13g2_nand2_1 _22373_ (.Y(_04763_),
    .A(\cpu.ex.r_stmp[12] ),
    .B(net457));
 sg13g2_o21ai_1 _22374_ (.B1(_04763_),
    .Y(_01020_),
    .A1(_04758_),
    .A2(_04762_));
 sg13g2_nor2_1 _22375_ (.A(_11444_),
    .B(net506),
    .Y(_04764_));
 sg13g2_a21oi_1 _22376_ (.A1(_10783_),
    .A2(net507),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nand2_1 _22377_ (.Y(_04766_),
    .A(\cpu.ex.r_stmp[13] ),
    .B(net457));
 sg13g2_o21ai_1 _22378_ (.B1(_04766_),
    .Y(_01021_),
    .A1(_04758_),
    .A2(_04765_));
 sg13g2_mux2_1 _22379_ (.A0(net598),
    .A1(_10861_),
    .S(net506),
    .X(_04767_));
 sg13g2_mux2_1 _22380_ (.A0(_04767_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net457),
    .X(_01022_));
 sg13g2_nor2_1 _22381_ (.A(_10749_),
    .B(net506),
    .Y(_04768_));
 sg13g2_a21oi_1 _22382_ (.A1(_10322_),
    .A2(_04747_),
    .Y(_04769_),
    .B1(_04768_));
 sg13g2_nand2_1 _22383_ (.Y(_04770_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(net457));
 sg13g2_o21ai_1 _22384_ (.B1(_04770_),
    .Y(_01023_),
    .A1(net456),
    .A2(_04769_));
 sg13g2_nor2_1 _22385_ (.A(_10204_),
    .B(net506),
    .Y(_04771_));
 sg13g2_a21oi_1 _22386_ (.A1(_10698_),
    .A2(net507),
    .Y(_04772_),
    .B1(_04771_));
 sg13g2_nand2_1 _22387_ (.Y(_04773_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net457));
 sg13g2_o21ai_1 _22388_ (.B1(_04773_),
    .Y(_01024_),
    .A1(net456),
    .A2(_04772_));
 sg13g2_nor2_1 _22389_ (.A(net654),
    .B(net506),
    .Y(_04774_));
 sg13g2_a21oi_1 _22390_ (.A1(_10443_),
    .A2(net507),
    .Y(_04775_),
    .B1(_04774_));
 sg13g2_nand2_1 _22391_ (.Y(_04776_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(_04753_));
 sg13g2_o21ai_1 _22392_ (.B1(_04776_),
    .Y(_01025_),
    .A1(net456),
    .A2(_04775_));
 sg13g2_nor2_1 _22393_ (.A(net796),
    .B(_04746_),
    .Y(_04777_));
 sg13g2_a21oi_1 _22394_ (.A1(_10515_),
    .A2(net507),
    .Y(_04778_),
    .B1(_04777_));
 sg13g2_nand2_1 _22395_ (.Y(_04779_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(_04753_));
 sg13g2_o21ai_1 _22396_ (.B1(_04779_),
    .Y(_01026_),
    .A1(net456),
    .A2(_04778_));
 sg13g2_nor2_1 _22397_ (.A(_03788_),
    .B(_04746_),
    .Y(_04780_));
 sg13g2_a21oi_1 _22398_ (.A1(_10582_),
    .A2(net507),
    .Y(_04781_),
    .B1(_04780_));
 sg13g2_nand2_1 _22399_ (.Y(_04782_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04753_));
 sg13g2_o21ai_1 _22400_ (.B1(_04782_),
    .Y(_01027_),
    .A1(net456),
    .A2(_04781_));
 sg13g2_nor2_1 _22401_ (.A(_12000_),
    .B(_04746_),
    .Y(_04783_));
 sg13g2_a21oi_1 _22402_ (.A1(_10547_),
    .A2(net507),
    .Y(_04784_),
    .B1(_04783_));
 sg13g2_nand2_1 _22403_ (.Y(_04785_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04753_));
 sg13g2_o21ai_1 _22404_ (.B1(_04785_),
    .Y(_01028_),
    .A1(net456),
    .A2(_04784_));
 sg13g2_nor2_1 _22405_ (.A(_03025_),
    .B(_04746_),
    .Y(_04786_));
 sg13g2_a21oi_1 _22406_ (.A1(\cpu.ex.r_sp[6] ),
    .A2(net507),
    .Y(_04787_),
    .B1(_04786_));
 sg13g2_nand2_1 _22407_ (.Y(_04788_),
    .A(\cpu.ex.r_stmp[6] ),
    .B(_04753_));
 sg13g2_o21ai_1 _22408_ (.B1(_04788_),
    .Y(_01029_),
    .A1(net456),
    .A2(_04787_));
 sg13g2_mux2_1 _22409_ (.A0(net1069),
    .A1(_10725_),
    .S(net506),
    .X(_04789_));
 sg13g2_mux2_1 _22410_ (.A0(_04789_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net457),
    .X(_01030_));
 sg13g2_mux2_1 _22411_ (.A0(net1070),
    .A1(_10802_),
    .S(net506),
    .X(_04790_));
 sg13g2_mux2_1 _22412_ (.A0(_04790_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(_04754_),
    .X(_01031_));
 sg13g2_mux2_1 _22413_ (.A0(_10819_),
    .A1(\cpu.ex.r_sp[9] ),
    .S(_04756_),
    .X(_04791_));
 sg13g2_mux2_1 _22414_ (.A0(_04791_),
    .A1(\cpu.ex.r_stmp[9] ),
    .S(_04754_),
    .X(_01032_));
 sg13g2_a21o_1 _22415_ (.A2(net340),
    .A1(_10246_),
    .B1(net178),
    .X(_04792_));
 sg13g2_nor2_1 _22416_ (.A(_11594_),
    .B(_04792_),
    .Y(_04793_));
 sg13g2_nor2_1 _22417_ (.A(net195),
    .B(net147),
    .Y(_04794_));
 sg13g2_nand2_1 _22418_ (.Y(_04795_),
    .A(_04205_),
    .B(net121));
 sg13g2_nand3_1 _22419_ (.B(_04393_),
    .C(_04795_),
    .A(_04317_),
    .Y(_04796_));
 sg13g2_nand2_1 _22420_ (.Y(_04797_),
    .A(_03705_),
    .B(_04142_));
 sg13g2_a22oi_1 _22421_ (.Y(_04798_),
    .B1(_04199_),
    .B2(net150),
    .A2(net179),
    .A1(_04176_));
 sg13g2_nand3_1 _22422_ (.B(_04797_),
    .C(_04798_),
    .A(_04653_),
    .Y(_04799_));
 sg13g2_nand2_1 _22423_ (.Y(_04800_),
    .A(net128),
    .B(_04197_));
 sg13g2_a22oi_1 _22424_ (.Y(_04801_),
    .B1(_04173_),
    .B2(net154),
    .A2(net122),
    .A1(_03743_));
 sg13g2_a22oi_1 _22425_ (.Y(_04802_),
    .B1(_04170_),
    .B2(_03681_),
    .A2(_04146_),
    .A1(_03672_));
 sg13g2_a22oi_1 _22426_ (.Y(_04803_),
    .B1(_04191_),
    .B2(_03766_),
    .A2(net123),
    .A1(_04166_));
 sg13g2_nand4_1 _22427_ (.B(_04801_),
    .C(_04802_),
    .A(_04800_),
    .Y(_04804_),
    .D(_04803_));
 sg13g2_nor3_1 _22428_ (.A(_04796_),
    .B(_04799_),
    .C(_04804_),
    .Y(_04805_));
 sg13g2_inv_1 _22429_ (.Y(_04806_),
    .A(_04805_));
 sg13g2_o21ai_1 _22430_ (.B1(_04805_),
    .Y(_04807_),
    .A1(net166),
    .A2(_11578_));
 sg13g2_a22oi_1 _22431_ (.Y(_04808_),
    .B1(_04807_),
    .B2(net1097),
    .A2(_04806_),
    .A1(net1135));
 sg13g2_nor2_1 _22432_ (.A(net1075),
    .B(net226),
    .Y(_04809_));
 sg13g2_nor2b_1 _22433_ (.A(_04112_),
    .B_N(_04113_),
    .Y(_04810_));
 sg13g2_a22oi_1 _22434_ (.Y(_04811_),
    .B1(_04810_),
    .B2(_11093_),
    .A2(_04809_),
    .A1(net159));
 sg13g2_or2_1 _22435_ (.X(_04812_),
    .B(_04811_),
    .A(net1059));
 sg13g2_nor2b_1 _22436_ (.A(net1059),
    .B_N(_04810_),
    .Y(_04813_));
 sg13g2_o21ai_1 _22437_ (.B1(_04103_),
    .Y(_04814_),
    .A1(_11093_),
    .A2(_04813_));
 sg13g2_a221oi_1 _22438_ (.B2(_04814_),
    .C1(_04099_),
    .B1(_04812_),
    .A1(net1076),
    .Y(_04815_),
    .A2(_11745_));
 sg13g2_o21ai_1 _22439_ (.B1(_04815_),
    .Y(_04816_),
    .A1(_04794_),
    .A2(_04808_));
 sg13g2_nand2_1 _22440_ (.Y(_04817_),
    .A(_11601_),
    .B(net196));
 sg13g2_nor2_1 _22441_ (.A(_03568_),
    .B(_04817_),
    .Y(_04818_));
 sg13g2_nand2_1 _22442_ (.Y(_04819_),
    .A(_04816_),
    .B(_04818_));
 sg13g2_buf_1 _22443_ (.A(_03568_),
    .X(_04820_));
 sg13g2_buf_1 _22444_ (.A(_03570_),
    .X(_04821_));
 sg13g2_buf_1 _22445_ (.A(net1025),
    .X(_04822_));
 sg13g2_nand2_1 _22446_ (.Y(_04823_),
    .A(_10619_),
    .B(_09231_));
 sg13g2_buf_2 _22447_ (.A(_04823_),
    .X(_04824_));
 sg13g2_inv_2 _22448_ (.Y(_04825_),
    .A(net1139));
 sg13g2_a21oi_1 _22449_ (.A1(_10089_),
    .A2(net774),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_nor3_1 _22450_ (.A(net1058),
    .B(net799),
    .C(_04826_),
    .Y(_04827_));
 sg13g2_nor2_1 _22451_ (.A(_10561_),
    .B(net796),
    .Y(_04828_));
 sg13g2_o21ai_1 _22452_ (.B1(net785),
    .Y(_04829_),
    .A1(_04827_),
    .A2(_04828_));
 sg13g2_nor3_1 _22453_ (.A(net1058),
    .B(net799),
    .C(net1139),
    .Y(_04830_));
 sg13g2_o21ai_1 _22454_ (.B1(net1067),
    .Y(_04831_),
    .A1(_09762_),
    .A2(_04830_));
 sg13g2_nand2_1 _22455_ (.Y(_04832_),
    .A(net909),
    .B(_04825_));
 sg13g2_o21ai_1 _22456_ (.B1(_04832_),
    .Y(_04833_),
    .A1(net796),
    .A2(_04825_));
 sg13g2_nand2_1 _22457_ (.Y(_04834_),
    .A(net798),
    .B(_10089_));
 sg13g2_buf_1 _22458_ (.A(_04834_),
    .X(_04835_));
 sg13g2_nand2_1 _22459_ (.Y(_04836_),
    .A(net774),
    .B(net1139));
 sg13g2_o21ai_1 _22460_ (.B1(_04832_),
    .Y(_04837_),
    .A1(net582),
    .A2(_04836_));
 sg13g2_a22oi_1 _22461_ (.Y(_04838_),
    .B1(_04837_),
    .B2(net1058),
    .A2(_04833_),
    .A1(net798));
 sg13g2_nand3_1 _22462_ (.B(_04831_),
    .C(_04838_),
    .A(_04829_),
    .Y(_04839_));
 sg13g2_buf_2 _22463_ (.A(_04839_),
    .X(_04840_));
 sg13g2_nand2_1 _22464_ (.Y(_04841_),
    .A(net785),
    .B(_10089_));
 sg13g2_buf_1 _22465_ (.A(_04841_),
    .X(_04842_));
 sg13g2_nand2_1 _22466_ (.Y(_04843_),
    .A(net904),
    .B(net919));
 sg13g2_buf_1 _22467_ (.A(_04843_),
    .X(_04844_));
 sg13g2_nor3_1 _22468_ (.A(net1058),
    .B(net581),
    .C(_04844_),
    .Y(_04845_));
 sg13g2_buf_1 _22469_ (.A(_04845_),
    .X(_04846_));
 sg13g2_a21o_1 _22470_ (.A2(_04840_),
    .A1(_09255_),
    .B1(net455),
    .X(_04847_));
 sg13g2_buf_2 _22471_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04848_));
 sg13g2_buf_1 _22472_ (.A(_09758_),
    .X(_04849_));
 sg13g2_nand2_1 _22473_ (.Y(_04850_),
    .A(net904),
    .B(net915));
 sg13g2_buf_2 _22474_ (.A(_04850_),
    .X(_04851_));
 sg13g2_nor3_2 _22475_ (.A(_04849_),
    .B(_04851_),
    .C(net582),
    .Y(_04852_));
 sg13g2_nor3_1 _22476_ (.A(net1058),
    .B(_04851_),
    .C(net582),
    .Y(_04853_));
 sg13g2_buf_2 _22477_ (.A(_04853_),
    .X(_04854_));
 sg13g2_a22oi_1 _22478_ (.Y(_04855_),
    .B1(_04854_),
    .B2(_09255_),
    .A2(_04852_),
    .A1(_04848_));
 sg13g2_nor3_1 _22479_ (.A(net785),
    .B(net1139),
    .C(_04844_),
    .Y(_04856_));
 sg13g2_buf_1 _22480_ (.A(_04856_),
    .X(_04857_));
 sg13g2_buf_2 _22481_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04858_));
 sg13g2_buf_2 _22482_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04859_));
 sg13g2_mux2_1 _22483_ (.A0(_04858_),
    .A1(_04859_),
    .S(net681),
    .X(_04860_));
 sg13g2_nor3_1 _22484_ (.A(net785),
    .B(net900),
    .C(_04851_),
    .Y(_04861_));
 sg13g2_buf_1 _22485_ (.A(_04861_),
    .X(_04862_));
 sg13g2_and2_1 _22486_ (.A(net871),
    .B(net504),
    .X(_04863_));
 sg13g2_buf_2 _22487_ (.A(_04863_),
    .X(_04864_));
 sg13g2_buf_2 _22488_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04865_));
 sg13g2_a22oi_1 _22489_ (.Y(_04866_),
    .B1(_04864_),
    .B2(_04865_),
    .A2(_04860_),
    .A1(net505));
 sg13g2_buf_2 _22490_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04867_));
 sg13g2_nor3_2 _22491_ (.A(_12008_),
    .B(net772),
    .C(_02764_),
    .Y(_04868_));
 sg13g2_buf_1 _22492_ (.A(net683),
    .X(_04869_));
 sg13g2_nand2_1 _22493_ (.Y(_04870_),
    .A(_09239_),
    .B(net580));
 sg13g2_nor2_1 _22494_ (.A(_04825_),
    .B(_04870_),
    .Y(_04871_));
 sg13g2_buf_2 _22495_ (.A(_04871_),
    .X(_04872_));
 sg13g2_buf_2 _22496_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04873_));
 sg13g2_a22oi_1 _22497_ (.Y(_04874_),
    .B1(_04872_),
    .B2(_04873_),
    .A2(_04868_),
    .A1(_04867_));
 sg13g2_nand3_1 _22498_ (.B(_04866_),
    .C(_04874_),
    .A(_04855_),
    .Y(_04875_));
 sg13g2_a21oi_1 _22499_ (.A1(\cpu.gpio.r_enable_in[0] ),
    .A2(_04847_),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_and2_1 _22500_ (.A(net1071),
    .B(_10028_),
    .X(_04877_));
 sg13g2_buf_1 _22501_ (.A(_04877_),
    .X(_04878_));
 sg13g2_mux2_1 _22502_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(\cpu.intr.r_timer_reload[16] ),
    .S(net772),
    .X(_04879_));
 sg13g2_mux2_1 _22503_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(net772),
    .X(_04880_));
 sg13g2_buf_1 _22504_ (.A(net580),
    .X(_04881_));
 sg13g2_buf_1 _22505_ (.A(net503),
    .X(_04882_));
 sg13g2_buf_1 _22506_ (.A(net454),
    .X(_04883_));
 sg13g2_a22oi_1 _22507_ (.Y(_04884_),
    .B1(_04880_),
    .B2(net416),
    .A2(_04879_),
    .A1(net485));
 sg13g2_buf_1 _22508_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04885_));
 sg13g2_nor2_1 _22509_ (.A(_04851_),
    .B(net582),
    .Y(_04886_));
 sg13g2_buf_1 _22510_ (.A(_04886_),
    .X(_04887_));
 sg13g2_buf_1 _22511_ (.A(_04887_),
    .X(_04888_));
 sg13g2_a22oi_1 _22512_ (.Y(_04889_),
    .B1(net415),
    .B2(_09280_),
    .A2(net426),
    .A1(_04885_));
 sg13g2_buf_1 _22513_ (.A(net619),
    .X(_04890_));
 sg13g2_buf_1 _22514_ (.A(net502),
    .X(_04891_));
 sg13g2_buf_1 _22515_ (.A(net453),
    .X(_04892_));
 sg13g2_a22oi_1 _22516_ (.Y(_04893_),
    .B1(net424),
    .B2(_10160_),
    .A2(net414),
    .A1(_09985_));
 sg13g2_buf_1 _22517_ (.A(net414),
    .X(_04894_));
 sg13g2_nand3_1 _22518_ (.B(_09989_),
    .C(net381),
    .A(net772),
    .Y(_04895_));
 sg13g2_o21ai_1 _22519_ (.B1(_04895_),
    .Y(_04896_),
    .A1(net681),
    .A2(_04893_));
 sg13g2_inv_1 _22520_ (.Y(_04897_),
    .A(_04896_));
 sg13g2_a21oi_1 _22521_ (.A1(_10152_),
    .A2(_04835_),
    .Y(_04898_),
    .B1(net799));
 sg13g2_nor2_1 _22522_ (.A(net909),
    .B(_04898_),
    .Y(_04899_));
 sg13g2_buf_2 _22523_ (.A(_04899_),
    .X(_04900_));
 sg13g2_nor2_1 _22524_ (.A(_04851_),
    .B(_10152_),
    .Y(_04901_));
 sg13g2_buf_2 _22525_ (.A(_04901_),
    .X(_04902_));
 sg13g2_buf_1 _22526_ (.A(_04902_),
    .X(_04903_));
 sg13g2_a21o_1 _22527_ (.A2(_04900_),
    .A1(_09280_),
    .B1(net413),
    .X(_04904_));
 sg13g2_o21ai_1 _22528_ (.B1(_04904_),
    .Y(_04905_),
    .A1(_09278_),
    .A2(_09279_));
 sg13g2_nand4_1 _22529_ (.B(_04889_),
    .C(_04897_),
    .A(_04884_),
    .Y(_04906_),
    .D(_04905_));
 sg13g2_nor2_1 _22530_ (.A(_09238_),
    .B(_02764_),
    .Y(_04907_));
 sg13g2_buf_2 _22531_ (.A(_04907_),
    .X(_04908_));
 sg13g2_nor2_1 _22532_ (.A(net798),
    .B(_04836_),
    .Y(_04909_));
 sg13g2_buf_2 _22533_ (.A(_00230_),
    .X(_04910_));
 sg13g2_nor2_1 _22534_ (.A(net799),
    .B(_04910_),
    .Y(_04911_));
 sg13g2_o21ai_1 _22535_ (.B1(net1067),
    .Y(_04912_),
    .A1(_04909_),
    .A2(_04911_));
 sg13g2_a21oi_1 _22536_ (.A1(net799),
    .A2(_04832_),
    .Y(_04913_),
    .B1(net798));
 sg13g2_o21ai_1 _22537_ (.B1(_10089_),
    .Y(_04914_),
    .A1(_10095_),
    .A2(_09451_));
 sg13g2_nor2b_1 _22538_ (.A(_04913_),
    .B_N(_04914_),
    .Y(_04915_));
 sg13g2_nor3_1 _22539_ (.A(net1058),
    .B(_10152_),
    .C(_04844_),
    .Y(_04916_));
 sg13g2_buf_2 _22540_ (.A(_04916_),
    .X(_04917_));
 sg13g2_a221oi_1 _22541_ (.B2(_04915_),
    .C1(_04917_),
    .B1(_04912_),
    .A1(_12000_),
    .Y(_04918_),
    .A2(_04908_));
 sg13g2_buf_2 _22542_ (.A(_04918_),
    .X(_04919_));
 sg13g2_nand2_1 _22543_ (.Y(_04920_),
    .A(_09343_),
    .B(_04919_));
 sg13g2_nor2_1 _22544_ (.A(_04842_),
    .B(_04844_),
    .Y(_04921_));
 sg13g2_buf_2 _22545_ (.A(_04921_),
    .X(_04922_));
 sg13g2_a22oi_1 _22546_ (.Y(_04923_),
    .B1(_04922_),
    .B2(_12033_),
    .A2(_04908_),
    .A1(\cpu.spi.r_mode[1][0] ));
 sg13g2_or2_1 _22547_ (.X(_04924_),
    .B(_04923_),
    .A(net747));
 sg13g2_buf_1 _22548_ (.A(_04922_),
    .X(_04925_));
 sg13g2_nand3_1 _22549_ (.B(\cpu.spi.r_mode[2][0] ),
    .C(_04925_),
    .A(net747),
    .Y(_04926_));
 sg13g2_a22oi_1 _22550_ (.Y(_04927_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net624),
    .A2(_04910_),
    .A1(_09275_));
 sg13g2_nand3_1 _22551_ (.B(net796),
    .C(\cpu.spi.r_ready ),
    .A(net771),
    .Y(_04928_));
 sg13g2_o21ai_1 _22552_ (.B1(_04928_),
    .Y(_04929_),
    .A1(net678),
    .A2(_04927_));
 sg13g2_nor3_1 _22553_ (.A(net1139),
    .B(net542),
    .C(_04844_),
    .Y(_04930_));
 sg13g2_buf_2 _22554_ (.A(_04930_),
    .X(_04931_));
 sg13g2_buf_1 _22555_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04932_));
 sg13g2_nand3_1 _22556_ (.B(net1139),
    .C(net619),
    .A(net1067),
    .Y(_04933_));
 sg13g2_buf_2 _22557_ (.A(_04933_),
    .X(_04934_));
 sg13g2_nand2b_1 _22558_ (.Y(_04935_),
    .B(_04917_),
    .A_N(_00316_));
 sg13g2_o21ai_1 _22559_ (.B1(_04935_),
    .Y(_04936_),
    .A1(_00315_),
    .A2(_04934_));
 sg13g2_a221oi_1 _22560_ (.B2(_04932_),
    .C1(_04936_),
    .B1(_04931_),
    .A1(net694),
    .Y(_04937_),
    .A2(_04929_));
 sg13g2_nand4_1 _22561_ (.B(_04924_),
    .C(_04926_),
    .A(_04920_),
    .Y(_04938_),
    .D(_04937_));
 sg13g2_inv_1 _22562_ (.Y(_04939_),
    .A(_09232_));
 sg13g2_nand2b_1 _22563_ (.Y(_04940_),
    .B(net679),
    .A_N(_09231_));
 sg13g2_buf_2 _22564_ (.A(_04940_),
    .X(_04941_));
 sg13g2_o21ai_1 _22565_ (.B1(net774),
    .Y(_04942_),
    .A1(net775),
    .A2(_09805_));
 sg13g2_buf_2 _22566_ (.A(_04942_),
    .X(_04943_));
 sg13g2_nor2_1 _22567_ (.A(net542),
    .B(_04844_),
    .Y(_04944_));
 sg13g2_buf_1 _22568_ (.A(_04944_),
    .X(_04945_));
 sg13g2_a22oi_1 _22569_ (.Y(_04946_),
    .B1(net411),
    .B2(\cpu.uart.r_div_value[8] ),
    .A2(net504),
    .A1(\cpu.uart.r_x_invert ));
 sg13g2_a22oi_1 _22570_ (.Y(_04947_),
    .B1(_04922_),
    .B2(\cpu.uart.r_div_value[0] ),
    .A2(net415),
    .A1(_09278_));
 sg13g2_nand2_1 _22571_ (.Y(_04948_),
    .A(_04946_),
    .B(_04947_));
 sg13g2_a21oi_1 _22572_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04943_),
    .Y(_04949_),
    .B1(_04948_));
 sg13g2_nor2_1 _22573_ (.A(_04941_),
    .B(_04949_),
    .Y(_04950_));
 sg13g2_a221oi_1 _22574_ (.B2(_04939_),
    .C1(_04950_),
    .B1(_04938_),
    .A1(_04878_),
    .Y(_04951_),
    .A2(_04906_));
 sg13g2_o21ai_1 _22575_ (.B1(_04951_),
    .Y(_04952_),
    .A1(_04824_),
    .A2(_04876_));
 sg13g2_nand2b_1 _22576_ (.Y(_04953_),
    .B(net1092),
    .A_N(_08350_));
 sg13g2_nor3_1 _22577_ (.A(net1030),
    .B(net1152),
    .C(_04953_),
    .Y(_04954_));
 sg13g2_buf_2 _22578_ (.A(_04954_),
    .X(_04955_));
 sg13g2_buf_1 _22579_ (.A(net621),
    .X(_04956_));
 sg13g2_buf_1 _22580_ (.A(net501),
    .X(_04957_));
 sg13g2_nand2_1 _22581_ (.Y(_04958_),
    .A(\cpu.dcache.r_data[0][0] ),
    .B(net452));
 sg13g2_buf_1 _22582_ (.A(net615),
    .X(_04959_));
 sg13g2_buf_1 _22583_ (.A(net620),
    .X(_04960_));
 sg13g2_buf_1 _22584_ (.A(net499),
    .X(_04961_));
 sg13g2_a22oi_1 _22585_ (.Y(_04962_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][0] ),
    .A2(net500),
    .A1(\cpu.dcache.r_data[3][0] ));
 sg13g2_buf_1 _22586_ (.A(net618),
    .X(_04963_));
 sg13g2_a22oi_1 _22587_ (.Y(_04964_),
    .B1(net498),
    .B2(\cpu.dcache.r_data[1][0] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][0] ));
 sg13g2_mux2_1 _22588_ (.A0(\cpu.dcache.r_data[5][0] ),
    .A1(\cpu.dcache.r_data[7][0] ),
    .S(net799),
    .X(_04965_));
 sg13g2_a22oi_1 _22589_ (.Y(_04966_),
    .B1(_04965_),
    .B2(net694),
    .A2(_09521_),
    .A1(\cpu.dcache.r_data[4][0] ));
 sg13g2_nand2b_1 _22590_ (.Y(_04967_),
    .B(net748),
    .A_N(_04966_));
 sg13g2_nand4_1 _22591_ (.B(_04962_),
    .C(_04964_),
    .A(_04958_),
    .Y(_04968_),
    .D(_04967_));
 sg13g2_nand2_1 _22592_ (.Y(_04969_),
    .A(\cpu.dcache.r_data[0][16] ),
    .B(net501));
 sg13g2_a22oi_1 _22593_ (.Y(_04970_),
    .B1(net471),
    .B2(\cpu.dcache.r_data[4][16] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][16] ));
 sg13g2_a22oi_1 _22594_ (.Y(_04971_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][16] ),
    .A2(net498),
    .A1(\cpu.dcache.r_data[1][16] ));
 sg13g2_mux2_1 _22595_ (.A0(\cpu.dcache.r_data[5][16] ),
    .A1(\cpu.dcache.r_data[7][16] ),
    .S(net799),
    .X(_04972_));
 sg13g2_a22oi_1 _22596_ (.Y(_04973_),
    .B1(_04972_),
    .B2(_09236_),
    .A2(net775),
    .A1(\cpu.dcache.r_data[6][16] ));
 sg13g2_nand2b_1 _22597_ (.Y(_04974_),
    .B(net909),
    .A_N(_04973_));
 sg13g2_nand4_1 _22598_ (.B(_04970_),
    .C(_04971_),
    .A(_04969_),
    .Y(_04975_),
    .D(_04974_));
 sg13g2_mux2_1 _22599_ (.A0(_04968_),
    .A1(_04975_),
    .S(net613),
    .X(_04976_));
 sg13g2_nor2_1 _22600_ (.A(net678),
    .B(net1119),
    .Y(_04977_));
 sg13g2_a21oi_2 _22601_ (.B1(_04953_),
    .Y(_04978_),
    .A2(_08402_),
    .A1(_10645_));
 sg13g2_buf_1 _22602_ (.A(_04978_),
    .X(_04979_));
 sg13g2_a221oi_1 _22603_ (.B2(_04977_),
    .C1(_04979_),
    .B1(_04975_),
    .A1(net1119),
    .Y(_04980_),
    .A2(_04968_));
 sg13g2_a21o_1 _22604_ (.A2(net1030),
    .A1(_10645_),
    .B1(_04953_),
    .X(_04981_));
 sg13g2_buf_1 _22605_ (.A(_04981_),
    .X(_04982_));
 sg13g2_a22oi_1 _22606_ (.Y(_04983_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(net502),
    .A1(\cpu.dcache.r_data[6][8] ));
 sg13g2_a22oi_1 _22607_ (.Y(_04984_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][8] ),
    .A2(net499),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_a22oi_1 _22608_ (.Y(_04985_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[5][8] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][8] ));
 sg13g2_nand3_1 _22609_ (.B(_04984_),
    .C(_04985_),
    .A(_04983_),
    .Y(_04986_));
 sg13g2_nand2_1 _22610_ (.Y(_04987_),
    .A(_00314_),
    .B(net912));
 sg13g2_o21ai_1 _22611_ (.B1(_04987_),
    .Y(_04988_),
    .A1(net912),
    .A2(_04986_));
 sg13g2_nor3_1 _22612_ (.A(\cpu.dcache.r_data[1][8] ),
    .B(net745),
    .C(_04986_),
    .Y(_04989_));
 sg13g2_a21o_1 _22613_ (.A2(_04988_),
    .A1(net745),
    .B1(_04989_),
    .X(_04990_));
 sg13g2_nor2_1 _22614_ (.A(_10019_),
    .B(_04990_),
    .Y(_04991_));
 sg13g2_inv_2 _22615_ (.Y(_04992_),
    .A(_12082_));
 sg13g2_a22oi_1 _22616_ (.Y(_04993_),
    .B1(net499),
    .B2(\cpu.dcache.r_data[2][24] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][24] ));
 sg13g2_a22oi_1 _22617_ (.Y(_04994_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net498),
    .A1(\cpu.dcache.r_data[1][24] ));
 sg13g2_inv_1 _22618_ (.Y(_04995_),
    .A(_00313_));
 sg13g2_a22oi_1 _22619_ (.Y(_04996_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][24] ),
    .A2(_04956_),
    .A1(_04995_));
 sg13g2_a22oi_1 _22620_ (.Y(_04997_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][24] ),
    .A2(net502),
    .A1(\cpu.dcache.r_data[6][24] ));
 sg13g2_nand4_1 _22621_ (.B(_04994_),
    .C(_04996_),
    .A(_04993_),
    .Y(_04998_),
    .D(_04997_));
 sg13g2_buf_1 _22622_ (.A(_04998_),
    .X(_04999_));
 sg13g2_and2_1 _22623_ (.A(_04992_),
    .B(_04999_),
    .X(_05000_));
 sg13g2_nor3_1 _22624_ (.A(net649),
    .B(_04991_),
    .C(_05000_),
    .Y(_05001_));
 sg13g2_nor3_1 _22625_ (.A(_04980_),
    .B(_05001_),
    .C(_04955_),
    .Y(_05002_));
 sg13g2_a21oi_1 _22626_ (.A1(_04955_),
    .A2(_04976_),
    .Y(_05003_),
    .B1(_05002_));
 sg13g2_nor2_1 _22627_ (.A(net1025),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_1 _22628_ (.A1(net846),
    .A2(_04952_),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_buf_1 _22629_ (.A(_03570_),
    .X(_05006_));
 sg13g2_nand2_1 _22630_ (.Y(_05007_),
    .A(_03517_),
    .B(net81));
 sg13g2_o21ai_1 _22631_ (.B1(_05007_),
    .Y(_05008_),
    .A1(net82),
    .A2(_05005_));
 sg13g2_buf_1 _22632_ (.A(_11610_),
    .X(_05009_));
 sg13g2_and3_1 _22633_ (.X(_05010_),
    .A(net734),
    .B(net80),
    .C(_04817_));
 sg13g2_a21oi_1 _22634_ (.A1(net83),
    .A2(_05008_),
    .Y(_05011_),
    .B1(_05010_));
 sg13g2_o21ai_1 _22635_ (.B1(_05011_),
    .Y(_01033_),
    .A1(_04793_),
    .A2(_04819_));
 sg13g2_nor2_1 _22636_ (.A(net679),
    .B(_04900_),
    .Y(_05012_));
 sg13g2_and2_1 _22637_ (.A(net1025),
    .B(_05012_),
    .X(_05013_));
 sg13g2_buf_2 _22638_ (.A(_05013_),
    .X(_05014_));
 sg13g2_nand2_2 _22639_ (.Y(_05015_),
    .A(_10090_),
    .B(net909));
 sg13g2_mux2_1 _22640_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(\cpu.intr.r_timer_reload[10] ),
    .S(net624),
    .X(_05016_));
 sg13g2_a22oi_1 _22641_ (.Y(_05017_),
    .B1(_05016_),
    .B2(_09237_),
    .A2(_09521_),
    .A1(_10212_));
 sg13g2_nor2_1 _22642_ (.A(net771),
    .B(_12717_),
    .Y(_05018_));
 sg13g2_buf_2 _22643_ (.A(_05018_),
    .X(_05019_));
 sg13g2_buf_1 _22644_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05020_));
 sg13g2_inv_1 _22645_ (.Y(_05021_),
    .A(_05020_));
 sg13g2_nor3_1 _22646_ (.A(_05021_),
    .B(_09463_),
    .C(net542),
    .Y(_05022_));
 sg13g2_a221oi_1 _22647_ (.B2(\cpu.intr.r_clock_cmp[26] ),
    .C1(_05022_),
    .B1(_05019_),
    .A1(_09990_),
    .Y(_05023_),
    .A2(_04908_));
 sg13g2_o21ai_1 _22648_ (.B1(_05023_),
    .Y(_05024_),
    .A1(_05015_),
    .A2(_05017_));
 sg13g2_inv_1 _22649_ (.Y(_05025_),
    .A(_00103_));
 sg13g2_buf_1 _22650_ (.A(net452),
    .X(_05026_));
 sg13g2_a22oi_1 _22651_ (.Y(_05027_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net410),
    .A1(_05025_));
 sg13g2_a22oi_1 _22652_ (.Y(_05028_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][10] ),
    .A2(net473),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_a22oi_1 _22653_ (.Y(_05029_),
    .B1(net414),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][10] ));
 sg13g2_buf_1 _22654_ (.A(net498),
    .X(_05030_));
 sg13g2_buf_1 _22655_ (.A(net450),
    .X(_05031_));
 sg13g2_buf_1 _22656_ (.A(_04961_),
    .X(_05032_));
 sg13g2_a22oi_1 _22657_ (.Y(_05033_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][10] ),
    .A2(net409),
    .A1(\cpu.dcache.r_data[1][10] ));
 sg13g2_nand4_1 _22658_ (.B(_05028_),
    .C(_05029_),
    .A(_05027_),
    .Y(_05034_),
    .D(_05033_));
 sg13g2_nand2_1 _22659_ (.Y(_05035_),
    .A(\cpu.dcache.r_data[4][26] ),
    .B(net529));
 sg13g2_a22oi_1 _22660_ (.Y(_05036_),
    .B1(net498),
    .B2(\cpu.dcache.r_data[1][26] ),
    .A2(net502),
    .A1(\cpu.dcache.r_data[6][26] ));
 sg13g2_a22oi_1 _22661_ (.Y(_05037_),
    .B1(_04869_),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_a22oi_1 _22662_ (.Y(_05038_),
    .B1(net499),
    .B2(\cpu.dcache.r_data[2][26] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][26] ));
 sg13g2_nand4_1 _22663_ (.B(_05036_),
    .C(_05037_),
    .A(_05035_),
    .Y(_05039_),
    .D(_05038_));
 sg13g2_nor2_1 _22664_ (.A(net452),
    .B(_05039_),
    .Y(_05040_));
 sg13g2_a21oi_1 _22665_ (.A1(_00102_),
    .A2(net410),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_buf_1 _22666_ (.A(_10019_),
    .X(_05042_));
 sg13g2_mux2_1 _22667_ (.A0(_05034_),
    .A1(_05041_),
    .S(net648),
    .X(_05043_));
 sg13g2_a22oi_1 _22668_ (.Y(_05044_),
    .B1(_05043_),
    .B2(_04955_),
    .A2(_05024_),
    .A1(_05014_));
 sg13g2_a21oi_2 _22669_ (.B1(net1152),
    .Y(_05045_),
    .A2(_08402_),
    .A1(net1151));
 sg13g2_nand2_2 _22670_ (.Y(_05046_),
    .A(_04978_),
    .B(_05045_));
 sg13g2_nand2_1 _22671_ (.Y(_05047_),
    .A(\cpu.dcache.r_data[2][23] ),
    .B(net620));
 sg13g2_a22oi_1 _22672_ (.Y(_05048_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[3][23] ),
    .A2(net619),
    .A1(\cpu.dcache.r_data[6][23] ));
 sg13g2_a22oi_1 _22673_ (.Y(_05049_),
    .B1(net617),
    .B2(\cpu.dcache.r_data[4][23] ),
    .A2(net580),
    .A1(\cpu.dcache.r_data[5][23] ));
 sg13g2_a22oi_1 _22674_ (.Y(_05050_),
    .B1(net618),
    .B2(\cpu.dcache.r_data[1][23] ),
    .A2(net786),
    .A1(\cpu.dcache.r_data[7][23] ));
 sg13g2_nand4_1 _22675_ (.B(_05048_),
    .C(_05049_),
    .A(_05047_),
    .Y(_05051_),
    .D(_05050_));
 sg13g2_nand2_1 _22676_ (.Y(_05052_),
    .A(_00153_),
    .B(net501));
 sg13g2_o21ai_1 _22677_ (.B1(_05052_),
    .Y(_05053_),
    .A1(net501),
    .A2(_05051_));
 sg13g2_or2_1 _22678_ (.X(_05054_),
    .B(_05053_),
    .A(_10090_));
 sg13g2_nand2_1 _22679_ (.Y(_05055_),
    .A(\cpu.dcache.r_data[2][7] ),
    .B(net620));
 sg13g2_a22oi_1 _22680_ (.Y(_05056_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[3][7] ),
    .A2(net619),
    .A1(\cpu.dcache.r_data[6][7] ));
 sg13g2_a22oi_1 _22681_ (.Y(_05057_),
    .B1(net617),
    .B2(\cpu.dcache.r_data[4][7] ),
    .A2(net580),
    .A1(\cpu.dcache.r_data[5][7] ));
 sg13g2_a22oi_1 _22682_ (.Y(_05058_),
    .B1(net618),
    .B2(\cpu.dcache.r_data[1][7] ),
    .A2(net786),
    .A1(\cpu.dcache.r_data[7][7] ));
 sg13g2_nand4_1 _22683_ (.B(_05056_),
    .C(_05057_),
    .A(_05055_),
    .Y(_05059_),
    .D(_05058_));
 sg13g2_nand2_1 _22684_ (.Y(_05060_),
    .A(_00152_),
    .B(net501));
 sg13g2_o21ai_1 _22685_ (.B1(_05060_),
    .Y(_05061_),
    .A1(net501),
    .A2(_05059_));
 sg13g2_mux2_1 _22686_ (.A0(_05054_),
    .A1(_05061_),
    .S(net1119),
    .X(_05062_));
 sg13g2_a22oi_1 _22687_ (.Y(_05063_),
    .B1(_09547_),
    .B2(\cpu.dcache.r_data[3][31] ),
    .A2(_09454_),
    .A1(\cpu.dcache.r_data[6][31] ));
 sg13g2_a22oi_1 _22688_ (.Y(_05064_),
    .B1(_09493_),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(_09447_),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_a22oi_1 _22689_ (.Y(_05065_),
    .B1(net683),
    .B2(\cpu.dcache.r_data[5][31] ),
    .A2(_09430_),
    .A1(\cpu.dcache.r_data[7][31] ));
 sg13g2_nand3_1 _22690_ (.B(_05064_),
    .C(_05065_),
    .A(_05063_),
    .Y(_05066_));
 sg13g2_nand2_1 _22691_ (.Y(_05067_),
    .A(_00154_),
    .B(net912));
 sg13g2_o21ai_1 _22692_ (.B1(_05067_),
    .Y(_05068_),
    .A1(net912),
    .A2(_05066_));
 sg13g2_nor3_1 _22693_ (.A(\cpu.dcache.r_data[1][31] ),
    .B(_09788_),
    .C(_05066_),
    .Y(_05069_));
 sg13g2_a21o_1 _22694_ (.A2(_05068_),
    .A1(_12188_),
    .B1(_05069_),
    .X(_05070_));
 sg13g2_buf_1 _22695_ (.A(_05070_),
    .X(_05071_));
 sg13g2_inv_1 _22696_ (.Y(_05072_),
    .A(_00155_));
 sg13g2_a22oi_1 _22697_ (.Y(_05073_),
    .B1(net620),
    .B2(\cpu.dcache.r_data[2][15] ),
    .A2(_04956_),
    .A1(_05072_));
 sg13g2_a22oi_1 _22698_ (.Y(_05074_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(_04869_),
    .A1(\cpu.dcache.r_data[5][15] ));
 sg13g2_a22oi_1 _22699_ (.Y(_05075_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[6][15] ),
    .A2(net786),
    .A1(\cpu.dcache.r_data[7][15] ));
 sg13g2_a22oi_1 _22700_ (.Y(_05076_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[3][15] ),
    .A2(net498),
    .A1(\cpu.dcache.r_data[1][15] ));
 sg13g2_nand4_1 _22701_ (.B(_05074_),
    .C(_05075_),
    .A(_05073_),
    .Y(_05077_),
    .D(_05076_));
 sg13g2_nand2_1 _22702_ (.Y(_05078_),
    .A(net900),
    .B(_05077_));
 sg13g2_o21ai_1 _22703_ (.B1(_05078_),
    .Y(_05079_),
    .A1(_00277_),
    .A2(_05071_));
 sg13g2_nand2_1 _22704_ (.Y(_05080_),
    .A(_04979_),
    .B(_05079_));
 sg13g2_o21ai_1 _22705_ (.B1(_05080_),
    .Y(_05081_),
    .A1(net650),
    .A2(_05062_));
 sg13g2_nand2b_1 _22706_ (.Y(_05082_),
    .B(net900),
    .A_N(_05061_));
 sg13g2_a21oi_1 _22707_ (.A1(_05054_),
    .A2(_05082_),
    .Y(_05083_),
    .B1(_05046_));
 sg13g2_a21oi_1 _22708_ (.A1(_05046_),
    .A2(_05081_),
    .Y(_05084_),
    .B1(_05083_));
 sg13g2_nor2_1 _22709_ (.A(net1067),
    .B(_10140_),
    .Y(_05085_));
 sg13g2_buf_2 _22710_ (.A(_05085_),
    .X(_05086_));
 sg13g2_nand2_1 _22711_ (.Y(_05087_),
    .A(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .B(_05086_));
 sg13g2_nor2_1 _22712_ (.A(net1067),
    .B(_12717_),
    .Y(_05088_));
 sg13g2_a22oi_1 _22713_ (.Y(_05089_),
    .B1(_05088_),
    .B2(net10),
    .A2(_10154_),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_a21oi_1 _22714_ (.A1(_09256_),
    .A2(_04902_),
    .Y(_05090_),
    .B1(_04861_));
 sg13g2_nand2b_1 _22715_ (.Y(_05091_),
    .B(_09257_),
    .A_N(_05090_));
 sg13g2_nand3_1 _22716_ (.B(_05089_),
    .C(_05091_),
    .A(_05087_),
    .Y(_05092_));
 sg13g2_a21o_1 _22717_ (.A2(_04840_),
    .A1(_09251_),
    .B1(_04854_),
    .X(_05093_));
 sg13g2_a221oi_1 _22718_ (.B2(_09256_),
    .C1(net1058),
    .B1(net411),
    .A1(_09251_),
    .Y(_05094_),
    .A2(_04922_));
 sg13g2_inv_1 _22719_ (.Y(_05095_),
    .A(_00159_));
 sg13g2_inv_1 _22720_ (.Y(_05096_),
    .A(_00161_));
 sg13g2_a221oi_1 _22721_ (.B2(_05096_),
    .C1(net872),
    .B1(_04902_),
    .A1(_05095_),
    .Y(_05097_),
    .A2(net504));
 sg13g2_inv_1 _22722_ (.Y(_05098_),
    .A(_00162_));
 sg13g2_nand2_2 _22723_ (.Y(_05099_),
    .A(_04825_),
    .B(_04887_));
 sg13g2_nor2_1 _22724_ (.A(net900),
    .B(_00158_),
    .Y(_05100_));
 sg13g2_buf_1 _22725_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05101_));
 sg13g2_nor2b_1 _22726_ (.A(_09239_),
    .B_N(_05101_),
    .Y(_05102_));
 sg13g2_o21ai_1 _22727_ (.B1(_04857_),
    .Y(_05103_),
    .A1(_05100_),
    .A2(_05102_));
 sg13g2_o21ai_1 _22728_ (.B1(_05103_),
    .Y(_05104_),
    .A1(_00160_),
    .A2(_05099_));
 sg13g2_a21oi_1 _22729_ (.A1(_05098_),
    .A2(_04872_),
    .Y(_05105_),
    .B1(_05104_));
 sg13g2_o21ai_1 _22730_ (.B1(_05105_),
    .Y(_05106_),
    .A1(_05094_),
    .A2(_05097_));
 sg13g2_a221oi_1 _22731_ (.B2(_09252_),
    .C1(_05106_),
    .B1(_05093_),
    .A1(net1139),
    .Y(_05107_),
    .A2(_05092_));
 sg13g2_inv_1 _22732_ (.Y(_05108_),
    .A(_00157_));
 sg13g2_buf_1 _22733_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05109_));
 sg13g2_a22oi_1 _22734_ (.Y(_05110_),
    .B1(_04931_),
    .B2(_05109_),
    .A2(_04917_),
    .A1(_05108_));
 sg13g2_nor3_1 _22735_ (.A(net654),
    .B(net900),
    .C(net796),
    .Y(_05111_));
 sg13g2_buf_2 _22736_ (.A(_05111_),
    .X(_05112_));
 sg13g2_nor2_1 _22737_ (.A(_00156_),
    .B(_04934_),
    .Y(_05113_));
 sg13g2_a21oi_1 _22738_ (.A1(\cpu.spi.r_timeout[7] ),
    .A2(_05112_),
    .Y(_05114_),
    .B1(_05113_));
 sg13g2_nand2b_1 _22739_ (.Y(_05115_),
    .B(_04919_),
    .A_N(_00224_));
 sg13g2_nand3_1 _22740_ (.B(_05114_),
    .C(_05115_),
    .A(_05110_),
    .Y(_05116_));
 sg13g2_a22oi_1 _22741_ (.Y(_05117_),
    .B1(_04943_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04922_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_a22oi_1 _22742_ (.Y(_05118_),
    .B1(net580),
    .B2(\cpu.intr.r_clock_cmp[23] ),
    .A2(net502),
    .A1(_10014_));
 sg13g2_nor2_1 _22743_ (.A(net900),
    .B(_05118_),
    .Y(_05119_));
 sg13g2_mux2_1 _22744_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(\cpu.intr.r_timer_reload[7] ),
    .S(net799),
    .X(_05120_));
 sg13g2_a22oi_1 _22745_ (.Y(_05121_),
    .B1(_05120_),
    .B2(net798),
    .A2(net775),
    .A1(_09991_));
 sg13g2_buf_2 _22746_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05122_));
 sg13g2_and3_1 _22747_ (.X(_05123_),
    .A(net1067),
    .B(\cpu.intr.r_timer_reload[23] ),
    .C(net680));
 sg13g2_a221oi_1 _22748_ (.B2(_10195_),
    .C1(_05123_),
    .B1(_05086_),
    .A1(_05122_),
    .Y(_05124_),
    .A2(_10154_));
 sg13g2_o21ai_1 _22749_ (.B1(_05124_),
    .Y(_05125_),
    .A1(_05015_),
    .A2(_05121_));
 sg13g2_o21ai_1 _22750_ (.B1(_05012_),
    .Y(_05126_),
    .A1(_05119_),
    .A2(_05125_));
 sg13g2_o21ai_1 _22751_ (.B1(_05126_),
    .Y(_05127_),
    .A1(_04941_),
    .A2(_05117_));
 sg13g2_a21oi_1 _22752_ (.A1(_04939_),
    .A2(_05116_),
    .Y(_05128_),
    .B1(_05127_));
 sg13g2_o21ai_1 _22753_ (.B1(_05128_),
    .Y(_05129_),
    .A1(_04824_),
    .A2(_05107_));
 sg13g2_nand2_1 _22754_ (.Y(_05130_),
    .A(_08350_),
    .B(_05129_));
 sg13g2_o21ai_1 _22755_ (.B1(_05130_),
    .Y(_05131_),
    .A1(_12080_),
    .A2(_05084_));
 sg13g2_a21oi_1 _22756_ (.A1(net1030),
    .A2(_05131_),
    .Y(_05132_),
    .B1(_11610_));
 sg13g2_buf_1 _22757_ (.A(_05132_),
    .X(_05133_));
 sg13g2_o21ai_1 _22758_ (.B1(_05133_),
    .Y(_05134_),
    .A1(net1030),
    .A2(_05044_));
 sg13g2_nand2b_1 _22759_ (.Y(_05135_),
    .B(net81),
    .A_N(_10903_));
 sg13g2_o21ai_1 _22760_ (.B1(_05135_),
    .Y(_05136_),
    .A1(net81),
    .A2(_05134_));
 sg13g2_buf_1 _22761_ (.A(_04216_),
    .X(_05137_));
 sg13g2_nand3_1 _22762_ (.B(net80),
    .C(net177),
    .A(net985),
    .Y(_05138_));
 sg13g2_o21ai_1 _22763_ (.B1(_05138_),
    .Y(_05139_),
    .A1(_11612_),
    .A2(_05136_));
 sg13g2_buf_1 _22764_ (.A(_11601_),
    .X(_05140_));
 sg13g2_a21oi_2 _22765_ (.B1(_04216_),
    .Y(_05141_),
    .A2(_03570_),
    .A1(_03568_));
 sg13g2_nand3_1 _22766_ (.B(_05134_),
    .C(_05141_),
    .A(net579),
    .Y(_05142_));
 sg13g2_a21oi_1 _22767_ (.A1(_04703_),
    .A2(_04731_),
    .Y(_05143_),
    .B1(_05142_));
 sg13g2_a21oi_1 _22768_ (.A1(_00260_),
    .A2(_11598_),
    .Y(_05144_),
    .B1(_11599_));
 sg13g2_buf_2 _22769_ (.A(_05144_),
    .X(_05145_));
 sg13g2_buf_1 _22770_ (.A(_05145_),
    .X(_05146_));
 sg13g2_and4_1 _22771_ (.A(net578),
    .B(_04735_),
    .C(_05134_),
    .D(_05141_),
    .X(_05147_));
 sg13g2_or3_1 _22772_ (.A(_05139_),
    .B(_05143_),
    .C(_05147_),
    .X(_01034_));
 sg13g2_nor3_1 _22773_ (.A(_04294_),
    .B(_04298_),
    .C(_04817_),
    .Y(_05148_));
 sg13g2_nor2_1 _22774_ (.A(\cpu.ex.pc[11] ),
    .B(_04095_),
    .Y(_05149_));
 sg13g2_nor3_1 _22775_ (.A(net579),
    .B(net177),
    .C(_04237_),
    .Y(_05150_));
 sg13g2_or3_1 _22776_ (.A(net83),
    .B(_05149_),
    .C(_05150_),
    .X(_05151_));
 sg13g2_nor2_1 _22777_ (.A(_11599_),
    .B(_05131_),
    .Y(_05152_));
 sg13g2_buf_1 _22778_ (.A(_04955_),
    .X(_05153_));
 sg13g2_nand2_1 _22779_ (.Y(_05154_),
    .A(\cpu.dcache.r_data[2][27] ),
    .B(net408));
 sg13g2_a22oi_1 _22780_ (.Y(_05155_),
    .B1(net500),
    .B2(\cpu.dcache.r_data[3][27] ),
    .A2(_04891_),
    .A1(\cpu.dcache.r_data[6][27] ));
 sg13g2_a22oi_1 _22781_ (.Y(_05156_),
    .B1(net471),
    .B2(\cpu.dcache.r_data[4][27] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[5][27] ));
 sg13g2_a22oi_1 _22782_ (.Y(_05157_),
    .B1(net450),
    .B2(\cpu.dcache.r_data[1][27] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][27] ));
 sg13g2_nand4_1 _22783_ (.B(_05155_),
    .C(_05156_),
    .A(_05154_),
    .Y(_05158_),
    .D(_05157_));
 sg13g2_nand2_1 _22784_ (.Y(_05159_),
    .A(_00112_),
    .B(net410));
 sg13g2_o21ai_1 _22785_ (.B1(_05159_),
    .Y(_05160_),
    .A1(net410),
    .A2(_05158_));
 sg13g2_inv_1 _22786_ (.Y(_05161_),
    .A(_00113_));
 sg13g2_a22oi_1 _22787_ (.Y(_05162_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[4][11] ),
    .A2(_05026_),
    .A1(_05161_));
 sg13g2_a22oi_1 _22788_ (.Y(_05163_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][11] ),
    .A2(net473),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_a22oi_1 _22789_ (.Y(_05164_),
    .B1(net414),
    .B2(\cpu.dcache.r_data[6][11] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][11] ));
 sg13g2_a22oi_1 _22790_ (.Y(_05165_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][11] ),
    .A2(net409),
    .A1(\cpu.dcache.r_data[1][11] ));
 sg13g2_nand4_1 _22791_ (.B(_05163_),
    .C(_05164_),
    .A(_05162_),
    .Y(_05166_),
    .D(_05165_));
 sg13g2_nand2_1 _22792_ (.Y(_05167_),
    .A(net611),
    .B(_05166_));
 sg13g2_o21ai_1 _22793_ (.B1(_05167_),
    .Y(_05168_),
    .A1(net544),
    .A2(_05160_));
 sg13g2_mux2_1 _22794_ (.A0(_10217_),
    .A1(\cpu.intr.r_timer_count[11] ),
    .S(net624),
    .X(_05169_));
 sg13g2_a22oi_1 _22795_ (.Y(_05170_),
    .B1(_05169_),
    .B2(net654),
    .A2(_10095_),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_buf_2 _22796_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05171_));
 sg13g2_mux2_1 _22797_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(\cpu.intr.r_clock_cmp[27] ),
    .S(net613),
    .X(_05172_));
 sg13g2_a22oi_1 _22798_ (.Y(_05173_),
    .B1(_05172_),
    .B2(net416),
    .A2(net384),
    .A1(_05171_));
 sg13g2_o21ai_1 _22799_ (.B1(_05173_),
    .Y(_05174_),
    .A1(_05015_),
    .A2(_05170_));
 sg13g2_a221oi_1 _22800_ (.B2(_05014_),
    .C1(net850),
    .B1(_05174_),
    .A1(net577),
    .Y(_05175_),
    .A2(_05168_));
 sg13g2_nor3_1 _22801_ (.A(net82),
    .B(_05152_),
    .C(_05175_),
    .Y(_05176_));
 sg13g2_and2_1 _22802_ (.A(_10925_),
    .B(net82),
    .X(_05177_));
 sg13g2_buf_1 _22803_ (.A(net83),
    .X(_05178_));
 sg13g2_o21ai_1 _22804_ (.B1(net74),
    .Y(_05179_),
    .A1(_05176_),
    .A2(_05177_));
 sg13g2_o21ai_1 _22805_ (.B1(_05179_),
    .Y(_01035_),
    .A1(_05148_),
    .A2(_05151_));
 sg13g2_nor3_1 _22806_ (.A(net579),
    .B(_05137_),
    .C(_04341_),
    .Y(_05180_));
 sg13g2_a21o_1 _22807_ (.A2(_05137_),
    .A1(_08373_),
    .B1(_05180_),
    .X(_05181_));
 sg13g2_buf_1 _22808_ (.A(net85),
    .X(_05182_));
 sg13g2_buf_1 _22809_ (.A(_05086_),
    .X(_05183_));
 sg13g2_buf_1 _22810_ (.A(_05088_),
    .X(_05184_));
 sg13g2_a22oi_1 _22811_ (.Y(_05185_),
    .B1(net448),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net449),
    .A1(_10224_));
 sg13g2_buf_2 _22812_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05186_));
 sg13g2_a22oi_1 _22813_ (.Y(_05187_),
    .B1(_05019_),
    .B2(\cpu.intr.r_clock_cmp[28] ),
    .A2(net384),
    .A1(_05186_));
 sg13g2_a22oi_1 _22814_ (.Y(_05188_),
    .B1(net381),
    .B2(\cpu.intr.r_timer_count[12] ),
    .A2(net485),
    .A1(\cpu.intr.r_timer_reload[12] ));
 sg13g2_or2_1 _22815_ (.X(_05189_),
    .B(_05188_),
    .A(net648));
 sg13g2_nand3_1 _22816_ (.B(_05187_),
    .C(_05189_),
    .A(_05185_),
    .Y(_05190_));
 sg13g2_a22oi_1 _22817_ (.Y(_05191_),
    .B1(_04960_),
    .B2(\cpu.dcache.r_data[2][28] ),
    .A2(_10023_),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_a22oi_1 _22818_ (.Y(_05192_),
    .B1(_12663_),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(_04963_),
    .A1(\cpu.dcache.r_data[1][28] ));
 sg13g2_inv_1 _22819_ (.Y(_05193_),
    .A(_00123_));
 sg13g2_a22oi_1 _22820_ (.Y(_05194_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(net501),
    .A1(_05193_));
 sg13g2_a22oi_1 _22821_ (.Y(_05195_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][28] ),
    .A2(_04890_),
    .A1(\cpu.dcache.r_data[6][28] ));
 sg13g2_nand4_1 _22822_ (.B(_05192_),
    .C(_05194_),
    .A(_05191_),
    .Y(_05196_),
    .D(_05195_));
 sg13g2_buf_1 _22823_ (.A(_05196_),
    .X(_05197_));
 sg13g2_a22oi_1 _22824_ (.Y(_05198_),
    .B1(_12534_),
    .B2(\cpu.dcache.r_data[3][12] ),
    .A2(_10023_),
    .A1(\cpu.dcache.r_data[7][12] ));
 sg13g2_o21ai_1 _22825_ (.B1(_05198_),
    .Y(_05199_),
    .A1(_00124_),
    .A2(net616));
 sg13g2_a221oi_1 _22826_ (.B2(\cpu.dcache.r_data[2][12] ),
    .C1(_05199_),
    .B1(net408),
    .A1(\cpu.dcache.r_data[1][12] ),
    .Y(_05200_),
    .A2(_05031_));
 sg13g2_mux2_1 _22827_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(\cpu.dcache.r_data[6][12] ),
    .S(_09222_),
    .X(_05201_));
 sg13g2_a22oi_1 _22828_ (.Y(_05202_),
    .B1(_05201_),
    .B2(_03785_),
    .A2(_09805_),
    .A1(\cpu.dcache.r_data[5][12] ));
 sg13g2_nand2b_1 _22829_ (.Y(_05203_),
    .B(net748),
    .A_N(_05202_));
 sg13g2_and2_1 _22830_ (.A(_05200_),
    .B(_05203_),
    .X(_05204_));
 sg13g2_nor2_1 _22831_ (.A(net648),
    .B(_05204_),
    .Y(_05205_));
 sg13g2_a21o_1 _22832_ (.A2(_05197_),
    .A1(net613),
    .B1(_05205_),
    .X(_05206_));
 sg13g2_a22oi_1 _22833_ (.Y(_05207_),
    .B1(_05206_),
    .B2(_05153_),
    .A2(_05190_),
    .A1(_05014_));
 sg13g2_o21ai_1 _22834_ (.B1(_05133_),
    .Y(_05208_),
    .A1(net1030),
    .A2(_05207_));
 sg13g2_nor2_1 _22835_ (.A(net81),
    .B(_05208_),
    .Y(_05209_));
 sg13g2_a21oi_1 _22836_ (.A1(_11946_),
    .A2(_04821_),
    .Y(_05210_),
    .B1(_05209_));
 sg13g2_nor2_1 _22837_ (.A(net85),
    .B(_05210_),
    .Y(_05211_));
 sg13g2_a221oi_1 _22838_ (.B2(net73),
    .C1(_05211_),
    .B1(_05181_),
    .A1(_04339_),
    .Y(_01036_),
    .A2(_04818_));
 sg13g2_mux2_1 _22839_ (.A0(_10230_),
    .A1(\cpu.intr.r_timer_count[13] ),
    .S(net695),
    .X(_05212_));
 sg13g2_a22oi_1 _22840_ (.Y(_05213_),
    .B1(_05212_),
    .B2(net654),
    .A2(_10095_),
    .A1(\cpu.intr.r_timer_reload[13] ));
 sg13g2_buf_1 _22841_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05214_));
 sg13g2_mux2_1 _22842_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(\cpu.intr.r_clock_cmp[29] ),
    .S(_10018_),
    .X(_05215_));
 sg13g2_a22oi_1 _22843_ (.Y(_05216_),
    .B1(_05215_),
    .B2(_04883_),
    .A2(net426),
    .A1(_05214_));
 sg13g2_o21ai_1 _22844_ (.B1(_05216_),
    .Y(_05217_),
    .A1(_05015_),
    .A2(_05213_));
 sg13g2_inv_1 _22845_ (.Y(_05218_),
    .A(_00130_));
 sg13g2_a22oi_1 _22846_ (.Y(_05219_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[4][29] ),
    .A2(net452),
    .A1(_05218_));
 sg13g2_a22oi_1 _22847_ (.Y(_05220_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][29] ),
    .A2(_04959_),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_a22oi_1 _22848_ (.Y(_05221_),
    .B1(net414),
    .B2(\cpu.dcache.r_data[6][29] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][29] ));
 sg13g2_a22oi_1 _22849_ (.Y(_05222_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][29] ),
    .A2(net450),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_nand4_1 _22850_ (.B(_05220_),
    .C(_05221_),
    .A(_05219_),
    .Y(_05223_),
    .D(_05222_));
 sg13g2_inv_1 _22851_ (.Y(_05224_),
    .A(_00131_));
 sg13g2_a22oi_1 _22852_ (.Y(_05225_),
    .B1(_05032_),
    .B2(\cpu.dcache.r_data[2][13] ),
    .A2(net452),
    .A1(_05224_));
 sg13g2_a22oi_1 _22853_ (.Y(_05226_),
    .B1(_12664_),
    .B2(\cpu.dcache.r_data[4][13] ),
    .A2(_04881_),
    .A1(\cpu.dcache.r_data[5][13] ));
 sg13g2_a22oi_1 _22854_ (.Y(_05227_),
    .B1(_04892_),
    .B2(\cpu.dcache.r_data[6][13] ),
    .A2(_10024_),
    .A1(\cpu.dcache.r_data[7][13] ));
 sg13g2_a22oi_1 _22855_ (.Y(_05228_),
    .B1(net473),
    .B2(\cpu.dcache.r_data[3][13] ),
    .A2(net450),
    .A1(\cpu.dcache.r_data[1][13] ));
 sg13g2_nand4_1 _22856_ (.B(_05226_),
    .C(_05227_),
    .A(_05225_),
    .Y(_05229_),
    .D(_05228_));
 sg13g2_mux2_1 _22857_ (.A0(_05223_),
    .A1(_05229_),
    .S(_10092_),
    .X(_05230_));
 sg13g2_a22oi_1 _22858_ (.Y(_05231_),
    .B1(_05230_),
    .B2(_04955_),
    .A2(_05217_),
    .A1(_05014_));
 sg13g2_nor2_1 _22859_ (.A(net1030),
    .B(_05231_),
    .Y(_05232_));
 sg13g2_nor2b_1 _22860_ (.A(_05232_),
    .B_N(_05133_),
    .Y(_05233_));
 sg13g2_nand2b_1 _22861_ (.Y(_05234_),
    .B(_05141_),
    .A_N(_05233_));
 sg13g2_nand2b_1 _22862_ (.Y(_05235_),
    .B(net579),
    .A_N(_05234_));
 sg13g2_nor2_1 _22863_ (.A(_03570_),
    .B(_05233_),
    .Y(_05236_));
 sg13g2_a21oi_1 _22864_ (.A1(net776),
    .A2(_05006_),
    .Y(_05237_),
    .B1(_05236_));
 sg13g2_nand3_1 _22865_ (.B(_05009_),
    .C(_04216_),
    .A(_08466_),
    .Y(_05238_));
 sg13g2_o21ai_1 _22866_ (.B1(_05238_),
    .Y(_05239_),
    .A1(_05009_),
    .A2(_05237_));
 sg13g2_nand2_1 _22867_ (.Y(_05240_),
    .A(net578),
    .B(_04380_));
 sg13g2_nor2_1 _22868_ (.A(_05234_),
    .B(_05240_),
    .Y(_05241_));
 sg13g2_nor2_1 _22869_ (.A(_05239_),
    .B(_05241_),
    .Y(_05242_));
 sg13g2_o21ai_1 _22870_ (.B1(_05242_),
    .Y(_01037_),
    .A1(_04378_),
    .A2(_05235_));
 sg13g2_buf_1 _22871_ (.A(_04095_),
    .X(_05243_));
 sg13g2_nand3b_1 _22872_ (.B(_05243_),
    .C(net578),
    .Y(_05244_),
    .A_N(_04418_));
 sg13g2_o21ai_1 _22873_ (.B1(_05244_),
    .Y(_05245_),
    .A1(_08476_),
    .A2(_05243_));
 sg13g2_nand2_1 _22874_ (.Y(_05246_),
    .A(\cpu.dcache.r_data[4][30] ),
    .B(_12663_));
 sg13g2_a22oi_1 _22875_ (.Y(_05247_),
    .B1(_04963_),
    .B2(\cpu.dcache.r_data[1][30] ),
    .A2(_04890_),
    .A1(\cpu.dcache.r_data[6][30] ));
 sg13g2_a22oi_1 _22876_ (.Y(_05248_),
    .B1(_04881_),
    .B2(\cpu.dcache.r_data[5][30] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_a22oi_1 _22877_ (.Y(_05249_),
    .B1(_04960_),
    .B2(\cpu.dcache.r_data[2][30] ),
    .A2(_10022_),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_nand4_1 _22878_ (.B(_05247_),
    .C(_05248_),
    .A(_05246_),
    .Y(_05250_),
    .D(_05249_));
 sg13g2_nand2_1 _22879_ (.Y(_05251_),
    .A(_00142_),
    .B(_04957_));
 sg13g2_o21ai_1 _22880_ (.B1(_05251_),
    .Y(_05252_),
    .A1(_04957_),
    .A2(_05250_));
 sg13g2_inv_1 _22881_ (.Y(_05253_),
    .A(_00143_));
 sg13g2_a22oi_1 _22882_ (.Y(_05254_),
    .B1(_12665_),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(_05026_),
    .A1(_05253_));
 sg13g2_a22oi_1 _22883_ (.Y(_05255_),
    .B1(_04882_),
    .B2(\cpu.dcache.r_data[5][14] ),
    .A2(_12535_),
    .A1(\cpu.dcache.r_data[3][14] ));
 sg13g2_a22oi_1 _22884_ (.Y(_05256_),
    .B1(_04892_),
    .B2(\cpu.dcache.r_data[6][14] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][14] ));
 sg13g2_a22oi_1 _22885_ (.Y(_05257_),
    .B1(_05032_),
    .B2(\cpu.dcache.r_data[2][14] ),
    .A2(net409),
    .A1(\cpu.dcache.r_data[1][14] ));
 sg13g2_nand4_1 _22886_ (.B(_05255_),
    .C(_05256_),
    .A(_05254_),
    .Y(_05258_),
    .D(_05257_));
 sg13g2_nand2_1 _22887_ (.Y(_05259_),
    .A(net611),
    .B(_05258_));
 sg13g2_o21ai_1 _22888_ (.B1(_05259_),
    .Y(_05260_),
    .A1(net544),
    .A2(_05252_));
 sg13g2_a22oi_1 _22889_ (.Y(_05261_),
    .B1(net448),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(net449),
    .A1(_10234_));
 sg13g2_buf_1 _22890_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05262_));
 sg13g2_a22oi_1 _22891_ (.Y(_05263_),
    .B1(_05019_),
    .B2(\cpu.intr.r_clock_cmp[30] ),
    .A2(net384),
    .A1(_05262_));
 sg13g2_a22oi_1 _22892_ (.Y(_05264_),
    .B1(net381),
    .B2(\cpu.intr.r_timer_count[14] ),
    .A2(net485),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_or2_1 _22893_ (.X(_05265_),
    .B(_05264_),
    .A(net613));
 sg13g2_nand3_1 _22894_ (.B(_05263_),
    .C(_05265_),
    .A(_05261_),
    .Y(_05266_));
 sg13g2_a221oi_1 _22895_ (.B2(_05014_),
    .C1(net850),
    .B1(_05266_),
    .A1(net577),
    .Y(_05267_),
    .A2(_05260_));
 sg13g2_nor3_1 _22896_ (.A(net82),
    .B(_05152_),
    .C(_05267_),
    .Y(_05268_));
 sg13g2_and2_1 _22897_ (.A(net598),
    .B(_04821_),
    .X(_05269_));
 sg13g2_nor3_1 _22898_ (.A(net85),
    .B(_05268_),
    .C(_05269_),
    .Y(_05270_));
 sg13g2_a221oi_1 _22899_ (.B2(net73),
    .C1(_05270_),
    .B1(_05245_),
    .A1(_04416_),
    .Y(_01038_),
    .A2(_04818_));
 sg13g2_o21ai_1 _22900_ (.B1(net196),
    .Y(_05271_),
    .A1(_11601_),
    .A2(_04452_));
 sg13g2_o21ai_1 _22901_ (.B1(_05271_),
    .Y(_05272_),
    .A1(_08474_),
    .A2(net196));
 sg13g2_nand2_1 _22902_ (.Y(_05273_),
    .A(net85),
    .B(_05272_));
 sg13g2_nor2_1 _22903_ (.A(_04449_),
    .B(_05273_),
    .Y(_05274_));
 sg13g2_a22oi_1 _22904_ (.Y(_05275_),
    .B1(net448),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net449),
    .A1(_10241_));
 sg13g2_buf_1 _22905_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05276_));
 sg13g2_a22oi_1 _22906_ (.Y(_05277_),
    .B1(_05019_),
    .B2(\cpu.intr.r_clock_cmp[31] ),
    .A2(_10156_),
    .A1(_05276_));
 sg13g2_a22oi_1 _22907_ (.Y(_05278_),
    .B1(_04894_),
    .B2(\cpu.intr.r_timer_count[15] ),
    .A2(net485),
    .A1(\cpu.intr.r_timer_reload[15] ));
 sg13g2_or2_1 _22908_ (.X(_05279_),
    .B(_05278_),
    .A(net613));
 sg13g2_nand3_1 _22909_ (.B(_05277_),
    .C(_05279_),
    .A(_05275_),
    .Y(_05280_));
 sg13g2_o21ai_1 _22910_ (.B1(_05078_),
    .Y(_05281_),
    .A1(net611),
    .A2(_05071_));
 sg13g2_a22oi_1 _22911_ (.Y(_05282_),
    .B1(_05281_),
    .B2(_05153_),
    .A2(_05280_),
    .A1(_05014_));
 sg13g2_o21ai_1 _22912_ (.B1(_05133_),
    .Y(_05283_),
    .A1(net850),
    .A2(_05282_));
 sg13g2_nand2_1 _22913_ (.Y(_05284_),
    .A(_10749_),
    .B(net81));
 sg13g2_o21ai_1 _22914_ (.B1(_05284_),
    .Y(_05285_),
    .A1(net82),
    .A2(_05283_));
 sg13g2_nand3_1 _22915_ (.B(_04817_),
    .C(_05272_),
    .A(net80),
    .Y(_05286_));
 sg13g2_o21ai_1 _22916_ (.B1(_05286_),
    .Y(_05287_),
    .A1(_11612_),
    .A2(_05285_));
 sg13g2_a21o_1 _22917_ (.A2(_05274_),
    .A1(_04448_),
    .B1(_05287_),
    .X(_01039_));
 sg13g2_mux2_1 _22918_ (.A0(_00200_),
    .A1(_04211_),
    .S(net579),
    .X(_05288_));
 sg13g2_nor2_1 _22919_ (.A(net1077),
    .B(net176),
    .Y(_05289_));
 sg13g2_a21oi_1 _22920_ (.A1(net176),
    .A2(_05288_),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_buf_1 _22921_ (.A(net80),
    .X(_05291_));
 sg13g2_buf_1 _22922_ (.A(net81),
    .X(_05292_));
 sg13g2_buf_1 _22923_ (.A(net1119),
    .X(_05293_));
 sg13g2_a22oi_1 _22924_ (.Y(_05294_),
    .B1(_12534_),
    .B2(\cpu.dcache.r_data[3][25] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_o21ai_1 _22925_ (.B1(_05294_),
    .Y(_05295_),
    .A1(_00092_),
    .A2(_09516_));
 sg13g2_a221oi_1 _22926_ (.B2(\cpu.dcache.r_data[2][25] ),
    .C1(_05295_),
    .B1(_04961_),
    .A1(\cpu.dcache.r_data[1][25] ),
    .Y(_05296_),
    .A2(_05030_));
 sg13g2_mux2_1 _22927_ (.A0(\cpu.dcache.r_data[4][25] ),
    .A1(\cpu.dcache.r_data[6][25] ),
    .S(_09222_),
    .X(_05297_));
 sg13g2_a22oi_1 _22928_ (.Y(_05298_),
    .B1(_05297_),
    .B2(_03785_),
    .A2(_09805_),
    .A1(\cpu.dcache.r_data[5][25] ));
 sg13g2_nand2b_1 _22929_ (.Y(_05299_),
    .B(_12001_),
    .A_N(_05298_));
 sg13g2_and2_1 _22930_ (.A(_05296_),
    .B(_05299_),
    .X(_05300_));
 sg13g2_buf_1 _22931_ (.A(_05300_),
    .X(_05301_));
 sg13g2_nand2_1 _22932_ (.Y(_05302_),
    .A(\cpu.dcache.r_data[2][9] ),
    .B(net499));
 sg13g2_o21ai_1 _22933_ (.B1(_05302_),
    .Y(_05303_),
    .A1(_00093_),
    .A2(net616));
 sg13g2_a221oi_1 _22934_ (.B2(\cpu.dcache.r_data[4][9] ),
    .C1(_05303_),
    .B1(_12664_),
    .A1(\cpu.dcache.r_data[5][9] ),
    .Y(_05304_),
    .A2(_04882_));
 sg13g2_a22oi_1 _22935_ (.Y(_05305_),
    .B1(_04891_),
    .B2(\cpu.dcache.r_data[6][9] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][9] ));
 sg13g2_a22oi_1 _22936_ (.Y(_05306_),
    .B1(_04959_),
    .B2(\cpu.dcache.r_data[3][9] ),
    .A2(_05030_),
    .A1(\cpu.dcache.r_data[1][9] ));
 sg13g2_and2_1 _22937_ (.A(_05305_),
    .B(_05306_),
    .X(_05307_));
 sg13g2_a21o_1 _22938_ (.A2(_05307_),
    .A1(_05304_),
    .B1(net681),
    .X(_05308_));
 sg13g2_o21ai_1 _22939_ (.B1(_05308_),
    .Y(_05309_),
    .A1(net983),
    .A2(_05301_));
 sg13g2_nand2_1 _22940_ (.Y(_05310_),
    .A(\cpu.dcache.r_data[4][1] ),
    .B(net424));
 sg13g2_a22oi_1 _22941_ (.Y(_05311_),
    .B1(net409),
    .B2(\cpu.dcache.r_data[1][1] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[6][1] ));
 sg13g2_a22oi_1 _22942_ (.Y(_05312_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][1] ),
    .A2(net473),
    .A1(\cpu.dcache.r_data[3][1] ));
 sg13g2_a22oi_1 _22943_ (.Y(_05313_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][1] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][1] ));
 sg13g2_nand4_1 _22944_ (.B(_05311_),
    .C(_05312_),
    .A(_05310_),
    .Y(_05314_),
    .D(_05313_));
 sg13g2_mux2_1 _22945_ (.A0(\cpu.dcache.r_data[0][1] ),
    .A1(_05314_),
    .S(net616),
    .X(_05315_));
 sg13g2_inv_1 _22946_ (.Y(_05316_),
    .A(_00091_));
 sg13g2_a22oi_1 _22947_ (.Y(_05317_),
    .B1(_12665_),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net410),
    .A1(_05316_));
 sg13g2_a22oi_1 _22948_ (.Y(_05318_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][17] ),
    .A2(_12535_),
    .A1(\cpu.dcache.r_data[3][17] ));
 sg13g2_a22oi_1 _22949_ (.Y(_05319_),
    .B1(net414),
    .B2(\cpu.dcache.r_data[6][17] ),
    .A2(_10024_),
    .A1(\cpu.dcache.r_data[7][17] ));
 sg13g2_a22oi_1 _22950_ (.Y(_05320_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][17] ),
    .A2(_05031_),
    .A1(\cpu.dcache.r_data[1][17] ));
 sg13g2_nand4_1 _22951_ (.B(_05318_),
    .C(_05319_),
    .A(_05317_),
    .Y(_05321_),
    .D(_05320_));
 sg13g2_buf_1 _22952_ (.A(_05321_),
    .X(_05322_));
 sg13g2_a22oi_1 _22953_ (.Y(_05323_),
    .B1(_05322_),
    .B2(_04977_),
    .A2(_05315_),
    .A1(net983));
 sg13g2_nor2_1 _22954_ (.A(net650),
    .B(_05323_),
    .Y(_05324_));
 sg13g2_a21oi_1 _22955_ (.A1(net650),
    .A2(_05309_),
    .Y(_05325_),
    .B1(_05324_));
 sg13g2_mux2_1 _22956_ (.A0(_05315_),
    .A1(_05322_),
    .S(net613),
    .X(_05326_));
 sg13g2_nand2_1 _22957_ (.Y(_05327_),
    .A(net577),
    .B(_05326_));
 sg13g2_o21ai_1 _22958_ (.B1(_05327_),
    .Y(_05328_),
    .A1(net577),
    .A2(_05325_));
 sg13g2_nand2_1 _22959_ (.Y(_05329_),
    .A(_09264_),
    .B(_04854_));
 sg13g2_o21ai_1 _22960_ (.B1(_05329_),
    .Y(_05330_),
    .A1(_00098_),
    .A2(_05099_));
 sg13g2_nand2_1 _22961_ (.Y(_05331_),
    .A(net871),
    .B(net504));
 sg13g2_nor2_1 _22962_ (.A(net771),
    .B(_00096_),
    .Y(_05332_));
 sg13g2_buf_2 _22963_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05333_));
 sg13g2_nor2b_1 _22964_ (.A(net772),
    .B_N(_05333_),
    .Y(_05334_));
 sg13g2_o21ai_1 _22965_ (.B1(net505),
    .Y(_05335_),
    .A1(_05332_),
    .A2(_05334_));
 sg13g2_o21ai_1 _22966_ (.B1(_05335_),
    .Y(_05336_),
    .A1(_00097_),
    .A2(_05331_));
 sg13g2_nand2_1 _22967_ (.Y(_05337_),
    .A(net872),
    .B(_04908_));
 sg13g2_nand2b_1 _22968_ (.Y(_05338_),
    .B(_04872_),
    .A_N(_00100_));
 sg13g2_o21ai_1 _22969_ (.B1(_05338_),
    .Y(_05339_),
    .A1(_00099_),
    .A2(_05337_));
 sg13g2_nor3_1 _22970_ (.A(_05330_),
    .B(_05336_),
    .C(_05339_),
    .Y(_05340_));
 sg13g2_a21oi_1 _22971_ (.A1(_09264_),
    .A2(_04840_),
    .Y(_05341_),
    .B1(net455));
 sg13g2_nand2b_1 _22972_ (.Y(_05342_),
    .B(\cpu.gpio.r_enable_in[1] ),
    .A_N(_05341_));
 sg13g2_a21oi_1 _22973_ (.A1(_05340_),
    .A2(_05342_),
    .Y(_05343_),
    .B1(_04824_));
 sg13g2_inv_1 _22974_ (.Y(_05344_),
    .A(_00095_));
 sg13g2_buf_1 _22975_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05345_));
 sg13g2_a22oi_1 _22976_ (.Y(_05346_),
    .B1(_04931_),
    .B2(_05345_),
    .A2(_04917_),
    .A1(_05344_));
 sg13g2_mux2_1 _22977_ (.A0(_11991_),
    .A1(_11996_),
    .S(net871),
    .X(_05347_));
 sg13g2_a22oi_1 _22978_ (.Y(_05348_),
    .B1(_05347_),
    .B2(_04922_),
    .A2(_05112_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_or2_1 _22979_ (.X(_05349_),
    .B(_04934_),
    .A(_00094_));
 sg13g2_nand3_1 _22980_ (.B(_05348_),
    .C(_05349_),
    .A(_05346_),
    .Y(_05350_));
 sg13g2_a221oi_1 _22981_ (.B2(_09342_),
    .C1(_05350_),
    .B1(_04919_),
    .A1(_11992_),
    .Y(_05351_),
    .A2(_04868_));
 sg13g2_nor2_1 _22982_ (.A(_09232_),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_a22oi_1 _22983_ (.Y(_05353_),
    .B1(net411),
    .B2(\cpu.uart.r_div_value[9] ),
    .A2(net504),
    .A1(\cpu.uart.r_r_invert ));
 sg13g2_a22oi_1 _22984_ (.Y(_05354_),
    .B1(net412),
    .B2(\cpu.uart.r_div_value[1] ),
    .A2(net415),
    .A1(_09279_));
 sg13g2_nand2_1 _22985_ (.Y(_05355_),
    .A(_05353_),
    .B(_05354_));
 sg13g2_a21oi_1 _22986_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04943_),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_nor2_1 _22987_ (.A(_04941_),
    .B(_05356_),
    .Y(_05357_));
 sg13g2_a22oi_1 _22988_ (.Y(_05358_),
    .B1(net416),
    .B2(\cpu.intr.r_clock_cmp[17] ),
    .A2(net381),
    .A1(_09988_));
 sg13g2_inv_1 _22989_ (.Y(_05359_),
    .A(_05358_));
 sg13g2_a22oi_1 _22990_ (.Y(_05360_),
    .B1(net416),
    .B2(\cpu.intr.r_clock_cmp[1] ),
    .A2(net381),
    .A1(_09993_));
 sg13g2_buf_1 _22991_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05361_));
 sg13g2_nand2_1 _22992_ (.Y(_05362_),
    .A(net902),
    .B(\cpu.intr.r_timer_reload[17] ));
 sg13g2_nand2_1 _22993_ (.Y(_05363_),
    .A(net771),
    .B(\cpu.intr.r_timer_reload[1] ));
 sg13g2_a21oi_1 _22994_ (.A1(_05362_),
    .A2(_05363_),
    .Y(_05364_),
    .B1(_10097_));
 sg13g2_a221oi_1 _22995_ (.B2(_09274_),
    .C1(_05364_),
    .B1(net413),
    .A1(_05361_),
    .Y(_05365_),
    .A2(net426));
 sg13g2_o21ai_1 _22996_ (.B1(_05365_),
    .Y(_05366_),
    .A1(net648),
    .A2(_05360_));
 sg13g2_a221oi_1 _22997_ (.B2(net648),
    .C1(_05366_),
    .B1(_05359_),
    .A1(_10161_),
    .Y(_05367_),
    .A2(net449));
 sg13g2_a21oi_1 _22998_ (.A1(_09274_),
    .A2(_04900_),
    .Y(_05368_),
    .B1(net415));
 sg13g2_nand2b_1 _22999_ (.Y(_05369_),
    .B(\cpu.intr.r_enable[1] ),
    .A_N(_05368_));
 sg13g2_a21oi_1 _23000_ (.A1(_05367_),
    .A2(_05369_),
    .Y(_05370_),
    .B1(net679));
 sg13g2_nor4_1 _23001_ (.A(_05343_),
    .B(_05352_),
    .C(_05357_),
    .D(_05370_),
    .Y(_05371_));
 sg13g2_nand2_1 _23002_ (.Y(_05372_),
    .A(net1025),
    .B(_05371_));
 sg13g2_o21ai_1 _23003_ (.B1(_05372_),
    .Y(_05373_),
    .A1(net846),
    .A2(_05328_));
 sg13g2_nand2_1 _23004_ (.Y(_05374_),
    .A(net543),
    .B(net82));
 sg13g2_o21ai_1 _23005_ (.B1(_05374_),
    .Y(_05375_),
    .A1(_05292_),
    .A2(_05373_));
 sg13g2_nor2_1 _23006_ (.A(net72),
    .B(_05375_),
    .Y(_05376_));
 sg13g2_a21oi_1 _23007_ (.A1(net73),
    .A2(_05290_),
    .Y(_01040_),
    .B1(_05376_));
 sg13g2_buf_1 _23008_ (.A(net83),
    .X(_05377_));
 sg13g2_a22oi_1 _23009_ (.Y(_05378_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][2] ),
    .A2(net499),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_a22oi_1 _23010_ (.Y(_05379_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[5][2] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][2] ));
 sg13g2_nand2_1 _23011_ (.Y(_05380_),
    .A(_05378_),
    .B(_05379_));
 sg13g2_a221oi_1 _23012_ (.B2(\cpu.dcache.r_data[3][2] ),
    .C1(_05380_),
    .B1(net500),
    .A1(\cpu.dcache.r_data[6][2] ),
    .Y(_05381_),
    .A2(net453));
 sg13g2_nor2_1 _23013_ (.A(\cpu.dcache.r_data[0][2] ),
    .B(_04851_),
    .Y(_05382_));
 sg13g2_a21oi_1 _23014_ (.A1(_04851_),
    .A2(_05381_),
    .Y(_05383_),
    .B1(_05382_));
 sg13g2_nand3b_1 _23015_ (.B(net409),
    .C(_05381_),
    .Y(_05384_),
    .A_N(\cpu.dcache.r_data[1][2] ));
 sg13g2_o21ai_1 _23016_ (.B1(_05384_),
    .Y(_05385_),
    .A1(net409),
    .A2(_05383_));
 sg13g2_a22oi_1 _23017_ (.Y(_05386_),
    .B1(net499),
    .B2(\cpu.dcache.r_data[2][18] ),
    .A2(net502),
    .A1(\cpu.dcache.r_data[6][18] ));
 sg13g2_a22oi_1 _23018_ (.Y(_05387_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][18] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][18] ));
 sg13g2_a22oi_1 _23019_ (.Y(_05388_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[5][18] ),
    .A2(_10022_),
    .A1(\cpu.dcache.r_data[7][18] ));
 sg13g2_nand3_1 _23020_ (.B(_05387_),
    .C(_05388_),
    .A(_05386_),
    .Y(_05389_));
 sg13g2_nand2_1 _23021_ (.Y(_05390_),
    .A(_00101_),
    .B(net912));
 sg13g2_o21ai_1 _23022_ (.B1(_05390_),
    .Y(_05391_),
    .A1(_09435_),
    .A2(_05389_));
 sg13g2_nor3_1 _23023_ (.A(\cpu.dcache.r_data[1][18] ),
    .B(net745),
    .C(_05389_),
    .Y(_05392_));
 sg13g2_a21o_1 _23024_ (.A2(_05391_),
    .A1(net745),
    .B1(_05392_),
    .X(_05393_));
 sg13g2_nand2b_1 _23025_ (.Y(_05394_),
    .B(net648),
    .A_N(_05393_));
 sg13g2_o21ai_1 _23026_ (.B1(_05394_),
    .Y(_05395_),
    .A1(net543),
    .A2(_05385_));
 sg13g2_mux2_1 _23027_ (.A0(_05394_),
    .A1(_05385_),
    .S(net983),
    .X(_05396_));
 sg13g2_a221oi_1 _23028_ (.B2(_04992_),
    .C1(net649),
    .B1(_05041_),
    .A1(net611),
    .Y(_05397_),
    .A2(_05034_));
 sg13g2_a21oi_1 _23029_ (.A1(net649),
    .A2(_05396_),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_mux2_1 _23030_ (.A0(_05395_),
    .A1(_05398_),
    .S(_05046_),
    .X(_05399_));
 sg13g2_nor2_1 _23031_ (.A(net678),
    .B(_00106_),
    .Y(_05400_));
 sg13g2_buf_1 _23032_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05401_));
 sg13g2_nor2b_1 _23033_ (.A(net681),
    .B_N(_05401_),
    .Y(_05402_));
 sg13g2_o21ai_1 _23034_ (.B1(net505),
    .Y(_05403_),
    .A1(_05400_),
    .A2(_05402_));
 sg13g2_o21ai_1 _23035_ (.B1(_05403_),
    .Y(_05404_),
    .A1(_00108_),
    .A2(_05099_));
 sg13g2_nand2_1 _23036_ (.Y(_05405_),
    .A(_09260_),
    .B(_04854_));
 sg13g2_o21ai_1 _23037_ (.B1(_05405_),
    .Y(_05406_),
    .A1(_00107_),
    .A2(_05331_));
 sg13g2_nand2b_1 _23038_ (.Y(_05407_),
    .B(_04872_),
    .A_N(_00110_));
 sg13g2_o21ai_1 _23039_ (.B1(_05407_),
    .Y(_05408_),
    .A1(_00109_),
    .A2(_05337_));
 sg13g2_a21oi_1 _23040_ (.A1(_09260_),
    .A2(_04840_),
    .Y(_05409_),
    .B1(net455));
 sg13g2_nor2b_1 _23041_ (.A(_05409_),
    .B_N(\cpu.gpio.r_enable_in[2] ),
    .Y(_05410_));
 sg13g2_nor4_1 _23042_ (.A(_05404_),
    .B(_05406_),
    .C(_05408_),
    .D(_05410_),
    .Y(_05411_));
 sg13g2_inv_1 _23043_ (.Y(_05412_),
    .A(_00105_));
 sg13g2_buf_1 _23044_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05413_));
 sg13g2_nand2_1 _23045_ (.Y(_05414_),
    .A(net871),
    .B(_11985_));
 sg13g2_o21ai_1 _23046_ (.B1(_05414_),
    .Y(_05415_),
    .A1(net871),
    .A2(_11981_));
 sg13g2_a22oi_1 _23047_ (.Y(_05416_),
    .B1(_05415_),
    .B2(_04922_),
    .A2(_05112_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _23048_ (.B1(_05416_),
    .Y(_05417_),
    .A1(_00104_),
    .A2(_04934_));
 sg13g2_a221oi_1 _23049_ (.B2(_05413_),
    .C1(_05417_),
    .B1(_04931_),
    .A1(_05412_),
    .Y(_05418_),
    .A2(_04917_));
 sg13g2_o21ai_1 _23050_ (.B1(_05418_),
    .Y(_05419_),
    .A1(_00285_),
    .A2(_05337_));
 sg13g2_a21o_1 _23051_ (.A2(_04919_),
    .A1(_09346_),
    .B1(_05419_),
    .X(_05420_));
 sg13g2_nand2_1 _23052_ (.Y(_05421_),
    .A(_10166_),
    .B(net449));
 sg13g2_a22oi_1 _23053_ (.Y(_05422_),
    .B1(net448),
    .B2(\cpu.intr.r_clock_cmp[2] ),
    .A2(_04908_),
    .A1(_09995_));
 sg13g2_a22oi_1 _23054_ (.Y(_05423_),
    .B1(net416),
    .B2(\cpu.intr.r_clock_cmp[18] ),
    .A2(net381),
    .A1(_09987_));
 sg13g2_nand2b_1 _23055_ (.Y(_05424_),
    .B(net681),
    .A_N(_05423_));
 sg13g2_mux2_1 _23056_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .S(net772),
    .X(_05425_));
 sg13g2_a22oi_1 _23057_ (.Y(_05426_),
    .B1(_05425_),
    .B2(net485),
    .A2(net415),
    .A1(_09271_));
 sg13g2_buf_2 _23058_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05427_));
 sg13g2_a22oi_1 _23059_ (.Y(_05428_),
    .B1(net413),
    .B2(_09270_),
    .A2(net426),
    .A1(_05427_));
 sg13g2_and3_1 _23060_ (.X(_05429_),
    .A(_05424_),
    .B(_05426_),
    .C(_05428_));
 sg13g2_nand3_1 _23061_ (.B(_09271_),
    .C(_04900_),
    .A(_09270_),
    .Y(_05430_));
 sg13g2_nand4_1 _23062_ (.B(_05422_),
    .C(_05429_),
    .A(_05421_),
    .Y(_05431_),
    .D(_05430_));
 sg13g2_and2_1 _23063_ (.A(\cpu.uart.r_in[2] ),
    .B(_04943_),
    .X(_05432_));
 sg13g2_a221oi_1 _23064_ (.B2(_09976_),
    .C1(_05432_),
    .B1(net411),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05433_),
    .A2(net412));
 sg13g2_o21ai_1 _23065_ (.B1(net1025),
    .Y(_05434_),
    .A1(_04941_),
    .A2(_05433_));
 sg13g2_a221oi_1 _23066_ (.B2(_04878_),
    .C1(_05434_),
    .B1(_05431_),
    .A1(_04939_),
    .Y(_05435_),
    .A2(_05420_));
 sg13g2_o21ai_1 _23067_ (.B1(_05435_),
    .Y(_05436_),
    .A1(_04824_),
    .A2(_05411_));
 sg13g2_o21ai_1 _23068_ (.B1(_05436_),
    .Y(_05437_),
    .A1(_04822_),
    .A2(_05399_));
 sg13g2_nor2_1 _23069_ (.A(net71),
    .B(_05437_),
    .Y(_05438_));
 sg13g2_a21oi_1 _23070_ (.A1(net590),
    .A2(net71),
    .Y(_05439_),
    .B1(_05438_));
 sg13g2_o21ai_1 _23071_ (.B1(net196),
    .Y(_05440_),
    .A1(net696),
    .A2(_05140_));
 sg13g2_nand2_1 _23072_ (.Y(_05441_),
    .A(_05145_),
    .B(_04486_));
 sg13g2_o21ai_1 _23073_ (.B1(_05441_),
    .Y(_05442_),
    .A1(net578),
    .A2(_04484_));
 sg13g2_a221oi_1 _23074_ (.B2(net176),
    .C1(net83),
    .B1(_05442_),
    .A1(net812),
    .Y(_05443_),
    .A2(_05440_));
 sg13g2_a21oi_1 _23075_ (.A1(net70),
    .A2(_05439_),
    .Y(_01041_),
    .B1(_05443_));
 sg13g2_o21ai_1 _23076_ (.B1(_05167_),
    .Y(_05444_),
    .A1(net983),
    .A2(_05160_));
 sg13g2_nand2_1 _23077_ (.Y(_05445_),
    .A(\cpu.dcache.r_data[4][3] ),
    .B(net471));
 sg13g2_a22oi_1 _23078_ (.Y(_05446_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][3] ),
    .A2(net498),
    .A1(\cpu.dcache.r_data[1][3] ));
 sg13g2_a22oi_1 _23079_ (.Y(_05447_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][3] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_a22oi_1 _23080_ (.Y(_05448_),
    .B1(net500),
    .B2(\cpu.dcache.r_data[3][3] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][3] ));
 sg13g2_nand4_1 _23081_ (.B(_05446_),
    .C(_05447_),
    .A(_05445_),
    .Y(_05449_),
    .D(_05448_));
 sg13g2_mux2_1 _23082_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(_05449_),
    .S(net616),
    .X(_05450_));
 sg13g2_a22oi_1 _23083_ (.Y(_05451_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][19] ));
 sg13g2_inv_1 _23084_ (.Y(_05452_),
    .A(_00111_));
 sg13g2_a22oi_1 _23085_ (.Y(_05453_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][19] ),
    .A2(net452),
    .A1(_05452_));
 sg13g2_a22oi_1 _23086_ (.Y(_05454_),
    .B1(net450),
    .B2(\cpu.dcache.r_data[1][19] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][19] ));
 sg13g2_a22oi_1 _23087_ (.Y(_05455_),
    .B1(net471),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net500),
    .A1(\cpu.dcache.r_data[3][19] ));
 sg13g2_nand4_1 _23088_ (.B(_05453_),
    .C(_05454_),
    .A(_05451_),
    .Y(_05456_),
    .D(_05455_));
 sg13g2_buf_1 _23089_ (.A(_05456_),
    .X(_05457_));
 sg13g2_a22oi_1 _23090_ (.Y(_05458_),
    .B1(_05457_),
    .B2(_04977_),
    .A2(_05450_),
    .A1(net983));
 sg13g2_nor2_1 _23091_ (.A(net650),
    .B(_05458_),
    .Y(_05459_));
 sg13g2_a21oi_1 _23092_ (.A1(net650),
    .A2(_05444_),
    .Y(_05460_),
    .B1(_05459_));
 sg13g2_mux2_1 _23093_ (.A0(_05450_),
    .A1(_05457_),
    .S(_10021_),
    .X(_05461_));
 sg13g2_nand2_1 _23094_ (.Y(_05462_),
    .A(net577),
    .B(_05461_));
 sg13g2_o21ai_1 _23095_ (.B1(_05462_),
    .Y(_05463_),
    .A1(net577),
    .A2(_05460_));
 sg13g2_a21o_1 _23096_ (.A2(_04840_),
    .A1(_09245_),
    .B1(_04846_),
    .X(_05464_));
 sg13g2_inv_1 _23097_ (.Y(_05465_),
    .A(_00119_));
 sg13g2_a22oi_1 _23098_ (.Y(_05466_),
    .B1(_05086_),
    .B2(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A2(_05019_),
    .A1(_05465_));
 sg13g2_inv_1 _23099_ (.Y(_05467_),
    .A(_00118_));
 sg13g2_nor2_1 _23100_ (.A(net900),
    .B(_00116_),
    .Y(_05468_));
 sg13g2_buf_1 _23101_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05469_));
 sg13g2_nor2b_1 _23102_ (.A(net902),
    .B_N(_05469_),
    .Y(_05470_));
 sg13g2_o21ai_1 _23103_ (.B1(net505),
    .Y(_05471_),
    .A1(_05468_),
    .A2(_05470_));
 sg13g2_o21ai_1 _23104_ (.B1(_05471_),
    .Y(_05472_),
    .A1(_00117_),
    .A2(_05331_));
 sg13g2_a221oi_1 _23105_ (.B2(_09245_),
    .C1(_05472_),
    .B1(_04854_),
    .A1(_05467_),
    .Y(_05473_),
    .A2(_04852_));
 sg13g2_o21ai_1 _23106_ (.B1(_05473_),
    .Y(_05474_),
    .A1(_04825_),
    .A2(_05466_));
 sg13g2_a21oi_1 _23107_ (.A1(\cpu.gpio.r_enable_in[3] ),
    .A2(_05464_),
    .Y(_05475_),
    .B1(_05474_));
 sg13g2_inv_1 _23108_ (.Y(_05476_),
    .A(_00115_));
 sg13g2_buf_1 _23109_ (.A(_04917_),
    .X(_05477_));
 sg13g2_buf_1 _23110_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05478_));
 sg13g2_a22oi_1 _23111_ (.Y(_05479_),
    .B1(_04931_),
    .B2(_05478_),
    .A2(net407),
    .A1(_05476_));
 sg13g2_nor2_1 _23112_ (.A(_00114_),
    .B(_04934_),
    .Y(_05480_));
 sg13g2_a21oi_1 _23113_ (.A1(\cpu.spi.r_timeout[3] ),
    .A2(_05112_),
    .Y(_05481_),
    .B1(_05480_));
 sg13g2_nand2_1 _23114_ (.Y(_05482_),
    .A(_09340_),
    .B(_04919_));
 sg13g2_and4_1 _23115_ (.A(net1071),
    .B(_05479_),
    .C(_05481_),
    .D(_05482_),
    .X(_05483_));
 sg13g2_a21oi_1 _23116_ (.A1(_10619_),
    .A2(_05475_),
    .Y(_05484_),
    .B1(_05483_));
 sg13g2_nand2_1 _23117_ (.Y(_05485_),
    .A(_10171_),
    .B(net449));
 sg13g2_buf_1 _23118_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05486_));
 sg13g2_a22oi_1 _23119_ (.Y(_05487_),
    .B1(net413),
    .B2(_09272_),
    .A2(net384),
    .A1(_05486_));
 sg13g2_a21oi_1 _23120_ (.A1(_09272_),
    .A2(_04900_),
    .Y(_05488_),
    .B1(net415));
 sg13g2_nand2b_1 _23121_ (.Y(_05489_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05488_));
 sg13g2_mux2_1 _23122_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(\cpu.intr.r_timer_reload[3] ),
    .S(net695),
    .X(_05490_));
 sg13g2_a22oi_1 _23123_ (.Y(_05491_),
    .B1(_05490_),
    .B2(net694),
    .A2(net775),
    .A1(\cpu.intr.r_timer_count[3] ));
 sg13g2_mux2_1 _23124_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .S(net695),
    .X(_05492_));
 sg13g2_a221oi_1 _23125_ (.B2(net694),
    .C1(net678),
    .B1(_05492_),
    .A1(_09986_),
    .Y(_05493_),
    .A2(net775));
 sg13g2_a21oi_1 _23126_ (.A1(net678),
    .A2(_05491_),
    .Y(_05494_),
    .B1(_05493_));
 sg13g2_nand2_1 _23127_ (.Y(_05495_),
    .A(net748),
    .B(_05494_));
 sg13g2_nand4_1 _23128_ (.B(_05487_),
    .C(_05489_),
    .A(_05485_),
    .Y(_05496_),
    .D(_05495_));
 sg13g2_nand2_1 _23129_ (.Y(_05497_),
    .A(\cpu.uart.r_div_value[11] ),
    .B(net411));
 sg13g2_a22oi_1 _23130_ (.Y(_05498_),
    .B1(_04943_),
    .B2(\cpu.uart.r_in[3] ),
    .A2(net412),
    .A1(\cpu.uart.r_div_value[3] ));
 sg13g2_a21oi_1 _23131_ (.A1(_05497_),
    .A2(_05498_),
    .Y(_05499_),
    .B1(_04941_));
 sg13g2_a221oi_1 _23132_ (.B2(_04878_),
    .C1(_05499_),
    .B1(_05496_),
    .A1(_09231_),
    .Y(_05500_),
    .A2(_05484_));
 sg13g2_nand2_1 _23133_ (.Y(_05501_),
    .A(net846),
    .B(_05500_));
 sg13g2_o21ai_1 _23134_ (.B1(_05501_),
    .Y(_05502_),
    .A1(net846),
    .A2(_05463_));
 sg13g2_nor2_1 _23135_ (.A(net71),
    .B(_05502_),
    .Y(_05503_));
 sg13g2_a21oi_1 _23136_ (.A1(_03534_),
    .A2(net71),
    .Y(_05504_),
    .B1(_05503_));
 sg13g2_a21o_1 _23137_ (.A2(_04516_),
    .A1(_05145_),
    .B1(net177),
    .X(_05505_));
 sg13g2_nand2_1 _23138_ (.Y(_05506_),
    .A(_05145_),
    .B(_04518_));
 sg13g2_o21ai_1 _23139_ (.B1(_05506_),
    .Y(_05507_),
    .A1(_05146_),
    .A2(_04515_));
 sg13g2_a221oi_1 _23140_ (.B2(net176),
    .C1(net83),
    .B1(_05507_),
    .A1(net698),
    .Y(_05508_),
    .A2(_05505_));
 sg13g2_a21oi_1 _23141_ (.A1(net70),
    .A2(_05504_),
    .Y(_01042_),
    .B1(_05508_));
 sg13g2_o21ai_1 _23142_ (.B1(net650),
    .Y(_05509_),
    .A1(_05045_),
    .A2(_05205_));
 sg13g2_inv_1 _23143_ (.Y(_05510_),
    .A(_00121_));
 sg13g2_a22oi_1 _23144_ (.Y(_05511_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[4][4] ),
    .A2(net410),
    .A1(_05510_));
 sg13g2_a22oi_1 _23145_ (.Y(_05512_),
    .B1(_04883_),
    .B2(\cpu.dcache.r_data[5][4] ),
    .A2(net473),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_a22oi_1 _23146_ (.Y(_05513_),
    .B1(_04894_),
    .B2(\cpu.dcache.r_data[6][4] ),
    .A2(_10025_),
    .A1(\cpu.dcache.r_data[7][4] ));
 sg13g2_a22oi_1 _23147_ (.Y(_05514_),
    .B1(net408),
    .B2(\cpu.dcache.r_data[2][4] ),
    .A2(net409),
    .A1(\cpu.dcache.r_data[1][4] ));
 sg13g2_and4_1 _23148_ (.A(_05511_),
    .B(_05512_),
    .C(_05513_),
    .D(_05514_),
    .X(_05515_));
 sg13g2_buf_1 _23149_ (.A(_05515_),
    .X(_05516_));
 sg13g2_nand2_1 _23150_ (.Y(_05517_),
    .A(net983),
    .B(net649));
 sg13g2_nor2_1 _23151_ (.A(_05516_),
    .B(_05517_),
    .Y(_05518_));
 sg13g2_nand2_1 _23152_ (.Y(_05519_),
    .A(net650),
    .B(_05197_));
 sg13g2_inv_1 _23153_ (.Y(_05520_),
    .A(_00122_));
 sg13g2_a22oi_1 _23154_ (.Y(_05521_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][20] ),
    .A2(net501),
    .A1(_05520_));
 sg13g2_a22oi_1 _23155_ (.Y(_05522_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][20] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][20] ));
 sg13g2_a22oi_1 _23156_ (.Y(_05523_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[6][20] ),
    .A2(net680),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_a22oi_1 _23157_ (.Y(_05524_),
    .B1(net499),
    .B2(\cpu.dcache.r_data[2][20] ),
    .A2(net498),
    .A1(\cpu.dcache.r_data[1][20] ));
 sg13g2_nand4_1 _23158_ (.B(_05522_),
    .C(_05523_),
    .A(_05521_),
    .Y(_05525_),
    .D(_05524_));
 sg13g2_buf_1 _23159_ (.A(_05525_),
    .X(_05526_));
 sg13g2_nand3_1 _23160_ (.B(net649),
    .C(_05526_),
    .A(_10021_),
    .Y(_05527_));
 sg13g2_a21oi_1 _23161_ (.A1(_05519_),
    .A2(_05527_),
    .Y(_05528_),
    .B1(net983));
 sg13g2_nor2_1 _23162_ (.A(_05518_),
    .B(_05528_),
    .Y(_05529_));
 sg13g2_nand2_1 _23163_ (.Y(_05530_),
    .A(net611),
    .B(_05516_));
 sg13g2_o21ai_1 _23164_ (.B1(_05530_),
    .Y(_05531_),
    .A1(net544),
    .A2(_05526_));
 sg13g2_a22oi_1 _23165_ (.Y(_05532_),
    .B1(_05531_),
    .B2(net577),
    .A2(_05529_),
    .A1(_05509_));
 sg13g2_nand3_1 _23166_ (.B(_09262_),
    .C(_04840_),
    .A(_09261_),
    .Y(_05533_));
 sg13g2_nand2_1 _23167_ (.Y(_05534_),
    .A(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .B(_10155_));
 sg13g2_a22oi_1 _23168_ (.Y(_05535_),
    .B1(_05184_),
    .B2(net7),
    .A2(_05086_),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_a21oi_1 _23169_ (.A1(_05534_),
    .A2(_05535_),
    .Y(_05536_),
    .B1(_04825_));
 sg13g2_and2_1 _23170_ (.A(_09253_),
    .B(net1139),
    .X(_05537_));
 sg13g2_a21oi_1 _23171_ (.A1(_04902_),
    .A2(_05537_),
    .Y(_05538_),
    .B1(_04917_));
 sg13g2_nand2b_1 _23172_ (.Y(_05539_),
    .B(\cpu.gpio.r_enable_io[4] ),
    .A_N(_05538_));
 sg13g2_buf_2 _23173_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05540_));
 sg13g2_buf_2 _23174_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05541_));
 sg13g2_mux2_1 _23175_ (.A0(_05540_),
    .A1(_05541_),
    .S(net902),
    .X(_05542_));
 sg13g2_and2_1 _23176_ (.A(net505),
    .B(_05542_),
    .X(_05543_));
 sg13g2_a221oi_1 _23177_ (.B2(_09261_),
    .C1(_05543_),
    .B1(net455),
    .A1(_09262_),
    .Y(_05544_),
    .A2(_04854_));
 sg13g2_buf_2 _23178_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05545_));
 sg13g2_a22oi_1 _23179_ (.Y(_05546_),
    .B1(net504),
    .B2(_05537_),
    .A2(_04852_),
    .A1(_05545_));
 sg13g2_buf_2 _23180_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05547_));
 sg13g2_buf_2 _23181_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05548_));
 sg13g2_buf_2 _23182_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05549_));
 sg13g2_a22oi_1 _23183_ (.Y(_05550_),
    .B1(_04902_),
    .B2(_05549_),
    .A2(net504),
    .A1(_05548_));
 sg13g2_inv_1 _23184_ (.Y(_05551_),
    .A(_05550_));
 sg13g2_a22oi_1 _23185_ (.Y(_05552_),
    .B1(_05551_),
    .B2(net871),
    .A2(_04872_),
    .A1(_05547_));
 sg13g2_nand4_1 _23186_ (.B(_05544_),
    .C(_05546_),
    .A(_05539_),
    .Y(_05553_),
    .D(_05552_));
 sg13g2_nor2_1 _23187_ (.A(_05536_),
    .B(_05553_),
    .Y(_05554_));
 sg13g2_a21oi_1 _23188_ (.A1(_05533_),
    .A2(_05554_),
    .Y(_05555_),
    .B1(_04824_));
 sg13g2_a22oi_1 _23189_ (.Y(_05556_),
    .B1(_04943_),
    .B2(\cpu.uart.r_in[4] ),
    .A2(net412),
    .A1(\cpu.uart.r_div_value[4] ));
 sg13g2_nor2_1 _23190_ (.A(_04941_),
    .B(_05556_),
    .Y(_05557_));
 sg13g2_buf_2 _23191_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05558_));
 sg13g2_mux2_1 _23192_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net902),
    .X(_05559_));
 sg13g2_mux2_1 _23193_ (.A0(\cpu.intr.r_timer_count[4] ),
    .A1(_10011_),
    .S(net902),
    .X(_05560_));
 sg13g2_a22oi_1 _23194_ (.Y(_05561_),
    .B1(_05560_),
    .B2(net381),
    .A2(_05559_),
    .A1(net485));
 sg13g2_mux2_1 _23195_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(\cpu.intr.r_clock_cmp[20] ),
    .S(_10018_),
    .X(_05562_));
 sg13g2_a22oi_1 _23196_ (.Y(_05563_),
    .B1(_05562_),
    .B2(net416),
    .A2(_04887_),
    .A1(_09244_));
 sg13g2_nand2_1 _23197_ (.Y(_05564_),
    .A(_05561_),
    .B(_05563_));
 sg13g2_a221oi_1 _23198_ (.B2(_10177_),
    .C1(_05564_),
    .B1(net449),
    .A1(_05558_),
    .Y(_05565_),
    .A2(net426));
 sg13g2_o21ai_1 _23199_ (.B1(_09269_),
    .Y(_05566_),
    .A1(net413),
    .A2(_04900_));
 sg13g2_a221oi_1 _23200_ (.B2(_05566_),
    .C1(net679),
    .B1(_05565_),
    .A1(_10381_),
    .Y(_05567_),
    .A2(_04900_));
 sg13g2_inv_1 _23201_ (.Y(_05568_),
    .A(_00126_));
 sg13g2_buf_1 _23202_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05569_));
 sg13g2_nand2_1 _23203_ (.Y(_05570_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(_05112_));
 sg13g2_o21ai_1 _23204_ (.B1(_05570_),
    .Y(_05571_),
    .A1(_00125_),
    .A2(_04934_));
 sg13g2_a221oi_1 _23205_ (.B2(_05569_),
    .C1(_05571_),
    .B1(_04931_),
    .A1(_05568_),
    .Y(_05572_),
    .A2(net407));
 sg13g2_nand2_1 _23206_ (.Y(_05573_),
    .A(_09348_),
    .B(_04919_));
 sg13g2_a21oi_1 _23207_ (.A1(_05572_),
    .A2(_05573_),
    .Y(_05574_),
    .B1(_09232_));
 sg13g2_nor4_1 _23208_ (.A(_05555_),
    .B(_05557_),
    .C(_05567_),
    .D(_05574_),
    .Y(_05575_));
 sg13g2_nand2_1 _23209_ (.Y(_05576_),
    .A(net846),
    .B(_05575_));
 sg13g2_o21ai_1 _23210_ (.B1(_05576_),
    .Y(_05577_),
    .A1(net846),
    .A2(_05532_));
 sg13g2_nor2_1 _23211_ (.A(net71),
    .B(_05577_),
    .Y(_05578_));
 sg13g2_a21oi_1 _23212_ (.A1(net517),
    .A2(net71),
    .Y(_05579_),
    .B1(_05578_));
 sg13g2_and2_1 _23213_ (.A(net696),
    .B(net810),
    .X(_05580_));
 sg13g2_o21ai_1 _23214_ (.B1(net196),
    .Y(_05581_),
    .A1(_05140_),
    .A2(_05580_));
 sg13g2_nand2_1 _23215_ (.Y(_05582_),
    .A(_05145_),
    .B(_04554_));
 sg13g2_o21ai_1 _23216_ (.B1(_05582_),
    .Y(_05583_),
    .A1(_05146_),
    .A2(_04552_));
 sg13g2_a221oi_1 _23217_ (.B2(net176),
    .C1(net83),
    .B1(_05583_),
    .A1(net1150),
    .Y(_05584_),
    .A2(_05581_));
 sg13g2_a21oi_1 _23218_ (.A1(_05377_),
    .A2(_05579_),
    .Y(_01043_),
    .B1(_05584_));
 sg13g2_nand2_1 _23219_ (.Y(_05585_),
    .A(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .B(net384));
 sg13g2_a22oi_1 _23220_ (.Y(_05586_),
    .B1(net448),
    .B2(net8),
    .A2(_05183_),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_nand2_1 _23221_ (.Y(_05587_),
    .A(_05585_),
    .B(_05586_));
 sg13g2_a21o_1 _23222_ (.A2(_04840_),
    .A1(_09248_),
    .B1(net455),
    .X(_05588_));
 sg13g2_nor2_1 _23223_ (.A(_00136_),
    .B(_05099_),
    .Y(_05589_));
 sg13g2_a221oi_1 _23224_ (.B2(_09265_),
    .C1(_05589_),
    .B1(net407),
    .A1(_09248_),
    .Y(_05590_),
    .A2(_04854_));
 sg13g2_nand2b_1 _23225_ (.Y(_05591_),
    .B(_04872_),
    .A_N(_00138_));
 sg13g2_nand3_1 _23226_ (.B(_09266_),
    .C(net984),
    .A(_09265_),
    .Y(_05592_));
 sg13g2_o21ai_1 _23227_ (.B1(_05592_),
    .Y(_05593_),
    .A1(net872),
    .A2(_00137_));
 sg13g2_nand2_1 _23228_ (.Y(_05594_),
    .A(_04903_),
    .B(_05593_));
 sg13g2_nand2_1 _23229_ (.Y(_05595_),
    .A(_09266_),
    .B(net984));
 sg13g2_o21ai_1 _23230_ (.B1(_05595_),
    .Y(_05596_),
    .A1(net872),
    .A2(_00135_));
 sg13g2_buf_2 _23231_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05597_));
 sg13g2_nand2_1 _23232_ (.Y(_05598_),
    .A(net678),
    .B(_05597_));
 sg13g2_o21ai_1 _23233_ (.B1(_05598_),
    .Y(_05599_),
    .A1(net678),
    .A2(_00134_));
 sg13g2_a22oi_1 _23234_ (.Y(_05600_),
    .B1(_05599_),
    .B2(_04857_),
    .A2(_05596_),
    .A1(_04862_));
 sg13g2_nand4_1 _23235_ (.B(_05591_),
    .C(_05594_),
    .A(_05590_),
    .Y(_05601_),
    .D(_05600_));
 sg13g2_a221oi_1 _23236_ (.B2(\cpu.gpio.r_enable_in[5] ),
    .C1(_05601_),
    .B1(_05588_),
    .A1(net984),
    .Y(_05602_),
    .A2(_05587_));
 sg13g2_inv_1 _23237_ (.Y(_05603_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_nor2_1 _23238_ (.A(_10091_),
    .B(_05603_),
    .Y(_05604_));
 sg13g2_a21oi_1 _23239_ (.A1(net771),
    .A2(\cpu.intr.r_timer_reload[5] ),
    .Y(_05605_),
    .B1(_05604_));
 sg13g2_buf_2 _23240_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05606_));
 sg13g2_a22oi_1 _23241_ (.Y(_05607_),
    .B1(_04887_),
    .B2(_09276_),
    .A2(net426),
    .A1(_05606_));
 sg13g2_o21ai_1 _23242_ (.B1(_05607_),
    .Y(_05608_),
    .A1(_10097_),
    .A2(_05605_));
 sg13g2_a221oi_1 _23243_ (.B2(_10183_),
    .C1(_05608_),
    .B1(net449),
    .A1(\cpu.intr.r_timer_count[5] ),
    .Y(_05609_),
    .A2(_04908_));
 sg13g2_a22oi_1 _23244_ (.Y(_05610_),
    .B1(net416),
    .B2(\cpu.intr.r_clock_cmp[21] ),
    .A2(net381),
    .A1(_10012_));
 sg13g2_inv_1 _23245_ (.Y(_05611_),
    .A(_05610_));
 sg13g2_a22oi_1 _23246_ (.Y(_05612_),
    .B1(_05611_),
    .B2(net648),
    .A2(net448),
    .A1(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_a21oi_1 _23247_ (.A1(_09276_),
    .A2(_04900_),
    .Y(_05613_),
    .B1(net413));
 sg13g2_nand2b_1 _23248_ (.Y(_05614_),
    .B(_09275_),
    .A_N(_05613_));
 sg13g2_nand3_1 _23249_ (.B(_05612_),
    .C(_05614_),
    .A(_05609_),
    .Y(_05615_));
 sg13g2_inv_1 _23250_ (.Y(_05616_),
    .A(_00133_));
 sg13g2_buf_1 _23251_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05617_));
 sg13g2_a22oi_1 _23252_ (.Y(_05618_),
    .B1(_04931_),
    .B2(_05617_),
    .A2(net407),
    .A1(_05616_));
 sg13g2_nor2_1 _23253_ (.A(_00132_),
    .B(_04934_),
    .Y(_05619_));
 sg13g2_a21oi_1 _23254_ (.A1(\cpu.spi.r_timeout[5] ),
    .A2(_05112_),
    .Y(_05620_),
    .B1(_05619_));
 sg13g2_nand2_1 _23255_ (.Y(_05621_),
    .A(_09347_),
    .B(_04919_));
 sg13g2_nand3_1 _23256_ (.B(_05620_),
    .C(_05621_),
    .A(_05618_),
    .Y(_05622_));
 sg13g2_a22oi_1 _23257_ (.Y(_05623_),
    .B1(_04943_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net412),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_nor2_1 _23258_ (.A(_04941_),
    .B(_05623_),
    .Y(_05624_));
 sg13g2_a221oi_1 _23259_ (.B2(_04939_),
    .C1(_05624_),
    .B1(_05622_),
    .A1(_04878_),
    .Y(_05625_),
    .A2(_05615_));
 sg13g2_o21ai_1 _23260_ (.B1(_05625_),
    .Y(_05626_),
    .A1(_04824_),
    .A2(_05602_));
 sg13g2_nand2_1 _23261_ (.Y(_05627_),
    .A(\cpu.dcache.r_data[4][5] ),
    .B(net471));
 sg13g2_a22oi_1 _23262_ (.Y(_05628_),
    .B1(net450),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][5] ));
 sg13g2_a22oi_1 _23263_ (.Y(_05629_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][5] ),
    .A2(net500),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_a22oi_1 _23264_ (.Y(_05630_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][5] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][5] ));
 sg13g2_nand4_1 _23265_ (.B(_05628_),
    .C(_05629_),
    .A(_05627_),
    .Y(_05631_),
    .D(_05630_));
 sg13g2_nor2_1 _23266_ (.A(net410),
    .B(_05631_),
    .Y(_05632_));
 sg13g2_a21oi_1 _23267_ (.A1(_00128_),
    .A2(net410),
    .Y(_05633_),
    .B1(_05632_));
 sg13g2_a22oi_1 _23268_ (.Y(_05634_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[5][21] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][21] ));
 sg13g2_inv_1 _23269_ (.Y(_05635_),
    .A(_00129_));
 sg13g2_a22oi_1 _23270_ (.Y(_05636_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][21] ),
    .A2(net452),
    .A1(_05635_));
 sg13g2_a22oi_1 _23271_ (.Y(_05637_),
    .B1(net450),
    .B2(\cpu.dcache.r_data[1][21] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][21] ));
 sg13g2_a22oi_1 _23272_ (.Y(_05638_),
    .B1(net471),
    .B2(\cpu.dcache.r_data[4][21] ),
    .A2(net500),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_nand4_1 _23273_ (.B(_05636_),
    .C(_05637_),
    .A(_05634_),
    .Y(_05639_),
    .D(_05638_));
 sg13g2_nand2_1 _23274_ (.Y(_05640_),
    .A(_10020_),
    .B(_05639_));
 sg13g2_nor2_1 _23275_ (.A(net1119),
    .B(_05640_),
    .Y(_05641_));
 sg13g2_a21oi_1 _23276_ (.A1(net1119),
    .A2(_05633_),
    .Y(_05642_),
    .B1(_05641_));
 sg13g2_a221oi_1 _23277_ (.B2(_10093_),
    .C1(_04982_),
    .B1(_05229_),
    .A1(_04992_),
    .Y(_05643_),
    .A2(_05223_));
 sg13g2_a21oi_1 _23278_ (.A1(net649),
    .A2(_05642_),
    .Y(_05644_),
    .B1(_05643_));
 sg13g2_nand2_1 _23279_ (.Y(_05645_),
    .A(net611),
    .B(_05633_));
 sg13g2_a21oi_1 _23280_ (.A1(_05640_),
    .A2(_05645_),
    .Y(_05646_),
    .B1(_05046_));
 sg13g2_a21oi_1 _23281_ (.A1(_05046_),
    .A2(_05644_),
    .Y(_05647_),
    .B1(_05646_));
 sg13g2_nor2_1 _23282_ (.A(_12080_),
    .B(_05647_),
    .Y(_05648_));
 sg13g2_a21oi_1 _23283_ (.A1(net846),
    .A2(_05626_),
    .Y(_05649_),
    .B1(_05648_));
 sg13g2_nor2_1 _23284_ (.A(net82),
    .B(_05649_),
    .Y(_05650_));
 sg13g2_a21oi_1 _23285_ (.A1(_12010_),
    .A2(net71),
    .Y(_05651_),
    .B1(_05650_));
 sg13g2_nand2b_1 _23286_ (.Y(_05652_),
    .B(net579),
    .A_N(_04580_));
 sg13g2_a21oi_1 _23287_ (.A1(_05145_),
    .A2(_04582_),
    .Y(_05653_),
    .B1(net177));
 sg13g2_and2_1 _23288_ (.A(net85),
    .B(_05653_),
    .X(_05654_));
 sg13g2_nor3_1 _23289_ (.A(net987),
    .B(net83),
    .C(net176),
    .Y(_05655_));
 sg13g2_a221oi_1 _23290_ (.B2(_05654_),
    .C1(_05655_),
    .B1(_05652_),
    .A1(net74),
    .Y(_01044_),
    .A2(_05651_));
 sg13g2_a21oi_1 _23291_ (.A1(_05145_),
    .A2(_04616_),
    .Y(_05656_),
    .B1(_04216_));
 sg13g2_o21ai_1 _23292_ (.B1(_05656_),
    .Y(_05657_),
    .A1(net578),
    .A2(_04613_));
 sg13g2_o21ai_1 _23293_ (.B1(_05657_),
    .Y(_05658_),
    .A1(net986),
    .A2(net176));
 sg13g2_a22oi_1 _23294_ (.Y(_05659_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[5][22] ),
    .A2(net453),
    .A1(\cpu.dcache.r_data[6][22] ));
 sg13g2_inv_1 _23295_ (.Y(_05660_),
    .A(_00141_));
 sg13g2_a22oi_1 _23296_ (.Y(_05661_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][22] ),
    .A2(net452),
    .A1(_05660_));
 sg13g2_a22oi_1 _23297_ (.Y(_05662_),
    .B1(net450),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[7][22] ));
 sg13g2_a22oi_1 _23298_ (.Y(_05663_),
    .B1(net471),
    .B2(\cpu.dcache.r_data[4][22] ),
    .A2(net500),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_and4_1 _23299_ (.A(_05659_),
    .B(_05661_),
    .C(_05662_),
    .D(_05663_),
    .X(_05664_));
 sg13g2_buf_1 _23300_ (.A(_05664_),
    .X(_05665_));
 sg13g2_a22oi_1 _23301_ (.Y(_05666_),
    .B1(net451),
    .B2(\cpu.dcache.r_data[2][6] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][6] ));
 sg13g2_o21ai_1 _23302_ (.B1(_05666_),
    .Y(_05667_),
    .A1(_00140_),
    .A2(net616));
 sg13g2_a221oi_1 _23303_ (.B2(\cpu.dcache.r_data[3][6] ),
    .C1(_05667_),
    .B1(net473),
    .A1(\cpu.dcache.r_data[1][6] ),
    .Y(_05668_),
    .A2(net409));
 sg13g2_mux2_1 _23304_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(\cpu.dcache.r_data[6][6] ),
    .S(net695),
    .X(_05669_));
 sg13g2_a22oi_1 _23305_ (.Y(_05670_),
    .B1(_05669_),
    .B2(net654),
    .A2(_09805_),
    .A1(\cpu.dcache.r_data[5][6] ));
 sg13g2_nand2b_1 _23306_ (.Y(_05671_),
    .B(_12001_),
    .A_N(_05670_));
 sg13g2_and2_1 _23307_ (.A(_05668_),
    .B(_05671_),
    .X(_05672_));
 sg13g2_buf_1 _23308_ (.A(_05672_),
    .X(_05673_));
 sg13g2_mux2_1 _23309_ (.A0(_05665_),
    .A1(_05673_),
    .S(net611),
    .X(_05674_));
 sg13g2_nand3b_1 _23310_ (.B(_05042_),
    .C(net649),
    .Y(_05675_),
    .A_N(_05665_));
 sg13g2_o21ai_1 _23311_ (.B1(_05675_),
    .Y(_05676_),
    .A1(net649),
    .A2(_05252_));
 sg13g2_nand2b_1 _23312_ (.Y(_05677_),
    .B(_05259_),
    .A_N(_05045_));
 sg13g2_nor2_1 _23313_ (.A(_05517_),
    .B(_05673_),
    .Y(_05678_));
 sg13g2_a221oi_1 _23314_ (.B2(net650),
    .C1(_05678_),
    .B1(_05677_),
    .A1(_04992_),
    .Y(_05679_),
    .A2(_05676_));
 sg13g2_a21oi_1 _23315_ (.A1(net577),
    .A2(_05674_),
    .Y(_05680_),
    .B1(_05679_));
 sg13g2_nand3b_1 _23316_ (.B(_04902_),
    .C(net871),
    .Y(_05681_),
    .A_N(_00149_));
 sg13g2_o21ai_1 _23317_ (.B1(_05681_),
    .Y(_05682_),
    .A1(_00148_),
    .A2(_05099_));
 sg13g2_a21oi_1 _23318_ (.A1(_09246_),
    .A2(_04854_),
    .Y(_05683_),
    .B1(_05682_));
 sg13g2_nand3_1 _23319_ (.B(net984),
    .C(_04902_),
    .A(_09249_),
    .Y(_05684_));
 sg13g2_nand2b_1 _23320_ (.Y(_05685_),
    .B(_05684_),
    .A_N(_04917_));
 sg13g2_nor2_1 _23321_ (.A(net771),
    .B(_00146_),
    .Y(_05686_));
 sg13g2_buf_1 _23322_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05687_));
 sg13g2_nor2b_1 _23323_ (.A(net902),
    .B_N(_05687_),
    .Y(_05688_));
 sg13g2_o21ai_1 _23324_ (.B1(net505),
    .Y(_05689_),
    .A1(_05686_),
    .A2(_05688_));
 sg13g2_o21ai_1 _23325_ (.B1(_05689_),
    .Y(_05690_),
    .A1(_00147_),
    .A2(_05331_));
 sg13g2_a21oi_1 _23326_ (.A1(\cpu.gpio.r_enable_io[6] ),
    .A2(_05685_),
    .Y(_05691_),
    .B1(_05690_));
 sg13g2_nor2_1 _23327_ (.A(net771),
    .B(_00150_),
    .Y(_05692_));
 sg13g2_nor2b_1 _23328_ (.A(net902),
    .B_N(net9),
    .Y(_05693_));
 sg13g2_o21ai_1 _23329_ (.B1(net416),
    .Y(_05694_),
    .A1(_05692_),
    .A2(_05693_));
 sg13g2_a22oi_1 _23330_ (.Y(_05695_),
    .B1(_04862_),
    .B2(_09249_),
    .A2(net426),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_nand2_1 _23331_ (.Y(_05696_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_05086_));
 sg13g2_nand3_1 _23332_ (.B(_05695_),
    .C(_05696_),
    .A(_05694_),
    .Y(_05697_));
 sg13g2_nand2_1 _23333_ (.Y(_05698_),
    .A(net984),
    .B(_05697_));
 sg13g2_a21oi_1 _23334_ (.A1(_09246_),
    .A2(_04840_),
    .Y(_05699_),
    .B1(net455));
 sg13g2_nand2b_1 _23335_ (.Y(_05700_),
    .B(\cpu.gpio.r_enable_in[6] ),
    .A_N(_05699_));
 sg13g2_and4_1 _23336_ (.A(_05683_),
    .B(_05691_),
    .C(_05698_),
    .D(_05700_),
    .X(_05701_));
 sg13g2_or2_1 _23337_ (.X(_05702_),
    .B(_05701_),
    .A(_04824_));
 sg13g2_a22oi_1 _23338_ (.Y(_05703_),
    .B1(_04943_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net412),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_or2_1 _23339_ (.X(_05704_),
    .B(_05703_),
    .A(_04941_));
 sg13g2_mux2_1 _23340_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .S(net624),
    .X(_05705_));
 sg13g2_a22oi_1 _23341_ (.Y(_05706_),
    .B1(_05705_),
    .B2(net694),
    .A2(net775),
    .A1(_10013_));
 sg13g2_mux2_1 _23342_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(\cpu.intr.r_timer_reload[6] ),
    .S(net695),
    .X(_05707_));
 sg13g2_a221oi_1 _23343_ (.B2(net694),
    .C1(net681),
    .B1(_05707_),
    .A1(_10189_),
    .Y(_05708_),
    .A2(_09521_));
 sg13g2_a21o_1 _23344_ (.A2(_05706_),
    .A1(net648),
    .B1(_05708_),
    .X(_05709_));
 sg13g2_buf_2 _23345_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05710_));
 sg13g2_a22oi_1 _23346_ (.Y(_05711_),
    .B1(_04908_),
    .B2(_09992_),
    .A2(_10156_),
    .A1(_05710_));
 sg13g2_o21ai_1 _23347_ (.B1(_05711_),
    .Y(_05712_),
    .A1(net774),
    .A2(_05709_));
 sg13g2_inv_1 _23348_ (.Y(_05713_),
    .A(_00145_));
 sg13g2_buf_1 _23349_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05714_));
 sg13g2_a22oi_1 _23350_ (.Y(_05715_),
    .B1(_04931_),
    .B2(_05714_),
    .A2(net407),
    .A1(_05713_));
 sg13g2_nor2_1 _23351_ (.A(_00144_),
    .B(_04934_),
    .Y(_05716_));
 sg13g2_a21oi_1 _23352_ (.A1(\cpu.spi.r_timeout[6] ),
    .A2(_05112_),
    .Y(_05717_),
    .B1(_05716_));
 sg13g2_nand2_1 _23353_ (.Y(_05718_),
    .A(_09341_),
    .B(_04919_));
 sg13g2_nand3_1 _23354_ (.B(_05717_),
    .C(_05718_),
    .A(_05715_),
    .Y(_05719_));
 sg13g2_a22oi_1 _23355_ (.Y(_05720_),
    .B1(_05719_),
    .B2(_04939_),
    .A2(_05712_),
    .A1(_05012_));
 sg13g2_nand4_1 _23356_ (.B(_05702_),
    .C(_05704_),
    .A(net1025),
    .Y(_05721_),
    .D(_05720_));
 sg13g2_o21ai_1 _23357_ (.B1(_05721_),
    .Y(_05722_),
    .A1(net846),
    .A2(_05680_));
 sg13g2_nand2_1 _23358_ (.Y(_05723_),
    .A(net1071),
    .B(net81));
 sg13g2_o21ai_1 _23359_ (.B1(_05723_),
    .Y(_05724_),
    .A1(net71),
    .A2(_05722_));
 sg13g2_nor2_1 _23360_ (.A(_05291_),
    .B(_05724_),
    .Y(_05725_));
 sg13g2_a21oi_1 _23361_ (.A1(net73),
    .A2(_05658_),
    .Y(_01045_),
    .B1(_05725_));
 sg13g2_mux2_1 _23362_ (.A0(_05131_),
    .A1(_09229_),
    .S(net82),
    .X(_05726_));
 sg13g2_nand3_1 _23363_ (.B(_04618_),
    .C(_04640_),
    .A(net579),
    .Y(_05727_));
 sg13g2_a21oi_1 _23364_ (.A1(_05145_),
    .A2(_04642_),
    .Y(_05728_),
    .B1(net177));
 sg13g2_a221oi_1 _23365_ (.B2(_05728_),
    .C1(_04820_),
    .B1(_05727_),
    .A1(net988),
    .Y(_05729_),
    .A2(net177));
 sg13g2_a21o_1 _23366_ (.A2(_05726_),
    .A1(_05377_),
    .B1(_05729_),
    .X(_01046_));
 sg13g2_mux2_1 _23367_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(\cpu.intr.r_timer_reload[8] ),
    .S(net695),
    .X(_05730_));
 sg13g2_a22oi_1 _23368_ (.Y(_05731_),
    .B1(_05730_),
    .B2(net694),
    .A2(_09521_),
    .A1(_10199_));
 sg13g2_inv_1 _23369_ (.Y(_05732_),
    .A(\cpu.intr.r_clock_count[24] ));
 sg13g2_nor3_1 _23370_ (.A(_05732_),
    .B(_09463_),
    .C(net542),
    .Y(_05733_));
 sg13g2_a221oi_1 _23371_ (.B2(\cpu.intr.r_clock_cmp[24] ),
    .C1(_05733_),
    .B1(_05019_),
    .A1(\cpu.intr.r_timer_count[8] ),
    .Y(_05734_),
    .A2(_04908_));
 sg13g2_o21ai_1 _23372_ (.B1(_05734_),
    .Y(_05735_),
    .A1(_05015_),
    .A2(_05731_));
 sg13g2_a21o_1 _23373_ (.A2(_04999_),
    .A1(_05042_),
    .B1(_04991_),
    .X(_05736_));
 sg13g2_a22oi_1 _23374_ (.Y(_05737_),
    .B1(_05736_),
    .B2(_04955_),
    .A2(_05735_),
    .A1(_05014_));
 sg13g2_nor2_1 _23375_ (.A(net1030),
    .B(_05737_),
    .Y(_05738_));
 sg13g2_nor2b_1 _23376_ (.A(_05738_),
    .B_N(_05133_),
    .Y(_05739_));
 sg13g2_nand2b_1 _23377_ (.Y(_05740_),
    .B(_05141_),
    .A_N(_05739_));
 sg13g2_nand2b_1 _23378_ (.Y(_05741_),
    .B(net579),
    .A_N(_05740_));
 sg13g2_nor2_1 _23379_ (.A(_03570_),
    .B(_05739_),
    .Y(_05742_));
 sg13g2_a21oi_1 _23380_ (.A1(_09227_),
    .A2(net81),
    .Y(_05743_),
    .B1(_05742_));
 sg13g2_nand3_1 _23381_ (.B(net80),
    .C(_04216_),
    .A(_08850_),
    .Y(_05744_));
 sg13g2_o21ai_1 _23382_ (.B1(_05744_),
    .Y(_05745_),
    .A1(net80),
    .A2(_05743_));
 sg13g2_nand2_1 _23383_ (.Y(_05746_),
    .A(net578),
    .B(_04670_));
 sg13g2_nor2_1 _23384_ (.A(_05740_),
    .B(_05746_),
    .Y(_05747_));
 sg13g2_nor2_1 _23385_ (.A(_05745_),
    .B(_05747_),
    .Y(_05748_));
 sg13g2_o21ai_1 _23386_ (.B1(_05748_),
    .Y(_01047_),
    .A1(_04669_),
    .A2(_05741_));
 sg13g2_nand2_1 _23387_ (.Y(_05749_),
    .A(_03571_),
    .B(net196));
 sg13g2_a22oi_1 _23388_ (.Y(_05750_),
    .B1(net448),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(_05086_),
    .A1(_10207_));
 sg13g2_buf_1 _23389_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05751_));
 sg13g2_a22oi_1 _23390_ (.Y(_05752_),
    .B1(_05019_),
    .B2(\cpu.intr.r_clock_cmp[25] ),
    .A2(net426),
    .A1(_05751_));
 sg13g2_a22oi_1 _23391_ (.Y(_05753_),
    .B1(net414),
    .B2(\cpu.intr.r_timer_count[9] ),
    .A2(net545),
    .A1(\cpu.intr.r_timer_reload[9] ));
 sg13g2_or2_1 _23392_ (.X(_05754_),
    .B(_05753_),
    .A(net681));
 sg13g2_nand3_1 _23393_ (.B(_05752_),
    .C(_05754_),
    .A(_05750_),
    .Y(_05755_));
 sg13g2_o21ai_1 _23394_ (.B1(_05308_),
    .Y(_05756_),
    .A1(_10092_),
    .A2(_05301_));
 sg13g2_a22oi_1 _23395_ (.Y(_05757_),
    .B1(_05756_),
    .B2(_04955_),
    .A2(_05755_),
    .A1(_05014_));
 sg13g2_nor2_1 _23396_ (.A(net1030),
    .B(_05757_),
    .Y(_05758_));
 sg13g2_nor2b_1 _23397_ (.A(_05758_),
    .B_N(_05133_),
    .Y(_05759_));
 sg13g2_or4_1 _23398_ (.A(net578),
    .B(_04699_),
    .C(_05749_),
    .D(_05759_),
    .X(_05760_));
 sg13g2_nor2_1 _23399_ (.A(_03570_),
    .B(_05759_),
    .Y(_05761_));
 sg13g2_a21oi_1 _23400_ (.A1(_10819_),
    .A2(_05006_),
    .Y(_05762_),
    .B1(_05761_));
 sg13g2_nand3_1 _23401_ (.B(net80),
    .C(_04216_),
    .A(_08824_),
    .Y(_05763_));
 sg13g2_o21ai_1 _23402_ (.B1(_05763_),
    .Y(_05764_),
    .A1(net80),
    .A2(_05762_));
 sg13g2_nand2_1 _23403_ (.Y(_05765_),
    .A(net578),
    .B(_04701_));
 sg13g2_nor3_1 _23404_ (.A(_05749_),
    .B(_05759_),
    .C(_05765_),
    .Y(_05766_));
 sg13g2_nor2_1 _23405_ (.A(_05764_),
    .B(_05766_),
    .Y(_05767_));
 sg13g2_o21ai_1 _23406_ (.B1(_05767_),
    .Y(_01048_),
    .A1(_04672_),
    .A2(_05760_));
 sg13g2_nand2b_1 _23407_ (.Y(_05768_),
    .B(\cpu.dec.r_rd[0] ),
    .A_N(_03476_));
 sg13g2_a21oi_1 _23408_ (.A1(net176),
    .A2(_05768_),
    .Y(_05769_),
    .B1(_04820_));
 sg13g2_a21o_1 _23409_ (.A2(_05178_),
    .A1(net1046),
    .B1(_05769_),
    .X(_01049_));
 sg13g2_nor2b_1 _23410_ (.A(_03476_),
    .B_N(\cpu.dec.r_rd[1] ),
    .Y(_05770_));
 sg13g2_o21ai_1 _23411_ (.B1(net72),
    .Y(_05771_),
    .A1(net177),
    .A2(_05770_));
 sg13g2_o21ai_1 _23412_ (.B1(_05771_),
    .Y(_01050_),
    .A1(_03546_),
    .A2(net73));
 sg13g2_nor3_1 _23413_ (.A(_03476_),
    .B(_09304_),
    .C(net177),
    .Y(_05772_));
 sg13g2_nand3_1 _23414_ (.B(net85),
    .C(_05772_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05773_));
 sg13g2_o21ai_1 _23415_ (.B1(_05773_),
    .Y(_01051_),
    .A1(_10261_),
    .A2(_05182_));
 sg13g2_inv_1 _23416_ (.Y(_05774_),
    .A(_10259_));
 sg13g2_nand3_1 _23417_ (.B(net85),
    .C(_05772_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05775_));
 sg13g2_o21ai_1 _23418_ (.B1(_05775_),
    .Y(_01052_),
    .A1(_05774_),
    .A2(_05182_));
 sg13g2_mux2_1 _23419_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05178_),
    .X(_01053_));
 sg13g2_mux2_1 _23420_ (.A0(net869),
    .A1(_11086_),
    .S(net73),
    .X(_01054_));
 sg13g2_nand2_1 _23421_ (.Y(_05776_),
    .A(net590),
    .B(net541));
 sg13g2_o21ai_1 _23422_ (.B1(_05776_),
    .Y(_05777_),
    .A1(net540),
    .A2(_11009_));
 sg13g2_a21oi_1 _23423_ (.A1(_11302_),
    .A2(_11303_),
    .Y(_05778_),
    .B1(net850));
 sg13g2_a21o_1 _23424_ (.A2(_05777_),
    .A1(net735),
    .B1(_05778_),
    .X(_05779_));
 sg13g2_mux2_1 _23425_ (.A0(_10215_),
    .A1(_05779_),
    .S(net73),
    .X(_01055_));
 sg13g2_nand2_1 _23426_ (.Y(_05780_),
    .A(_09223_),
    .B(net541));
 sg13g2_o21ai_1 _23427_ (.B1(_05780_),
    .Y(_05781_),
    .A1(net540),
    .A2(_10970_));
 sg13g2_a21oi_1 _23428_ (.A1(_11464_),
    .A2(_11483_),
    .Y(_05782_),
    .B1(net850));
 sg13g2_a21oi_1 _23429_ (.A1(net735),
    .A2(_05781_),
    .Y(_05783_),
    .B1(_05782_));
 sg13g2_nand2_1 _23430_ (.Y(_05784_),
    .A(_10222_),
    .B(net74));
 sg13g2_o21ai_1 _23431_ (.B1(_05784_),
    .Y(_01056_),
    .A1(net70),
    .A2(_05783_));
 sg13g2_nand2_1 _23432_ (.Y(_05785_),
    .A(_03535_),
    .B(_10292_));
 sg13g2_o21ai_1 _23433_ (.B1(net601),
    .Y(_05786_),
    .A1(_11135_),
    .A2(_11148_));
 sg13g2_nand2_2 _23434_ (.Y(_05787_),
    .A(_05785_),
    .B(_05786_));
 sg13g2_a21oi_1 _23435_ (.A1(_11412_),
    .A2(_11414_),
    .Y(_05788_),
    .B1(net850));
 sg13g2_a21oi_1 _23436_ (.A1(net735),
    .A2(_05787_),
    .Y(_05789_),
    .B1(_05788_));
 sg13g2_nand2_1 _23437_ (.Y(_05790_),
    .A(_10227_),
    .B(net74));
 sg13g2_o21ai_1 _23438_ (.B1(_05790_),
    .Y(_01057_),
    .A1(net70),
    .A2(_05789_));
 sg13g2_nor3_1 _23439_ (.A(net850),
    .B(_11443_),
    .C(_11445_),
    .Y(_05791_));
 sg13g2_a21o_1 _23440_ (.A2(_11119_),
    .A1(net735),
    .B1(_05791_),
    .X(_05792_));
 sg13g2_nand2_1 _23441_ (.Y(_05793_),
    .A(_10229_),
    .B(net74));
 sg13g2_o21ai_1 _23442_ (.B1(_05793_),
    .Y(_01058_),
    .A1(net70),
    .A2(_05792_));
 sg13g2_nand2_1 _23443_ (.Y(_05794_),
    .A(_03099_),
    .B(_11211_));
 sg13g2_o21ai_1 _23444_ (.B1(_05794_),
    .Y(_05795_),
    .A1(net735),
    .A2(_11541_));
 sg13g2_mux2_1 _23445_ (.A0(_10239_),
    .A1(_05795_),
    .S(net73),
    .X(_01059_));
 sg13g2_and2_1 _23446_ (.A(_03098_),
    .B(_11184_),
    .X(_05796_));
 sg13g2_a21oi_1 _23447_ (.A1(_11599_),
    .A2(_10360_),
    .Y(_05797_),
    .B1(_05796_));
 sg13g2_nand2_1 _23448_ (.Y(_05798_),
    .A(_10244_),
    .B(net74));
 sg13g2_o21ai_1 _23449_ (.B1(_05798_),
    .Y(_01060_),
    .A1(net70),
    .A2(_05797_));
 sg13g2_nand2_1 _23450_ (.Y(_05799_),
    .A(net543),
    .B(net541));
 sg13g2_o21ai_1 _23451_ (.B1(_05799_),
    .Y(_05800_),
    .A1(_10358_),
    .A2(_11050_));
 sg13g2_mux2_1 _23452_ (.A0(_10145_),
    .A1(_05800_),
    .S(net72),
    .X(_01061_));
 sg13g2_mux2_1 _23453_ (.A0(_10165_),
    .A1(_05777_),
    .S(net72),
    .X(_01062_));
 sg13g2_mux2_1 _23454_ (.A0(net896),
    .A1(_05781_),
    .S(net72),
    .X(_01063_));
 sg13g2_mux2_1 _23455_ (.A0(net1047),
    .A1(_05787_),
    .S(net72),
    .X(_01064_));
 sg13g2_nand2_1 _23456_ (.Y(_05801_),
    .A(net1011),
    .B(net74));
 sg13g2_o21ai_1 _23457_ (.B1(_05801_),
    .Y(_01065_),
    .A1(_11119_),
    .A2(net70));
 sg13g2_nand2_1 _23458_ (.Y(_05802_),
    .A(net1010),
    .B(net74));
 sg13g2_o21ai_1 _23459_ (.B1(_05802_),
    .Y(_01066_),
    .A1(_11212_),
    .A2(net70));
 sg13g2_mux2_1 _23460_ (.A0(net899),
    .A1(_11184_),
    .S(net72),
    .X(_01067_));
 sg13g2_a22oi_1 _23461_ (.Y(_05803_),
    .B1(net601),
    .B2(_11375_),
    .A2(net541),
    .A1(net1070));
 sg13g2_nand2_1 _23462_ (.Y(_05804_),
    .A(net735),
    .B(_11086_));
 sg13g2_o21ai_1 _23463_ (.B1(_05804_),
    .Y(_05805_),
    .A1(net735),
    .A2(_05803_));
 sg13g2_mux2_1 _23464_ (.A0(_10205_),
    .A1(_05805_),
    .S(net72),
    .X(_01068_));
 sg13g2_a21oi_1 _23465_ (.A1(_11335_),
    .A2(_11336_),
    .Y(_05806_),
    .B1(_03098_));
 sg13g2_a21o_1 _23466_ (.A2(_05800_),
    .A1(net735),
    .B1(_05806_),
    .X(_05807_));
 sg13g2_mux2_1 _23467_ (.A0(_10210_),
    .A1(_05807_),
    .S(_05291_),
    .X(_01069_));
 sg13g2_buf_1 _23468_ (.A(net916),
    .X(_05808_));
 sg13g2_buf_1 _23469_ (.A(net275),
    .X(_05809_));
 sg13g2_nor2_1 _23470_ (.A(net664),
    .B(_10595_),
    .Y(_05810_));
 sg13g2_a21oi_1 _23471_ (.A1(_08373_),
    .A2(_10595_),
    .Y(_05811_),
    .B1(_05810_));
 sg13g2_or3_1 _23472_ (.A(_11088_),
    .B(_11010_),
    .C(\cpu.dec.imm[3] ),
    .X(_05812_));
 sg13g2_buf_1 _23473_ (.A(_05812_),
    .X(_05813_));
 sg13g2_o21ai_1 _23474_ (.B1(_03356_),
    .Y(_05814_),
    .A1(_11051_),
    .A2(_05813_));
 sg13g2_buf_1 _23475_ (.A(_05814_),
    .X(_05815_));
 sg13g2_nor4_2 _23476_ (.A(_08308_),
    .B(_04737_),
    .C(_10263_),
    .Y(_05816_),
    .D(_03547_));
 sg13g2_and2_1 _23477_ (.A(_05815_),
    .B(_05816_),
    .X(_05817_));
 sg13g2_buf_1 _23478_ (.A(_05817_),
    .X(_05818_));
 sg13g2_buf_1 _23479_ (.A(_00290_),
    .X(_05819_));
 sg13g2_nand2b_1 _23480_ (.Y(_05820_),
    .B(net990),
    .A_N(net1107));
 sg13g2_o21ai_1 _23481_ (.B1(_05820_),
    .Y(_05821_),
    .A1(net990),
    .A2(net664));
 sg13g2_nand3_1 _23482_ (.B(_05818_),
    .C(_05821_),
    .A(net275),
    .Y(_05822_));
 sg13g2_o21ai_1 _23483_ (.B1(_05822_),
    .Y(_05823_),
    .A1(_05809_),
    .A2(_05811_));
 sg13g2_o21ai_1 _23484_ (.B1(net916),
    .Y(_05824_),
    .A1(_08457_),
    .A2(_05818_));
 sg13g2_buf_1 _23485_ (.A(_05824_),
    .X(_05825_));
 sg13g2_inv_1 _23486_ (.Y(_05826_),
    .A(_10851_));
 sg13g2_a22oi_1 _23487_ (.Y(_01072_),
    .B1(_05825_),
    .B2(_05826_),
    .A2(_05823_),
    .A1(net728));
 sg13g2_inv_2 _23488_ (.Y(_05827_),
    .A(net1126));
 sg13g2_nor2_1 _23489_ (.A(_08466_),
    .B(net490),
    .Y(_05828_));
 sg13g2_a21oi_1 _23490_ (.A1(_11444_),
    .A2(net490),
    .Y(_05829_),
    .B1(_05828_));
 sg13g2_nor2_1 _23491_ (.A(_05826_),
    .B(_05827_),
    .Y(_05830_));
 sg13g2_buf_2 _23492_ (.A(_05830_),
    .X(_05831_));
 sg13g2_buf_1 _23493_ (.A(_10851_),
    .X(_05832_));
 sg13g2_nor2_2 _23494_ (.A(net982),
    .B(net1126),
    .Y(_05833_));
 sg13g2_o21ai_1 _23495_ (.B1(net990),
    .Y(_05834_),
    .A1(_05831_),
    .A2(_05833_));
 sg13g2_o21ai_1 _23496_ (.B1(_05834_),
    .Y(_05835_),
    .A1(net990),
    .A2(net776));
 sg13g2_nand3_1 _23497_ (.B(_05818_),
    .C(_05835_),
    .A(net210),
    .Y(_05836_));
 sg13g2_o21ai_1 _23498_ (.B1(_05836_),
    .Y(_05837_),
    .A1(net210),
    .A2(_05829_));
 sg13g2_buf_2 _23499_ (.A(net797),
    .X(_05838_));
 sg13g2_a22oi_1 _23500_ (.Y(_01073_),
    .B1(_05837_),
    .B2(net647),
    .A2(_05825_),
    .A1(_05827_));
 sg13g2_inv_2 _23501_ (.Y(_05839_),
    .A(_10872_));
 sg13g2_mux2_1 _23502_ (.A0(_08476_),
    .A1(net598),
    .S(net490),
    .X(_05840_));
 sg13g2_buf_1 _23503_ (.A(_10872_),
    .X(_05841_));
 sg13g2_nand2_1 _23504_ (.Y(_05842_),
    .A(_10851_),
    .B(net1126));
 sg13g2_buf_1 _23505_ (.A(_05842_),
    .X(_05843_));
 sg13g2_nor2_1 _23506_ (.A(_05841_),
    .B(net845),
    .Y(_05844_));
 sg13g2_buf_1 _23507_ (.A(net981),
    .X(_05845_));
 sg13g2_nand2_1 _23508_ (.Y(_05846_),
    .A(net844),
    .B(net845));
 sg13g2_nand3b_1 _23509_ (.B(_05846_),
    .C(_08403_),
    .Y(_05847_),
    .A_N(_05844_));
 sg13g2_o21ai_1 _23510_ (.B1(_05847_),
    .Y(_05848_),
    .A1(net990),
    .A2(net598));
 sg13g2_nand3_1 _23511_ (.B(_05818_),
    .C(_05848_),
    .A(net275),
    .Y(_05849_));
 sg13g2_o21ai_1 _23512_ (.B1(_05849_),
    .Y(_05850_),
    .A1(net210),
    .A2(_05840_));
 sg13g2_a22oi_1 _23513_ (.Y(_01074_),
    .B1(_05850_),
    .B2(_05838_),
    .A2(_05825_),
    .A1(_05839_));
 sg13g2_inv_1 _23514_ (.Y(_05851_),
    .A(_10308_));
 sg13g2_nor2_1 _23515_ (.A(net907),
    .B(_10595_),
    .Y(_05852_));
 sg13g2_a21oi_1 _23516_ (.A1(_08474_),
    .A2(_10595_),
    .Y(_05853_),
    .B1(_05852_));
 sg13g2_nand2_1 _23517_ (.Y(_05854_),
    .A(_10872_),
    .B(_05831_));
 sg13g2_buf_2 _23518_ (.A(_05854_),
    .X(_05855_));
 sg13g2_xnor2_1 _23519_ (.Y(_05856_),
    .A(net980),
    .B(_05855_));
 sg13g2_nand2_1 _23520_ (.Y(_05857_),
    .A(net990),
    .B(_05856_));
 sg13g2_o21ai_1 _23521_ (.B1(_05857_),
    .Y(_05858_),
    .A1(net990),
    .A2(net907));
 sg13g2_nand3_1 _23522_ (.B(_05818_),
    .C(_05858_),
    .A(net275),
    .Y(_05859_));
 sg13g2_o21ai_1 _23523_ (.B1(_05859_),
    .Y(_05860_),
    .A1(net210),
    .A2(_05853_));
 sg13g2_a22oi_1 _23524_ (.Y(_01075_),
    .B1(_05860_),
    .B2(_05808_),
    .A2(_05825_),
    .A1(net980));
 sg13g2_buf_2 _23525_ (.A(_00188_),
    .X(_05861_));
 sg13g2_nor2_1 _23526_ (.A(_10419_),
    .B(_10308_),
    .Y(_05862_));
 sg13g2_buf_2 _23527_ (.A(_05862_),
    .X(_05863_));
 sg13g2_nand2_1 _23528_ (.Y(_05864_),
    .A(_05861_),
    .B(_05863_));
 sg13g2_nand3b_1 _23529_ (.B(_05816_),
    .C(_08403_),
    .Y(_05865_),
    .A_N(_10503_));
 sg13g2_buf_1 _23530_ (.A(_05865_),
    .X(_05866_));
 sg13g2_nand3b_1 _23531_ (.B(_05827_),
    .C(_05826_),
    .Y(_05867_),
    .A_N(_05866_));
 sg13g2_buf_1 _23532_ (.A(_05867_),
    .X(_05868_));
 sg13g2_nor2_1 _23533_ (.A(_05864_),
    .B(_05868_),
    .Y(_05869_));
 sg13g2_buf_1 _23534_ (.A(_05869_),
    .X(_05870_));
 sg13g2_buf_1 _23535_ (.A(_05870_),
    .X(_05871_));
 sg13g2_mux2_1 _23536_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(_03536_),
    .S(_05871_),
    .X(_01143_));
 sg13g2_mux2_1 _23537_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net512),
    .S(net255),
    .X(_01144_));
 sg13g2_mux2_1 _23538_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(_03530_),
    .S(net255),
    .X(_01145_));
 sg13g2_mux2_1 _23539_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net514),
    .S(net255),
    .X(_01146_));
 sg13g2_mux2_1 _23540_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net732),
    .S(net255),
    .X(_01147_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net730),
    .S(net255),
    .X(_01148_));
 sg13g2_mux2_1 _23542_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net729),
    .S(net255),
    .X(_01149_));
 sg13g2_buf_1 _23543_ (.A(_10819_),
    .X(_05872_));
 sg13g2_mux2_1 _23544_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net979),
    .S(net255),
    .X(_01150_));
 sg13g2_buf_1 _23545_ (.A(net992),
    .X(_05873_));
 sg13g2_mux2_1 _23546_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net843),
    .S(_05871_),
    .X(_01151_));
 sg13g2_buf_1 _23547_ (.A(net991),
    .X(_05874_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net842),
    .S(net255),
    .X(_01152_));
 sg13g2_mux2_1 _23549_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(_03526_),
    .S(_05870_),
    .X(_01153_));
 sg13g2_mux2_1 _23550_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(_03527_),
    .S(_05870_),
    .X(_01154_));
 sg13g2_buf_1 _23551_ (.A(net517),
    .X(_05875_));
 sg13g2_buf_1 _23552_ (.A(_05866_),
    .X(_05876_));
 sg13g2_nand2_1 _23553_ (.Y(_05877_),
    .A(_05826_),
    .B(net1126));
 sg13g2_buf_1 _23554_ (.A(_05877_),
    .X(_05878_));
 sg13g2_nand2_1 _23555_ (.Y(_05879_),
    .A(_10420_),
    .B(_10308_));
 sg13g2_buf_2 _23556_ (.A(_05879_),
    .X(_05880_));
 sg13g2_nor3_2 _23557_ (.A(net981),
    .B(net727),
    .C(_05880_),
    .Y(_05881_));
 sg13g2_nor2b_1 _23558_ (.A(net446),
    .B_N(_05881_),
    .Y(_05882_));
 sg13g2_buf_1 _23559_ (.A(_05882_),
    .X(_05883_));
 sg13g2_buf_1 _23560_ (.A(_05883_),
    .X(_05884_));
 sg13g2_mux2_1 _23561_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net447),
    .S(net330),
    .X(_01155_));
 sg13g2_mux2_1 _23562_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net512),
    .S(net330),
    .X(_01156_));
 sg13g2_buf_1 _23563_ (.A(net907),
    .X(_05885_));
 sg13g2_mux2_1 _23564_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net726),
    .S(net330),
    .X(_01157_));
 sg13g2_mux2_1 _23565_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net514),
    .S(_05884_),
    .X(_01158_));
 sg13g2_mux2_1 _23566_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net732),
    .S(net330),
    .X(_01159_));
 sg13g2_mux2_1 _23567_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net730),
    .S(net330),
    .X(_01160_));
 sg13g2_mux2_1 _23568_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net729),
    .S(net330),
    .X(_01161_));
 sg13g2_mux2_1 _23569_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net979),
    .S(_05884_),
    .X(_01162_));
 sg13g2_mux2_1 _23570_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net843),
    .S(net330),
    .X(_01163_));
 sg13g2_mux2_1 _23571_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net842),
    .S(net330),
    .X(_01164_));
 sg13g2_buf_1 _23572_ (.A(net664),
    .X(_05886_));
 sg13g2_mux2_1 _23573_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(_05886_),
    .S(_05883_),
    .X(_01165_));
 sg13g2_buf_1 _23574_ (.A(net776),
    .X(_05887_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(_05887_),
    .S(_05883_),
    .X(_01166_));
 sg13g2_nor3_1 _23576_ (.A(net981),
    .B(net845),
    .C(_05880_),
    .Y(_05888_));
 sg13g2_buf_2 _23577_ (.A(_05888_),
    .X(_05889_));
 sg13g2_nor2b_1 _23578_ (.A(net446),
    .B_N(_05889_),
    .Y(_05890_));
 sg13g2_buf_1 _23579_ (.A(_05890_),
    .X(_05891_));
 sg13g2_buf_1 _23580_ (.A(_05891_),
    .X(_05892_));
 sg13g2_mux2_1 _23581_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net447),
    .S(net329),
    .X(_01167_));
 sg13g2_mux2_1 _23582_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net512),
    .S(net329),
    .X(_01168_));
 sg13g2_mux2_1 _23583_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(_05885_),
    .S(net329),
    .X(_01169_));
 sg13g2_mux2_1 _23584_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net514),
    .S(_05892_),
    .X(_01170_));
 sg13g2_mux2_1 _23585_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net732),
    .S(net329),
    .X(_01171_));
 sg13g2_mux2_1 _23586_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(_04742_),
    .S(net329),
    .X(_01172_));
 sg13g2_mux2_1 _23587_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net729),
    .S(net329),
    .X(_01173_));
 sg13g2_mux2_1 _23588_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(_05872_),
    .S(_05892_),
    .X(_01174_));
 sg13g2_mux2_1 _23589_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net843),
    .S(net329),
    .X(_01175_));
 sg13g2_mux2_1 _23590_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net842),
    .S(net329),
    .X(_01176_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(_05886_),
    .S(_05891_),
    .X(_01177_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(_05887_),
    .S(_05891_),
    .X(_01178_));
 sg13g2_nor2_2 _23593_ (.A(_10419_),
    .B(net980),
    .Y(_05893_));
 sg13g2_nand2b_1 _23594_ (.Y(_05894_),
    .B(_05893_),
    .A_N(_05861_));
 sg13g2_buf_1 _23595_ (.A(_05894_),
    .X(_05895_));
 sg13g2_nor2_1 _23596_ (.A(_05868_),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_buf_1 _23597_ (.A(_05896_),
    .X(_05897_));
 sg13g2_buf_1 _23598_ (.A(_05897_),
    .X(_05898_));
 sg13g2_mux2_1 _23599_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net447),
    .S(net254),
    .X(_01179_));
 sg13g2_mux2_1 _23600_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net512),
    .S(net254),
    .X(_01180_));
 sg13g2_mux2_1 _23601_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(_05885_),
    .S(net254),
    .X(_01181_));
 sg13g2_mux2_1 _23602_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(_03555_),
    .S(net254),
    .X(_01182_));
 sg13g2_mux2_1 _23603_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net732),
    .S(net254),
    .X(_01183_));
 sg13g2_mux2_1 _23604_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net730),
    .S(net254),
    .X(_01184_));
 sg13g2_mux2_1 _23605_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net729),
    .S(net254),
    .X(_01185_));
 sg13g2_mux2_1 _23606_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(_05872_),
    .S(net254),
    .X(_01186_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net843),
    .S(_05898_),
    .X(_01187_));
 sg13g2_mux2_1 _23608_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net842),
    .S(_05898_),
    .X(_01188_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net576),
    .S(_05897_),
    .X(_01189_));
 sg13g2_mux2_1 _23610_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net646),
    .S(_05897_),
    .X(_01190_));
 sg13g2_nand2_1 _23611_ (.Y(_05899_),
    .A(_10851_),
    .B(_05827_));
 sg13g2_buf_2 _23612_ (.A(_05899_),
    .X(_05900_));
 sg13g2_or2_1 _23613_ (.X(_05901_),
    .B(_05866_),
    .A(_05900_));
 sg13g2_buf_2 _23614_ (.A(_05901_),
    .X(_05902_));
 sg13g2_nor2_1 _23615_ (.A(_05895_),
    .B(_05902_),
    .Y(_05903_));
 sg13g2_buf_1 _23616_ (.A(_05903_),
    .X(_05904_));
 sg13g2_buf_1 _23617_ (.A(_05904_),
    .X(_05905_));
 sg13g2_mux2_1 _23618_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net447),
    .S(net253),
    .X(_01191_));
 sg13g2_mux2_1 _23619_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net512),
    .S(net253),
    .X(_01192_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net726),
    .S(net253),
    .X(_01193_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(_03555_),
    .S(net253),
    .X(_01194_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(_03556_),
    .S(net253),
    .X(_01195_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net730),
    .S(net253),
    .X(_01196_));
 sg13g2_mux2_1 _23624_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net729),
    .S(net253),
    .X(_01197_));
 sg13g2_mux2_1 _23625_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net979),
    .S(_05905_),
    .X(_01198_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net843),
    .S(_05905_),
    .X(_01199_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net842),
    .S(net253),
    .X(_01200_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net576),
    .S(_05904_),
    .X(_01201_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net646),
    .S(_05904_),
    .X(_01202_));
 sg13g2_buf_1 _23630_ (.A(_05866_),
    .X(_05906_));
 sg13g2_nor3_1 _23631_ (.A(net727),
    .B(_05906_),
    .C(_05895_),
    .Y(_05907_));
 sg13g2_buf_1 _23632_ (.A(_05907_),
    .X(_05908_));
 sg13g2_buf_1 _23633_ (.A(_05908_),
    .X(_05909_));
 sg13g2_mux2_1 _23634_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(_05875_),
    .S(net328),
    .X(_01203_));
 sg13g2_mux2_1 _23635_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(_03563_),
    .S(net328),
    .X(_01204_));
 sg13g2_mux2_1 _23636_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net726),
    .S(net328),
    .X(_01205_));
 sg13g2_buf_1 _23637_ (.A(net662),
    .X(_05910_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_05910_),
    .S(net328),
    .X(_01206_));
 sg13g2_mux2_1 _23639_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(_03556_),
    .S(net328),
    .X(_01207_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net730),
    .S(net328),
    .X(_01208_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net729),
    .S(net328),
    .X(_01209_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net979),
    .S(_05909_),
    .X(_01210_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(_05873_),
    .S(_05909_),
    .X(_01211_));
 sg13g2_mux2_1 _23644_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(_05874_),
    .S(net328),
    .X(_01212_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(net576),
    .S(_05908_),
    .X(_01213_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(net646),
    .S(_05908_),
    .X(_01214_));
 sg13g2_nor3_1 _23647_ (.A(net845),
    .B(net445),
    .C(_05895_),
    .Y(_05911_));
 sg13g2_buf_1 _23648_ (.A(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _23649_ (.A(_05912_),
    .X(_05913_));
 sg13g2_mux2_1 _23650_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05875_),
    .S(net327),
    .X(_01215_));
 sg13g2_mux2_1 _23651_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(_03563_),
    .S(net327),
    .X(_01216_));
 sg13g2_mux2_1 _23652_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(net726),
    .S(net327),
    .X(_01217_));
 sg13g2_mux2_1 _23653_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(net575),
    .S(net327),
    .X(_01218_));
 sg13g2_buf_1 _23654_ (.A(net857),
    .X(_05914_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(_05914_),
    .S(net327),
    .X(_01219_));
 sg13g2_mux2_1 _23656_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(net730),
    .S(net327),
    .X(_01220_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(_04743_),
    .S(net327),
    .X(_01221_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(net979),
    .S(_05913_),
    .X(_01222_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(_05873_),
    .S(_05913_),
    .X(_01223_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(_05874_),
    .S(net327),
    .X(_01224_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(net576),
    .S(_05912_),
    .X(_01225_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(net646),
    .S(_05912_),
    .X(_01226_));
 sg13g2_nand2_1 _23663_ (.Y(_05915_),
    .A(_10419_),
    .B(net980));
 sg13g2_buf_2 _23664_ (.A(_05915_),
    .X(_05916_));
 sg13g2_nand2_2 _23665_ (.Y(_05917_),
    .A(_05839_),
    .B(_05833_));
 sg13g2_nor3_1 _23666_ (.A(net445),
    .B(_05916_),
    .C(_05917_),
    .Y(_05918_));
 sg13g2_buf_1 _23667_ (.A(_05918_),
    .X(_05919_));
 sg13g2_buf_1 _23668_ (.A(_05919_),
    .X(_05920_));
 sg13g2_mux2_1 _23669_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net447),
    .S(net326),
    .X(_01227_));
 sg13g2_buf_1 _23670_ (.A(_11523_),
    .X(_05921_));
 sg13g2_mux2_1 _23671_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net497),
    .S(net326),
    .X(_01228_));
 sg13g2_mux2_1 _23672_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net726),
    .S(net326),
    .X(_01229_));
 sg13g2_mux2_1 _23673_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net575),
    .S(net326),
    .X(_01230_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net725),
    .S(net326),
    .X(_01231_));
 sg13g2_mux2_1 _23675_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net730),
    .S(net326),
    .X(_01232_));
 sg13g2_mux2_1 _23676_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net729),
    .S(net326),
    .X(_01233_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net979),
    .S(_05920_),
    .X(_01234_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net843),
    .S(_05920_),
    .X(_01235_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net842),
    .S(net326),
    .X(_01236_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net576),
    .S(_05919_),
    .X(_01237_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net646),
    .S(_05919_),
    .X(_01238_));
 sg13g2_nor3_1 _23682_ (.A(_05845_),
    .B(_05902_),
    .C(_05916_),
    .Y(_05922_));
 sg13g2_buf_1 _23683_ (.A(_05922_),
    .X(_05923_));
 sg13g2_buf_1 _23684_ (.A(_05923_),
    .X(_05924_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net447),
    .S(net252),
    .X(_01239_));
 sg13g2_mux2_1 _23686_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net497),
    .S(net252),
    .X(_01240_));
 sg13g2_mux2_1 _23687_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net726),
    .S(net252),
    .X(_01241_));
 sg13g2_mux2_1 _23688_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net575),
    .S(net252),
    .X(_01242_));
 sg13g2_mux2_1 _23689_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net725),
    .S(net252),
    .X(_01243_));
 sg13g2_mux2_1 _23690_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net730),
    .S(net252),
    .X(_01244_));
 sg13g2_mux2_1 _23691_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net729),
    .S(net252),
    .X(_01245_));
 sg13g2_mux2_1 _23692_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net979),
    .S(_05924_),
    .X(_01246_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net843),
    .S(net252),
    .X(_01247_));
 sg13g2_mux2_1 _23694_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net842),
    .S(_05924_),
    .X(_01248_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net576),
    .S(_05923_),
    .X(_01249_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net646),
    .S(_05923_),
    .X(_01250_));
 sg13g2_buf_1 _23697_ (.A(_10308_),
    .X(_05925_));
 sg13g2_nor2_1 _23698_ (.A(_10420_),
    .B(_10851_),
    .Y(_05926_));
 sg13g2_nand3_1 _23699_ (.B(_05839_),
    .C(_05926_),
    .A(_11433_),
    .Y(_05927_));
 sg13g2_nor2_2 _23700_ (.A(net978),
    .B(_05927_),
    .Y(_05928_));
 sg13g2_nor2b_1 _23701_ (.A(net446),
    .B_N(_05928_),
    .Y(_05929_));
 sg13g2_buf_1 _23702_ (.A(_05929_),
    .X(_05930_));
 sg13g2_buf_1 _23703_ (.A(_05930_),
    .X(_05931_));
 sg13g2_mux2_1 _23704_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net447),
    .S(net325),
    .X(_01251_));
 sg13g2_mux2_1 _23705_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net497),
    .S(net325),
    .X(_01252_));
 sg13g2_mux2_1 _23706_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net726),
    .S(net325),
    .X(_01253_));
 sg13g2_mux2_1 _23707_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net575),
    .S(net325),
    .X(_01254_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net725),
    .S(net325),
    .X(_01255_));
 sg13g2_buf_1 _23709_ (.A(net1069),
    .X(_05932_));
 sg13g2_mux2_1 _23710_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net841),
    .S(net325),
    .X(_01256_));
 sg13g2_buf_1 _23711_ (.A(_09227_),
    .X(_05933_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(_05933_),
    .S(net325),
    .X(_01257_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net979),
    .S(_05931_),
    .X(_01258_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net843),
    .S(net325),
    .X(_01259_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net842),
    .S(_05931_),
    .X(_01260_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net576),
    .S(_05930_),
    .X(_01261_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net646),
    .S(_05930_),
    .X(_01262_));
 sg13g2_nor3_1 _23718_ (.A(net981),
    .B(net845),
    .C(_05916_),
    .Y(_05934_));
 sg13g2_buf_2 _23719_ (.A(_05934_),
    .X(_05935_));
 sg13g2_nor2b_1 _23720_ (.A(net446),
    .B_N(_05935_),
    .Y(_05936_));
 sg13g2_buf_1 _23721_ (.A(_05936_),
    .X(_05937_));
 sg13g2_buf_1 _23722_ (.A(_05937_),
    .X(_05938_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(net447),
    .S(net324),
    .X(_01263_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(_05921_),
    .S(net324),
    .X(_01264_));
 sg13g2_mux2_1 _23725_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net726),
    .S(net324),
    .X(_01265_));
 sg13g2_mux2_1 _23726_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net575),
    .S(net324),
    .X(_01266_));
 sg13g2_mux2_1 _23727_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(net725),
    .S(net324),
    .X(_01267_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(_05932_),
    .S(net324),
    .X(_01268_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(_05933_),
    .S(net324),
    .X(_01269_));
 sg13g2_buf_1 _23730_ (.A(_10819_),
    .X(_05939_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(_05939_),
    .S(_05938_),
    .X(_01270_));
 sg13g2_buf_1 _23732_ (.A(_10903_),
    .X(_05940_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(_05940_),
    .S(net324),
    .X(_01271_));
 sg13g2_buf_1 _23734_ (.A(_10925_),
    .X(_05941_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(_05941_),
    .S(_05938_),
    .X(_01272_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net576),
    .S(_05937_),
    .X(_01273_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net646),
    .S(_05937_),
    .X(_01274_));
 sg13g2_buf_1 _23738_ (.A(net517),
    .X(_05942_));
 sg13g2_nor2_1 _23739_ (.A(_05864_),
    .B(_05902_),
    .Y(_05943_));
 sg13g2_buf_1 _23740_ (.A(_05943_),
    .X(_05944_));
 sg13g2_buf_1 _23741_ (.A(_05944_),
    .X(_05945_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(net444),
    .S(net251),
    .X(_01275_));
 sg13g2_mux2_1 _23743_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(_05921_),
    .S(net251),
    .X(_01276_));
 sg13g2_buf_1 _23744_ (.A(net907),
    .X(_05946_));
 sg13g2_mux2_1 _23745_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05946_),
    .S(net251),
    .X(_01277_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05910_),
    .S(net251),
    .X(_01278_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(_05914_),
    .S(net251),
    .X(_01279_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(_05932_),
    .S(net251),
    .X(_01280_));
 sg13g2_mux2_1 _23749_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(net840),
    .S(_05945_),
    .X(_01281_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05939_),
    .S(_05945_),
    .X(_01282_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05940_),
    .S(net251),
    .X(_01283_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(_05941_),
    .S(net251),
    .X(_01284_));
 sg13g2_buf_1 _23753_ (.A(net664),
    .X(_05947_));
 sg13g2_mux2_1 _23754_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(_05947_),
    .S(_05944_),
    .X(_01285_));
 sg13g2_buf_1 _23755_ (.A(net776),
    .X(_05948_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05948_),
    .S(_05944_),
    .X(_01286_));
 sg13g2_or2_1 _23757_ (.X(_05949_),
    .B(_05916_),
    .A(_05861_));
 sg13g2_buf_1 _23758_ (.A(_05949_),
    .X(_05950_));
 sg13g2_nor2_1 _23759_ (.A(_05868_),
    .B(_05950_),
    .Y(_05951_));
 sg13g2_buf_1 _23760_ (.A(_05951_),
    .X(_05952_));
 sg13g2_buf_1 _23761_ (.A(_05952_),
    .X(_05953_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net444),
    .S(net250),
    .X(_01287_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net497),
    .S(net250),
    .X(_01288_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net724),
    .S(net250),
    .X(_01289_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net575),
    .S(net250),
    .X(_01290_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net725),
    .S(net250),
    .X(_01291_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net841),
    .S(net250),
    .X(_01292_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net840),
    .S(net250),
    .X(_01293_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net977),
    .S(_05953_),
    .X(_01294_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net976),
    .S(net250),
    .X(_01295_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net975),
    .S(_05953_),
    .X(_01296_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(_05947_),
    .S(_05952_),
    .X(_01297_));
 sg13g2_mux2_1 _23773_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net645),
    .S(_05952_),
    .X(_01298_));
 sg13g2_nor2_1 _23774_ (.A(_05902_),
    .B(_05950_),
    .Y(_05954_));
 sg13g2_buf_1 _23775_ (.A(_05954_),
    .X(_05955_));
 sg13g2_buf_1 _23776_ (.A(_05955_),
    .X(_05956_));
 sg13g2_mux2_1 _23777_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net444),
    .S(net249),
    .X(_01299_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net497),
    .S(net249),
    .X(_01300_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net724),
    .S(net249),
    .X(_01301_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net575),
    .S(net249),
    .X(_01302_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net725),
    .S(net249),
    .X(_01303_));
 sg13g2_mux2_1 _23782_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net841),
    .S(net249),
    .X(_01304_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net840),
    .S(net249),
    .X(_01305_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net977),
    .S(_05956_),
    .X(_01306_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net976),
    .S(net249),
    .X(_01307_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net975),
    .S(_05956_),
    .X(_01308_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net574),
    .S(_05955_),
    .X(_01309_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net645),
    .S(_05955_),
    .X(_01310_));
 sg13g2_nor3_1 _23789_ (.A(net727),
    .B(net445),
    .C(_05950_),
    .Y(_05957_));
 sg13g2_buf_1 _23790_ (.A(_05957_),
    .X(_05958_));
 sg13g2_buf_1 _23791_ (.A(_05958_),
    .X(_05959_));
 sg13g2_mux2_1 _23792_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net444),
    .S(net323),
    .X(_01311_));
 sg13g2_mux2_1 _23793_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net497),
    .S(net323),
    .X(_01312_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net724),
    .S(net323),
    .X(_01313_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net575),
    .S(net323),
    .X(_01314_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net725),
    .S(net323),
    .X(_01315_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net841),
    .S(net323),
    .X(_01316_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net840),
    .S(_05959_),
    .X(_01317_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net977),
    .S(_05959_),
    .X(_01318_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net976),
    .S(net323),
    .X(_01319_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net975),
    .S(net323),
    .X(_01320_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net574),
    .S(_05958_),
    .X(_01321_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net645),
    .S(_05958_),
    .X(_01322_));
 sg13g2_nor3_1 _23804_ (.A(net845),
    .B(net445),
    .C(_05950_),
    .Y(_05960_));
 sg13g2_buf_1 _23805_ (.A(_05960_),
    .X(_05961_));
 sg13g2_buf_1 _23806_ (.A(_05961_),
    .X(_05962_));
 sg13g2_mux2_1 _23807_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net444),
    .S(net322),
    .X(_01323_));
 sg13g2_mux2_1 _23808_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net497),
    .S(net322),
    .X(_01324_));
 sg13g2_mux2_1 _23809_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net724),
    .S(net322),
    .X(_01325_));
 sg13g2_buf_1 _23810_ (.A(_12010_),
    .X(_05963_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(_05963_),
    .S(net322),
    .X(_01326_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net725),
    .S(net322),
    .X(_01327_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net841),
    .S(net322),
    .X(_01328_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net840),
    .S(_05962_),
    .X(_01329_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net977),
    .S(_05962_),
    .X(_01330_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net976),
    .S(net322),
    .X(_01331_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net975),
    .S(net322),
    .X(_01332_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net574),
    .S(_05961_),
    .X(_01333_));
 sg13g2_mux2_1 _23819_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net645),
    .S(_05961_),
    .X(_01334_));
 sg13g2_buf_1 _23820_ (.A(_10419_),
    .X(_05964_));
 sg13g2_nand2_2 _23821_ (.Y(_05965_),
    .A(net974),
    .B(net978));
 sg13g2_nor3_1 _23822_ (.A(net445),
    .B(_05917_),
    .C(_05965_),
    .Y(_05966_));
 sg13g2_buf_1 _23823_ (.A(_05966_),
    .X(_05967_));
 sg13g2_buf_1 _23824_ (.A(_05967_),
    .X(_05968_));
 sg13g2_mux2_1 _23825_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net444),
    .S(net321),
    .X(_01335_));
 sg13g2_mux2_1 _23826_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net497),
    .S(net321),
    .X(_01336_));
 sg13g2_mux2_1 _23827_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net724),
    .S(net321),
    .X(_01337_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net573),
    .S(net321),
    .X(_01338_));
 sg13g2_buf_1 _23829_ (.A(_09225_),
    .X(_05969_));
 sg13g2_mux2_1 _23830_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net839),
    .S(net321),
    .X(_01339_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net841),
    .S(net321),
    .X(_01340_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net840),
    .S(net321),
    .X(_01341_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net977),
    .S(_05968_),
    .X(_01342_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net976),
    .S(_05968_),
    .X(_01343_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net975),
    .S(net321),
    .X(_01344_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net574),
    .S(_05967_),
    .X(_01345_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net645),
    .S(_05967_),
    .X(_01346_));
 sg13g2_nor3_1 _23838_ (.A(_05845_),
    .B(_05902_),
    .C(_05965_),
    .Y(_05970_));
 sg13g2_buf_1 _23839_ (.A(_05970_),
    .X(_05971_));
 sg13g2_buf_1 _23840_ (.A(_05971_),
    .X(_05972_));
 sg13g2_mux2_1 _23841_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net444),
    .S(net248),
    .X(_01347_));
 sg13g2_buf_1 _23842_ (.A(_11523_),
    .X(_05973_));
 sg13g2_mux2_1 _23843_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net496),
    .S(net248),
    .X(_01348_));
 sg13g2_mux2_1 _23844_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net724),
    .S(net248),
    .X(_01349_));
 sg13g2_mux2_1 _23845_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net573),
    .S(net248),
    .X(_01350_));
 sg13g2_mux2_1 _23846_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net839),
    .S(net248),
    .X(_01351_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net841),
    .S(net248),
    .X(_01352_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net840),
    .S(net248),
    .X(_01353_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net977),
    .S(_05972_),
    .X(_01354_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net976),
    .S(_05972_),
    .X(_01355_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net975),
    .S(net248),
    .X(_01356_));
 sg13g2_mux2_1 _23852_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net574),
    .S(_05971_),
    .X(_01357_));
 sg13g2_mux2_1 _23853_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net645),
    .S(_05971_),
    .X(_01358_));
 sg13g2_nor2_2 _23854_ (.A(net980),
    .B(_05927_),
    .Y(_05974_));
 sg13g2_nor2b_1 _23855_ (.A(net446),
    .B_N(_05974_),
    .Y(_05975_));
 sg13g2_buf_1 _23856_ (.A(_05975_),
    .X(_05976_));
 sg13g2_buf_1 _23857_ (.A(_05976_),
    .X(_05977_));
 sg13g2_mux2_1 _23858_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(_05942_),
    .S(net320),
    .X(_01359_));
 sg13g2_mux2_1 _23859_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net496),
    .S(net320),
    .X(_01360_));
 sg13g2_mux2_1 _23860_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net724),
    .S(net320),
    .X(_01361_));
 sg13g2_mux2_1 _23861_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net573),
    .S(net320),
    .X(_01362_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net839),
    .S(net320),
    .X(_01363_));
 sg13g2_mux2_1 _23863_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net841),
    .S(net320),
    .X(_01364_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net840),
    .S(net320),
    .X(_01365_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net977),
    .S(_05977_),
    .X(_01366_));
 sg13g2_mux2_1 _23866_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net976),
    .S(_05977_),
    .X(_01367_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net975),
    .S(net320),
    .X(_01368_));
 sg13g2_mux2_1 _23868_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net574),
    .S(_05976_),
    .X(_01369_));
 sg13g2_mux2_1 _23869_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net645),
    .S(_05976_),
    .X(_01370_));
 sg13g2_nor3_1 _23870_ (.A(net981),
    .B(net845),
    .C(_05965_),
    .Y(_05978_));
 sg13g2_buf_2 _23871_ (.A(_05978_),
    .X(_05979_));
 sg13g2_nor2b_1 _23872_ (.A(net446),
    .B_N(_05979_),
    .Y(_05980_));
 sg13g2_buf_1 _23873_ (.A(_05980_),
    .X(_05981_));
 sg13g2_buf_1 _23874_ (.A(_05981_),
    .X(_05982_));
 sg13g2_mux2_1 _23875_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(_05942_),
    .S(net319),
    .X(_01371_));
 sg13g2_mux2_1 _23876_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net496),
    .S(net319),
    .X(_01372_));
 sg13g2_mux2_1 _23877_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net724),
    .S(net319),
    .X(_01373_));
 sg13g2_mux2_1 _23878_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net573),
    .S(net319),
    .X(_01374_));
 sg13g2_mux2_1 _23879_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net839),
    .S(net319),
    .X(_01375_));
 sg13g2_buf_1 _23880_ (.A(net1069),
    .X(_05983_));
 sg13g2_mux2_1 _23881_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net838),
    .S(net319),
    .X(_01376_));
 sg13g2_buf_1 _23882_ (.A(net1070),
    .X(_05984_));
 sg13g2_mux2_1 _23883_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net837),
    .S(net319),
    .X(_01377_));
 sg13g2_mux2_1 _23884_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net977),
    .S(_05982_),
    .X(_01378_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net976),
    .S(_05982_),
    .X(_01379_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net975),
    .S(net319),
    .X(_01380_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net574),
    .S(_05981_),
    .X(_01381_));
 sg13g2_mux2_1 _23888_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net645),
    .S(_05981_),
    .X(_01382_));
 sg13g2_or2_1 _23889_ (.X(_05985_),
    .B(_05965_),
    .A(_05861_));
 sg13g2_buf_1 _23890_ (.A(_05985_),
    .X(_05986_));
 sg13g2_nor2_1 _23891_ (.A(_05868_),
    .B(_05986_),
    .Y(_05987_));
 sg13g2_buf_1 _23892_ (.A(_05987_),
    .X(_05988_));
 sg13g2_buf_1 _23893_ (.A(_05988_),
    .X(_05989_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net444),
    .S(net247),
    .X(_01383_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net496),
    .S(net247),
    .X(_01384_));
 sg13g2_mux2_1 _23896_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(_05946_),
    .S(net247),
    .X(_01385_));
 sg13g2_mux2_1 _23897_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net573),
    .S(net247),
    .X(_01386_));
 sg13g2_mux2_1 _23898_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net839),
    .S(net247),
    .X(_01387_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net838),
    .S(net247),
    .X(_01388_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net837),
    .S(net247),
    .X(_01389_));
 sg13g2_buf_1 _23901_ (.A(_10819_),
    .X(_05990_));
 sg13g2_mux2_1 _23902_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net973),
    .S(_05989_),
    .X(_01390_));
 sg13g2_buf_1 _23903_ (.A(_10903_),
    .X(_05991_));
 sg13g2_mux2_1 _23904_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net972),
    .S(_05989_),
    .X(_01391_));
 sg13g2_buf_1 _23905_ (.A(_10925_),
    .X(_05992_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net971),
    .S(net247),
    .X(_01392_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net574),
    .S(_05988_),
    .X(_01393_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(_05948_),
    .S(_05988_),
    .X(_01394_));
 sg13g2_buf_1 _23909_ (.A(net517),
    .X(_05993_));
 sg13g2_nor2_1 _23910_ (.A(_05902_),
    .B(_05986_),
    .Y(_05994_));
 sg13g2_buf_1 _23911_ (.A(_05994_),
    .X(_05995_));
 sg13g2_buf_1 _23912_ (.A(_05995_),
    .X(_05996_));
 sg13g2_mux2_1 _23913_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net443),
    .S(net246),
    .X(_01395_));
 sg13g2_mux2_1 _23914_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net496),
    .S(net246),
    .X(_01396_));
 sg13g2_buf_1 _23915_ (.A(_09558_),
    .X(_05997_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net723),
    .S(net246),
    .X(_01397_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net573),
    .S(net246),
    .X(_01398_));
 sg13g2_mux2_1 _23918_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net839),
    .S(net246),
    .X(_01399_));
 sg13g2_mux2_1 _23919_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net838),
    .S(net246),
    .X(_01400_));
 sg13g2_mux2_1 _23920_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net837),
    .S(net246),
    .X(_01401_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net973),
    .S(_05996_),
    .X(_01402_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net972),
    .S(_05996_),
    .X(_01403_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net971),
    .S(net246),
    .X(_01404_));
 sg13g2_buf_1 _23924_ (.A(_11413_),
    .X(_05998_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net572),
    .S(_05995_),
    .X(_01405_));
 sg13g2_buf_1 _23926_ (.A(_09710_),
    .X(_05999_));
 sg13g2_mux2_1 _23927_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net644),
    .S(_05995_),
    .X(_01406_));
 sg13g2_nor3_1 _23928_ (.A(net727),
    .B(_05864_),
    .C(_05876_),
    .Y(_06000_));
 sg13g2_buf_1 _23929_ (.A(_06000_),
    .X(_06001_));
 sg13g2_buf_1 _23930_ (.A(_06001_),
    .X(_06002_));
 sg13g2_mux2_1 _23931_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net443),
    .S(net318),
    .X(_01407_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(_05973_),
    .S(net318),
    .X(_01408_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(net723),
    .S(net318),
    .X(_01409_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05963_),
    .S(net318),
    .X(_01410_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(_05969_),
    .S(net318),
    .X(_01411_));
 sg13g2_mux2_1 _23936_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net838),
    .S(net318),
    .X(_01412_));
 sg13g2_mux2_1 _23937_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net837),
    .S(_06002_),
    .X(_01413_));
 sg13g2_mux2_1 _23938_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(net973),
    .S(net318),
    .X(_01414_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(net972),
    .S(_06002_),
    .X(_01415_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net971),
    .S(net318),
    .X(_01416_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(net572),
    .S(_06001_),
    .X(_01417_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net644),
    .S(_06001_),
    .X(_01418_));
 sg13g2_nor3_1 _23943_ (.A(_05878_),
    .B(net445),
    .C(_05986_),
    .Y(_06003_));
 sg13g2_buf_1 _23944_ (.A(_06003_),
    .X(_06004_));
 sg13g2_buf_1 _23945_ (.A(_06004_),
    .X(_06005_));
 sg13g2_mux2_1 _23946_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net443),
    .S(net317),
    .X(_01419_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net496),
    .S(net317),
    .X(_01420_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net723),
    .S(net317),
    .X(_01421_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(net573),
    .S(net317),
    .X(_01422_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net839),
    .S(net317),
    .X(_01423_));
 sg13g2_mux2_1 _23951_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net838),
    .S(net317),
    .X(_01424_));
 sg13g2_mux2_1 _23952_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net837),
    .S(net317),
    .X(_01425_));
 sg13g2_mux2_1 _23953_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net973),
    .S(_06005_),
    .X(_01426_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(net972),
    .S(_06005_),
    .X(_01427_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net971),
    .S(net317),
    .X(_01428_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net572),
    .S(_06004_),
    .X(_01429_));
 sg13g2_mux2_1 _23957_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net644),
    .S(_06004_),
    .X(_01430_));
 sg13g2_nor3_1 _23958_ (.A(net845),
    .B(net445),
    .C(_05986_),
    .Y(_06006_));
 sg13g2_buf_1 _23959_ (.A(_06006_),
    .X(_06007_));
 sg13g2_buf_1 _23960_ (.A(_06007_),
    .X(_06008_));
 sg13g2_mux2_1 _23961_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net443),
    .S(net316),
    .X(_01431_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net496),
    .S(net316),
    .X(_01432_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net723),
    .S(net316),
    .X(_01433_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(net573),
    .S(net316),
    .X(_01434_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net839),
    .S(net316),
    .X(_01435_));
 sg13g2_mux2_1 _23966_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net838),
    .S(net316),
    .X(_01436_));
 sg13g2_mux2_1 _23967_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net837),
    .S(net316),
    .X(_01437_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net973),
    .S(_06008_),
    .X(_01438_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net972),
    .S(_06008_),
    .X(_01439_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net971),
    .S(net316),
    .X(_01440_));
 sg13g2_mux2_1 _23971_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net572),
    .S(_06007_),
    .X(_01441_));
 sg13g2_mux2_1 _23972_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net644),
    .S(_06007_),
    .X(_01442_));
 sg13g2_nor3_1 _23973_ (.A(_05843_),
    .B(_05864_),
    .C(_05906_),
    .Y(_06009_));
 sg13g2_buf_1 _23974_ (.A(_06009_),
    .X(_06010_));
 sg13g2_buf_1 _23975_ (.A(_06010_),
    .X(_06011_));
 sg13g2_mux2_1 _23976_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net443),
    .S(net315),
    .X(_01443_));
 sg13g2_mux2_1 _23977_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net496),
    .S(net315),
    .X(_01444_));
 sg13g2_mux2_1 _23978_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(net723),
    .S(net315),
    .X(_01445_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net592),
    .S(_06011_),
    .X(_01446_));
 sg13g2_mux2_1 _23980_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(_05969_),
    .S(net315),
    .X(_01447_));
 sg13g2_mux2_1 _23981_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net838),
    .S(net315),
    .X(_01448_));
 sg13g2_mux2_1 _23982_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net837),
    .S(net315),
    .X(_01449_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net973),
    .S(net315),
    .X(_01450_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net972),
    .S(_06011_),
    .X(_01451_));
 sg13g2_mux2_1 _23985_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net971),
    .S(net315),
    .X(_01452_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net572),
    .S(_06010_),
    .X(_01453_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(net644),
    .S(_06010_),
    .X(_01454_));
 sg13g2_nand2_2 _23988_ (.Y(_06012_),
    .A(_10872_),
    .B(_05863_));
 sg13g2_nor2_1 _23989_ (.A(_05868_),
    .B(_06012_),
    .Y(_06013_));
 sg13g2_buf_1 _23990_ (.A(_06013_),
    .X(_06014_));
 sg13g2_buf_1 _23991_ (.A(_06014_),
    .X(_06015_));
 sg13g2_mux2_1 _23992_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net443),
    .S(net245),
    .X(_01455_));
 sg13g2_mux2_1 _23993_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(_05973_),
    .S(net245),
    .X(_01456_));
 sg13g2_mux2_1 _23994_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net723),
    .S(net245),
    .X(_01457_));
 sg13g2_mux2_1 _23995_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net592),
    .S(_06015_),
    .X(_01458_));
 sg13g2_mux2_1 _23996_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net857),
    .S(net245),
    .X(_01459_));
 sg13g2_mux2_1 _23997_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(_05983_),
    .S(net245),
    .X(_01460_));
 sg13g2_mux2_1 _23998_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net837),
    .S(net245),
    .X(_01461_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net973),
    .S(net245),
    .X(_01462_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net972),
    .S(_06015_),
    .X(_01463_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net971),
    .S(net245),
    .X(_01464_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net572),
    .S(_06014_),
    .X(_01465_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05999_),
    .S(_06014_),
    .X(_01466_));
 sg13g2_nor2_1 _24004_ (.A(_05900_),
    .B(_06012_),
    .Y(_06016_));
 sg13g2_buf_2 _24005_ (.A(_06016_),
    .X(_06017_));
 sg13g2_nor2b_1 _24006_ (.A(_05876_),
    .B_N(_06017_),
    .Y(_06018_));
 sg13g2_buf_1 _24007_ (.A(_06018_),
    .X(_06019_));
 sg13g2_buf_1 _24008_ (.A(_06019_),
    .X(_06020_));
 sg13g2_mux2_1 _24009_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net443),
    .S(net314),
    .X(_01467_));
 sg13g2_mux2_1 _24010_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net520),
    .S(net314),
    .X(_01468_));
 sg13g2_mux2_1 _24011_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net723),
    .S(net314),
    .X(_01469_));
 sg13g2_mux2_1 _24012_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net592),
    .S(net314),
    .X(_01470_));
 sg13g2_mux2_1 _24013_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net857),
    .S(net314),
    .X(_01471_));
 sg13g2_mux2_1 _24014_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net838),
    .S(net314),
    .X(_01472_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(_05984_),
    .S(net314),
    .X(_01473_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net973),
    .S(_06020_),
    .X(_01474_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net972),
    .S(_06020_),
    .X(_01475_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net971),
    .S(net314),
    .X(_01476_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(_05998_),
    .S(_06019_),
    .X(_01477_));
 sg13g2_mux2_1 _24020_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net644),
    .S(_06019_),
    .X(_01478_));
 sg13g2_nor2_2 _24021_ (.A(net982),
    .B(_05827_),
    .Y(_06021_));
 sg13g2_nand2_2 _24022_ (.Y(_06022_),
    .A(net981),
    .B(_06021_));
 sg13g2_nor3_2 _24023_ (.A(net974),
    .B(net978),
    .C(_06022_),
    .Y(_06023_));
 sg13g2_nor2b_1 _24024_ (.A(net446),
    .B_N(_06023_),
    .Y(_06024_));
 sg13g2_buf_1 _24025_ (.A(_06024_),
    .X(_06025_));
 sg13g2_buf_1 _24026_ (.A(_06025_),
    .X(_06026_));
 sg13g2_mux2_1 _24027_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(_05993_),
    .S(net313),
    .X(_01479_));
 sg13g2_mux2_1 _24028_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(net520),
    .S(net313),
    .X(_01480_));
 sg13g2_mux2_1 _24029_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(_05997_),
    .S(net313),
    .X(_01481_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net592),
    .S(net313),
    .X(_01482_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net857),
    .S(net313),
    .X(_01483_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(_05983_),
    .S(net313),
    .X(_01484_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(_05984_),
    .S(net313),
    .X(_01485_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_05990_),
    .S(_06026_),
    .X(_01486_));
 sg13g2_mux2_1 _24035_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(_05991_),
    .S(_06026_),
    .X(_01487_));
 sg13g2_mux2_1 _24036_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(_05992_),
    .S(net313),
    .X(_01488_));
 sg13g2_mux2_1 _24037_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net572),
    .S(_06025_),
    .X(_01489_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net644),
    .S(_06025_),
    .X(_01490_));
 sg13g2_nor2b_1 _24039_ (.A(_05855_),
    .B_N(_05863_),
    .Y(_06027_));
 sg13g2_buf_2 _24040_ (.A(_06027_),
    .X(_06028_));
 sg13g2_nor2b_1 _24041_ (.A(net446),
    .B_N(_06028_),
    .Y(_06029_));
 sg13g2_buf_1 _24042_ (.A(_06029_),
    .X(_06030_));
 sg13g2_buf_1 _24043_ (.A(_06030_),
    .X(_06031_));
 sg13g2_mux2_1 _24044_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_05993_),
    .S(net312),
    .X(_01491_));
 sg13g2_mux2_1 _24045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net520),
    .S(net312),
    .X(_01492_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net723),
    .S(net312),
    .X(_01493_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net592),
    .S(net312),
    .X(_01494_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net857),
    .S(net312),
    .X(_01495_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net862),
    .S(net312),
    .X(_01496_));
 sg13g2_mux2_1 _24050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net861),
    .S(_06031_),
    .X(_01497_));
 sg13g2_mux2_1 _24051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(_05990_),
    .S(net312),
    .X(_01498_));
 sg13g2_mux2_1 _24052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(_05991_),
    .S(_06031_),
    .X(_01499_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(_05992_),
    .S(net312),
    .X(_01500_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net572),
    .S(_06030_),
    .X(_01501_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net644),
    .S(_06030_),
    .X(_01502_));
 sg13g2_nor3_1 _24056_ (.A(net445),
    .B(_05880_),
    .C(_05917_),
    .Y(_06032_));
 sg13g2_buf_1 _24057_ (.A(_06032_),
    .X(_06033_));
 sg13g2_buf_1 _24058_ (.A(_06033_),
    .X(_06034_));
 sg13g2_mux2_1 _24059_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(net443),
    .S(net311),
    .X(_01503_));
 sg13g2_mux2_1 _24060_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(_03528_),
    .S(net311),
    .X(_01504_));
 sg13g2_mux2_1 _24061_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_05997_),
    .S(net311),
    .X(_01505_));
 sg13g2_mux2_1 _24062_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_03038_),
    .S(net311),
    .X(_01506_));
 sg13g2_mux2_1 _24063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(_03042_),
    .S(net311),
    .X(_01507_));
 sg13g2_mux2_1 _24064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(net862),
    .S(net311),
    .X(_01508_));
 sg13g2_mux2_1 _24065_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net861),
    .S(net311),
    .X(_01509_));
 sg13g2_mux2_1 _24066_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net993),
    .S(net311),
    .X(_01510_));
 sg13g2_mux2_1 _24067_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net992),
    .S(_06034_),
    .X(_01511_));
 sg13g2_mux2_1 _24068_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net991),
    .S(_06034_),
    .X(_01512_));
 sg13g2_mux2_1 _24069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(_05998_),
    .S(_06033_),
    .X(_01513_));
 sg13g2_mux2_1 _24070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_05999_),
    .S(_06033_),
    .X(_01514_));
 sg13g2_nor3_1 _24071_ (.A(net844),
    .B(_05880_),
    .C(_05902_),
    .Y(_06035_));
 sg13g2_buf_1 _24072_ (.A(_06035_),
    .X(_06036_));
 sg13g2_buf_1 _24073_ (.A(_06036_),
    .X(_06037_));
 sg13g2_mux2_1 _24074_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(_03535_),
    .S(net244),
    .X(_01515_));
 sg13g2_mux2_1 _24075_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_03528_),
    .S(net244),
    .X(_01516_));
 sg13g2_mux2_1 _24076_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(net907),
    .S(net244),
    .X(_01517_));
 sg13g2_mux2_1 _24077_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_03038_),
    .S(net244),
    .X(_01518_));
 sg13g2_mux2_1 _24078_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(_03042_),
    .S(net244),
    .X(_01519_));
 sg13g2_mux2_1 _24079_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_03028_),
    .S(net244),
    .X(_01520_));
 sg13g2_mux2_1 _24080_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(_03030_),
    .S(net244),
    .X(_01521_));
 sg13g2_mux2_1 _24081_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(_03032_),
    .S(_06037_),
    .X(_01522_));
 sg13g2_mux2_1 _24082_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_03034_),
    .S(net244),
    .X(_01523_));
 sg13g2_mux2_1 _24083_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_03036_),
    .S(_06037_),
    .X(_01524_));
 sg13g2_mux2_1 _24084_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_11413_),
    .S(_06036_),
    .X(_01525_));
 sg13g2_mux2_1 _24085_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(net776),
    .S(_06036_),
    .X(_01526_));
 sg13g2_and2_1 _24086_ (.A(_05861_),
    .B(_05863_),
    .X(_06038_));
 sg13g2_buf_1 _24087_ (.A(_06038_),
    .X(_06039_));
 sg13g2_and3_1 _24088_ (.X(_06040_),
    .A(net1151),
    .B(_10503_),
    .C(_05816_));
 sg13g2_buf_1 _24089_ (.A(_06040_),
    .X(_06041_));
 sg13g2_and2_1 _24090_ (.A(_05833_),
    .B(_06041_),
    .X(_06042_));
 sg13g2_buf_1 _24091_ (.A(_06042_),
    .X(_06043_));
 sg13g2_nand2_1 _24092_ (.Y(_06044_),
    .A(_06039_),
    .B(_06043_));
 sg13g2_buf_1 _24093_ (.A(_06044_),
    .X(_06045_));
 sg13g2_buf_1 _24094_ (.A(net310),
    .X(_06046_));
 sg13g2_nand2_1 _24095_ (.Y(_06047_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(net310));
 sg13g2_o21ai_1 _24096_ (.B1(_06047_),
    .Y(_01527_),
    .A1(net583),
    .A2(net243));
 sg13g2_mux2_1 _24097_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(_06046_),
    .X(_01528_));
 sg13g2_nand2_1 _24098_ (.Y(_06048_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(net310));
 sg13g2_o21ai_1 _24099_ (.B1(_06048_),
    .Y(_01529_),
    .A1(net584),
    .A2(net243));
 sg13g2_nand2_1 _24100_ (.Y(_06049_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(net310));
 sg13g2_o21ai_1 _24101_ (.B1(_06049_),
    .Y(_01530_),
    .A1(net657),
    .A2(net243));
 sg13g2_nand2_1 _24102_ (.Y(_06050_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .B(net310));
 sg13g2_o21ai_1 _24103_ (.B1(_06050_),
    .Y(_01531_),
    .A1(net743),
    .A2(net243));
 sg13g2_mux2_1 _24104_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .S(net243),
    .X(_01532_));
 sg13g2_mux2_1 _24105_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net243),
    .X(_01533_));
 sg13g2_mux2_1 _24106_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net243),
    .X(_01534_));
 sg13g2_mux2_1 _24107_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(_06045_),
    .X(_01535_));
 sg13g2_mux2_1 _24108_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net310),
    .X(_01536_));
 sg13g2_nand2_1 _24109_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .B(net310));
 sg13g2_o21ai_1 _24110_ (.B1(_06051_),
    .Y(_01537_),
    .A1(net655),
    .A2(_06046_));
 sg13g2_nand2_1 _24111_ (.Y(_06052_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .B(net310));
 sg13g2_o21ai_1 _24112_ (.B1(_06052_),
    .Y(_01538_),
    .A1(net731),
    .A2(net243));
 sg13g2_buf_1 _24113_ (.A(_06041_),
    .X(_06053_));
 sg13g2_nand2_1 _24114_ (.Y(_06054_),
    .A(_05881_),
    .B(net442));
 sg13g2_buf_1 _24115_ (.A(_06054_),
    .X(_06055_));
 sg13g2_buf_1 _24116_ (.A(net380),
    .X(_06056_));
 sg13g2_nand2_1 _24117_ (.Y(_06057_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(net380));
 sg13g2_o21ai_1 _24118_ (.B1(_06057_),
    .Y(_01539_),
    .A1(net583),
    .A2(net309));
 sg13g2_mux2_1 _24119_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(_06056_),
    .X(_01540_));
 sg13g2_nand2_1 _24120_ (.Y(_06058_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(net380));
 sg13g2_o21ai_1 _24121_ (.B1(_06058_),
    .Y(_01541_),
    .A1(net584),
    .A2(_06056_));
 sg13g2_nand2_1 _24122_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(net380));
 sg13g2_o21ai_1 _24123_ (.B1(_06059_),
    .Y(_01542_),
    .A1(net657),
    .A2(net309));
 sg13g2_nand2_1 _24124_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .B(net380));
 sg13g2_o21ai_1 _24125_ (.B1(_06060_),
    .Y(_01543_),
    .A1(net743),
    .A2(net309));
 sg13g2_mux2_1 _24126_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .S(net309),
    .X(_01544_));
 sg13g2_mux2_1 _24127_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net309),
    .X(_01545_));
 sg13g2_mux2_1 _24128_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net309),
    .X(_01546_));
 sg13g2_mux2_1 _24129_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net380),
    .X(_01547_));
 sg13g2_mux2_1 _24130_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net380),
    .X(_01548_));
 sg13g2_nand2_1 _24131_ (.Y(_06061_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .B(_06055_));
 sg13g2_o21ai_1 _24132_ (.B1(_06061_),
    .Y(_01549_),
    .A1(net655),
    .A2(net309));
 sg13g2_nand2_1 _24133_ (.Y(_06062_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .B(net380));
 sg13g2_o21ai_1 _24134_ (.B1(_06062_),
    .Y(_01550_),
    .A1(net731),
    .A2(net309));
 sg13g2_nand2_1 _24135_ (.Y(_06063_),
    .A(_05889_),
    .B(net442));
 sg13g2_buf_1 _24136_ (.A(_06063_),
    .X(_06064_));
 sg13g2_buf_1 _24137_ (.A(net379),
    .X(_06065_));
 sg13g2_nand2_1 _24138_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(net379));
 sg13g2_o21ai_1 _24139_ (.B1(_06066_),
    .Y(_01551_),
    .A1(net583),
    .A2(net308));
 sg13g2_mux2_1 _24140_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(_06065_),
    .X(_01552_));
 sg13g2_nand2_1 _24141_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(net379));
 sg13g2_o21ai_1 _24142_ (.B1(_06067_),
    .Y(_01553_),
    .A1(net584),
    .A2(_06065_));
 sg13g2_nand2_1 _24143_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(net379));
 sg13g2_o21ai_1 _24144_ (.B1(_06068_),
    .Y(_01554_),
    .A1(net657),
    .A2(net308));
 sg13g2_nand2_1 _24145_ (.Y(_06069_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .B(net379));
 sg13g2_o21ai_1 _24146_ (.B1(_06069_),
    .Y(_01555_),
    .A1(net743),
    .A2(net308));
 sg13g2_mux2_1 _24147_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S(net308),
    .X(_01556_));
 sg13g2_mux2_1 _24148_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net308),
    .X(_01557_));
 sg13g2_mux2_1 _24149_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net308),
    .X(_01558_));
 sg13g2_mux2_1 _24150_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net379),
    .X(_01559_));
 sg13g2_mux2_1 _24151_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net379),
    .X(_01560_));
 sg13g2_nand2_1 _24152_ (.Y(_06070_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .B(_06064_));
 sg13g2_o21ai_1 _24153_ (.B1(_06070_),
    .Y(_01561_),
    .A1(net655),
    .A2(net308));
 sg13g2_nand2_1 _24154_ (.Y(_06071_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .B(net379));
 sg13g2_o21ai_1 _24155_ (.B1(_06071_),
    .Y(_01562_),
    .A1(net731),
    .A2(net308));
 sg13g2_nor2_2 _24156_ (.A(_05861_),
    .B(_05880_),
    .Y(_06072_));
 sg13g2_nand2_1 _24157_ (.Y(_06073_),
    .A(_06072_),
    .B(_06043_));
 sg13g2_buf_1 _24158_ (.A(_06073_),
    .X(_06074_));
 sg13g2_buf_1 _24159_ (.A(net307),
    .X(_06075_));
 sg13g2_nand2_1 _24160_ (.Y(_06076_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(net307));
 sg13g2_o21ai_1 _24161_ (.B1(_06076_),
    .Y(_01563_),
    .A1(net583),
    .A2(net242));
 sg13g2_mux2_1 _24162_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net242),
    .X(_01564_));
 sg13g2_nand2_1 _24163_ (.Y(_06077_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(net307));
 sg13g2_o21ai_1 _24164_ (.B1(_06077_),
    .Y(_01565_),
    .A1(net584),
    .A2(net242));
 sg13g2_nand2_1 _24165_ (.Y(_06078_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(net307));
 sg13g2_o21ai_1 _24166_ (.B1(_06078_),
    .Y(_01566_),
    .A1(net657),
    .A2(net242));
 sg13g2_nand2_1 _24167_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .B(net307));
 sg13g2_o21ai_1 _24168_ (.B1(_06079_),
    .Y(_01567_),
    .A1(net743),
    .A2(net242));
 sg13g2_mux2_1 _24169_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .S(net242),
    .X(_01568_));
 sg13g2_mux2_1 _24170_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net242),
    .X(_01569_));
 sg13g2_mux2_1 _24171_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net242),
    .X(_01570_));
 sg13g2_mux2_1 _24172_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net307),
    .X(_01571_));
 sg13g2_mux2_1 _24173_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net307),
    .X(_01572_));
 sg13g2_nand2_1 _24174_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .B(_06074_));
 sg13g2_o21ai_1 _24175_ (.B1(_06080_),
    .Y(_01573_),
    .A1(net655),
    .A2(_06075_));
 sg13g2_nand2_1 _24176_ (.Y(_06081_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .B(net307));
 sg13g2_o21ai_1 _24177_ (.B1(_06081_),
    .Y(_01574_),
    .A1(net731),
    .A2(_06075_));
 sg13g2_nor2b_1 _24178_ (.A(_05900_),
    .B_N(_06041_),
    .Y(_06082_));
 sg13g2_buf_2 _24179_ (.A(_06082_),
    .X(_06083_));
 sg13g2_nand2_1 _24180_ (.Y(_06084_),
    .A(_06072_),
    .B(_06083_));
 sg13g2_buf_1 _24181_ (.A(_06084_),
    .X(_06085_));
 sg13g2_buf_1 _24182_ (.A(net306),
    .X(_06086_));
 sg13g2_nand2_1 _24183_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(net306));
 sg13g2_o21ai_1 _24184_ (.B1(_06087_),
    .Y(_01575_),
    .A1(net583),
    .A2(net241));
 sg13g2_mux2_1 _24185_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net241),
    .X(_01576_));
 sg13g2_nand2_1 _24186_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(net306));
 sg13g2_o21ai_1 _24187_ (.B1(_06088_),
    .Y(_01577_),
    .A1(net584),
    .A2(net241));
 sg13g2_nand2_1 _24188_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(net306));
 sg13g2_o21ai_1 _24189_ (.B1(_06089_),
    .Y(_01578_),
    .A1(net657),
    .A2(net241));
 sg13g2_nand2_1 _24190_ (.Y(_06090_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .B(net306));
 sg13g2_o21ai_1 _24191_ (.B1(_06090_),
    .Y(_01579_),
    .A1(net743),
    .A2(net241));
 sg13g2_mux2_1 _24192_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .S(net241),
    .X(_01580_));
 sg13g2_mux2_1 _24193_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net241),
    .X(_01581_));
 sg13g2_mux2_1 _24194_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net241),
    .X(_01582_));
 sg13g2_mux2_1 _24195_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net306),
    .X(_01583_));
 sg13g2_mux2_1 _24196_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net306),
    .X(_01584_));
 sg13g2_nand2_1 _24197_ (.Y(_06091_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .B(_06085_));
 sg13g2_o21ai_1 _24198_ (.B1(_06091_),
    .Y(_01585_),
    .A1(net655),
    .A2(_06086_));
 sg13g2_nand2_1 _24199_ (.Y(_06092_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .B(net306));
 sg13g2_o21ai_1 _24200_ (.B1(_06092_),
    .Y(_01586_),
    .A1(net731),
    .A2(_06086_));
 sg13g2_nand3_1 _24201_ (.B(_06072_),
    .C(_06053_),
    .A(_06021_),
    .Y(_06093_));
 sg13g2_buf_1 _24202_ (.A(_06093_),
    .X(_06094_));
 sg13g2_buf_1 _24203_ (.A(net378),
    .X(_06095_));
 sg13g2_nand2_1 _24204_ (.Y(_06096_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(net378));
 sg13g2_o21ai_1 _24205_ (.B1(_06096_),
    .Y(_01587_),
    .A1(net583),
    .A2(net305));
 sg13g2_mux2_1 _24206_ (.A0(_03782_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net305),
    .X(_01588_));
 sg13g2_nand2_1 _24207_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(net378));
 sg13g2_o21ai_1 _24208_ (.B1(_06097_),
    .Y(_01589_),
    .A1(net584),
    .A2(net305));
 sg13g2_nand2_1 _24209_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(net378));
 sg13g2_o21ai_1 _24210_ (.B1(_06098_),
    .Y(_01590_),
    .A1(net657),
    .A2(net305));
 sg13g2_nand2_1 _24211_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .B(net378));
 sg13g2_o21ai_1 _24212_ (.B1(_06099_),
    .Y(_01591_),
    .A1(net743),
    .A2(net305));
 sg13g2_mux2_1 _24213_ (.A0(net742),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .S(net305),
    .X(_01592_));
 sg13g2_mux2_1 _24214_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net305),
    .X(_01593_));
 sg13g2_mux2_1 _24215_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net305),
    .X(_01594_));
 sg13g2_mux2_1 _24216_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net378),
    .X(_01595_));
 sg13g2_mux2_1 _24217_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net378),
    .X(_01596_));
 sg13g2_nand2_1 _24218_ (.Y(_06100_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .B(_06094_));
 sg13g2_o21ai_1 _24219_ (.B1(_06100_),
    .Y(_01597_),
    .A1(net655),
    .A2(_06095_));
 sg13g2_nand2_1 _24220_ (.Y(_06101_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .B(net378));
 sg13g2_o21ai_1 _24221_ (.B1(_06101_),
    .Y(_01598_),
    .A1(_03780_),
    .A2(_06095_));
 sg13g2_buf_1 _24222_ (.A(_06041_),
    .X(_06102_));
 sg13g2_nand3_1 _24223_ (.B(_06072_),
    .C(net441),
    .A(_05831_),
    .Y(_06103_));
 sg13g2_buf_1 _24224_ (.A(_06103_),
    .X(_06104_));
 sg13g2_buf_1 _24225_ (.A(net377),
    .X(_06105_));
 sg13g2_nand2_1 _24226_ (.Y(_06106_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(net377));
 sg13g2_o21ai_1 _24227_ (.B1(_06106_),
    .Y(_01599_),
    .A1(net583),
    .A2(net304));
 sg13g2_mux2_1 _24228_ (.A0(_03782_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net304),
    .X(_01600_));
 sg13g2_nand2_1 _24229_ (.Y(_06107_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(net377));
 sg13g2_o21ai_1 _24230_ (.B1(_06107_),
    .Y(_01601_),
    .A1(net584),
    .A2(net304));
 sg13g2_buf_1 _24231_ (.A(_03019_),
    .X(_06108_));
 sg13g2_nand2_1 _24232_ (.Y(_06109_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(net377));
 sg13g2_o21ai_1 _24233_ (.B1(_06109_),
    .Y(_01602_),
    .A1(_06108_),
    .A2(net304));
 sg13g2_buf_1 _24234_ (.A(net863),
    .X(_06110_));
 sg13g2_nand2_1 _24235_ (.Y(_06111_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .B(net377));
 sg13g2_o21ai_1 _24236_ (.B1(_06111_),
    .Y(_01603_),
    .A1(_06110_),
    .A2(net304));
 sg13g2_buf_1 _24237_ (.A(net862),
    .X(_06112_));
 sg13g2_mux2_1 _24238_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S(net304),
    .X(_01604_));
 sg13g2_buf_1 _24239_ (.A(net861),
    .X(_06113_));
 sg13g2_mux2_1 _24240_ (.A0(_06113_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net304),
    .X(_01605_));
 sg13g2_buf_1 _24241_ (.A(net993),
    .X(_06114_));
 sg13g2_mux2_1 _24242_ (.A0(_06114_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net304),
    .X(_01606_));
 sg13g2_buf_1 _24243_ (.A(net992),
    .X(_06115_));
 sg13g2_mux2_1 _24244_ (.A0(_06115_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(net377),
    .X(_01607_));
 sg13g2_buf_1 _24245_ (.A(net991),
    .X(_06116_));
 sg13g2_mux2_1 _24246_ (.A0(_06116_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net377),
    .X(_01608_));
 sg13g2_nand2_1 _24247_ (.Y(_06117_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .B(net377));
 sg13g2_o21ai_1 _24248_ (.B1(_06117_),
    .Y(_01609_),
    .A1(net655),
    .A2(_06105_));
 sg13g2_nand2_1 _24249_ (.Y(_06118_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .B(_06104_));
 sg13g2_o21ai_1 _24250_ (.B1(_06118_),
    .Y(_01610_),
    .A1(_03780_),
    .A2(_06105_));
 sg13g2_nor3_2 _24251_ (.A(net982),
    .B(net1126),
    .C(_05841_),
    .Y(_06119_));
 sg13g2_nand4_1 _24252_ (.B(net980),
    .C(_06119_),
    .A(net974),
    .Y(_06120_),
    .D(net441));
 sg13g2_buf_1 _24253_ (.A(_06120_),
    .X(_06121_));
 sg13g2_buf_1 _24254_ (.A(_06121_),
    .X(_06122_));
 sg13g2_nand2_1 _24255_ (.Y(_06123_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(net376));
 sg13g2_o21ai_1 _24256_ (.B1(_06123_),
    .Y(_01611_),
    .A1(net583),
    .A2(net303));
 sg13g2_mux2_1 _24257_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(_06122_),
    .X(_01612_));
 sg13g2_nand2_1 _24258_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(net376));
 sg13g2_o21ai_1 _24259_ (.B1(_06124_),
    .Y(_01613_),
    .A1(net584),
    .A2(net303));
 sg13g2_nand2_1 _24260_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(net376));
 sg13g2_o21ai_1 _24261_ (.B1(_06125_),
    .Y(_01614_),
    .A1(net643),
    .A2(net303));
 sg13g2_nand2_1 _24262_ (.Y(_06126_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .B(net376));
 sg13g2_o21ai_1 _24263_ (.B1(_06126_),
    .Y(_01615_),
    .A1(net722),
    .A2(net303));
 sg13g2_mux2_1 _24264_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .S(net303),
    .X(_01616_));
 sg13g2_mux2_1 _24265_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net303),
    .X(_01617_));
 sg13g2_mux2_1 _24266_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net303),
    .X(_01618_));
 sg13g2_mux2_1 _24267_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net376),
    .X(_01619_));
 sg13g2_mux2_1 _24268_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(net376),
    .X(_01620_));
 sg13g2_nand2_1 _24269_ (.Y(_06127_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .B(net376));
 sg13g2_o21ai_1 _24270_ (.B1(_06127_),
    .Y(_01621_),
    .A1(net655),
    .A2(_06122_));
 sg13g2_nand2_1 _24271_ (.Y(_06128_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .B(net376));
 sg13g2_o21ai_1 _24272_ (.B1(_06128_),
    .Y(_01622_),
    .A1(net731),
    .A2(net303));
 sg13g2_buf_1 _24273_ (.A(net653),
    .X(_06129_));
 sg13g2_nand4_1 _24274_ (.B(_05839_),
    .C(net980),
    .A(net974),
    .Y(_06130_),
    .D(_06083_));
 sg13g2_buf_1 _24275_ (.A(_06130_),
    .X(_06131_));
 sg13g2_buf_1 _24276_ (.A(net302),
    .X(_06132_));
 sg13g2_nand2_1 _24277_ (.Y(_06133_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(net302));
 sg13g2_o21ai_1 _24278_ (.B1(_06133_),
    .Y(_01623_),
    .A1(net571),
    .A2(net240));
 sg13g2_buf_1 _24279_ (.A(net520),
    .X(_06134_));
 sg13g2_mux2_1 _24280_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(_06132_),
    .X(_01624_));
 sg13g2_buf_1 _24281_ (.A(net666),
    .X(_06135_));
 sg13g2_nand2_1 _24282_ (.Y(_06136_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(_06131_));
 sg13g2_o21ai_1 _24283_ (.B1(_06136_),
    .Y(_01625_),
    .A1(net570),
    .A2(_06132_));
 sg13g2_nand2_1 _24284_ (.Y(_06137_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(net302));
 sg13g2_o21ai_1 _24285_ (.B1(_06137_),
    .Y(_01626_),
    .A1(net643),
    .A2(net240));
 sg13g2_nand2_1 _24286_ (.Y(_06138_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .B(net302));
 sg13g2_o21ai_1 _24287_ (.B1(_06138_),
    .Y(_01627_),
    .A1(net722),
    .A2(net240));
 sg13g2_mux2_1 _24288_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .S(net240),
    .X(_01628_));
 sg13g2_mux2_1 _24289_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net240),
    .X(_01629_));
 sg13g2_mux2_1 _24290_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net240),
    .X(_01630_));
 sg13g2_mux2_1 _24291_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net302),
    .X(_01631_));
 sg13g2_mux2_1 _24292_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(net302),
    .X(_01632_));
 sg13g2_buf_1 _24293_ (.A(net749),
    .X(_06139_));
 sg13g2_nand2_1 _24294_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .B(net302));
 sg13g2_o21ai_1 _24295_ (.B1(_06140_),
    .Y(_01633_),
    .A1(net642),
    .A2(net240));
 sg13g2_buf_1 _24296_ (.A(net875),
    .X(_06141_));
 sg13g2_nand2_1 _24297_ (.Y(_06142_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .B(net302));
 sg13g2_o21ai_1 _24298_ (.B1(_06142_),
    .Y(_01634_),
    .A1(net719),
    .A2(net240));
 sg13g2_nand2_1 _24299_ (.Y(_06143_),
    .A(_05928_),
    .B(net442));
 sg13g2_buf_1 _24300_ (.A(_06143_),
    .X(_06144_));
 sg13g2_buf_1 _24301_ (.A(net375),
    .X(_06145_));
 sg13g2_nand2_1 _24302_ (.Y(_06146_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(net375));
 sg13g2_o21ai_1 _24303_ (.B1(_06146_),
    .Y(_01635_),
    .A1(net571),
    .A2(net301));
 sg13g2_mux2_1 _24304_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(_06145_),
    .X(_01636_));
 sg13g2_nand2_1 _24305_ (.Y(_06147_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24306_ (.B1(_06147_),
    .Y(_01637_),
    .A1(net570),
    .A2(_06145_));
 sg13g2_nand2_1 _24307_ (.Y(_06148_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(net375));
 sg13g2_o21ai_1 _24308_ (.B1(_06148_),
    .Y(_01638_),
    .A1(net643),
    .A2(net301));
 sg13g2_nand2_1 _24309_ (.Y(_06149_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .B(net375));
 sg13g2_o21ai_1 _24310_ (.B1(_06149_),
    .Y(_01639_),
    .A1(net722),
    .A2(net301));
 sg13g2_mux2_1 _24311_ (.A0(_06112_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .S(net301),
    .X(_01640_));
 sg13g2_mux2_1 _24312_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net301),
    .X(_01641_));
 sg13g2_mux2_1 _24313_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net301),
    .X(_01642_));
 sg13g2_mux2_1 _24314_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net375),
    .X(_01643_));
 sg13g2_mux2_1 _24315_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(net375),
    .X(_01644_));
 sg13g2_nand2_1 _24316_ (.Y(_06150_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .B(net375));
 sg13g2_o21ai_1 _24317_ (.B1(_06150_),
    .Y(_01645_),
    .A1(net642),
    .A2(net301));
 sg13g2_nand2_1 _24318_ (.Y(_06151_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .B(net375));
 sg13g2_o21ai_1 _24319_ (.B1(_06151_),
    .Y(_01646_),
    .A1(net719),
    .A2(net301));
 sg13g2_nand2_1 _24320_ (.Y(_06152_),
    .A(_05935_),
    .B(net442));
 sg13g2_buf_1 _24321_ (.A(_06152_),
    .X(_06153_));
 sg13g2_buf_1 _24322_ (.A(_06153_),
    .X(_06154_));
 sg13g2_nand2_1 _24323_ (.Y(_06155_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(net374));
 sg13g2_o21ai_1 _24324_ (.B1(_06155_),
    .Y(_01647_),
    .A1(_06129_),
    .A2(net300));
 sg13g2_mux2_1 _24325_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(_06154_),
    .X(_01648_));
 sg13g2_nand2_1 _24326_ (.Y(_06156_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(net374));
 sg13g2_o21ai_1 _24327_ (.B1(_06156_),
    .Y(_01649_),
    .A1(_06135_),
    .A2(_06154_));
 sg13g2_nand2_1 _24328_ (.Y(_06157_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(net374));
 sg13g2_o21ai_1 _24329_ (.B1(_06157_),
    .Y(_01650_),
    .A1(net643),
    .A2(net300));
 sg13g2_nand2_1 _24330_ (.Y(_06158_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .B(net374));
 sg13g2_o21ai_1 _24331_ (.B1(_06158_),
    .Y(_01651_),
    .A1(net722),
    .A2(net300));
 sg13g2_mux2_1 _24332_ (.A0(_06112_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S(net300),
    .X(_01652_));
 sg13g2_mux2_1 _24333_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net300),
    .X(_01653_));
 sg13g2_mux2_1 _24334_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net300),
    .X(_01654_));
 sg13g2_mux2_1 _24335_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net374),
    .X(_01655_));
 sg13g2_mux2_1 _24336_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net374),
    .X(_01656_));
 sg13g2_nand2_1 _24337_ (.Y(_06159_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .B(net374));
 sg13g2_o21ai_1 _24338_ (.B1(_06159_),
    .Y(_01657_),
    .A1(_06139_),
    .A2(net300));
 sg13g2_nand2_1 _24339_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .B(net374));
 sg13g2_o21ai_1 _24340_ (.B1(_06160_),
    .Y(_01658_),
    .A1(_06141_),
    .A2(net300));
 sg13g2_nand2_1 _24341_ (.Y(_06161_),
    .A(_06039_),
    .B(_06083_));
 sg13g2_buf_1 _24342_ (.A(_06161_),
    .X(_06162_));
 sg13g2_buf_1 _24343_ (.A(net299),
    .X(_06163_));
 sg13g2_nand2_1 _24344_ (.Y(_06164_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(net299));
 sg13g2_o21ai_1 _24345_ (.B1(_06164_),
    .Y(_01659_),
    .A1(_06129_),
    .A2(net239));
 sg13g2_mux2_1 _24346_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(_06163_),
    .X(_01660_));
 sg13g2_nand2_1 _24347_ (.Y(_06165_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(net299));
 sg13g2_o21ai_1 _24348_ (.B1(_06165_),
    .Y(_01661_),
    .A1(_06135_),
    .A2(net239));
 sg13g2_nand2_1 _24349_ (.Y(_06166_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(net299));
 sg13g2_o21ai_1 _24350_ (.B1(_06166_),
    .Y(_01662_),
    .A1(_06108_),
    .A2(net239));
 sg13g2_nand2_1 _24351_ (.Y(_06167_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .B(net299));
 sg13g2_o21ai_1 _24352_ (.B1(_06167_),
    .Y(_01663_),
    .A1(_06110_),
    .A2(net239));
 sg13g2_mux2_1 _24353_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .S(net239),
    .X(_01664_));
 sg13g2_mux2_1 _24354_ (.A0(_06113_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net239),
    .X(_01665_));
 sg13g2_mux2_1 _24355_ (.A0(_06114_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net239),
    .X(_01666_));
 sg13g2_mux2_1 _24356_ (.A0(_06115_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net299),
    .X(_01667_));
 sg13g2_mux2_1 _24357_ (.A0(_06116_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(_06162_),
    .X(_01668_));
 sg13g2_nand2_1 _24358_ (.Y(_06168_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .B(net299));
 sg13g2_o21ai_1 _24359_ (.B1(_06168_),
    .Y(_01669_),
    .A1(_06139_),
    .A2(_06163_));
 sg13g2_nand2_1 _24360_ (.Y(_06169_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .B(net299));
 sg13g2_o21ai_1 _24361_ (.B1(_06169_),
    .Y(_01670_),
    .A1(_06141_),
    .A2(net239));
 sg13g2_nor2_2 _24362_ (.A(_05861_),
    .B(_05916_),
    .Y(_06170_));
 sg13g2_nand2_1 _24363_ (.Y(_06171_),
    .A(_06170_),
    .B(_06043_));
 sg13g2_buf_1 _24364_ (.A(_06171_),
    .X(_06172_));
 sg13g2_buf_1 _24365_ (.A(net298),
    .X(_06173_));
 sg13g2_nand2_1 _24366_ (.Y(_06174_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(net298));
 sg13g2_o21ai_1 _24367_ (.B1(_06174_),
    .Y(_01671_),
    .A1(net571),
    .A2(net238));
 sg13g2_mux2_1 _24368_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(_06173_),
    .X(_01672_));
 sg13g2_nand2_1 _24369_ (.Y(_06175_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(net298));
 sg13g2_o21ai_1 _24370_ (.B1(_06175_),
    .Y(_01673_),
    .A1(net570),
    .A2(_06173_));
 sg13g2_nand2_1 _24371_ (.Y(_06176_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(net298));
 sg13g2_o21ai_1 _24372_ (.B1(_06176_),
    .Y(_01674_),
    .A1(net643),
    .A2(net238));
 sg13g2_nand2_1 _24373_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .B(net298));
 sg13g2_o21ai_1 _24374_ (.B1(_06177_),
    .Y(_01675_),
    .A1(net722),
    .A2(net238));
 sg13g2_mux2_1 _24375_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .S(net238),
    .X(_01676_));
 sg13g2_mux2_1 _24376_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net238),
    .X(_01677_));
 sg13g2_mux2_1 _24377_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(net238),
    .X(_01678_));
 sg13g2_mux2_1 _24378_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net298),
    .X(_01679_));
 sg13g2_mux2_1 _24379_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(_06172_),
    .X(_01680_));
 sg13g2_nand2_1 _24380_ (.Y(_06178_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .B(net298));
 sg13g2_o21ai_1 _24381_ (.B1(_06178_),
    .Y(_01681_),
    .A1(net642),
    .A2(net238));
 sg13g2_nand2_1 _24382_ (.Y(_06179_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .B(net298));
 sg13g2_o21ai_1 _24383_ (.B1(_06179_),
    .Y(_01682_),
    .A1(net719),
    .A2(net238));
 sg13g2_nand2_1 _24384_ (.Y(_06180_),
    .A(_06170_),
    .B(_06083_));
 sg13g2_buf_1 _24385_ (.A(_06180_),
    .X(_06181_));
 sg13g2_buf_1 _24386_ (.A(net297),
    .X(_06182_));
 sg13g2_nand2_1 _24387_ (.Y(_06183_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(net297));
 sg13g2_o21ai_1 _24388_ (.B1(_06183_),
    .Y(_01683_),
    .A1(net571),
    .A2(net237));
 sg13g2_mux2_1 _24389_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(_06182_),
    .X(_01684_));
 sg13g2_nand2_1 _24390_ (.Y(_06184_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(net297));
 sg13g2_o21ai_1 _24391_ (.B1(_06184_),
    .Y(_01685_),
    .A1(net570),
    .A2(_06182_));
 sg13g2_nand2_1 _24392_ (.Y(_06185_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(net297));
 sg13g2_o21ai_1 _24393_ (.B1(_06185_),
    .Y(_01686_),
    .A1(net643),
    .A2(net237));
 sg13g2_nand2_1 _24394_ (.Y(_06186_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .B(net297));
 sg13g2_o21ai_1 _24395_ (.B1(_06186_),
    .Y(_01687_),
    .A1(net722),
    .A2(net237));
 sg13g2_mux2_1 _24396_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .S(net237),
    .X(_01688_));
 sg13g2_mux2_1 _24397_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net237),
    .X(_01689_));
 sg13g2_mux2_1 _24398_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(net237),
    .X(_01690_));
 sg13g2_mux2_1 _24399_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net297),
    .X(_01691_));
 sg13g2_mux2_1 _24400_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(_06181_),
    .X(_01692_));
 sg13g2_nand2_1 _24401_ (.Y(_06187_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .B(net297));
 sg13g2_o21ai_1 _24402_ (.B1(_06187_),
    .Y(_01693_),
    .A1(net642),
    .A2(net237));
 sg13g2_nand2_1 _24403_ (.Y(_06188_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .B(net297));
 sg13g2_o21ai_1 _24404_ (.B1(_06188_),
    .Y(_01694_),
    .A1(net719),
    .A2(net237));
 sg13g2_nand3_1 _24405_ (.B(_06170_),
    .C(net441),
    .A(_06021_),
    .Y(_06189_));
 sg13g2_buf_1 _24406_ (.A(_06189_),
    .X(_06190_));
 sg13g2_buf_1 _24407_ (.A(net373),
    .X(_06191_));
 sg13g2_nand2_1 _24408_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(net373));
 sg13g2_o21ai_1 _24409_ (.B1(_06192_),
    .Y(_01695_),
    .A1(net571),
    .A2(net296));
 sg13g2_mux2_1 _24410_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(_06191_),
    .X(_01696_));
 sg13g2_nand2_1 _24411_ (.Y(_06193_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(net373));
 sg13g2_o21ai_1 _24412_ (.B1(_06193_),
    .Y(_01697_),
    .A1(net570),
    .A2(_06191_));
 sg13g2_nand2_1 _24413_ (.Y(_06194_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(net373));
 sg13g2_o21ai_1 _24414_ (.B1(_06194_),
    .Y(_01698_),
    .A1(net643),
    .A2(net296));
 sg13g2_nand2_1 _24415_ (.Y(_06195_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .B(net373));
 sg13g2_o21ai_1 _24416_ (.B1(_06195_),
    .Y(_01699_),
    .A1(net722),
    .A2(net296));
 sg13g2_mux2_1 _24417_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .S(net296),
    .X(_01700_));
 sg13g2_mux2_1 _24418_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net296),
    .X(_01701_));
 sg13g2_mux2_1 _24419_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(net296),
    .X(_01702_));
 sg13g2_mux2_1 _24420_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net373),
    .X(_01703_));
 sg13g2_mux2_1 _24421_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(_06190_),
    .X(_01704_));
 sg13g2_nand2_1 _24422_ (.Y(_06196_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .B(net373));
 sg13g2_o21ai_1 _24423_ (.B1(_06196_),
    .Y(_01705_),
    .A1(net642),
    .A2(net296));
 sg13g2_nand2_1 _24424_ (.Y(_06197_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .B(net373));
 sg13g2_o21ai_1 _24425_ (.B1(_06197_),
    .Y(_01706_),
    .A1(net719),
    .A2(net296));
 sg13g2_nand3_1 _24426_ (.B(_06170_),
    .C(net441),
    .A(_05831_),
    .Y(_06198_));
 sg13g2_buf_1 _24427_ (.A(_06198_),
    .X(_06199_));
 sg13g2_buf_1 _24428_ (.A(net372),
    .X(_06200_));
 sg13g2_nand2_1 _24429_ (.Y(_06201_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(net372));
 sg13g2_o21ai_1 _24430_ (.B1(_06201_),
    .Y(_01707_),
    .A1(net571),
    .A2(net295));
 sg13g2_mux2_1 _24431_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(_06200_),
    .X(_01708_));
 sg13g2_nand2_1 _24432_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(net372));
 sg13g2_o21ai_1 _24433_ (.B1(_06202_),
    .Y(_01709_),
    .A1(net570),
    .A2(_06200_));
 sg13g2_nand2_1 _24434_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(net372));
 sg13g2_o21ai_1 _24435_ (.B1(_06203_),
    .Y(_01710_),
    .A1(net643),
    .A2(net295));
 sg13g2_nand2_1 _24436_ (.Y(_06204_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .B(_06199_));
 sg13g2_o21ai_1 _24437_ (.B1(_06204_),
    .Y(_01711_),
    .A1(net722),
    .A2(net295));
 sg13g2_mux2_1 _24438_ (.A0(net721),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S(net295),
    .X(_01712_));
 sg13g2_mux2_1 _24439_ (.A0(net720),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net295),
    .X(_01713_));
 sg13g2_mux2_1 _24440_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(net295),
    .X(_01714_));
 sg13g2_mux2_1 _24441_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net372),
    .X(_01715_));
 sg13g2_mux2_1 _24442_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net372),
    .X(_01716_));
 sg13g2_nand2_1 _24443_ (.Y(_06205_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .B(net372));
 sg13g2_o21ai_1 _24444_ (.B1(_06205_),
    .Y(_01717_),
    .A1(net642),
    .A2(net295));
 sg13g2_nand2_1 _24445_ (.Y(_06206_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .B(net372));
 sg13g2_o21ai_1 _24446_ (.B1(_06206_),
    .Y(_01718_),
    .A1(net719),
    .A2(net295));
 sg13g2_nand4_1 _24447_ (.B(net978),
    .C(_06119_),
    .A(net974),
    .Y(_06207_),
    .D(_06102_));
 sg13g2_buf_1 _24448_ (.A(_06207_),
    .X(_06208_));
 sg13g2_buf_1 _24449_ (.A(net371),
    .X(_06209_));
 sg13g2_nand2_1 _24450_ (.Y(_06210_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(net371));
 sg13g2_o21ai_1 _24451_ (.B1(_06210_),
    .Y(_01719_),
    .A1(net571),
    .A2(net294));
 sg13g2_mux2_1 _24452_ (.A0(_06134_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net294),
    .X(_01720_));
 sg13g2_nand2_1 _24453_ (.Y(_06211_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(net371));
 sg13g2_o21ai_1 _24454_ (.B1(_06211_),
    .Y(_01721_),
    .A1(net570),
    .A2(_06209_));
 sg13g2_buf_1 _24455_ (.A(net744),
    .X(_06212_));
 sg13g2_nand2_1 _24456_ (.Y(_06213_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(net371));
 sg13g2_o21ai_1 _24457_ (.B1(_06213_),
    .Y(_01722_),
    .A1(net641),
    .A2(net294));
 sg13g2_buf_1 _24458_ (.A(net863),
    .X(_06214_));
 sg13g2_nand2_1 _24459_ (.Y(_06215_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .B(_06208_));
 sg13g2_o21ai_1 _24460_ (.B1(_06215_),
    .Y(_01723_),
    .A1(net718),
    .A2(_06209_));
 sg13g2_buf_1 _24461_ (.A(net862),
    .X(_06216_));
 sg13g2_mux2_1 _24462_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .S(net294),
    .X(_01724_));
 sg13g2_buf_1 _24463_ (.A(net861),
    .X(_06217_));
 sg13g2_mux2_1 _24464_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net294),
    .X(_01725_));
 sg13g2_buf_1 _24465_ (.A(net993),
    .X(_06218_));
 sg13g2_mux2_1 _24466_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(net294),
    .X(_01726_));
 sg13g2_buf_1 _24467_ (.A(net992),
    .X(_06219_));
 sg13g2_mux2_1 _24468_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net371),
    .X(_01727_));
 sg13g2_buf_1 _24469_ (.A(net991),
    .X(_06220_));
 sg13g2_mux2_1 _24470_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net371),
    .X(_01728_));
 sg13g2_nand2_1 _24471_ (.Y(_06221_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .B(net371));
 sg13g2_o21ai_1 _24472_ (.B1(_06221_),
    .Y(_01729_),
    .A1(net642),
    .A2(net294));
 sg13g2_nand2_1 _24473_ (.Y(_06222_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .B(net371));
 sg13g2_o21ai_1 _24474_ (.B1(_06222_),
    .Y(_01730_),
    .A1(net719),
    .A2(net294));
 sg13g2_nand4_1 _24475_ (.B(_05839_),
    .C(net978),
    .A(net974),
    .Y(_06223_),
    .D(_06083_));
 sg13g2_buf_1 _24476_ (.A(_06223_),
    .X(_06224_));
 sg13g2_buf_1 _24477_ (.A(net293),
    .X(_06225_));
 sg13g2_nand2_1 _24478_ (.Y(_06226_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(net293));
 sg13g2_o21ai_1 _24479_ (.B1(_06226_),
    .Y(_01731_),
    .A1(net571),
    .A2(net236));
 sg13g2_mux2_1 _24480_ (.A0(_06134_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net236),
    .X(_01732_));
 sg13g2_nand2_1 _24481_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(net293));
 sg13g2_o21ai_1 _24482_ (.B1(_06227_),
    .Y(_01733_),
    .A1(net570),
    .A2(_06225_));
 sg13g2_nand2_1 _24483_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(net293));
 sg13g2_o21ai_1 _24484_ (.B1(_06228_),
    .Y(_01734_),
    .A1(net641),
    .A2(net236));
 sg13g2_nand2_1 _24485_ (.Y(_06229_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .B(_06224_));
 sg13g2_o21ai_1 _24486_ (.B1(_06229_),
    .Y(_01735_),
    .A1(net718),
    .A2(_06225_));
 sg13g2_mux2_1 _24487_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .S(net236),
    .X(_01736_));
 sg13g2_mux2_1 _24488_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net236),
    .X(_01737_));
 sg13g2_mux2_1 _24489_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(net236),
    .X(_01738_));
 sg13g2_mux2_1 _24490_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net293),
    .X(_01739_));
 sg13g2_mux2_1 _24491_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net293),
    .X(_01740_));
 sg13g2_nand2_1 _24492_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .B(net293));
 sg13g2_o21ai_1 _24493_ (.B1(_06230_),
    .Y(_01741_),
    .A1(net642),
    .A2(net236));
 sg13g2_nand2_1 _24494_ (.Y(_06231_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .B(net293));
 sg13g2_o21ai_1 _24495_ (.B1(_06231_),
    .Y(_01742_),
    .A1(net719),
    .A2(net236));
 sg13g2_buf_1 _24496_ (.A(net653),
    .X(_06232_));
 sg13g2_nand2_1 _24497_ (.Y(_06233_),
    .A(_05974_),
    .B(net442));
 sg13g2_buf_1 _24498_ (.A(_06233_),
    .X(_06234_));
 sg13g2_buf_1 _24499_ (.A(net370),
    .X(_06235_));
 sg13g2_nand2_1 _24500_ (.Y(_06236_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(net370));
 sg13g2_o21ai_1 _24501_ (.B1(_06236_),
    .Y(_01743_),
    .A1(net569),
    .A2(net292));
 sg13g2_buf_1 _24502_ (.A(net520),
    .X(_06237_));
 sg13g2_mux2_1 _24503_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net292),
    .X(_01744_));
 sg13g2_buf_1 _24504_ (.A(net666),
    .X(_06238_));
 sg13g2_nand2_1 _24505_ (.Y(_06239_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(net370));
 sg13g2_o21ai_1 _24506_ (.B1(_06239_),
    .Y(_01745_),
    .A1(net568),
    .A2(net292));
 sg13g2_nand2_1 _24507_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(net370));
 sg13g2_o21ai_1 _24508_ (.B1(_06240_),
    .Y(_01746_),
    .A1(net641),
    .A2(net292));
 sg13g2_nand2_1 _24509_ (.Y(_06241_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .B(_06234_));
 sg13g2_o21ai_1 _24510_ (.B1(_06241_),
    .Y(_01747_),
    .A1(_06214_),
    .A2(_06235_));
 sg13g2_mux2_1 _24511_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .S(net292),
    .X(_01748_));
 sg13g2_mux2_1 _24512_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net292),
    .X(_01749_));
 sg13g2_mux2_1 _24513_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(net292),
    .X(_01750_));
 sg13g2_mux2_1 _24514_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(net370),
    .X(_01751_));
 sg13g2_mux2_1 _24515_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net370),
    .X(_01752_));
 sg13g2_buf_1 _24516_ (.A(net749),
    .X(_06242_));
 sg13g2_nand2_1 _24517_ (.Y(_06243_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .B(net370));
 sg13g2_o21ai_1 _24518_ (.B1(_06243_),
    .Y(_01753_),
    .A1(net640),
    .A2(net292));
 sg13g2_buf_1 _24519_ (.A(net875),
    .X(_06244_));
 sg13g2_nand2_1 _24520_ (.Y(_06245_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .B(net370));
 sg13g2_o21ai_1 _24521_ (.B1(_06245_),
    .Y(_01754_),
    .A1(net715),
    .A2(_06235_));
 sg13g2_nand2_1 _24522_ (.Y(_06246_),
    .A(_05979_),
    .B(net442));
 sg13g2_buf_1 _24523_ (.A(_06246_),
    .X(_06247_));
 sg13g2_buf_1 _24524_ (.A(net369),
    .X(_06248_));
 sg13g2_nand2_1 _24525_ (.Y(_06249_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(net369));
 sg13g2_o21ai_1 _24526_ (.B1(_06249_),
    .Y(_01755_),
    .A1(_06232_),
    .A2(net291));
 sg13g2_mux2_1 _24527_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net291),
    .X(_01756_));
 sg13g2_nand2_1 _24528_ (.Y(_06250_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(net369));
 sg13g2_o21ai_1 _24529_ (.B1(_06250_),
    .Y(_01757_),
    .A1(net568),
    .A2(net291));
 sg13g2_nand2_1 _24530_ (.Y(_06251_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(net369));
 sg13g2_o21ai_1 _24531_ (.B1(_06251_),
    .Y(_01758_),
    .A1(net641),
    .A2(net291));
 sg13g2_nand2_1 _24532_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .B(_06247_));
 sg13g2_o21ai_1 _24533_ (.B1(_06252_),
    .Y(_01759_),
    .A1(_06214_),
    .A2(_06248_));
 sg13g2_mux2_1 _24534_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S(net291),
    .X(_01760_));
 sg13g2_mux2_1 _24535_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net291),
    .X(_01761_));
 sg13g2_mux2_1 _24536_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(net291),
    .X(_01762_));
 sg13g2_mux2_1 _24537_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(net369),
    .X(_01763_));
 sg13g2_mux2_1 _24538_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net369),
    .X(_01764_));
 sg13g2_nand2_1 _24539_ (.Y(_06253_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .B(net369));
 sg13g2_o21ai_1 _24540_ (.B1(_06253_),
    .Y(_01765_),
    .A1(net640),
    .A2(net291));
 sg13g2_nand2_1 _24541_ (.Y(_06254_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .B(net369));
 sg13g2_o21ai_1 _24542_ (.B1(_06254_),
    .Y(_01766_),
    .A1(net715),
    .A2(_06248_));
 sg13g2_nor2_2 _24543_ (.A(_05861_),
    .B(_05965_),
    .Y(_06255_));
 sg13g2_nand2_1 _24544_ (.Y(_06256_),
    .A(_06255_),
    .B(_06043_));
 sg13g2_buf_1 _24545_ (.A(_06256_),
    .X(_06257_));
 sg13g2_buf_1 _24546_ (.A(net290),
    .X(_06258_));
 sg13g2_nand2_1 _24547_ (.Y(_06259_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(net290));
 sg13g2_o21ai_1 _24548_ (.B1(_06259_),
    .Y(_01767_),
    .A1(net569),
    .A2(net235));
 sg13g2_mux2_1 _24549_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(_06258_),
    .X(_01768_));
 sg13g2_nand2_1 _24550_ (.Y(_06260_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(net290));
 sg13g2_o21ai_1 _24551_ (.B1(_06260_),
    .Y(_01769_),
    .A1(net568),
    .A2(net235));
 sg13g2_nand2_1 _24552_ (.Y(_06261_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(net290));
 sg13g2_o21ai_1 _24553_ (.B1(_06261_),
    .Y(_01770_),
    .A1(net641),
    .A2(net235));
 sg13g2_nand2_1 _24554_ (.Y(_06262_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .B(net290));
 sg13g2_o21ai_1 _24555_ (.B1(_06262_),
    .Y(_01771_),
    .A1(net718),
    .A2(net235));
 sg13g2_mux2_1 _24556_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .S(net235),
    .X(_01772_));
 sg13g2_mux2_1 _24557_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net235),
    .X(_01773_));
 sg13g2_mux2_1 _24558_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(net235),
    .X(_01774_));
 sg13g2_mux2_1 _24559_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(net290),
    .X(_01775_));
 sg13g2_mux2_1 _24560_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(_06257_),
    .X(_01776_));
 sg13g2_nand2_1 _24561_ (.Y(_06263_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .B(net290));
 sg13g2_o21ai_1 _24562_ (.B1(_06263_),
    .Y(_01777_),
    .A1(net640),
    .A2(net235));
 sg13g2_nand2_1 _24563_ (.Y(_06264_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .B(net290));
 sg13g2_o21ai_1 _24564_ (.B1(_06264_),
    .Y(_01778_),
    .A1(net715),
    .A2(_06258_));
 sg13g2_nand2_1 _24565_ (.Y(_06265_),
    .A(_06255_),
    .B(_06083_));
 sg13g2_buf_1 _24566_ (.A(_06265_),
    .X(_06266_));
 sg13g2_buf_1 _24567_ (.A(net289),
    .X(_06267_));
 sg13g2_nand2_1 _24568_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(net289));
 sg13g2_o21ai_1 _24569_ (.B1(_06268_),
    .Y(_01779_),
    .A1(net569),
    .A2(net234));
 sg13g2_mux2_1 _24570_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(_06267_),
    .X(_01780_));
 sg13g2_nand2_1 _24571_ (.Y(_06269_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(net289));
 sg13g2_o21ai_1 _24572_ (.B1(_06269_),
    .Y(_01781_),
    .A1(net568),
    .A2(net234));
 sg13g2_nand2_1 _24573_ (.Y(_06270_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(net289));
 sg13g2_o21ai_1 _24574_ (.B1(_06270_),
    .Y(_01782_),
    .A1(net641),
    .A2(net234));
 sg13g2_nand2_1 _24575_ (.Y(_06271_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .B(net289));
 sg13g2_o21ai_1 _24576_ (.B1(_06271_),
    .Y(_01783_),
    .A1(net718),
    .A2(net234));
 sg13g2_mux2_1 _24577_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .S(net234),
    .X(_01784_));
 sg13g2_mux2_1 _24578_ (.A0(_06217_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net234),
    .X(_01785_));
 sg13g2_mux2_1 _24579_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(net234),
    .X(_01786_));
 sg13g2_mux2_1 _24580_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(net289),
    .X(_01787_));
 sg13g2_mux2_1 _24581_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(_06266_),
    .X(_01788_));
 sg13g2_nand2_1 _24582_ (.Y(_06272_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .B(net289));
 sg13g2_o21ai_1 _24583_ (.B1(_06272_),
    .Y(_01789_),
    .A1(net640),
    .A2(net234));
 sg13g2_nand2_1 _24584_ (.Y(_06273_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .B(net289));
 sg13g2_o21ai_1 _24585_ (.B1(_06273_),
    .Y(_01790_),
    .A1(net715),
    .A2(_06267_));
 sg13g2_nand3_1 _24586_ (.B(_06039_),
    .C(net441),
    .A(_06021_),
    .Y(_06274_));
 sg13g2_buf_1 _24587_ (.A(_06274_),
    .X(_06275_));
 sg13g2_buf_1 _24588_ (.A(net368),
    .X(_06276_));
 sg13g2_nand2_1 _24589_ (.Y(_06277_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(net368));
 sg13g2_o21ai_1 _24590_ (.B1(_06277_),
    .Y(_01791_),
    .A1(net569),
    .A2(net288));
 sg13g2_mux2_1 _24591_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(_06276_),
    .X(_01792_));
 sg13g2_nand2_1 _24592_ (.Y(_06278_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(net368));
 sg13g2_o21ai_1 _24593_ (.B1(_06278_),
    .Y(_01793_),
    .A1(_06238_),
    .A2(net288));
 sg13g2_nand2_1 _24594_ (.Y(_06279_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(net368));
 sg13g2_o21ai_1 _24595_ (.B1(_06279_),
    .Y(_01794_),
    .A1(_06212_),
    .A2(net288));
 sg13g2_nand2_1 _24596_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .B(net368));
 sg13g2_o21ai_1 _24597_ (.B1(_06280_),
    .Y(_01795_),
    .A1(net718),
    .A2(net288));
 sg13g2_mux2_1 _24598_ (.A0(_06216_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .S(net288),
    .X(_01796_));
 sg13g2_mux2_1 _24599_ (.A0(_06217_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net288),
    .X(_01797_));
 sg13g2_mux2_1 _24600_ (.A0(_06218_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(net288),
    .X(_01798_));
 sg13g2_mux2_1 _24601_ (.A0(_06219_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net368),
    .X(_01799_));
 sg13g2_mux2_1 _24602_ (.A0(_06220_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(_06275_),
    .X(_01800_));
 sg13g2_nand2_1 _24603_ (.Y(_06281_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .B(net368));
 sg13g2_o21ai_1 _24604_ (.B1(_06281_),
    .Y(_01801_),
    .A1(_06242_),
    .A2(_06276_));
 sg13g2_nand2_1 _24605_ (.Y(_06282_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .B(net368));
 sg13g2_o21ai_1 _24606_ (.B1(_06282_),
    .Y(_01802_),
    .A1(_06244_),
    .A2(net288));
 sg13g2_nand3_1 _24607_ (.B(_06255_),
    .C(net441),
    .A(_06021_),
    .Y(_06283_));
 sg13g2_buf_1 _24608_ (.A(_06283_),
    .X(_06284_));
 sg13g2_buf_1 _24609_ (.A(net367),
    .X(_06285_));
 sg13g2_nand2_1 _24610_ (.Y(_06286_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(net367));
 sg13g2_o21ai_1 _24611_ (.B1(_06286_),
    .Y(_01803_),
    .A1(net569),
    .A2(net287));
 sg13g2_mux2_1 _24612_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(_06285_),
    .X(_01804_));
 sg13g2_nand2_1 _24613_ (.Y(_06287_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(net367));
 sg13g2_o21ai_1 _24614_ (.B1(_06287_),
    .Y(_01805_),
    .A1(net568),
    .A2(net287));
 sg13g2_nand2_1 _24615_ (.Y(_06288_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(net367));
 sg13g2_o21ai_1 _24616_ (.B1(_06288_),
    .Y(_01806_),
    .A1(net641),
    .A2(net287));
 sg13g2_nand2_1 _24617_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .B(net367));
 sg13g2_o21ai_1 _24618_ (.B1(_06289_),
    .Y(_01807_),
    .A1(net718),
    .A2(net287));
 sg13g2_mux2_1 _24619_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .S(net287),
    .X(_01808_));
 sg13g2_mux2_1 _24620_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net287),
    .X(_01809_));
 sg13g2_mux2_1 _24621_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(net287),
    .X(_01810_));
 sg13g2_mux2_1 _24622_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(net367),
    .X(_01811_));
 sg13g2_mux2_1 _24623_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(_06284_),
    .X(_01812_));
 sg13g2_nand2_1 _24624_ (.Y(_06290_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .B(net367));
 sg13g2_o21ai_1 _24625_ (.B1(_06290_),
    .Y(_01813_),
    .A1(net640),
    .A2(net287));
 sg13g2_nand2_1 _24626_ (.Y(_06291_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .B(net367));
 sg13g2_o21ai_1 _24627_ (.B1(_06291_),
    .Y(_01814_),
    .A1(net715),
    .A2(_06285_));
 sg13g2_nand3_1 _24628_ (.B(_06255_),
    .C(net441),
    .A(_05831_),
    .Y(_06292_));
 sg13g2_buf_1 _24629_ (.A(_06292_),
    .X(_06293_));
 sg13g2_buf_1 _24630_ (.A(net366),
    .X(_06294_));
 sg13g2_nand2_1 _24631_ (.Y(_06295_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(net366));
 sg13g2_o21ai_1 _24632_ (.B1(_06295_),
    .Y(_01815_),
    .A1(net569),
    .A2(net286));
 sg13g2_mux2_1 _24633_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(_06294_),
    .X(_01816_));
 sg13g2_nand2_1 _24634_ (.Y(_06296_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(net366));
 sg13g2_o21ai_1 _24635_ (.B1(_06296_),
    .Y(_01817_),
    .A1(net568),
    .A2(net286));
 sg13g2_nand2_1 _24636_ (.Y(_06297_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(net366));
 sg13g2_o21ai_1 _24637_ (.B1(_06297_),
    .Y(_01818_),
    .A1(net641),
    .A2(net286));
 sg13g2_nand2_1 _24638_ (.Y(_06298_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .B(net366));
 sg13g2_o21ai_1 _24639_ (.B1(_06298_),
    .Y(_01819_),
    .A1(net718),
    .A2(net286));
 sg13g2_mux2_1 _24640_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S(net286),
    .X(_01820_));
 sg13g2_mux2_1 _24641_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net286),
    .X(_01821_));
 sg13g2_mux2_1 _24642_ (.A0(net833),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(net286),
    .X(_01822_));
 sg13g2_mux2_1 _24643_ (.A0(net832),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(net366),
    .X(_01823_));
 sg13g2_mux2_1 _24644_ (.A0(net831),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(_06293_),
    .X(_01824_));
 sg13g2_nand2_1 _24645_ (.Y(_06299_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .B(net366));
 sg13g2_o21ai_1 _24646_ (.B1(_06299_),
    .Y(_01825_),
    .A1(net640),
    .A2(net286));
 sg13g2_nand2_1 _24647_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .B(net366));
 sg13g2_o21ai_1 _24648_ (.B1(_06300_),
    .Y(_01826_),
    .A1(net715),
    .A2(_06294_));
 sg13g2_nand3_1 _24649_ (.B(_06039_),
    .C(net441),
    .A(_05831_),
    .Y(_06301_));
 sg13g2_buf_1 _24650_ (.A(_06301_),
    .X(_06302_));
 sg13g2_buf_1 _24651_ (.A(net365),
    .X(_06303_));
 sg13g2_nand2_1 _24652_ (.Y(_06304_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(net365));
 sg13g2_o21ai_1 _24653_ (.B1(_06304_),
    .Y(_01827_),
    .A1(_06232_),
    .A2(net285));
 sg13g2_mux2_1 _24654_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(_06303_),
    .X(_01828_));
 sg13g2_nand2_1 _24655_ (.Y(_06305_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(net365));
 sg13g2_o21ai_1 _24656_ (.B1(_06305_),
    .Y(_01829_),
    .A1(_06238_),
    .A2(net285));
 sg13g2_nand2_1 _24657_ (.Y(_06306_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(net365));
 sg13g2_o21ai_1 _24658_ (.B1(_06306_),
    .Y(_01830_),
    .A1(_06212_),
    .A2(net285));
 sg13g2_nand2_1 _24659_ (.Y(_06307_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .B(net365));
 sg13g2_o21ai_1 _24660_ (.B1(_06307_),
    .Y(_01831_),
    .A1(net718),
    .A2(net285));
 sg13g2_mux2_1 _24661_ (.A0(_06216_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S(net285),
    .X(_01832_));
 sg13g2_mux2_1 _24662_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net285),
    .X(_01833_));
 sg13g2_mux2_1 _24663_ (.A0(_06218_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(net285),
    .X(_01834_));
 sg13g2_mux2_1 _24664_ (.A0(_06219_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net365),
    .X(_01835_));
 sg13g2_mux2_1 _24665_ (.A0(_06220_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(_06302_),
    .X(_01836_));
 sg13g2_nand2_1 _24666_ (.Y(_06308_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .B(net365));
 sg13g2_o21ai_1 _24667_ (.B1(_06308_),
    .Y(_01837_),
    .A1(_06242_),
    .A2(_06303_));
 sg13g2_nand2_1 _24668_ (.Y(_06309_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .B(net365));
 sg13g2_o21ai_1 _24669_ (.B1(_06309_),
    .Y(_01838_),
    .A1(_06244_),
    .A2(net285));
 sg13g2_nand2b_1 _24670_ (.Y(_06310_),
    .B(_06043_),
    .A_N(_06012_));
 sg13g2_buf_1 _24671_ (.A(_06310_),
    .X(_06311_));
 sg13g2_buf_1 _24672_ (.A(net284),
    .X(_06312_));
 sg13g2_nand2_1 _24673_ (.Y(_06313_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(net284));
 sg13g2_o21ai_1 _24674_ (.B1(_06313_),
    .Y(_01839_),
    .A1(net569),
    .A2(net233));
 sg13g2_mux2_1 _24675_ (.A0(_06237_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net233),
    .X(_01840_));
 sg13g2_nand2_1 _24676_ (.Y(_06314_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(net284));
 sg13g2_o21ai_1 _24677_ (.B1(_06314_),
    .Y(_01841_),
    .A1(net568),
    .A2(net233));
 sg13g2_nand2_1 _24678_ (.Y(_06315_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(net284));
 sg13g2_o21ai_1 _24679_ (.B1(_06315_),
    .Y(_01842_),
    .A1(net744),
    .A2(net233));
 sg13g2_nand2_1 _24680_ (.Y(_06316_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .B(net284));
 sg13g2_o21ai_1 _24681_ (.B1(_06316_),
    .Y(_01843_),
    .A1(net863),
    .A2(net233));
 sg13g2_mux2_1 _24682_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .S(net233),
    .X(_01844_));
 sg13g2_mux2_1 _24683_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net233),
    .X(_01845_));
 sg13g2_mux2_1 _24684_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net233),
    .X(_01846_));
 sg13g2_mux2_1 _24685_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net284),
    .X(_01847_));
 sg13g2_mux2_1 _24686_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(_06311_),
    .X(_01848_));
 sg13g2_nand2_1 _24687_ (.Y(_06317_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .B(net284));
 sg13g2_o21ai_1 _24688_ (.B1(_06317_),
    .Y(_01849_),
    .A1(net640),
    .A2(_06312_));
 sg13g2_nand2_1 _24689_ (.Y(_06318_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .B(net284));
 sg13g2_o21ai_1 _24690_ (.B1(_06318_),
    .Y(_01850_),
    .A1(net715),
    .A2(_06312_));
 sg13g2_nand2_1 _24691_ (.Y(_06319_),
    .A(_06017_),
    .B(net442));
 sg13g2_buf_1 _24692_ (.A(_06319_),
    .X(_06320_));
 sg13g2_buf_1 _24693_ (.A(net364),
    .X(_06321_));
 sg13g2_nand2_1 _24694_ (.Y(_06322_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(net364));
 sg13g2_o21ai_1 _24695_ (.B1(_06322_),
    .Y(_01851_),
    .A1(net569),
    .A2(net283));
 sg13g2_mux2_1 _24696_ (.A0(_06237_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net283),
    .X(_01852_));
 sg13g2_nand2_1 _24697_ (.Y(_06323_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(net364));
 sg13g2_o21ai_1 _24698_ (.B1(_06323_),
    .Y(_01853_),
    .A1(net568),
    .A2(net283));
 sg13g2_nand2_1 _24699_ (.Y(_06324_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(net364));
 sg13g2_o21ai_1 _24700_ (.B1(_06324_),
    .Y(_01854_),
    .A1(net744),
    .A2(net283));
 sg13g2_nand2_1 _24701_ (.Y(_06325_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .B(net364));
 sg13g2_o21ai_1 _24702_ (.B1(_06325_),
    .Y(_01855_),
    .A1(net863),
    .A2(net283));
 sg13g2_mux2_1 _24703_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .S(net283),
    .X(_01856_));
 sg13g2_mux2_1 _24704_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net283),
    .X(_01857_));
 sg13g2_mux2_1 _24705_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net283),
    .X(_01858_));
 sg13g2_mux2_1 _24706_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net364),
    .X(_01859_));
 sg13g2_mux2_1 _24707_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net364),
    .X(_01860_));
 sg13g2_nand2_1 _24708_ (.Y(_06326_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .B(net364));
 sg13g2_o21ai_1 _24709_ (.B1(_06326_),
    .Y(_01861_),
    .A1(net640),
    .A2(_06321_));
 sg13g2_nand2_1 _24710_ (.Y(_06327_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .B(_06320_));
 sg13g2_o21ai_1 _24711_ (.B1(_06327_),
    .Y(_01862_),
    .A1(net715),
    .A2(_06321_));
 sg13g2_nand2_1 _24712_ (.Y(_06328_),
    .A(_06023_),
    .B(_06053_));
 sg13g2_buf_1 _24713_ (.A(_06328_),
    .X(_06329_));
 sg13g2_buf_1 _24714_ (.A(net363),
    .X(_06330_));
 sg13g2_nand2_1 _24715_ (.Y(_06331_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(net363));
 sg13g2_o21ai_1 _24716_ (.B1(_06331_),
    .Y(_01863_),
    .A1(net653),
    .A2(net282));
 sg13g2_mux2_1 _24717_ (.A0(net462),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net282),
    .X(_01864_));
 sg13g2_nand2_1 _24718_ (.Y(_06332_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(net363));
 sg13g2_o21ai_1 _24719_ (.B1(_06332_),
    .Y(_01865_),
    .A1(net666),
    .A2(net282));
 sg13g2_nand2_1 _24720_ (.Y(_06333_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(net363));
 sg13g2_o21ai_1 _24721_ (.B1(_06333_),
    .Y(_01866_),
    .A1(net744),
    .A2(net282));
 sg13g2_nand2_1 _24722_ (.Y(_06334_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .B(net363));
 sg13g2_o21ai_1 _24723_ (.B1(_06334_),
    .Y(_01867_),
    .A1(net863),
    .A2(net282));
 sg13g2_mux2_1 _24724_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .S(net282),
    .X(_01868_));
 sg13g2_mux2_1 _24725_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net282),
    .X(_01869_));
 sg13g2_mux2_1 _24726_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net282),
    .X(_01870_));
 sg13g2_mux2_1 _24727_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net363),
    .X(_01871_));
 sg13g2_mux2_1 _24728_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(_06329_),
    .X(_01872_));
 sg13g2_nand2_1 _24729_ (.Y(_06335_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .B(net363));
 sg13g2_o21ai_1 _24730_ (.B1(_06335_),
    .Y(_01873_),
    .A1(net749),
    .A2(_06330_));
 sg13g2_nand2_1 _24731_ (.Y(_06336_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .B(net363));
 sg13g2_o21ai_1 _24732_ (.B1(_06336_),
    .Y(_01874_),
    .A1(net875),
    .A2(_06330_));
 sg13g2_nand2_1 _24733_ (.Y(_06337_),
    .A(_06028_),
    .B(net442));
 sg13g2_buf_1 _24734_ (.A(_06337_),
    .X(_06338_));
 sg13g2_buf_1 _24735_ (.A(net362),
    .X(_06339_));
 sg13g2_nand2_1 _24736_ (.Y(_06340_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(net362));
 sg13g2_o21ai_1 _24737_ (.B1(_06340_),
    .Y(_01875_),
    .A1(net653),
    .A2(net281));
 sg13g2_mux2_1 _24738_ (.A0(net462),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net281),
    .X(_01876_));
 sg13g2_nand2_1 _24739_ (.Y(_06341_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(net362));
 sg13g2_o21ai_1 _24740_ (.B1(_06341_),
    .Y(_01877_),
    .A1(net666),
    .A2(_06339_));
 sg13g2_nand2_1 _24741_ (.Y(_06342_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(net362));
 sg13g2_o21ai_1 _24742_ (.B1(_06342_),
    .Y(_01878_),
    .A1(net744),
    .A2(net281));
 sg13g2_nand2_1 _24743_ (.Y(_06343_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .B(net362));
 sg13g2_o21ai_1 _24744_ (.B1(_06343_),
    .Y(_01879_),
    .A1(net863),
    .A2(net281));
 sg13g2_mux2_1 _24745_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S(net281),
    .X(_01880_));
 sg13g2_mux2_1 _24746_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net281),
    .X(_01881_));
 sg13g2_mux2_1 _24747_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net281),
    .X(_01882_));
 sg13g2_mux2_1 _24748_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net362),
    .X(_01883_));
 sg13g2_mux2_1 _24749_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(_06338_),
    .X(_01884_));
 sg13g2_nand2_1 _24750_ (.Y(_06344_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .B(net362));
 sg13g2_o21ai_1 _24751_ (.B1(_06344_),
    .Y(_01885_),
    .A1(net749),
    .A2(net281));
 sg13g2_nand2_1 _24752_ (.Y(_06345_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .B(net362));
 sg13g2_o21ai_1 _24753_ (.B1(_06345_),
    .Y(_01886_),
    .A1(net875),
    .A2(_06339_));
 sg13g2_nand3_1 _24754_ (.B(_06119_),
    .C(_06102_),
    .A(_05893_),
    .Y(_06346_));
 sg13g2_buf_1 _24755_ (.A(_06346_),
    .X(_06347_));
 sg13g2_buf_1 _24756_ (.A(net361),
    .X(_06348_));
 sg13g2_nand2_1 _24757_ (.Y(_06349_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(net361));
 sg13g2_o21ai_1 _24758_ (.B1(_06349_),
    .Y(_01887_),
    .A1(net653),
    .A2(net280));
 sg13g2_mux2_1 _24759_ (.A0(net462),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(net280),
    .X(_01888_));
 sg13g2_nand2_1 _24760_ (.Y(_06350_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(net361));
 sg13g2_o21ai_1 _24761_ (.B1(_06350_),
    .Y(_01889_),
    .A1(net666),
    .A2(net280));
 sg13g2_nand2_1 _24762_ (.Y(_06351_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(net361));
 sg13g2_o21ai_1 _24763_ (.B1(_06351_),
    .Y(_01890_),
    .A1(net744),
    .A2(net280));
 sg13g2_nand2_1 _24764_ (.Y(_06352_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .B(net361));
 sg13g2_o21ai_1 _24765_ (.B1(_06352_),
    .Y(_01891_),
    .A1(net863),
    .A2(net280));
 sg13g2_mux2_1 _24766_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .S(net280),
    .X(_01892_));
 sg13g2_mux2_1 _24767_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net280),
    .X(_01893_));
 sg13g2_mux2_1 _24768_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net280),
    .X(_01894_));
 sg13g2_mux2_1 _24769_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net361),
    .X(_01895_));
 sg13g2_mux2_1 _24770_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net361),
    .X(_01896_));
 sg13g2_nand2_1 _24771_ (.Y(_06353_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .B(_06347_));
 sg13g2_o21ai_1 _24772_ (.B1(_06353_),
    .Y(_01897_),
    .A1(net749),
    .A2(_06348_));
 sg13g2_nand2_1 _24773_ (.Y(_06354_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .B(net361));
 sg13g2_o21ai_1 _24774_ (.B1(_06354_),
    .Y(_01898_),
    .A1(net875),
    .A2(_06348_));
 sg13g2_nand3_1 _24775_ (.B(_05893_),
    .C(_06083_),
    .A(_05839_),
    .Y(_06355_));
 sg13g2_buf_1 _24776_ (.A(_06355_),
    .X(_06356_));
 sg13g2_buf_1 _24777_ (.A(net279),
    .X(_06357_));
 sg13g2_nand2_1 _24778_ (.Y(_06358_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(net279));
 sg13g2_o21ai_1 _24779_ (.B1(_06358_),
    .Y(_01899_),
    .A1(net653),
    .A2(net232));
 sg13g2_mux2_1 _24780_ (.A0(net462),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(net232),
    .X(_01900_));
 sg13g2_nand2_1 _24781_ (.Y(_06359_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(net279));
 sg13g2_o21ai_1 _24782_ (.B1(_06359_),
    .Y(_01901_),
    .A1(net666),
    .A2(net232));
 sg13g2_nand2_1 _24783_ (.Y(_06360_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(net279));
 sg13g2_o21ai_1 _24784_ (.B1(_06360_),
    .Y(_01902_),
    .A1(net744),
    .A2(net232));
 sg13g2_nand2_1 _24785_ (.Y(_06361_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .B(net279));
 sg13g2_o21ai_1 _24786_ (.B1(_06361_),
    .Y(_01903_),
    .A1(net863),
    .A2(net232));
 sg13g2_mux2_1 _24787_ (.A0(net739),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .S(net232),
    .X(_01904_));
 sg13g2_mux2_1 _24788_ (.A0(net738),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net232),
    .X(_01905_));
 sg13g2_mux2_1 _24789_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net232),
    .X(_01906_));
 sg13g2_mux2_1 _24790_ (.A0(net854),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net279),
    .X(_01907_));
 sg13g2_mux2_1 _24791_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net279),
    .X(_01908_));
 sg13g2_nand2_1 _24792_ (.Y(_06362_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .B(_06356_));
 sg13g2_o21ai_1 _24793_ (.B1(_06362_),
    .Y(_01909_),
    .A1(net749),
    .A2(_06357_));
 sg13g2_nand2_1 _24794_ (.Y(_06363_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .B(net279));
 sg13g2_o21ai_1 _24795_ (.B1(_06363_),
    .Y(_01910_),
    .A1(net875),
    .A2(_06357_));
 sg13g2_mux2_1 _24796_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(_03533_),
    .S(_05870_),
    .X(_01911_));
 sg13g2_mux2_1 _24797_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(_03533_),
    .S(_05883_),
    .X(_01912_));
 sg13g2_buf_1 _24798_ (.A(net590),
    .X(_06364_));
 sg13g2_mux2_1 _24799_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net495),
    .S(_05891_),
    .X(_01913_));
 sg13g2_mux2_1 _24800_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net495),
    .S(_05897_),
    .X(_01914_));
 sg13g2_mux2_1 _24801_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(_06364_),
    .S(_05904_),
    .X(_01915_));
 sg13g2_mux2_1 _24802_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(net495),
    .S(_05908_),
    .X(_01916_));
 sg13g2_mux2_1 _24803_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(net495),
    .S(_05912_),
    .X(_01917_));
 sg13g2_mux2_1 _24804_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net495),
    .S(_05919_),
    .X(_01918_));
 sg13g2_mux2_1 _24805_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net495),
    .S(_05923_),
    .X(_01919_));
 sg13g2_mux2_1 _24806_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net495),
    .S(_05930_),
    .X(_01920_));
 sg13g2_mux2_1 _24807_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net495),
    .S(_05937_),
    .X(_01921_));
 sg13g2_mux2_1 _24808_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(_06364_),
    .S(_05944_),
    .X(_01922_));
 sg13g2_buf_1 _24809_ (.A(net590),
    .X(_06365_));
 sg13g2_mux2_1 _24810_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net494),
    .S(_05952_),
    .X(_01923_));
 sg13g2_mux2_1 _24811_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net494),
    .S(_05955_),
    .X(_01924_));
 sg13g2_mux2_1 _24812_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(_06365_),
    .S(_05958_),
    .X(_01925_));
 sg13g2_mux2_1 _24813_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net494),
    .S(_05961_),
    .X(_01926_));
 sg13g2_mux2_1 _24814_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net494),
    .S(_05967_),
    .X(_01927_));
 sg13g2_mux2_1 _24815_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net494),
    .S(_05971_),
    .X(_01928_));
 sg13g2_mux2_1 _24816_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net494),
    .S(_05976_),
    .X(_01929_));
 sg13g2_mux2_1 _24817_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(_06365_),
    .S(_05981_),
    .X(_01930_));
 sg13g2_mux2_1 _24818_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net494),
    .S(_05988_),
    .X(_01931_));
 sg13g2_mux2_1 _24819_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net494),
    .S(_05995_),
    .X(_01932_));
 sg13g2_buf_1 _24820_ (.A(net590),
    .X(_06366_));
 sg13g2_mux2_1 _24821_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(net493),
    .S(_06001_),
    .X(_01933_));
 sg13g2_mux2_1 _24822_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net493),
    .S(_06004_),
    .X(_01934_));
 sg13g2_mux2_1 _24823_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net493),
    .S(_06007_),
    .X(_01935_));
 sg13g2_mux2_1 _24824_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net493),
    .S(_06010_),
    .X(_01936_));
 sg13g2_mux2_1 _24825_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net493),
    .S(_06014_),
    .X(_01937_));
 sg13g2_mux2_1 _24826_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net493),
    .S(_06019_),
    .X(_01938_));
 sg13g2_mux2_1 _24827_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net493),
    .S(_06025_),
    .X(_01939_));
 sg13g2_mux2_1 _24828_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(net493),
    .S(_06030_),
    .X(_01940_));
 sg13g2_mux2_1 _24829_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(_06366_),
    .S(_06033_),
    .X(_01941_));
 sg13g2_mux2_1 _24830_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_06366_),
    .S(_06036_),
    .X(_01942_));
 sg13g2_nor2_1 _24831_ (.A(net1071),
    .B(_09292_),
    .Y(_06367_));
 sg13g2_and3_1 _24832_ (.X(_06368_),
    .A(net1069),
    .B(_00237_),
    .C(_06367_));
 sg13g2_buf_2 _24833_ (.A(_06368_),
    .X(_06369_));
 sg13g2_and2_1 _24834_ (.A(net1066),
    .B(_06369_),
    .X(_06370_));
 sg13g2_buf_2 _24835_ (.A(_06370_),
    .X(_06371_));
 sg13g2_and3_1 _24836_ (.X(_06372_),
    .A(net984),
    .B(net384),
    .C(_06371_));
 sg13g2_buf_1 _24837_ (.A(_06372_),
    .X(_06373_));
 sg13g2_mux2_1 _24838_ (.A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net865),
    .S(_06373_),
    .X(_01959_));
 sg13g2_mux2_1 _24839_ (.A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1014),
    .S(_06373_),
    .X(_01960_));
 sg13g2_mux2_1 _24840_ (.A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1013),
    .S(_06373_),
    .X(_01961_));
 sg13g2_mux2_1 _24841_ (.A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1005),
    .S(_06373_),
    .X(_01962_));
 sg13g2_nand3_1 _24842_ (.B(_05183_),
    .C(_06371_),
    .A(net984),
    .Y(_06374_));
 sg13g2_buf_2 _24843_ (.A(_06374_),
    .X(_06375_));
 sg13g2_mux2_1 _24844_ (.A0(net896),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06375_),
    .X(_01963_));
 sg13g2_mux2_1 _24845_ (.A0(net1047),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06375_),
    .X(_01964_));
 sg13g2_mux2_1 _24846_ (.A0(net895),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06375_),
    .X(_01965_));
 sg13g2_mux2_1 _24847_ (.A0(net894),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .S(_06375_),
    .X(_01966_));
 sg13g2_mux2_1 _24848_ (.A0(net899),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .S(_06375_),
    .X(_01967_));
 sg13g2_nand2_1 _24849_ (.Y(_06376_),
    .A(_04872_),
    .B(_06371_));
 sg13g2_buf_4 _24850_ (.X(_06377_),
    .A(_06376_));
 sg13g2_mux2_1 _24851_ (.A0(net869),
    .A1(_04873_),
    .S(_06377_),
    .X(_01968_));
 sg13g2_buf_1 _24852_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06378_));
 sg13g2_mux2_1 _24853_ (.A0(net898),
    .A1(_06378_),
    .S(_06377_),
    .X(_01969_));
 sg13g2_mux2_1 _24854_ (.A0(net897),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(_06377_),
    .X(_01970_));
 sg13g2_mux2_1 _24855_ (.A0(net896),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .S(_06377_),
    .X(_01971_));
 sg13g2_mux2_1 _24856_ (.A0(net1047),
    .A1(_05547_),
    .S(_06377_),
    .X(_01972_));
 sg13g2_buf_1 _24857_ (.A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .X(_06379_));
 sg13g2_mux2_1 _24858_ (.A0(net895),
    .A1(_06379_),
    .S(_06377_),
    .X(_01973_));
 sg13g2_mux2_1 _24859_ (.A0(_10188_),
    .A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .S(_06377_),
    .X(_01974_));
 sg13g2_mux2_1 _24860_ (.A0(net899),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .S(_06377_),
    .X(_01975_));
 sg13g2_and3_1 _24861_ (.X(_06380_),
    .A(net544),
    .B(net505),
    .C(_06371_));
 sg13g2_buf_4 _24862_ (.X(_06381_),
    .A(_06380_));
 sg13g2_mux2_1 _24863_ (.A0(_04858_),
    .A1(net869),
    .S(_06381_),
    .X(_01976_));
 sg13g2_mux2_1 _24864_ (.A0(_05333_),
    .A1(net898),
    .S(_06381_),
    .X(_01977_));
 sg13g2_mux2_1 _24865_ (.A0(_05401_),
    .A1(net897),
    .S(_06381_),
    .X(_01978_));
 sg13g2_mux2_1 _24866_ (.A0(_05469_),
    .A1(net896),
    .S(_06381_),
    .X(_01979_));
 sg13g2_mux2_1 _24867_ (.A0(_05540_),
    .A1(net865),
    .S(_06381_),
    .X(_01980_));
 sg13g2_mux2_1 _24868_ (.A0(_05597_),
    .A1(net1014),
    .S(_06381_),
    .X(_01981_));
 sg13g2_mux2_1 _24869_ (.A0(_05687_),
    .A1(net1013),
    .S(_06381_),
    .X(_01982_));
 sg13g2_mux2_1 _24870_ (.A0(_05101_),
    .A1(net1005),
    .S(_06381_),
    .X(_01983_));
 sg13g2_nand3_1 _24871_ (.B(net505),
    .C(_06371_),
    .A(net543),
    .Y(_06382_));
 sg13g2_buf_4 _24872_ (.X(_06383_),
    .A(_06382_));
 sg13g2_mux2_1 _24873_ (.A0(net869),
    .A1(_04859_),
    .S(_06383_),
    .X(_01984_));
 sg13g2_buf_1 _24874_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06384_));
 sg13g2_mux2_1 _24875_ (.A0(net898),
    .A1(_06384_),
    .S(_06383_),
    .X(_01985_));
 sg13g2_mux2_1 _24876_ (.A0(net897),
    .A1(\cpu.gpio.r_src_io[6][2] ),
    .S(_06383_),
    .X(_01986_));
 sg13g2_mux2_1 _24877_ (.A0(net896),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .S(_06383_),
    .X(_01987_));
 sg13g2_mux2_1 _24878_ (.A0(net1047),
    .A1(_05541_),
    .S(_06383_),
    .X(_01988_));
 sg13g2_buf_1 _24879_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06385_));
 sg13g2_mux2_1 _24880_ (.A0(net895),
    .A1(_06385_),
    .S(_06383_),
    .X(_01989_));
 sg13g2_mux2_1 _24881_ (.A0(net894),
    .A1(\cpu.gpio.r_src_io[7][2] ),
    .S(_06383_),
    .X(_01990_));
 sg13g2_mux2_1 _24882_ (.A0(net899),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .S(_06383_),
    .X(_01991_));
 sg13g2_and3_1 _24883_ (.X(_06386_),
    .A(net662),
    .B(_04903_),
    .C(_06371_));
 sg13g2_buf_1 _24884_ (.A(_06386_),
    .X(_06387_));
 sg13g2_mux2_1 _24885_ (.A0(_05549_),
    .A1(net865),
    .S(_06387_),
    .X(_01992_));
 sg13g2_buf_1 _24886_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06388_));
 sg13g2_mux2_1 _24887_ (.A0(_06388_),
    .A1(net1014),
    .S(_06387_),
    .X(_01993_));
 sg13g2_mux2_1 _24888_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(net1013),
    .S(_06387_),
    .X(_01994_));
 sg13g2_mux2_1 _24889_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net1005),
    .S(_06387_),
    .X(_01995_));
 sg13g2_nand2_1 _24890_ (.Y(_06389_),
    .A(_04852_),
    .B(_06371_));
 sg13g2_buf_4 _24891_ (.X(_06390_),
    .A(_06389_));
 sg13g2_mux2_1 _24892_ (.A0(net869),
    .A1(_04848_),
    .S(_06390_),
    .X(_01996_));
 sg13g2_buf_1 _24893_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06391_));
 sg13g2_mux2_1 _24894_ (.A0(net898),
    .A1(_06391_),
    .S(_06390_),
    .X(_01997_));
 sg13g2_mux2_1 _24895_ (.A0(net897),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(_06390_),
    .X(_01998_));
 sg13g2_mux2_1 _24896_ (.A0(net896),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(_06390_),
    .X(_01999_));
 sg13g2_mux2_1 _24897_ (.A0(net1047),
    .A1(_05545_),
    .S(_06390_),
    .X(_02000_));
 sg13g2_buf_1 _24898_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06392_));
 sg13g2_mux2_1 _24899_ (.A0(net895),
    .A1(_06392_),
    .S(_06390_),
    .X(_02001_));
 sg13g2_mux2_1 _24900_ (.A0(net894),
    .A1(\cpu.gpio.r_src_o[5][2] ),
    .S(_06390_),
    .X(_02002_));
 sg13g2_mux2_1 _24901_ (.A0(net899),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .S(_06390_),
    .X(_02003_));
 sg13g2_nand2_2 _24902_ (.Y(_06393_),
    .A(_04864_),
    .B(_06371_));
 sg13g2_mux2_1 _24903_ (.A0(net1047),
    .A1(_05548_),
    .S(_06393_),
    .X(_02008_));
 sg13g2_buf_1 _24904_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06394_));
 sg13g2_mux2_1 _24905_ (.A0(net895),
    .A1(_06394_),
    .S(_06393_),
    .X(_02009_));
 sg13g2_mux2_1 _24906_ (.A0(net894),
    .A1(\cpu.gpio.r_src_o[7][2] ),
    .S(_06393_),
    .X(_02010_));
 sg13g2_mux2_1 _24907_ (.A0(net899),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .S(_06393_),
    .X(_02011_));
 sg13g2_buf_1 _24908_ (.A(net1111),
    .X(_06395_));
 sg13g2_and2_1 _24909_ (.A(net815),
    .B(_08856_),
    .X(_06396_));
 sg13g2_buf_4 _24910_ (.X(_06397_),
    .A(_06396_));
 sg13g2_buf_1 _24911_ (.A(\cpu.icache.r_offset[2] ),
    .X(_06398_));
 sg13g2_buf_2 _24912_ (.A(_00255_),
    .X(_06399_));
 sg13g2_buf_1 _24913_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06400_));
 sg13g2_buf_1 _24914_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06401_));
 sg13g2_nand2b_1 _24915_ (.Y(_06402_),
    .B(_06401_),
    .A_N(_06400_));
 sg13g2_nor3_1 _24916_ (.A(_06398_),
    .B(_06399_),
    .C(_06402_),
    .Y(_06403_));
 sg13g2_buf_2 _24917_ (.A(_06403_),
    .X(_06404_));
 sg13g2_nand2_2 _24918_ (.Y(_06405_),
    .A(_06397_),
    .B(_06404_));
 sg13g2_mux2_1 _24919_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06405_),
    .X(_02015_));
 sg13g2_buf_1 _24920_ (.A(net1110),
    .X(_06406_));
 sg13g2_buf_1 _24921_ (.A(_00256_),
    .X(_06407_));
 sg13g2_inv_1 _24922_ (.Y(_06408_),
    .A(_06407_));
 sg13g2_nand2_1 _24923_ (.Y(_06409_),
    .A(_06400_),
    .B(_06401_));
 sg13g2_nor3_1 _24924_ (.A(_06399_),
    .B(_06408_),
    .C(_06409_),
    .Y(_06410_));
 sg13g2_buf_2 _24925_ (.A(_06410_),
    .X(_06411_));
 sg13g2_nand2_2 _24926_ (.Y(_06412_),
    .A(_06397_),
    .B(_06411_));
 sg13g2_mux2_1 _24927_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06412_),
    .X(_02016_));
 sg13g2_buf_1 _24928_ (.A(net1109),
    .X(_06413_));
 sg13g2_mux2_1 _24929_ (.A0(_06413_),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06412_),
    .X(_02017_));
 sg13g2_nand2b_1 _24930_ (.Y(_06414_),
    .B(_06400_),
    .A_N(_06401_));
 sg13g2_nor3_1 _24931_ (.A(_06398_),
    .B(_06399_),
    .C(_06414_),
    .Y(_06415_));
 sg13g2_buf_2 _24932_ (.A(_06415_),
    .X(_06416_));
 sg13g2_nand2_2 _24933_ (.Y(_06417_),
    .A(_06397_),
    .B(_06416_));
 sg13g2_mux2_1 _24934_ (.A0(_06395_),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06417_),
    .X(_02018_));
 sg13g2_buf_1 _24935_ (.A(net1108),
    .X(_06418_));
 sg13g2_mux2_1 _24936_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06417_),
    .X(_02019_));
 sg13g2_mux2_1 _24937_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06417_),
    .X(_02020_));
 sg13g2_mux2_1 _24938_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06417_),
    .X(_02021_));
 sg13g2_nor3_1 _24939_ (.A(_06399_),
    .B(_06407_),
    .C(_06402_),
    .Y(_06419_));
 sg13g2_buf_4 _24940_ (.X(_06420_),
    .A(_06419_));
 sg13g2_nand2_2 _24941_ (.Y(_06421_),
    .A(_06397_),
    .B(_06420_));
 sg13g2_mux2_1 _24942_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06421_),
    .X(_02022_));
 sg13g2_mux2_1 _24943_ (.A0(_06418_),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06421_),
    .X(_02023_));
 sg13g2_mux2_1 _24944_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06421_),
    .X(_02024_));
 sg13g2_mux2_1 _24945_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06421_),
    .X(_02025_));
 sg13g2_mux2_1 _24946_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06405_),
    .X(_02026_));
 sg13g2_nor4_1 _24947_ (.A(_06400_),
    .B(_06401_),
    .C(_06399_),
    .D(_06407_),
    .Y(_06422_));
 sg13g2_buf_2 _24948_ (.A(_06422_),
    .X(_06423_));
 sg13g2_nand2_2 _24949_ (.Y(_06424_),
    .A(_06397_),
    .B(_06423_));
 sg13g2_mux2_1 _24950_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06424_),
    .X(_02027_));
 sg13g2_mux2_1 _24951_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06424_),
    .X(_02028_));
 sg13g2_mux2_1 _24952_ (.A0(_06406_),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06424_),
    .X(_02029_));
 sg13g2_mux2_1 _24953_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06424_),
    .X(_02030_));
 sg13g2_inv_1 _24954_ (.Y(_06425_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_1 _24955_ (.A(_06407_),
    .B(_06425_),
    .C(_06409_),
    .Y(_06426_));
 sg13g2_buf_2 _24956_ (.A(_06426_),
    .X(_06427_));
 sg13g2_nand2_1 _24957_ (.Y(_06428_),
    .A(_06397_),
    .B(_06427_));
 sg13g2_buf_1 _24958_ (.A(_06428_),
    .X(_06429_));
 sg13g2_buf_1 _24959_ (.A(_06429_),
    .X(_06430_));
 sg13g2_mux2_1 _24960_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(_06430_),
    .X(_02031_));
 sg13g2_mux2_1 _24961_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(_06430_),
    .X(_02032_));
 sg13g2_mux2_1 _24962_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net406),
    .X(_02033_));
 sg13g2_buf_1 _24963_ (.A(_06429_),
    .X(_06431_));
 sg13g2_mux2_1 _24964_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net405),
    .X(_02034_));
 sg13g2_nor3_1 _24965_ (.A(_06399_),
    .B(_06407_),
    .C(_06414_),
    .Y(_06432_));
 sg13g2_buf_4 _24966_ (.X(_06433_),
    .A(_06432_));
 sg13g2_nand2_2 _24967_ (.Y(_06434_),
    .A(_06397_),
    .B(_06433_));
 sg13g2_mux2_1 _24968_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06434_),
    .X(_02035_));
 sg13g2_mux2_1 _24969_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06434_),
    .X(_02036_));
 sg13g2_mux2_1 _24970_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06405_),
    .X(_02037_));
 sg13g2_mux2_1 _24971_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06434_),
    .X(_02038_));
 sg13g2_mux2_1 _24972_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06434_),
    .X(_02039_));
 sg13g2_mux2_1 _24973_ (.A0(_06413_),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06405_),
    .X(_02040_));
 sg13g2_nor4_1 _24974_ (.A(_06400_),
    .B(_06401_),
    .C(_06398_),
    .D(_06399_),
    .Y(_06435_));
 sg13g2_buf_2 _24975_ (.A(_06435_),
    .X(_06436_));
 sg13g2_nand2_2 _24976_ (.Y(_06437_),
    .A(_06397_),
    .B(_06436_));
 sg13g2_mux2_1 _24977_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06437_),
    .X(_02041_));
 sg13g2_mux2_1 _24978_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06437_),
    .X(_02042_));
 sg13g2_mux2_1 _24979_ (.A0(net969),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06437_),
    .X(_02043_));
 sg13g2_mux2_1 _24980_ (.A0(net968),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06437_),
    .X(_02044_));
 sg13g2_mux2_1 _24981_ (.A0(net970),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06412_),
    .X(_02045_));
 sg13g2_mux2_1 _24982_ (.A0(net967),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06412_),
    .X(_02046_));
 sg13g2_buf_1 _24983_ (.A(net1111),
    .X(_06438_));
 sg13g2_and2_1 _24984_ (.A(net524),
    .B(_06404_),
    .X(_06439_));
 sg13g2_buf_1 _24985_ (.A(_06439_),
    .X(_06440_));
 sg13g2_mux2_1 _24986_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(_06438_),
    .S(_06440_),
    .X(_02047_));
 sg13g2_buf_1 _24987_ (.A(net1110),
    .X(_06441_));
 sg13g2_and2_1 _24988_ (.A(net524),
    .B(_06411_),
    .X(_06442_));
 sg13g2_buf_1 _24989_ (.A(_06442_),
    .X(_06443_));
 sg13g2_mux2_1 _24990_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net965),
    .S(_06443_),
    .X(_02048_));
 sg13g2_buf_1 _24991_ (.A(net1109),
    .X(_06444_));
 sg13g2_mux2_1 _24992_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net964),
    .S(_06443_),
    .X(_02049_));
 sg13g2_and2_1 _24993_ (.A(net524),
    .B(_06416_),
    .X(_06445_));
 sg13g2_buf_1 _24994_ (.A(_06445_),
    .X(_06446_));
 sg13g2_mux2_1 _24995_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net966),
    .S(_06446_),
    .X(_02050_));
 sg13g2_buf_1 _24996_ (.A(net1108),
    .X(_06447_));
 sg13g2_mux2_1 _24997_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net963),
    .S(_06446_),
    .X(_02051_));
 sg13g2_mux2_1 _24998_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net965),
    .S(_06446_),
    .X(_02052_));
 sg13g2_mux2_1 _24999_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net964),
    .S(_06446_),
    .X(_02053_));
 sg13g2_and2_1 _25000_ (.A(net524),
    .B(_06420_),
    .X(_06448_));
 sg13g2_buf_1 _25001_ (.A(_06448_),
    .X(_06449_));
 sg13g2_mux2_1 _25002_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net966),
    .S(_06449_),
    .X(_02054_));
 sg13g2_mux2_1 _25003_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net963),
    .S(_06449_),
    .X(_02055_));
 sg13g2_mux2_1 _25004_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net965),
    .S(_06449_),
    .X(_02056_));
 sg13g2_mux2_1 _25005_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(_06444_),
    .S(_06449_),
    .X(_02057_));
 sg13g2_mux2_1 _25006_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net963),
    .S(_06440_),
    .X(_02058_));
 sg13g2_buf_1 _25007_ (.A(net1111),
    .X(_06450_));
 sg13g2_and2_1 _25008_ (.A(_03114_),
    .B(_06423_),
    .X(_06451_));
 sg13g2_buf_1 _25009_ (.A(_06451_),
    .X(_06452_));
 sg13g2_mux2_1 _25010_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net962),
    .S(_06452_),
    .X(_02059_));
 sg13g2_buf_1 _25011_ (.A(net1108),
    .X(_06453_));
 sg13g2_mux2_1 _25012_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net961),
    .S(_06452_),
    .X(_02060_));
 sg13g2_buf_1 _25013_ (.A(net1110),
    .X(_06454_));
 sg13g2_mux2_1 _25014_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(_06454_),
    .S(_06452_),
    .X(_02061_));
 sg13g2_buf_1 _25015_ (.A(net1109),
    .X(_06455_));
 sg13g2_mux2_1 _25016_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net959),
    .S(_06452_),
    .X(_02062_));
 sg13g2_and2_1 _25017_ (.A(net524),
    .B(_06427_),
    .X(_06456_));
 sg13g2_buf_2 _25018_ (.A(_06456_),
    .X(_06457_));
 sg13g2_mux2_1 _25019_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net962),
    .S(_06457_),
    .X(_02063_));
 sg13g2_mux2_1 _25020_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net961),
    .S(_06457_),
    .X(_02064_));
 sg13g2_mux2_1 _25021_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(net960),
    .S(_06457_),
    .X(_02065_));
 sg13g2_mux2_1 _25022_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net959),
    .S(_06457_),
    .X(_02066_));
 sg13g2_and2_1 _25023_ (.A(_03114_),
    .B(_06433_),
    .X(_06458_));
 sg13g2_buf_1 _25024_ (.A(_06458_),
    .X(_06459_));
 sg13g2_mux2_1 _25025_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net962),
    .S(_06459_),
    .X(_02067_));
 sg13g2_mux2_1 _25026_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(_06453_),
    .S(_06459_),
    .X(_02068_));
 sg13g2_mux2_1 _25027_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net960),
    .S(_06440_),
    .X(_02069_));
 sg13g2_mux2_1 _25028_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net960),
    .S(_06459_),
    .X(_02070_));
 sg13g2_mux2_1 _25029_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net959),
    .S(_06459_),
    .X(_02071_));
 sg13g2_mux2_1 _25030_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net959),
    .S(_06440_),
    .X(_02072_));
 sg13g2_and2_1 _25031_ (.A(net524),
    .B(_06436_),
    .X(_06460_));
 sg13g2_buf_1 _25032_ (.A(_06460_),
    .X(_06461_));
 sg13g2_mux2_1 _25033_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net962),
    .S(_06461_),
    .X(_02073_));
 sg13g2_mux2_1 _25034_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net961),
    .S(_06461_),
    .X(_02074_));
 sg13g2_mux2_1 _25035_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net960),
    .S(_06461_),
    .X(_02075_));
 sg13g2_mux2_1 _25036_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net959),
    .S(_06461_),
    .X(_02076_));
 sg13g2_mux2_1 _25037_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(_06450_),
    .S(_06443_),
    .X(_02077_));
 sg13g2_mux2_1 _25038_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(_06453_),
    .S(_06443_),
    .X(_02078_));
 sg13g2_and2_1 _25039_ (.A(net463),
    .B(_06404_),
    .X(_06462_));
 sg13g2_buf_2 _25040_ (.A(_06462_),
    .X(_06463_));
 sg13g2_mux2_1 _25041_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(_06450_),
    .S(_06463_),
    .X(_02079_));
 sg13g2_and2_1 _25042_ (.A(_03115_),
    .B(_06411_),
    .X(_06464_));
 sg13g2_buf_1 _25043_ (.A(_06464_),
    .X(_06465_));
 sg13g2_mux2_1 _25044_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net960),
    .S(_06465_),
    .X(_02080_));
 sg13g2_mux2_1 _25045_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(_06455_),
    .S(_06465_),
    .X(_02081_));
 sg13g2_and2_1 _25046_ (.A(net463),
    .B(_06416_),
    .X(_06466_));
 sg13g2_buf_1 _25047_ (.A(_06466_),
    .X(_06467_));
 sg13g2_mux2_1 _25048_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net962),
    .S(_06467_),
    .X(_02082_));
 sg13g2_mux2_1 _25049_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net961),
    .S(_06467_),
    .X(_02083_));
 sg13g2_mux2_1 _25050_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net960),
    .S(_06467_),
    .X(_02084_));
 sg13g2_mux2_1 _25051_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net959),
    .S(_06467_),
    .X(_02085_));
 sg13g2_and2_1 _25052_ (.A(net463),
    .B(_06420_),
    .X(_06468_));
 sg13g2_buf_1 _25053_ (.A(_06468_),
    .X(_06469_));
 sg13g2_mux2_1 _25054_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net962),
    .S(_06469_),
    .X(_02086_));
 sg13g2_mux2_1 _25055_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net961),
    .S(_06469_),
    .X(_02087_));
 sg13g2_mux2_1 _25056_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(_06454_),
    .S(_06469_),
    .X(_02088_));
 sg13g2_mux2_1 _25057_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(_06455_),
    .S(_06469_),
    .X(_02089_));
 sg13g2_mux2_1 _25058_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net961),
    .S(_06463_),
    .X(_02090_));
 sg13g2_and2_1 _25059_ (.A(net463),
    .B(_06423_),
    .X(_06470_));
 sg13g2_buf_1 _25060_ (.A(_06470_),
    .X(_06471_));
 sg13g2_mux2_1 _25061_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net962),
    .S(_06471_),
    .X(_02091_));
 sg13g2_mux2_1 _25062_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net961),
    .S(_06471_),
    .X(_02092_));
 sg13g2_mux2_1 _25063_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net960),
    .S(_06471_),
    .X(_02093_));
 sg13g2_mux2_1 _25064_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net959),
    .S(_06471_),
    .X(_02094_));
 sg13g2_and2_1 _25065_ (.A(net463),
    .B(_06427_),
    .X(_06472_));
 sg13g2_buf_2 _25066_ (.A(_06472_),
    .X(_06473_));
 sg13g2_mux2_1 _25067_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net962),
    .S(_06473_),
    .X(_02095_));
 sg13g2_mux2_1 _25068_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net961),
    .S(_06473_),
    .X(_02096_));
 sg13g2_mux2_1 _25069_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net960),
    .S(_06473_),
    .X(_02097_));
 sg13g2_mux2_1 _25070_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net959),
    .S(_06473_),
    .X(_02098_));
 sg13g2_buf_1 _25071_ (.A(_12052_),
    .X(_06474_));
 sg13g2_and2_1 _25072_ (.A(_03115_),
    .B(_06433_),
    .X(_06475_));
 sg13g2_buf_1 _25073_ (.A(_06475_),
    .X(_06476_));
 sg13g2_mux2_1 _25074_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net958),
    .S(_06476_),
    .X(_02099_));
 sg13g2_buf_1 _25075_ (.A(_12119_),
    .X(_06477_));
 sg13g2_mux2_1 _25076_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net957),
    .S(_06476_),
    .X(_02100_));
 sg13g2_buf_1 _25077_ (.A(_12087_),
    .X(_06478_));
 sg13g2_mux2_1 _25078_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net956),
    .S(_06463_),
    .X(_02101_));
 sg13g2_mux2_1 _25079_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net956),
    .S(_06476_),
    .X(_02102_));
 sg13g2_buf_2 _25080_ (.A(net1117),
    .X(_06479_));
 sg13g2_mux2_1 _25081_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net955),
    .S(_06476_),
    .X(_02103_));
 sg13g2_mux2_1 _25082_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net955),
    .S(_06463_),
    .X(_02104_));
 sg13g2_and2_1 _25083_ (.A(net463),
    .B(_06436_),
    .X(_06480_));
 sg13g2_buf_1 _25084_ (.A(_06480_),
    .X(_06481_));
 sg13g2_mux2_1 _25085_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net958),
    .S(_06481_),
    .X(_02105_));
 sg13g2_mux2_1 _25086_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net957),
    .S(_06481_),
    .X(_02106_));
 sg13g2_mux2_1 _25087_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net956),
    .S(_06481_),
    .X(_02107_));
 sg13g2_mux2_1 _25088_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net955),
    .S(_06481_),
    .X(_02108_));
 sg13g2_mux2_1 _25089_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net958),
    .S(_06465_),
    .X(_02109_));
 sg13g2_mux2_1 _25090_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net957),
    .S(_06465_),
    .X(_02110_));
 sg13g2_nand2_2 _25091_ (.Y(_06482_),
    .A(net546),
    .B(_06404_));
 sg13g2_mux2_1 _25092_ (.A0(_06395_),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06482_),
    .X(_02111_));
 sg13g2_and2_1 _25093_ (.A(_09021_),
    .B(_06411_),
    .X(_06483_));
 sg13g2_buf_1 _25094_ (.A(_06483_),
    .X(_06484_));
 sg13g2_mux2_1 _25095_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net956),
    .S(_06484_),
    .X(_02112_));
 sg13g2_mux2_1 _25096_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net955),
    .S(_06484_),
    .X(_02113_));
 sg13g2_nand2_2 _25097_ (.Y(_06485_),
    .A(net546),
    .B(_06416_));
 sg13g2_mux2_1 _25098_ (.A0(net970),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06485_),
    .X(_02114_));
 sg13g2_mux2_1 _25099_ (.A0(net967),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06485_),
    .X(_02115_));
 sg13g2_mux2_1 _25100_ (.A0(net969),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06485_),
    .X(_02116_));
 sg13g2_mux2_1 _25101_ (.A0(net968),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06485_),
    .X(_02117_));
 sg13g2_buf_1 _25102_ (.A(_02909_),
    .X(_06486_));
 sg13g2_nand2_2 _25103_ (.Y(_06487_),
    .A(net546),
    .B(_06420_));
 sg13g2_mux2_1 _25104_ (.A0(net954),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06487_),
    .X(_02118_));
 sg13g2_mux2_1 _25105_ (.A0(_06418_),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06487_),
    .X(_02119_));
 sg13g2_mux2_1 _25106_ (.A0(_06406_),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06487_),
    .X(_02120_));
 sg13g2_mux2_1 _25107_ (.A0(net968),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06487_),
    .X(_02121_));
 sg13g2_buf_1 _25108_ (.A(_02933_),
    .X(_06488_));
 sg13g2_mux2_1 _25109_ (.A0(net953),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06482_),
    .X(_02122_));
 sg13g2_nand2_2 _25110_ (.Y(_06489_),
    .A(_09021_),
    .B(_06423_));
 sg13g2_mux2_1 _25111_ (.A0(_06486_),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06489_),
    .X(_02123_));
 sg13g2_mux2_1 _25112_ (.A0(_06488_),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06489_),
    .X(_02124_));
 sg13g2_buf_1 _25113_ (.A(_02918_),
    .X(_06490_));
 sg13g2_mux2_1 _25114_ (.A0(net952),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06489_),
    .X(_02125_));
 sg13g2_buf_1 _25115_ (.A(_02922_),
    .X(_06491_));
 sg13g2_mux2_1 _25116_ (.A0(_06491_),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06489_),
    .X(_02126_));
 sg13g2_nand2_1 _25117_ (.Y(_06492_),
    .A(net546),
    .B(_06427_));
 sg13g2_buf_1 _25118_ (.A(_06492_),
    .X(_06493_));
 sg13g2_buf_1 _25119_ (.A(_06493_),
    .X(_06494_));
 sg13g2_mux2_1 _25120_ (.A0(net954),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net360),
    .X(_02127_));
 sg13g2_mux2_1 _25121_ (.A0(net953),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(_06494_),
    .X(_02128_));
 sg13g2_mux2_1 _25122_ (.A0(net952),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net360),
    .X(_02129_));
 sg13g2_buf_1 _25123_ (.A(_06493_),
    .X(_06495_));
 sg13g2_mux2_1 _25124_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(_06495_),
    .X(_02130_));
 sg13g2_nand2_2 _25125_ (.Y(_06496_),
    .A(net546),
    .B(_06433_));
 sg13g2_mux2_1 _25126_ (.A0(_06486_),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06496_),
    .X(_02131_));
 sg13g2_mux2_1 _25127_ (.A0(net953),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06496_),
    .X(_02132_));
 sg13g2_mux2_1 _25128_ (.A0(_06490_),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06482_),
    .X(_02133_));
 sg13g2_mux2_1 _25129_ (.A0(net952),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06496_),
    .X(_02134_));
 sg13g2_mux2_1 _25130_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06496_),
    .X(_02135_));
 sg13g2_mux2_1 _25131_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06482_),
    .X(_02136_));
 sg13g2_nand2_2 _25132_ (.Y(_06497_),
    .A(net546),
    .B(_06436_));
 sg13g2_mux2_1 _25133_ (.A0(net954),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06497_),
    .X(_02137_));
 sg13g2_mux2_1 _25134_ (.A0(_06488_),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06497_),
    .X(_02138_));
 sg13g2_mux2_1 _25135_ (.A0(_06490_),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06497_),
    .X(_02139_));
 sg13g2_mux2_1 _25136_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06497_),
    .X(_02140_));
 sg13g2_mux2_1 _25137_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net958),
    .S(_06484_),
    .X(_02141_));
 sg13g2_mux2_1 _25138_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net957),
    .S(_06484_),
    .X(_02142_));
 sg13g2_nand2_2 _25139_ (.Y(_06498_),
    .A(net522),
    .B(_06404_));
 sg13g2_mux2_1 _25140_ (.A0(net954),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06498_),
    .X(_02143_));
 sg13g2_and2_1 _25141_ (.A(net522),
    .B(_06411_),
    .X(_06499_));
 sg13g2_buf_1 _25142_ (.A(_06499_),
    .X(_06500_));
 sg13g2_mux2_1 _25143_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net956),
    .S(_06500_),
    .X(_02144_));
 sg13g2_mux2_1 _25144_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net955),
    .S(_06500_),
    .X(_02145_));
 sg13g2_nand2_2 _25145_ (.Y(_06501_),
    .A(net522),
    .B(_06416_));
 sg13g2_mux2_1 _25146_ (.A0(net954),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06501_),
    .X(_02146_));
 sg13g2_mux2_1 _25147_ (.A0(net953),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06501_),
    .X(_02147_));
 sg13g2_mux2_1 _25148_ (.A0(net952),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06501_),
    .X(_02148_));
 sg13g2_mux2_1 _25149_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06501_),
    .X(_02149_));
 sg13g2_nand2_2 _25150_ (.Y(_06502_),
    .A(net522),
    .B(_06420_));
 sg13g2_mux2_1 _25151_ (.A0(net954),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06502_),
    .X(_02150_));
 sg13g2_mux2_1 _25152_ (.A0(net953),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06502_),
    .X(_02151_));
 sg13g2_mux2_1 _25153_ (.A0(net952),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06502_),
    .X(_02152_));
 sg13g2_mux2_1 _25154_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06502_),
    .X(_02153_));
 sg13g2_mux2_1 _25155_ (.A0(net953),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06498_),
    .X(_02154_));
 sg13g2_nand2_2 _25156_ (.Y(_06503_),
    .A(_03118_),
    .B(_06423_));
 sg13g2_mux2_1 _25157_ (.A0(net954),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06503_),
    .X(_02155_));
 sg13g2_mux2_1 _25158_ (.A0(net953),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06503_),
    .X(_02156_));
 sg13g2_mux2_1 _25159_ (.A0(net952),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06503_),
    .X(_02157_));
 sg13g2_mux2_1 _25160_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06503_),
    .X(_02158_));
 sg13g2_and2_1 _25161_ (.A(net522),
    .B(_06427_),
    .X(_06504_));
 sg13g2_buf_2 _25162_ (.A(_06504_),
    .X(_06505_));
 sg13g2_mux2_1 _25163_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net958),
    .S(_06505_),
    .X(_02159_));
 sg13g2_mux2_1 _25164_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net957),
    .S(_06505_),
    .X(_02160_));
 sg13g2_mux2_1 _25165_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net956),
    .S(_06505_),
    .X(_02161_));
 sg13g2_mux2_1 _25166_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(net955),
    .S(_06505_),
    .X(_02162_));
 sg13g2_nand2_2 _25167_ (.Y(_06506_),
    .A(_03118_),
    .B(_06433_));
 sg13g2_mux2_1 _25168_ (.A0(net954),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06506_),
    .X(_02163_));
 sg13g2_mux2_1 _25169_ (.A0(net953),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06506_),
    .X(_02164_));
 sg13g2_mux2_1 _25170_ (.A0(net952),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06498_),
    .X(_02165_));
 sg13g2_mux2_1 _25171_ (.A0(net952),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06506_),
    .X(_02166_));
 sg13g2_mux2_1 _25172_ (.A0(_06491_),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06506_),
    .X(_02167_));
 sg13g2_mux2_1 _25173_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06498_),
    .X(_02168_));
 sg13g2_buf_1 _25174_ (.A(_02909_),
    .X(_06507_));
 sg13g2_nand2_2 _25175_ (.Y(_06508_),
    .A(net522),
    .B(_06436_));
 sg13g2_mux2_1 _25176_ (.A0(net950),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06508_),
    .X(_02169_));
 sg13g2_buf_1 _25177_ (.A(_02933_),
    .X(_06509_));
 sg13g2_mux2_1 _25178_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06508_),
    .X(_02170_));
 sg13g2_buf_1 _25179_ (.A(_02918_),
    .X(_06510_));
 sg13g2_mux2_1 _25180_ (.A0(net948),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06508_),
    .X(_02171_));
 sg13g2_buf_1 _25181_ (.A(_02922_),
    .X(_06511_));
 sg13g2_mux2_1 _25182_ (.A0(net947),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06508_),
    .X(_02172_));
 sg13g2_mux2_1 _25183_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net958),
    .S(_06500_),
    .X(_02173_));
 sg13g2_mux2_1 _25184_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(net957),
    .S(_06500_),
    .X(_02174_));
 sg13g2_nand2_2 _25185_ (.Y(_06512_),
    .A(net625),
    .B(_06404_));
 sg13g2_mux2_1 _25186_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][0] ),
    .S(_06512_),
    .X(_02175_));
 sg13g2_nand2_2 _25187_ (.Y(_06513_),
    .A(net625),
    .B(_06411_));
 sg13g2_mux2_1 _25188_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][10] ),
    .S(_06513_),
    .X(_02176_));
 sg13g2_mux2_1 _25189_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][11] ),
    .S(_06513_),
    .X(_02177_));
 sg13g2_nand2_2 _25190_ (.Y(_06514_),
    .A(net625),
    .B(_06416_));
 sg13g2_mux2_1 _25191_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][12] ),
    .S(_06514_),
    .X(_02178_));
 sg13g2_mux2_1 _25192_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][13] ),
    .S(_06514_),
    .X(_02179_));
 sg13g2_mux2_1 _25193_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][14] ),
    .S(_06514_),
    .X(_02180_));
 sg13g2_mux2_1 _25194_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][15] ),
    .S(_06514_),
    .X(_02181_));
 sg13g2_nand2_2 _25195_ (.Y(_06515_),
    .A(_09002_),
    .B(_06420_));
 sg13g2_mux2_1 _25196_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][16] ),
    .S(_06515_),
    .X(_02182_));
 sg13g2_mux2_1 _25197_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][17] ),
    .S(_06515_),
    .X(_02183_));
 sg13g2_mux2_1 _25198_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][18] ),
    .S(_06515_),
    .X(_02184_));
 sg13g2_mux2_1 _25199_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][19] ),
    .S(_06515_),
    .X(_02185_));
 sg13g2_mux2_1 _25200_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][1] ),
    .S(_06512_),
    .X(_02186_));
 sg13g2_nand2_2 _25201_ (.Y(_06516_),
    .A(_09002_),
    .B(_06423_));
 sg13g2_mux2_1 _25202_ (.A0(_06507_),
    .A1(\cpu.icache.r_data[5][20] ),
    .S(_06516_),
    .X(_02187_));
 sg13g2_mux2_1 _25203_ (.A0(_06509_),
    .A1(\cpu.icache.r_data[5][21] ),
    .S(_06516_),
    .X(_02188_));
 sg13g2_mux2_1 _25204_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[5][22] ),
    .S(_06516_),
    .X(_02189_));
 sg13g2_mux2_1 _25205_ (.A0(_06511_),
    .A1(\cpu.icache.r_data[5][23] ),
    .S(_06516_),
    .X(_02190_));
 sg13g2_nand2_1 _25206_ (.Y(_06517_),
    .A(net625),
    .B(_06427_));
 sg13g2_buf_2 _25207_ (.A(_06517_),
    .X(_06518_));
 sg13g2_mux2_1 _25208_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][24] ),
    .S(_06518_),
    .X(_02191_));
 sg13g2_mux2_1 _25209_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][25] ),
    .S(_06518_),
    .X(_02192_));
 sg13g2_mux2_1 _25210_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][26] ),
    .S(_06518_),
    .X(_02193_));
 sg13g2_mux2_1 _25211_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][27] ),
    .S(_06518_),
    .X(_02194_));
 sg13g2_nand2_2 _25212_ (.Y(_06519_),
    .A(net625),
    .B(_06433_));
 sg13g2_mux2_1 _25213_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][28] ),
    .S(_06519_),
    .X(_02195_));
 sg13g2_mux2_1 _25214_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][29] ),
    .S(_06519_),
    .X(_02196_));
 sg13g2_mux2_1 _25215_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][2] ),
    .S(_06512_),
    .X(_02197_));
 sg13g2_mux2_1 _25216_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[5][30] ),
    .S(_06519_),
    .X(_02198_));
 sg13g2_mux2_1 _25217_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][31] ),
    .S(_06519_),
    .X(_02199_));
 sg13g2_mux2_1 _25218_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][3] ),
    .S(_06512_),
    .X(_02200_));
 sg13g2_nand2_2 _25219_ (.Y(_06520_),
    .A(net625),
    .B(_06436_));
 sg13g2_mux2_1 _25220_ (.A0(net950),
    .A1(\cpu.icache.r_data[5][4] ),
    .S(_06520_),
    .X(_02201_));
 sg13g2_mux2_1 _25221_ (.A0(net949),
    .A1(\cpu.icache.r_data[5][5] ),
    .S(_06520_),
    .X(_02202_));
 sg13g2_mux2_1 _25222_ (.A0(net948),
    .A1(\cpu.icache.r_data[5][6] ),
    .S(_06520_),
    .X(_02203_));
 sg13g2_mux2_1 _25223_ (.A0(net947),
    .A1(\cpu.icache.r_data[5][7] ),
    .S(_06520_),
    .X(_02204_));
 sg13g2_mux2_1 _25224_ (.A0(_06507_),
    .A1(\cpu.icache.r_data[5][8] ),
    .S(_06513_),
    .X(_02205_));
 sg13g2_mux2_1 _25225_ (.A0(_06509_),
    .A1(\cpu.icache.r_data[5][9] ),
    .S(_06513_),
    .X(_02206_));
 sg13g2_nand2_2 _25226_ (.Y(_06521_),
    .A(net523),
    .B(_06404_));
 sg13g2_mux2_1 _25227_ (.A0(net950),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06521_),
    .X(_02207_));
 sg13g2_nand2_2 _25228_ (.Y(_06522_),
    .A(net523),
    .B(_06411_));
 sg13g2_mux2_1 _25229_ (.A0(net948),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06522_),
    .X(_02208_));
 sg13g2_mux2_1 _25230_ (.A0(_06511_),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06522_),
    .X(_02209_));
 sg13g2_nand2_2 _25231_ (.Y(_06523_),
    .A(net523),
    .B(_06416_));
 sg13g2_mux2_1 _25232_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06523_),
    .X(_02210_));
 sg13g2_mux2_1 _25233_ (.A0(net949),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06523_),
    .X(_02211_));
 sg13g2_mux2_1 _25234_ (.A0(net965),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06523_),
    .X(_02212_));
 sg13g2_mux2_1 _25235_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06523_),
    .X(_02213_));
 sg13g2_nand2_2 _25236_ (.Y(_06524_),
    .A(net523),
    .B(_06420_));
 sg13g2_mux2_1 _25237_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06524_),
    .X(_02214_));
 sg13g2_mux2_1 _25238_ (.A0(net963),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06524_),
    .X(_02215_));
 sg13g2_mux2_1 _25239_ (.A0(net965),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06524_),
    .X(_02216_));
 sg13g2_mux2_1 _25240_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06524_),
    .X(_02217_));
 sg13g2_mux2_1 _25241_ (.A0(net963),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06521_),
    .X(_02218_));
 sg13g2_nand2_2 _25242_ (.Y(_06525_),
    .A(_03117_),
    .B(_06423_));
 sg13g2_mux2_1 _25243_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06525_),
    .X(_02219_));
 sg13g2_mux2_1 _25244_ (.A0(_06447_),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06525_),
    .X(_02220_));
 sg13g2_mux2_1 _25245_ (.A0(_06441_),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06525_),
    .X(_02221_));
 sg13g2_mux2_1 _25246_ (.A0(_06444_),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06525_),
    .X(_02222_));
 sg13g2_nand2_1 _25247_ (.Y(_06526_),
    .A(net523),
    .B(_06427_));
 sg13g2_buf_2 _25248_ (.A(_06526_),
    .X(_06527_));
 sg13g2_mux2_1 _25249_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06527_),
    .X(_02223_));
 sg13g2_mux2_1 _25250_ (.A0(net963),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06527_),
    .X(_02224_));
 sg13g2_mux2_1 _25251_ (.A0(net965),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06527_),
    .X(_02225_));
 sg13g2_mux2_1 _25252_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06527_),
    .X(_02226_));
 sg13g2_nand2_2 _25253_ (.Y(_06528_),
    .A(_03117_),
    .B(_06433_));
 sg13g2_mux2_1 _25254_ (.A0(_06438_),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06528_),
    .X(_02227_));
 sg13g2_mux2_1 _25255_ (.A0(net963),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06528_),
    .X(_02228_));
 sg13g2_mux2_1 _25256_ (.A0(net965),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06521_),
    .X(_02229_));
 sg13g2_mux2_1 _25257_ (.A0(_06441_),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06528_),
    .X(_02230_));
 sg13g2_mux2_1 _25258_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06528_),
    .X(_02231_));
 sg13g2_mux2_1 _25259_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06521_),
    .X(_02232_));
 sg13g2_nand2_2 _25260_ (.Y(_06529_),
    .A(net523),
    .B(_06436_));
 sg13g2_mux2_1 _25261_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06529_),
    .X(_02233_));
 sg13g2_mux2_1 _25262_ (.A0(net963),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06529_),
    .X(_02234_));
 sg13g2_mux2_1 _25263_ (.A0(net965),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06529_),
    .X(_02235_));
 sg13g2_mux2_1 _25264_ (.A0(net964),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06529_),
    .X(_02236_));
 sg13g2_mux2_1 _25265_ (.A0(net966),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06522_),
    .X(_02237_));
 sg13g2_mux2_1 _25266_ (.A0(_06447_),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06522_),
    .X(_02238_));
 sg13g2_and2_1 _25267_ (.A(net626),
    .B(_06404_),
    .X(_06530_));
 sg13g2_buf_1 _25268_ (.A(_06530_),
    .X(_06531_));
 sg13g2_mux2_1 _25269_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net958),
    .S(_06531_),
    .X(_02239_));
 sg13g2_and2_1 _25270_ (.A(_08956_),
    .B(_06411_),
    .X(_06532_));
 sg13g2_buf_1 _25271_ (.A(_06532_),
    .X(_06533_));
 sg13g2_mux2_1 _25272_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net956),
    .S(_06533_),
    .X(_02240_));
 sg13g2_mux2_1 _25273_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net955),
    .S(_06533_),
    .X(_02241_));
 sg13g2_and2_1 _25274_ (.A(net626),
    .B(_06416_),
    .X(_06534_));
 sg13g2_buf_1 _25275_ (.A(_06534_),
    .X(_06535_));
 sg13g2_mux2_1 _25276_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(net958),
    .S(_06535_),
    .X(_02242_));
 sg13g2_mux2_1 _25277_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net957),
    .S(_06535_),
    .X(_02243_));
 sg13g2_mux2_1 _25278_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net956),
    .S(_06535_),
    .X(_02244_));
 sg13g2_mux2_1 _25279_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net955),
    .S(_06535_),
    .X(_02245_));
 sg13g2_and2_1 _25280_ (.A(_08956_),
    .B(_06420_),
    .X(_06536_));
 sg13g2_buf_1 _25281_ (.A(_06536_),
    .X(_06537_));
 sg13g2_mux2_1 _25282_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(_06474_),
    .S(_06537_),
    .X(_02246_));
 sg13g2_mux2_1 _25283_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(_06477_),
    .S(_06537_),
    .X(_02247_));
 sg13g2_mux2_1 _25284_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(_06478_),
    .S(_06537_),
    .X(_02248_));
 sg13g2_mux2_1 _25285_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(_06479_),
    .S(_06537_),
    .X(_02249_));
 sg13g2_mux2_1 _25286_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net957),
    .S(_06531_),
    .X(_02250_));
 sg13g2_and2_1 _25287_ (.A(net626),
    .B(_06423_),
    .X(_06538_));
 sg13g2_buf_1 _25288_ (.A(_06538_),
    .X(_06539_));
 sg13g2_mux2_1 _25289_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(_06474_),
    .S(_06539_),
    .X(_02251_));
 sg13g2_mux2_1 _25290_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(_06477_),
    .S(_06539_),
    .X(_02252_));
 sg13g2_mux2_1 _25291_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(_06478_),
    .S(_06539_),
    .X(_02253_));
 sg13g2_mux2_1 _25292_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(_06479_),
    .S(_06539_),
    .X(_02254_));
 sg13g2_and2_1 _25293_ (.A(net626),
    .B(_06427_),
    .X(_06540_));
 sg13g2_buf_2 _25294_ (.A(_06540_),
    .X(_06541_));
 sg13g2_mux2_1 _25295_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1021),
    .S(_06541_),
    .X(_02255_));
 sg13g2_mux2_1 _25296_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net1020),
    .S(_06541_),
    .X(_02256_));
 sg13g2_mux2_1 _25297_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net1023),
    .S(_06541_),
    .X(_02257_));
 sg13g2_mux2_1 _25298_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net1022),
    .S(_06541_),
    .X(_02258_));
 sg13g2_and2_1 _25299_ (.A(net626),
    .B(_06433_),
    .X(_06542_));
 sg13g2_buf_1 _25300_ (.A(_06542_),
    .X(_06543_));
 sg13g2_mux2_1 _25301_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1021),
    .S(_06543_),
    .X(_02259_));
 sg13g2_mux2_1 _25302_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net1020),
    .S(_06543_),
    .X(_02260_));
 sg13g2_mux2_1 _25303_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net1023),
    .S(_06531_),
    .X(_02261_));
 sg13g2_mux2_1 _25304_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12209_),
    .S(_06543_),
    .X(_02262_));
 sg13g2_mux2_1 _25305_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net1022),
    .S(_06543_),
    .X(_02263_));
 sg13g2_mux2_1 _25306_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12216_),
    .S(_06531_),
    .X(_02264_));
 sg13g2_and2_1 _25307_ (.A(net626),
    .B(_06436_),
    .X(_06544_));
 sg13g2_buf_1 _25308_ (.A(_06544_),
    .X(_06545_));
 sg13g2_mux2_1 _25309_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12220_),
    .S(_06545_),
    .X(_02265_));
 sg13g2_mux2_1 _25310_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12227_),
    .S(_06545_),
    .X(_02266_));
 sg13g2_mux2_1 _25311_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12209_),
    .S(_06545_),
    .X(_02267_));
 sg13g2_mux2_1 _25312_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12216_),
    .S(_06545_),
    .X(_02268_));
 sg13g2_mux2_1 _25313_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12220_),
    .S(_06533_),
    .X(_02269_));
 sg13g2_mux2_1 _25314_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12227_),
    .S(_06533_),
    .X(_02270_));
 sg13g2_mux2_1 _25315_ (.A0(net987),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(_06431_),
    .X(_02274_));
 sg13g2_buf_1 _25316_ (.A(_06429_),
    .X(_06546_));
 sg13g2_nand2_1 _25317_ (.Y(_06547_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net405));
 sg13g2_o21ai_1 _25318_ (.B1(_06547_),
    .Y(_02275_),
    .A1(net392),
    .A2(net404));
 sg13g2_nand2_1 _25319_ (.Y(_06548_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net405));
 sg13g2_o21ai_1 _25320_ (.B1(_06548_),
    .Y(_02276_),
    .A1(net393),
    .A2(net404));
 sg13g2_nand2_1 _25321_ (.Y(_06549_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net405));
 sg13g2_o21ai_1 _25322_ (.B1(_06549_),
    .Y(_02277_),
    .A1(net394),
    .A2(_06546_));
 sg13g2_nand2_1 _25323_ (.Y(_06550_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net405));
 sg13g2_o21ai_1 _25324_ (.B1(_06550_),
    .Y(_02278_),
    .A1(net344),
    .A2(net404));
 sg13g2_nand2_1 _25325_ (.Y(_06551_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(net405));
 sg13g2_o21ai_1 _25326_ (.B1(_06551_),
    .Y(_02279_),
    .A1(net395),
    .A2(net404));
 sg13g2_nand2_1 _25327_ (.Y(_06552_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net405));
 sg13g2_o21ai_1 _25328_ (.B1(_06552_),
    .Y(_02280_),
    .A1(net391),
    .A2(net404));
 sg13g2_buf_1 _25329_ (.A(_06429_),
    .X(_06553_));
 sg13g2_nand2_1 _25330_ (.Y(_06554_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net403));
 sg13g2_o21ai_1 _25331_ (.B1(_06554_),
    .Y(_02281_),
    .A1(net396),
    .A2(net404));
 sg13g2_nand2_1 _25332_ (.Y(_06555_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net403));
 sg13g2_o21ai_1 _25333_ (.B1(_06555_),
    .Y(_02282_),
    .A1(net436),
    .A2(net404));
 sg13g2_nand2_1 _25334_ (.Y(_06556_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net403));
 sg13g2_o21ai_1 _25335_ (.B1(_06556_),
    .Y(_02283_),
    .A1(net487),
    .A2(net404));
 sg13g2_mux2_1 _25336_ (.A0(net986),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net405),
    .X(_02284_));
 sg13g2_nand2_1 _25337_ (.Y(_06557_),
    .A(\cpu.icache.r_tag[0][7] ),
    .B(net403));
 sg13g2_o21ai_1 _25338_ (.B1(_06557_),
    .Y(_02285_),
    .A1(net988),
    .A2(net406));
 sg13g2_nand2_1 _25339_ (.Y(_06558_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(net403));
 sg13g2_o21ai_1 _25340_ (.B1(_06558_),
    .Y(_02286_),
    .A1(net922),
    .A2(net406));
 sg13g2_nand2_1 _25341_ (.Y(_06559_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(_06553_));
 sg13g2_o21ai_1 _25342_ (.B1(_06559_),
    .Y(_02287_),
    .A1(net1080),
    .A2(net406));
 sg13g2_mux2_1 _25343_ (.A0(net985),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(_06431_),
    .X(_02288_));
 sg13g2_nand2_1 _25344_ (.Y(_06560_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net403));
 sg13g2_o21ai_1 _25345_ (.B1(_06560_),
    .Y(_02289_),
    .A1(net1079),
    .A2(net406));
 sg13g2_nand2_1 _25346_ (.Y(_06561_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(_06553_));
 sg13g2_o21ai_1 _25347_ (.B1(_06561_),
    .Y(_02290_),
    .A1(net488),
    .A2(net406));
 sg13g2_nand2_1 _25348_ (.Y(_06562_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(net403));
 sg13g2_o21ai_1 _25349_ (.B1(_06562_),
    .Y(_02291_),
    .A1(net437),
    .A2(net406));
 sg13g2_nand2_1 _25350_ (.Y(_06563_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net403));
 sg13g2_o21ai_1 _25351_ (.B1(_06563_),
    .Y(_02292_),
    .A1(net486),
    .A2(net406));
 sg13g2_nor3_1 _25352_ (.A(_06399_),
    .B(_06407_),
    .C(_06409_),
    .Y(_06564_));
 sg13g2_buf_1 _25353_ (.A(_06564_),
    .X(_06565_));
 sg13g2_nand2_1 _25354_ (.Y(_06566_),
    .A(net524),
    .B(_06565_));
 sg13g2_buf_2 _25355_ (.A(_06566_),
    .X(_06567_));
 sg13g2_buf_1 _25356_ (.A(_06567_),
    .X(_06568_));
 sg13g2_mux2_1 _25357_ (.A0(net987),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net358),
    .X(_02293_));
 sg13g2_buf_1 _25358_ (.A(_06567_),
    .X(_06569_));
 sg13g2_nand2_1 _25359_ (.Y(_06570_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(_06568_));
 sg13g2_o21ai_1 _25360_ (.B1(_06570_),
    .Y(_02294_),
    .A1(net392),
    .A2(net357));
 sg13g2_buf_1 _25361_ (.A(_06567_),
    .X(_06571_));
 sg13g2_nand2_1 _25362_ (.Y(_06572_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net356));
 sg13g2_o21ai_1 _25363_ (.B1(_06572_),
    .Y(_02295_),
    .A1(net393),
    .A2(net357));
 sg13g2_nand2_1 _25364_ (.Y(_06573_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net356));
 sg13g2_o21ai_1 _25365_ (.B1(_06573_),
    .Y(_02296_),
    .A1(net394),
    .A2(net357));
 sg13g2_nand2_1 _25366_ (.Y(_06574_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net356));
 sg13g2_o21ai_1 _25367_ (.B1(_06574_),
    .Y(_02297_),
    .A1(net344),
    .A2(net357));
 sg13g2_nand2_1 _25368_ (.Y(_06575_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net356));
 sg13g2_o21ai_1 _25369_ (.B1(_06575_),
    .Y(_02298_),
    .A1(net395),
    .A2(net357));
 sg13g2_nand2_1 _25370_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net356));
 sg13g2_o21ai_1 _25371_ (.B1(_06576_),
    .Y(_02299_),
    .A1(net391),
    .A2(net357));
 sg13g2_nand2_1 _25372_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net356));
 sg13g2_o21ai_1 _25373_ (.B1(_06577_),
    .Y(_02300_),
    .A1(net396),
    .A2(net357));
 sg13g2_nand2_1 _25374_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25375_ (.B1(_06578_),
    .Y(_02301_),
    .A1(net436),
    .A2(_06569_));
 sg13g2_nand2_1 _25376_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25377_ (.B1(_06579_),
    .Y(_02302_),
    .A1(net487),
    .A2(_06569_));
 sg13g2_mux2_1 _25378_ (.A0(net986),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net358),
    .X(_02303_));
 sg13g2_nand2_1 _25379_ (.Y(_06580_),
    .A(\cpu.icache.r_tag[1][7] ),
    .B(net356));
 sg13g2_o21ai_1 _25380_ (.B1(_06580_),
    .Y(_02304_),
    .A1(net988),
    .A2(net357));
 sg13g2_nand2_1 _25381_ (.Y(_06581_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net356));
 sg13g2_o21ai_1 _25382_ (.B1(_06581_),
    .Y(_02305_),
    .A1(net922),
    .A2(net358));
 sg13g2_nand2_1 _25383_ (.Y(_06582_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25384_ (.B1(_06582_),
    .Y(_02306_),
    .A1(net1080),
    .A2(net358));
 sg13g2_mux2_1 _25385_ (.A0(net985),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net358),
    .X(_02307_));
 sg13g2_nand2_1 _25386_ (.Y(_06583_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25387_ (.B1(_06583_),
    .Y(_02308_),
    .A1(net1079),
    .A2(net358));
 sg13g2_nand2_1 _25388_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25389_ (.B1(_06584_),
    .Y(_02309_),
    .A1(net488),
    .A2(net358));
 sg13g2_nand2_1 _25390_ (.Y(_06585_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25391_ (.B1(_06585_),
    .Y(_02310_),
    .A1(net437),
    .A2(net358));
 sg13g2_nand2_1 _25392_ (.Y(_06586_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25393_ (.B1(_06586_),
    .Y(_02311_),
    .A1(net486),
    .A2(_06568_));
 sg13g2_nand2_1 _25394_ (.Y(_06587_),
    .A(net463),
    .B(_06565_));
 sg13g2_buf_2 _25395_ (.A(_06587_),
    .X(_06588_));
 sg13g2_buf_1 _25396_ (.A(_06588_),
    .X(_06589_));
 sg13g2_mux2_1 _25397_ (.A0(net987),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net278),
    .X(_02312_));
 sg13g2_buf_1 _25398_ (.A(_06588_),
    .X(_06590_));
 sg13g2_nand2_1 _25399_ (.Y(_06591_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net278));
 sg13g2_o21ai_1 _25400_ (.B1(_06591_),
    .Y(_02313_),
    .A1(net392),
    .A2(net277));
 sg13g2_buf_1 _25401_ (.A(_06588_),
    .X(_06592_));
 sg13g2_nand2_1 _25402_ (.Y(_06593_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net276));
 sg13g2_o21ai_1 _25403_ (.B1(_06593_),
    .Y(_02314_),
    .A1(net393),
    .A2(net277));
 sg13g2_nand2_1 _25404_ (.Y(_06594_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net276));
 sg13g2_o21ai_1 _25405_ (.B1(_06594_),
    .Y(_02315_),
    .A1(net394),
    .A2(net277));
 sg13g2_nand2_1 _25406_ (.Y(_06595_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net276));
 sg13g2_o21ai_1 _25407_ (.B1(_06595_),
    .Y(_02316_),
    .A1(net344),
    .A2(net277));
 sg13g2_nand2_1 _25408_ (.Y(_06596_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net276));
 sg13g2_o21ai_1 _25409_ (.B1(_06596_),
    .Y(_02317_),
    .A1(net395),
    .A2(net277));
 sg13g2_nand2_1 _25410_ (.Y(_06597_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net276));
 sg13g2_o21ai_1 _25411_ (.B1(_06597_),
    .Y(_02318_),
    .A1(net391),
    .A2(net277));
 sg13g2_nand2_1 _25412_ (.Y(_06598_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net276));
 sg13g2_o21ai_1 _25413_ (.B1(_06598_),
    .Y(_02319_),
    .A1(net396),
    .A2(net277));
 sg13g2_nand2_1 _25414_ (.Y(_06599_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(_06592_));
 sg13g2_o21ai_1 _25415_ (.B1(_06599_),
    .Y(_02320_),
    .A1(_08670_),
    .A2(_06590_));
 sg13g2_nand2_1 _25416_ (.Y(_06600_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net276));
 sg13g2_o21ai_1 _25417_ (.B1(_06600_),
    .Y(_02321_),
    .A1(net487),
    .A2(net277));
 sg13g2_mux2_1 _25418_ (.A0(net986),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net278),
    .X(_02322_));
 sg13g2_nand2_1 _25419_ (.Y(_06601_),
    .A(\cpu.icache.r_tag[2][7] ),
    .B(net276));
 sg13g2_o21ai_1 _25420_ (.B1(_06601_),
    .Y(_02323_),
    .A1(net988),
    .A2(_06590_));
 sg13g2_nand2_1 _25421_ (.Y(_06602_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(_06592_));
 sg13g2_o21ai_1 _25422_ (.B1(_06602_),
    .Y(_02324_),
    .A1(net922),
    .A2(net278));
 sg13g2_nand2_1 _25423_ (.Y(_06603_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25424_ (.B1(_06603_),
    .Y(_02325_),
    .A1(_08825_),
    .A2(_06589_));
 sg13g2_mux2_1 _25425_ (.A0(net985),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net278),
    .X(_02326_));
 sg13g2_nand2_1 _25426_ (.Y(_06604_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25427_ (.B1(_06604_),
    .Y(_02327_),
    .A1(net1079),
    .A2(_06589_));
 sg13g2_nand2_1 _25428_ (.Y(_06605_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25429_ (.B1(_06605_),
    .Y(_02328_),
    .A1(net488),
    .A2(net278));
 sg13g2_nand2_1 _25430_ (.Y(_06606_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25431_ (.B1(_06606_),
    .Y(_02329_),
    .A1(net437),
    .A2(net278));
 sg13g2_nand2_1 _25432_ (.Y(_06607_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25433_ (.B1(_06607_),
    .Y(_02330_),
    .A1(_08691_),
    .A2(net278));
 sg13g2_mux2_1 _25434_ (.A0(net987),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net359),
    .X(_02331_));
 sg13g2_buf_1 _25435_ (.A(_06493_),
    .X(_06608_));
 sg13g2_nand2_1 _25436_ (.Y(_06609_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net359));
 sg13g2_o21ai_1 _25437_ (.B1(_06609_),
    .Y(_02332_),
    .A1(_08784_),
    .A2(_06608_));
 sg13g2_nand2_1 _25438_ (.Y(_06610_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net359));
 sg13g2_o21ai_1 _25439_ (.B1(_06610_),
    .Y(_02333_),
    .A1(net393),
    .A2(net355));
 sg13g2_nand2_1 _25440_ (.Y(_06611_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net359));
 sg13g2_o21ai_1 _25441_ (.B1(_06611_),
    .Y(_02334_),
    .A1(net394),
    .A2(net355));
 sg13g2_nand2_1 _25442_ (.Y(_06612_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net359));
 sg13g2_o21ai_1 _25443_ (.B1(_06612_),
    .Y(_02335_),
    .A1(net344),
    .A2(net355));
 sg13g2_nand2_1 _25444_ (.Y(_06613_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net359));
 sg13g2_o21ai_1 _25445_ (.B1(_06613_),
    .Y(_02336_),
    .A1(net395),
    .A2(net355));
 sg13g2_nand2_1 _25446_ (.Y(_06614_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net359));
 sg13g2_o21ai_1 _25447_ (.B1(_06614_),
    .Y(_02337_),
    .A1(net391),
    .A2(net355));
 sg13g2_buf_1 _25448_ (.A(_06493_),
    .X(_06615_));
 sg13g2_nand2_1 _25449_ (.Y(_06616_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net354));
 sg13g2_o21ai_1 _25450_ (.B1(_06616_),
    .Y(_02338_),
    .A1(net396),
    .A2(net355));
 sg13g2_nand2_1 _25451_ (.Y(_06617_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net354));
 sg13g2_o21ai_1 _25452_ (.B1(_06617_),
    .Y(_02339_),
    .A1(net436),
    .A2(net355));
 sg13g2_nand2_1 _25453_ (.Y(_06618_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net354));
 sg13g2_o21ai_1 _25454_ (.B1(_06618_),
    .Y(_02340_),
    .A1(net487),
    .A2(net355));
 sg13g2_mux2_1 _25455_ (.A0(net986),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net359),
    .X(_02341_));
 sg13g2_nand2_1 _25456_ (.Y(_06619_),
    .A(\cpu.icache.r_tag[3][7] ),
    .B(net354));
 sg13g2_o21ai_1 _25457_ (.B1(_06619_),
    .Y(_02342_),
    .A1(net988),
    .A2(net360));
 sg13g2_nand2_1 _25458_ (.Y(_06620_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net354));
 sg13g2_o21ai_1 _25459_ (.B1(_06620_),
    .Y(_02343_),
    .A1(net922),
    .A2(net360));
 sg13g2_nand2_1 _25460_ (.Y(_06621_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(net354));
 sg13g2_o21ai_1 _25461_ (.B1(_06621_),
    .Y(_02344_),
    .A1(net1080),
    .A2(net360));
 sg13g2_mux2_1 _25462_ (.A0(net985),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(_06495_),
    .X(_02345_));
 sg13g2_nand2_1 _25463_ (.Y(_06622_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net354));
 sg13g2_o21ai_1 _25464_ (.B1(_06622_),
    .Y(_02346_),
    .A1(net1079),
    .A2(net360));
 sg13g2_nand2_1 _25465_ (.Y(_06623_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(_06615_));
 sg13g2_o21ai_1 _25466_ (.B1(_06623_),
    .Y(_02347_),
    .A1(net488),
    .A2(net360));
 sg13g2_nand2_1 _25467_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(_06615_));
 sg13g2_o21ai_1 _25468_ (.B1(_06624_),
    .Y(_02348_),
    .A1(net437),
    .A2(net360));
 sg13g2_nand2_1 _25469_ (.Y(_06625_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net354));
 sg13g2_o21ai_1 _25470_ (.B1(_06625_),
    .Y(_02349_),
    .A1(net486),
    .A2(_06494_));
 sg13g2_nand2_1 _25471_ (.Y(_06626_),
    .A(net522),
    .B(_06565_));
 sg13g2_buf_2 _25472_ (.A(_06626_),
    .X(_06627_));
 sg13g2_buf_1 _25473_ (.A(_06627_),
    .X(_06628_));
 sg13g2_mux2_1 _25474_ (.A0(net987),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net353),
    .X(_02350_));
 sg13g2_buf_1 _25475_ (.A(_06627_),
    .X(_06629_));
 sg13g2_nand2_1 _25476_ (.Y(_06630_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net353));
 sg13g2_o21ai_1 _25477_ (.B1(_06630_),
    .Y(_02351_),
    .A1(net392),
    .A2(net352));
 sg13g2_buf_1 _25478_ (.A(_06627_),
    .X(_06631_));
 sg13g2_nand2_1 _25479_ (.Y(_06632_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net351));
 sg13g2_o21ai_1 _25480_ (.B1(_06632_),
    .Y(_02352_),
    .A1(net393),
    .A2(net352));
 sg13g2_nand2_1 _25481_ (.Y(_06633_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net351));
 sg13g2_o21ai_1 _25482_ (.B1(_06633_),
    .Y(_02353_),
    .A1(net394),
    .A2(net352));
 sg13g2_nand2_1 _25483_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net351));
 sg13g2_o21ai_1 _25484_ (.B1(_06634_),
    .Y(_02354_),
    .A1(net344),
    .A2(net352));
 sg13g2_nand2_1 _25485_ (.Y(_06635_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net351));
 sg13g2_o21ai_1 _25486_ (.B1(_06635_),
    .Y(_02355_),
    .A1(net395),
    .A2(net352));
 sg13g2_nand2_1 _25487_ (.Y(_06636_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net351));
 sg13g2_o21ai_1 _25488_ (.B1(_06636_),
    .Y(_02356_),
    .A1(net391),
    .A2(net352));
 sg13g2_nand2_1 _25489_ (.Y(_06637_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net351));
 sg13g2_o21ai_1 _25490_ (.B1(_06637_),
    .Y(_02357_),
    .A1(net396),
    .A2(net352));
 sg13g2_nand2_1 _25491_ (.Y(_06638_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(_06631_));
 sg13g2_o21ai_1 _25492_ (.B1(_06638_),
    .Y(_02358_),
    .A1(net436),
    .A2(_06629_));
 sg13g2_nand2_1 _25493_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net351));
 sg13g2_o21ai_1 _25494_ (.B1(_06639_),
    .Y(_02359_),
    .A1(_08615_),
    .A2(net352));
 sg13g2_mux2_1 _25495_ (.A0(net986),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net353),
    .X(_02360_));
 sg13g2_nand2_1 _25496_ (.Y(_06640_),
    .A(\cpu.icache.r_tag[4][7] ),
    .B(_06631_));
 sg13g2_o21ai_1 _25497_ (.B1(_06640_),
    .Y(_02361_),
    .A1(net988),
    .A2(_06629_));
 sg13g2_nand2_1 _25498_ (.Y(_06641_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(net351));
 sg13g2_o21ai_1 _25499_ (.B1(_06641_),
    .Y(_02362_),
    .A1(net922),
    .A2(net353));
 sg13g2_nand2_1 _25500_ (.Y(_06642_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(_06627_));
 sg13g2_o21ai_1 _25501_ (.B1(_06642_),
    .Y(_02363_),
    .A1(net1080),
    .A2(_06628_));
 sg13g2_mux2_1 _25502_ (.A0(net985),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net353),
    .X(_02364_));
 sg13g2_nand2_1 _25503_ (.Y(_06643_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(_06627_));
 sg13g2_o21ai_1 _25504_ (.B1(_06643_),
    .Y(_02365_),
    .A1(net1079),
    .A2(net353));
 sg13g2_nand2_1 _25505_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06627_));
 sg13g2_o21ai_1 _25506_ (.B1(_06644_),
    .Y(_02366_),
    .A1(net488),
    .A2(net353));
 sg13g2_nand2_1 _25507_ (.Y(_06645_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06627_));
 sg13g2_o21ai_1 _25508_ (.B1(_06645_),
    .Y(_02367_),
    .A1(net437),
    .A2(_06628_));
 sg13g2_nand2_1 _25509_ (.Y(_06646_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06627_));
 sg13g2_o21ai_1 _25510_ (.B1(_06646_),
    .Y(_02368_),
    .A1(net486),
    .A2(net353));
 sg13g2_nand2_1 _25511_ (.Y(_06647_),
    .A(net625),
    .B(_06565_));
 sg13g2_buf_2 _25512_ (.A(_06647_),
    .X(_06648_));
 sg13g2_buf_1 _25513_ (.A(_06648_),
    .X(_06649_));
 sg13g2_mux2_1 _25514_ (.A0(net987),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net402),
    .X(_02369_));
 sg13g2_buf_1 _25515_ (.A(_06648_),
    .X(_06650_));
 sg13g2_nand2_1 _25516_ (.Y(_06651_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net402));
 sg13g2_o21ai_1 _25517_ (.B1(_06651_),
    .Y(_02370_),
    .A1(net392),
    .A2(net401));
 sg13g2_buf_1 _25518_ (.A(_06648_),
    .X(_06652_));
 sg13g2_nand2_1 _25519_ (.Y(_06653_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net400));
 sg13g2_o21ai_1 _25520_ (.B1(_06653_),
    .Y(_02371_),
    .A1(net393),
    .A2(net401));
 sg13g2_nand2_1 _25521_ (.Y(_06654_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net400));
 sg13g2_o21ai_1 _25522_ (.B1(_06654_),
    .Y(_02372_),
    .A1(net394),
    .A2(net401));
 sg13g2_nand2_1 _25523_ (.Y(_06655_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net400));
 sg13g2_o21ai_1 _25524_ (.B1(_06655_),
    .Y(_02373_),
    .A1(net344),
    .A2(net401));
 sg13g2_nand2_1 _25525_ (.Y(_06656_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net400));
 sg13g2_o21ai_1 _25526_ (.B1(_06656_),
    .Y(_02374_),
    .A1(net395),
    .A2(net401));
 sg13g2_nand2_1 _25527_ (.Y(_06657_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net400));
 sg13g2_o21ai_1 _25528_ (.B1(_06657_),
    .Y(_02375_),
    .A1(net391),
    .A2(net401));
 sg13g2_nand2_1 _25529_ (.Y(_06658_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(_06652_));
 sg13g2_o21ai_1 _25530_ (.B1(_06658_),
    .Y(_02376_),
    .A1(net396),
    .A2(_06650_));
 sg13g2_nand2_1 _25531_ (.Y(_06659_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(_06652_));
 sg13g2_o21ai_1 _25532_ (.B1(_06659_),
    .Y(_02377_),
    .A1(net436),
    .A2(_06650_));
 sg13g2_nand2_1 _25533_ (.Y(_06660_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net400));
 sg13g2_o21ai_1 _25534_ (.B1(_06660_),
    .Y(_02378_),
    .A1(net487),
    .A2(net401));
 sg13g2_mux2_1 _25535_ (.A0(net986),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(net402),
    .X(_02379_));
 sg13g2_nand2_1 _25536_ (.Y(_06661_),
    .A(\cpu.icache.r_tag[5][7] ),
    .B(net400));
 sg13g2_o21ai_1 _25537_ (.B1(_06661_),
    .Y(_02380_),
    .A1(net988),
    .A2(net401));
 sg13g2_nand2_1 _25538_ (.Y(_06662_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net400));
 sg13g2_o21ai_1 _25539_ (.B1(_06662_),
    .Y(_02381_),
    .A1(net922),
    .A2(net402));
 sg13g2_nand2_1 _25540_ (.Y(_06663_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(_06648_));
 sg13g2_o21ai_1 _25541_ (.B1(_06663_),
    .Y(_02382_),
    .A1(net1080),
    .A2(net402));
 sg13g2_mux2_1 _25542_ (.A0(net985),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net402),
    .X(_02383_));
 sg13g2_nand2_1 _25543_ (.Y(_06664_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(_06648_));
 sg13g2_o21ai_1 _25544_ (.B1(_06664_),
    .Y(_02384_),
    .A1(_08883_),
    .A2(net402));
 sg13g2_nand2_1 _25545_ (.Y(_06665_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06648_));
 sg13g2_o21ai_1 _25546_ (.B1(_06665_),
    .Y(_02385_),
    .A1(_08556_),
    .A2(_06649_));
 sg13g2_nand2_1 _25547_ (.Y(_06666_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06648_));
 sg13g2_o21ai_1 _25548_ (.B1(_06666_),
    .Y(_02386_),
    .A1(_08587_),
    .A2(net402));
 sg13g2_nand2_1 _25549_ (.Y(_06667_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06648_));
 sg13g2_o21ai_1 _25550_ (.B1(_06667_),
    .Y(_02387_),
    .A1(net486),
    .A2(_06649_));
 sg13g2_nand2_1 _25551_ (.Y(_06668_),
    .A(net523),
    .B(_06565_));
 sg13g2_buf_2 _25552_ (.A(_06668_),
    .X(_06669_));
 sg13g2_buf_1 _25553_ (.A(_06669_),
    .X(_06670_));
 sg13g2_mux2_1 _25554_ (.A0(_04581_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net350),
    .X(_02388_));
 sg13g2_buf_1 _25555_ (.A(_06669_),
    .X(_06671_));
 sg13g2_nand2_1 _25556_ (.Y(_06672_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net350));
 sg13g2_o21ai_1 _25557_ (.B1(_06672_),
    .Y(_02389_),
    .A1(net392),
    .A2(_06671_));
 sg13g2_buf_1 _25558_ (.A(_06669_),
    .X(_06673_));
 sg13g2_nand2_1 _25559_ (.Y(_06674_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net348));
 sg13g2_o21ai_1 _25560_ (.B1(_06674_),
    .Y(_02390_),
    .A1(net393),
    .A2(net349));
 sg13g2_nand2_1 _25561_ (.Y(_06675_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net348));
 sg13g2_o21ai_1 _25562_ (.B1(_06675_),
    .Y(_02391_),
    .A1(net394),
    .A2(net349));
 sg13g2_nand2_1 _25563_ (.Y(_06676_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net348));
 sg13g2_o21ai_1 _25564_ (.B1(_06676_),
    .Y(_02392_),
    .A1(_09046_),
    .A2(net349));
 sg13g2_nand2_1 _25565_ (.Y(_06677_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net348));
 sg13g2_o21ai_1 _25566_ (.B1(_06677_),
    .Y(_02393_),
    .A1(net395),
    .A2(net349));
 sg13g2_nand2_1 _25567_ (.Y(_06678_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net348));
 sg13g2_o21ai_1 _25568_ (.B1(_06678_),
    .Y(_02394_),
    .A1(net391),
    .A2(net349));
 sg13g2_nand2_1 _25569_ (.Y(_06679_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net348));
 sg13g2_o21ai_1 _25570_ (.B1(_06679_),
    .Y(_02395_),
    .A1(net396),
    .A2(net349));
 sg13g2_nand2_1 _25571_ (.Y(_06680_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net348));
 sg13g2_o21ai_1 _25572_ (.B1(_06680_),
    .Y(_02396_),
    .A1(net436),
    .A2(net349));
 sg13g2_nand2_1 _25573_ (.Y(_06681_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net348));
 sg13g2_o21ai_1 _25574_ (.B1(_06681_),
    .Y(_02397_),
    .A1(net487),
    .A2(net349));
 sg13g2_mux2_1 _25575_ (.A0(_04614_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net350),
    .X(_02398_));
 sg13g2_nand2_1 _25576_ (.Y(_06682_),
    .A(\cpu.icache.r_tag[6][7] ),
    .B(_06673_));
 sg13g2_o21ai_1 _25577_ (.B1(_06682_),
    .Y(_02399_),
    .A1(_04229_),
    .A2(_06671_));
 sg13g2_nand2_1 _25578_ (.Y(_06683_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(_06673_));
 sg13g2_o21ai_1 _25579_ (.B1(_06683_),
    .Y(_02400_),
    .A1(net922),
    .A2(net350));
 sg13g2_nand2_1 _25580_ (.Y(_06684_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(_06669_));
 sg13g2_o21ai_1 _25581_ (.B1(_06684_),
    .Y(_02401_),
    .A1(net1080),
    .A2(_06670_));
 sg13g2_mux2_1 _25582_ (.A0(_04733_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net350),
    .X(_02402_));
 sg13g2_nand2_1 _25583_ (.Y(_06685_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06669_));
 sg13g2_o21ai_1 _25584_ (.B1(_06685_),
    .Y(_02403_),
    .A1(net1079),
    .A2(net350));
 sg13g2_nand2_1 _25585_ (.Y(_06686_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06669_));
 sg13g2_o21ai_1 _25586_ (.B1(_06686_),
    .Y(_02404_),
    .A1(net488),
    .A2(net350));
 sg13g2_nand2_1 _25587_ (.Y(_06687_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06669_));
 sg13g2_o21ai_1 _25588_ (.B1(_06687_),
    .Y(_02405_),
    .A1(net437),
    .A2(net350));
 sg13g2_nand2_1 _25589_ (.Y(_06688_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06669_));
 sg13g2_o21ai_1 _25590_ (.B1(_06688_),
    .Y(_02406_),
    .A1(net486),
    .A2(_06670_));
 sg13g2_nand2_1 _25591_ (.Y(_06689_),
    .A(net626),
    .B(_06565_));
 sg13g2_buf_2 _25592_ (.A(_06689_),
    .X(_06690_));
 sg13g2_buf_1 _25593_ (.A(_06690_),
    .X(_06691_));
 sg13g2_mux2_1 _25594_ (.A0(_04581_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net399),
    .X(_02407_));
 sg13g2_buf_1 _25595_ (.A(_06690_),
    .X(_06692_));
 sg13g2_nand2_1 _25596_ (.Y(_06693_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net399));
 sg13g2_o21ai_1 _25597_ (.B1(_06693_),
    .Y(_02408_),
    .A1(net392),
    .A2(net398));
 sg13g2_buf_1 _25598_ (.A(_06690_),
    .X(_06694_));
 sg13g2_nand2_1 _25599_ (.Y(_06695_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net397));
 sg13g2_o21ai_1 _25600_ (.B1(_06695_),
    .Y(_02409_),
    .A1(net393),
    .A2(net398));
 sg13g2_nand2_1 _25601_ (.Y(_06696_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net397));
 sg13g2_o21ai_1 _25602_ (.B1(_06696_),
    .Y(_02410_),
    .A1(_08738_),
    .A2(net398));
 sg13g2_nand2_1 _25603_ (.Y(_06697_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net397));
 sg13g2_o21ai_1 _25604_ (.B1(_06697_),
    .Y(_02411_),
    .A1(net344),
    .A2(net398));
 sg13g2_nand2_1 _25605_ (.Y(_06698_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net397));
 sg13g2_o21ai_1 _25606_ (.B1(_06698_),
    .Y(_02412_),
    .A1(net395),
    .A2(net398));
 sg13g2_nand2_1 _25607_ (.Y(_06699_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net397));
 sg13g2_o21ai_1 _25608_ (.B1(_06699_),
    .Y(_02413_),
    .A1(net391),
    .A2(net398));
 sg13g2_nand2_1 _25609_ (.Y(_06700_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(_06694_));
 sg13g2_o21ai_1 _25610_ (.B1(_06700_),
    .Y(_02414_),
    .A1(_08487_),
    .A2(_06692_));
 sg13g2_nand2_1 _25611_ (.Y(_06701_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(_06694_));
 sg13g2_o21ai_1 _25612_ (.B1(_06701_),
    .Y(_02415_),
    .A1(net436),
    .A2(_06692_));
 sg13g2_nand2_1 _25613_ (.Y(_06702_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net397));
 sg13g2_o21ai_1 _25614_ (.B1(_06702_),
    .Y(_02416_),
    .A1(net487),
    .A2(net398));
 sg13g2_mux2_1 _25615_ (.A0(_04614_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net399),
    .X(_02417_));
 sg13g2_nand2_1 _25616_ (.Y(_06703_),
    .A(\cpu.icache.r_tag[7][7] ),
    .B(net397));
 sg13g2_o21ai_1 _25617_ (.B1(_06703_),
    .Y(_02418_),
    .A1(_04229_),
    .A2(net398));
 sg13g2_nand2_1 _25618_ (.Y(_06704_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net397));
 sg13g2_o21ai_1 _25619_ (.B1(_06704_),
    .Y(_02419_),
    .A1(_08852_),
    .A2(net399));
 sg13g2_nand2_1 _25620_ (.Y(_06705_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(_06690_));
 sg13g2_o21ai_1 _25621_ (.B1(_06705_),
    .Y(_02420_),
    .A1(net1080),
    .A2(_06691_));
 sg13g2_mux2_1 _25622_ (.A0(_04733_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net399),
    .X(_02421_));
 sg13g2_nand2_1 _25623_ (.Y(_06706_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06690_));
 sg13g2_o21ai_1 _25624_ (.B1(_06706_),
    .Y(_02422_),
    .A1(net1079),
    .A2(net399));
 sg13g2_nand2_1 _25625_ (.Y(_06707_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06690_));
 sg13g2_o21ai_1 _25626_ (.B1(_06707_),
    .Y(_02423_),
    .A1(net488),
    .A2(_06691_));
 sg13g2_nand2_1 _25627_ (.Y(_06708_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06690_));
 sg13g2_o21ai_1 _25628_ (.B1(_06708_),
    .Y(_02424_),
    .A1(net437),
    .A2(net399));
 sg13g2_nand2_1 _25629_ (.Y(_06709_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06690_));
 sg13g2_o21ai_1 _25630_ (.B1(_06709_),
    .Y(_02425_),
    .A1(net486),
    .A2(net399));
 sg13g2_and2_1 _25631_ (.A(net193),
    .B(net448),
    .X(_06710_));
 sg13g2_buf_2 _25632_ (.A(_06710_),
    .X(_06711_));
 sg13g2_buf_1 _25633_ (.A(_06711_),
    .X(_06712_));
 sg13g2_mux2_1 _25634_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(net869),
    .S(net97),
    .X(_02435_));
 sg13g2_mux2_1 _25635_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(_10215_),
    .S(net97),
    .X(_02436_));
 sg13g2_mux2_1 _25636_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(_10222_),
    .S(net97),
    .X(_02437_));
 sg13g2_mux2_1 _25637_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(_10227_),
    .S(net97),
    .X(_02438_));
 sg13g2_mux2_1 _25638_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(_10229_),
    .S(net97),
    .X(_02439_));
 sg13g2_mux2_1 _25639_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(_10239_),
    .S(_06712_),
    .X(_02440_));
 sg13g2_mux2_1 _25640_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(_10244_),
    .S(_06712_),
    .X(_02441_));
 sg13g2_nor3_1 _25641_ (.A(_09292_),
    .B(_10030_),
    .C(_04870_),
    .Y(_06713_));
 sg13g2_buf_2 _25642_ (.A(_06713_),
    .X(_06714_));
 sg13g2_buf_1 _25643_ (.A(_06714_),
    .X(_06715_));
 sg13g2_mux2_1 _25644_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(net869),
    .S(net146),
    .X(_02442_));
 sg13g2_mux2_1 _25645_ (.A0(\cpu.intr.r_clock_cmp[17] ),
    .A1(net898),
    .S(net146),
    .X(_02443_));
 sg13g2_mux2_1 _25646_ (.A0(\cpu.intr.r_clock_cmp[18] ),
    .A1(net897),
    .S(net146),
    .X(_02444_));
 sg13g2_mux2_1 _25647_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(net896),
    .S(net146),
    .X(_02445_));
 sg13g2_mux2_1 _25648_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(net898),
    .S(net97),
    .X(_02446_));
 sg13g2_mux2_1 _25649_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(net865),
    .S(net146),
    .X(_02447_));
 sg13g2_mux2_1 _25650_ (.A0(\cpu.intr.r_clock_cmp[21] ),
    .A1(net1014),
    .S(net146),
    .X(_02448_));
 sg13g2_mux2_1 _25651_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(net1013),
    .S(_06715_),
    .X(_02449_));
 sg13g2_mux2_1 _25652_ (.A0(\cpu.intr.r_clock_cmp[23] ),
    .A1(_12541_),
    .S(_06715_),
    .X(_02450_));
 sg13g2_mux2_1 _25653_ (.A0(\cpu.intr.r_clock_cmp[24] ),
    .A1(_10205_),
    .S(net146),
    .X(_02451_));
 sg13g2_mux2_1 _25654_ (.A0(\cpu.intr.r_clock_cmp[25] ),
    .A1(_10210_),
    .S(net146),
    .X(_02452_));
 sg13g2_mux2_1 _25655_ (.A0(\cpu.intr.r_clock_cmp[26] ),
    .A1(_10215_),
    .S(_06714_),
    .X(_02453_));
 sg13g2_mux2_1 _25656_ (.A0(\cpu.intr.r_clock_cmp[27] ),
    .A1(_10222_),
    .S(_06714_),
    .X(_02454_));
 sg13g2_mux2_1 _25657_ (.A0(\cpu.intr.r_clock_cmp[28] ),
    .A1(_10227_),
    .S(_06714_),
    .X(_02455_));
 sg13g2_mux2_1 _25658_ (.A0(\cpu.intr.r_clock_cmp[29] ),
    .A1(_10229_),
    .S(_06714_),
    .X(_02456_));
 sg13g2_mux2_1 _25659_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(net897),
    .S(net97),
    .X(_02457_));
 sg13g2_mux2_1 _25660_ (.A0(\cpu.intr.r_clock_cmp[30] ),
    .A1(_10239_),
    .S(_06714_),
    .X(_02458_));
 sg13g2_mux2_1 _25661_ (.A0(\cpu.intr.r_clock_cmp[31] ),
    .A1(_10244_),
    .S(_06714_),
    .X(_02459_));
 sg13g2_mux2_1 _25662_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(net1016),
    .S(net97),
    .X(_02460_));
 sg13g2_mux2_1 _25663_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(_12581_),
    .S(_06711_),
    .X(_02461_));
 sg13g2_mux2_1 _25664_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(net1014),
    .S(_06711_),
    .X(_02462_));
 sg13g2_mux2_1 _25665_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(_12279_),
    .S(_06711_),
    .X(_02463_));
 sg13g2_mux2_1 _25666_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(net1005),
    .S(_06711_),
    .X(_02464_));
 sg13g2_mux2_1 _25667_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(_10205_),
    .S(_06711_),
    .X(_02465_));
 sg13g2_mux2_1 _25668_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(_10210_),
    .S(_06711_),
    .X(_02466_));
 sg13g2_nor4_1 _25669_ (.A(net543),
    .B(_09292_),
    .C(_10097_),
    .D(net679),
    .Y(_06716_));
 sg13g2_buf_2 _25670_ (.A(_06716_),
    .X(_06717_));
 sg13g2_buf_1 _25671_ (.A(_06717_),
    .X(_06718_));
 sg13g2_mux2_1 _25672_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net869),
    .S(net145),
    .X(_02490_));
 sg13g2_mux2_1 _25673_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10215_),
    .S(net145),
    .X(_02491_));
 sg13g2_mux2_1 _25674_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10222_),
    .S(net145),
    .X(_02492_));
 sg13g2_mux2_1 _25675_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10227_),
    .S(net145),
    .X(_02493_));
 sg13g2_mux2_1 _25676_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10229_),
    .S(net145),
    .X(_02494_));
 sg13g2_mux2_1 _25677_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10239_),
    .S(_06718_),
    .X(_02495_));
 sg13g2_mux2_1 _25678_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10244_),
    .S(_06718_),
    .X(_02496_));
 sg13g2_mux2_1 _25679_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net868),
    .S(net171),
    .X(_02497_));
 sg13g2_inv_1 _25680_ (.Y(_06719_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_o21ai_1 _25681_ (.B1(_10101_),
    .Y(_02498_),
    .A1(_06719_),
    .A2(net171));
 sg13g2_inv_1 _25682_ (.Y(_06720_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_o21ai_1 _25683_ (.B1(_10107_),
    .Y(_02499_),
    .A1(_06720_),
    .A2(net171));
 sg13g2_inv_1 _25684_ (.Y(_06721_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25685_ (.B1(_10112_),
    .Y(_02500_),
    .A1(_06721_),
    .A2(net171));
 sg13g2_mux2_1 _25686_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(_12250_),
    .S(net145),
    .X(_02501_));
 sg13g2_mux2_1 _25687_ (.A0(\cpu.intr.r_timer_reload[20] ),
    .A1(net865),
    .S(_10100_),
    .X(_02502_));
 sg13g2_o21ai_1 _25688_ (.B1(_10124_),
    .Y(_02503_),
    .A1(_05603_),
    .A2(_10100_));
 sg13g2_inv_1 _25689_ (.Y(_06722_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25690_ (.B1(_10130_),
    .Y(_02504_),
    .A1(_06722_),
    .A2(net171));
 sg13g2_mux2_1 _25691_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net1005),
    .S(net171),
    .X(_02505_));
 sg13g2_mux2_1 _25692_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(net866),
    .S(net145),
    .X(_02506_));
 sg13g2_mux2_1 _25693_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(net1016),
    .S(net145),
    .X(_02507_));
 sg13g2_mux2_1 _25694_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(net865),
    .S(_06717_),
    .X(_02508_));
 sg13g2_mux2_1 _25695_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(net1014),
    .S(_06717_),
    .X(_02509_));
 sg13g2_mux2_1 _25696_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net1013),
    .S(_06717_),
    .X(_02510_));
 sg13g2_mux2_1 _25697_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(_12283_),
    .S(_06717_),
    .X(_02511_));
 sg13g2_mux2_1 _25698_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10205_),
    .S(_06717_),
    .X(_02512_));
 sg13g2_mux2_1 _25699_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10210_),
    .S(_06717_),
    .X(_02513_));
 sg13g2_inv_1 _25700_ (.Y(_06723_),
    .A(_09842_));
 sg13g2_nor4_1 _25701_ (.A(_11968_),
    .B(_09859_),
    .C(_11965_),
    .D(_11938_),
    .Y(_06724_));
 sg13g2_nand2b_1 _25702_ (.Y(_06725_),
    .B(_06724_),
    .A_N(_11967_));
 sg13g2_nor3_1 _25703_ (.A(_11937_),
    .B(_11935_),
    .C(_06725_),
    .Y(_06726_));
 sg13g2_inv_1 _25704_ (.Y(_06727_),
    .A(_06726_));
 sg13g2_nor4_1 _25705_ (.A(_09848_),
    .B(_09840_),
    .C(_09838_),
    .D(_06727_),
    .Y(_06728_));
 sg13g2_o21ai_1 _25706_ (.B1(_06728_),
    .Y(_06729_),
    .A1(_09881_),
    .A2(_09882_));
 sg13g2_buf_1 _25707_ (.A(_06729_),
    .X(_06730_));
 sg13g2_and2_1 _25708_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_09873_),
    .X(_06731_));
 sg13g2_a221oi_1 _25709_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06731_),
    .B1(_09878_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06732_),
    .A2(_09876_));
 sg13g2_or4_1 _25710_ (.A(_09847_),
    .B(_09858_),
    .C(_09862_),
    .D(_09851_),
    .X(_06733_));
 sg13g2_buf_1 _25711_ (.A(_06733_),
    .X(_06734_));
 sg13g2_a221oi_1 _25712_ (.B2(_06734_),
    .C1(net1138),
    .B1(_00178_),
    .A1(net1136),
    .Y(_06735_),
    .A2(_06723_));
 sg13g2_o21ai_1 _25713_ (.B1(_06735_),
    .Y(_06736_),
    .A1(_09934_),
    .A2(_06732_));
 sg13g2_nor2_1 _25714_ (.A(_06730_),
    .B(_06736_),
    .Y(_06737_));
 sg13g2_a21oi_1 _25715_ (.A1(_06723_),
    .A2(net29),
    .Y(_02514_),
    .B1(_06737_));
 sg13g2_inv_1 _25716_ (.Y(_06738_),
    .A(_09843_));
 sg13g2_a22oi_1 _25717_ (.Y(_06739_),
    .B1(_09873_),
    .B2(\cpu.qspi.r_read_delay[1][1] ),
    .A2(_09876_),
    .A1(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_nand2_1 _25718_ (.Y(_06740_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_09878_));
 sg13g2_a21oi_1 _25719_ (.A1(_06739_),
    .A2(_06740_),
    .Y(_06741_),
    .B1(_09934_));
 sg13g2_xnor2_1 _25720_ (.Y(_06742_),
    .A(_09842_),
    .B(_09843_));
 sg13g2_nor2_1 _25721_ (.A(net1136),
    .B(_06734_),
    .Y(_06743_));
 sg13g2_mux2_1 _25722_ (.A0(_06742_),
    .A1(_09934_),
    .S(_06743_),
    .X(_06744_));
 sg13g2_nor4_1 _25723_ (.A(net1138),
    .B(net29),
    .C(_06741_),
    .D(_06744_),
    .Y(_06745_));
 sg13g2_a21oi_1 _25724_ (.A1(_06738_),
    .A2(net29),
    .Y(_02515_),
    .B1(_06745_));
 sg13g2_inv_1 _25725_ (.Y(_06746_),
    .A(\cpu.qspi.r_count[2] ));
 sg13g2_nor2_1 _25726_ (.A(_09842_),
    .B(_09843_),
    .Y(_06747_));
 sg13g2_xor2_1 _25727_ (.B(_06747_),
    .A(_00179_),
    .X(_06748_));
 sg13g2_nor4_1 _25728_ (.A(_09847_),
    .B(_09858_),
    .C(net1137),
    .D(_09851_),
    .Y(_06749_));
 sg13g2_o21ai_1 _25729_ (.B1(_09935_),
    .Y(_06750_),
    .A1(net1136),
    .A2(_06749_));
 sg13g2_a22oi_1 _25730_ (.Y(_06751_),
    .B1(_06748_),
    .B2(_06750_),
    .A2(_06743_),
    .A1(_09933_));
 sg13g2_a22oi_1 _25731_ (.Y(_06752_),
    .B1(_09873_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09876_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25732_ (.Y(_06753_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09878_));
 sg13g2_a21oi_1 _25733_ (.A1(_06752_),
    .A2(_06753_),
    .Y(_06754_),
    .B1(_09934_));
 sg13g2_nor4_1 _25734_ (.A(net1138),
    .B(net29),
    .C(_06751_),
    .D(_06754_),
    .Y(_06755_));
 sg13g2_a21oi_1 _25735_ (.A1(_06746_),
    .A2(net29),
    .Y(_02516_),
    .B1(_06755_));
 sg13g2_a21oi_1 _25736_ (.A1(net1136),
    .A2(net773),
    .Y(_06756_),
    .B1(_06734_));
 sg13g2_inv_1 _25737_ (.Y(_06757_),
    .A(_06756_));
 sg13g2_a22oi_1 _25738_ (.Y(_06758_),
    .B1(_09873_),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(_09876_),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_nand2_1 _25739_ (.Y(_06759_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_09878_));
 sg13g2_nand2_1 _25740_ (.Y(_06760_),
    .A(_06758_),
    .B(_06759_));
 sg13g2_a22oi_1 _25741_ (.Y(_06761_),
    .B1(_06760_),
    .B2(_09933_),
    .A2(_06757_),
    .A1(_09844_));
 sg13g2_a21oi_1 _25742_ (.A1(_06746_),
    .A2(_06747_),
    .Y(_06762_),
    .B1(_06756_));
 sg13g2_o21ai_1 _25743_ (.B1(\cpu.qspi.r_count[3] ),
    .Y(_06763_),
    .A1(net29),
    .A2(_06762_));
 sg13g2_o21ai_1 _25744_ (.B1(_06763_),
    .Y(_02517_),
    .A1(net29),
    .A2(_06761_));
 sg13g2_or2_1 _25745_ (.X(_06764_),
    .B(_09844_),
    .A(_00254_));
 sg13g2_a21oi_1 _25746_ (.A1(net773),
    .A2(_06764_),
    .Y(_06765_),
    .B1(_06756_));
 sg13g2_mux2_1 _25747_ (.A0(_06765_),
    .A1(\cpu.qspi.r_count[4] ),
    .S(net29),
    .X(_02518_));
 sg13g2_nand2_1 _25748_ (.Y(_06766_),
    .A(_10028_),
    .B(_06367_));
 sg13g2_nor2_1 _25749_ (.A(net581),
    .B(_06766_),
    .Y(_06767_));
 sg13g2_buf_1 _25750_ (.A(_06767_),
    .X(_06768_));
 sg13g2_nand2_1 _25751_ (.Y(_06769_),
    .A(net901),
    .B(_06768_));
 sg13g2_and2_1 _25752_ (.A(_10028_),
    .B(_06367_),
    .X(_06770_));
 sg13g2_buf_1 _25753_ (.A(_06770_),
    .X(_06771_));
 sg13g2_nand2_1 _25754_ (.Y(_06772_),
    .A(_09240_),
    .B(_06771_));
 sg13g2_buf_1 _25755_ (.A(_06772_),
    .X(_06773_));
 sg13g2_nand2_1 _25756_ (.Y(_06774_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06773_));
 sg13g2_a21oi_1 _25757_ (.A1(_06769_),
    .A2(_06774_),
    .Y(_02529_),
    .B1(net623));
 sg13g2_nand2_1 _25758_ (.Y(_06775_),
    .A(net999),
    .B(_06768_));
 sg13g2_nand2_1 _25759_ (.Y(_06776_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06773_));
 sg13g2_a21oi_1 _25760_ (.A1(_06775_),
    .A2(_06776_),
    .Y(_02530_),
    .B1(net623));
 sg13g2_nand2_1 _25761_ (.Y(_06777_),
    .A(net864),
    .B(_06768_));
 sg13g2_nand2_1 _25762_ (.Y(_06778_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06773_));
 sg13g2_nand3_1 _25763_ (.B(_06777_),
    .C(_06778_),
    .A(net728),
    .Y(_02531_));
 sg13g2_nand2_1 _25764_ (.Y(_06779_),
    .A(_12694_),
    .B(_06768_));
 sg13g2_nand2_1 _25765_ (.Y(_06780_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06773_));
 sg13g2_a21oi_1 _25766_ (.A1(_06779_),
    .A2(_06780_),
    .Y(_02532_),
    .B1(_09369_));
 sg13g2_buf_1 _25767_ (.A(_10153_),
    .X(_06781_));
 sg13g2_nor2_1 _25768_ (.A(_06781_),
    .B(_06766_),
    .Y(_06782_));
 sg13g2_nand2_1 _25769_ (.Y(_06783_),
    .A(net901),
    .B(_06782_));
 sg13g2_nand2b_1 _25770_ (.Y(_06784_),
    .B(_06771_),
    .A_N(_06781_));
 sg13g2_buf_1 _25771_ (.A(_06784_),
    .X(_06785_));
 sg13g2_nand2_1 _25772_ (.Y(_06786_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06785_));
 sg13g2_a21oi_1 _25773_ (.A1(_06783_),
    .A2(_06786_),
    .Y(_02533_),
    .B1(_09369_));
 sg13g2_nand2_1 _25774_ (.Y(_06787_),
    .A(net999),
    .B(_06782_));
 sg13g2_nand2_1 _25775_ (.Y(_06788_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06785_));
 sg13g2_buf_1 _25776_ (.A(_09368_),
    .X(_06789_));
 sg13g2_a21oi_1 _25777_ (.A1(_06787_),
    .A2(_06788_),
    .Y(_02534_),
    .B1(net567));
 sg13g2_nand2_1 _25778_ (.Y(_06790_),
    .A(net864),
    .B(_06782_));
 sg13g2_nand2_1 _25779_ (.Y(_06791_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06785_));
 sg13g2_nand3_1 _25780_ (.B(_06790_),
    .C(_06791_),
    .A(net728),
    .Y(_02535_));
 sg13g2_nand2_1 _25781_ (.Y(_06792_),
    .A(net1000),
    .B(_06782_));
 sg13g2_nand2_1 _25782_ (.Y(_06793_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06785_));
 sg13g2_a21oi_1 _25783_ (.A1(_06792_),
    .A2(_06793_),
    .Y(_02536_),
    .B1(net567));
 sg13g2_buf_1 _25784_ (.A(_10080_),
    .X(_06794_));
 sg13g2_nor2_1 _25785_ (.A(net582),
    .B(_06766_),
    .Y(_06795_));
 sg13g2_buf_1 _25786_ (.A(_06795_),
    .X(_06796_));
 sg13g2_nand2_1 _25787_ (.Y(_06797_),
    .A(_06794_),
    .B(_06796_));
 sg13g2_nand2b_1 _25788_ (.Y(_06798_),
    .B(_06771_),
    .A_N(net582));
 sg13g2_buf_1 _25789_ (.A(_06798_),
    .X(_06799_));
 sg13g2_nand2_1 _25790_ (.Y(_06800_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06799_));
 sg13g2_a21oi_1 _25791_ (.A1(_06797_),
    .A2(_06800_),
    .Y(_02537_),
    .B1(net567));
 sg13g2_nand2_1 _25792_ (.Y(_06801_),
    .A(net999),
    .B(_06796_));
 sg13g2_nand2_1 _25793_ (.Y(_06802_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06799_));
 sg13g2_a21oi_1 _25794_ (.A1(_06801_),
    .A2(_06802_),
    .Y(_02538_),
    .B1(net567));
 sg13g2_nand2_1 _25795_ (.Y(_06803_),
    .A(net864),
    .B(_06796_));
 sg13g2_nand2_1 _25796_ (.Y(_06804_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06799_));
 sg13g2_nand3_1 _25797_ (.B(_06803_),
    .C(_06804_),
    .A(net728),
    .Y(_02539_));
 sg13g2_nand2_1 _25798_ (.Y(_06805_),
    .A(net1054),
    .B(_06796_));
 sg13g2_nand2_1 _25799_ (.Y(_06806_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06799_));
 sg13g2_a21oi_1 _25800_ (.A1(_06805_),
    .A2(_06806_),
    .Y(_02540_),
    .B1(net567));
 sg13g2_or3_1 _25801_ (.A(_09933_),
    .B(\cpu.qspi.r_state[14] ),
    .C(_09838_),
    .X(_06807_));
 sg13g2_and2_1 _25802_ (.A(\cpu.qspi.r_mask[1] ),
    .B(_09873_),
    .X(_06808_));
 sg13g2_a221oi_1 _25803_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06808_),
    .B1(_09878_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06809_),
    .A2(_09876_));
 sg13g2_nand2_1 _25804_ (.Y(_06810_),
    .A(_11937_),
    .B(_06809_));
 sg13g2_nor3_2 _25805_ (.A(_09847_),
    .B(_09848_),
    .C(_09840_),
    .Y(_06811_));
 sg13g2_nand3b_1 _25806_ (.B(_06810_),
    .C(_06811_),
    .Y(_06812_),
    .A_N(_06807_));
 sg13g2_buf_2 _25807_ (.A(_06812_),
    .X(_06813_));
 sg13g2_nor4_1 _25808_ (.A(_09858_),
    .B(net1138),
    .C(_09862_),
    .D(_09851_),
    .Y(_06814_));
 sg13g2_and2_1 _25809_ (.A(_06726_),
    .B(_06814_),
    .X(_06815_));
 sg13g2_buf_1 _25810_ (.A(_06815_),
    .X(_06816_));
 sg13g2_nand2_1 _25811_ (.Y(_06817_),
    .A(_09861_),
    .B(_06816_));
 sg13g2_xor2_1 _25812_ (.B(_09881_),
    .A(net172),
    .X(_06818_));
 sg13g2_buf_1 _25813_ (.A(_09397_),
    .X(_06819_));
 sg13g2_mux2_1 _25814_ (.A0(_09686_),
    .A1(net429),
    .S(net139),
    .X(_06820_));
 sg13g2_nand2_1 _25815_ (.Y(_06821_),
    .A(net830),
    .B(_06820_));
 sg13g2_o21ai_1 _25816_ (.B1(_06821_),
    .Y(_06822_),
    .A1(net830),
    .A2(_08762_));
 sg13g2_nand2b_1 _25817_ (.Y(_06823_),
    .B(_09859_),
    .A_N(net172));
 sg13g2_buf_1 _25818_ (.A(net1026),
    .X(_06824_));
 sg13g2_nand3_1 _25819_ (.B(net829),
    .C(net1027),
    .A(_12059_),
    .Y(_06825_));
 sg13g2_mux4_1 _25820_ (.S0(_12059_),
    .A0(_05526_),
    .A1(_05197_),
    .A2(_04975_),
    .A3(_04999_),
    .S1(net1026),
    .X(_06826_));
 sg13g2_nand3_1 _25821_ (.B(_12056_),
    .C(_04968_),
    .A(net1026),
    .Y(_06827_));
 sg13g2_o21ai_1 _25822_ (.B1(_06827_),
    .Y(_06828_),
    .A1(net1026),
    .A2(net994));
 sg13g2_nor2_1 _25823_ (.A(_12060_),
    .B(_12061_),
    .Y(_06829_));
 sg13g2_nand2_1 _25824_ (.Y(_06830_),
    .A(_12056_),
    .B(_06829_));
 sg13g2_or2_1 _25825_ (.X(_06831_),
    .B(_12056_),
    .A(_12071_));
 sg13g2_buf_1 _25826_ (.A(_06831_),
    .X(_06832_));
 sg13g2_o21ai_1 _25827_ (.B1(_06832_),
    .Y(_06833_),
    .A1(_05204_),
    .A2(_06830_));
 sg13g2_a221oi_1 _25828_ (.B2(_12060_),
    .C1(_06833_),
    .B1(_06828_),
    .A1(net994),
    .Y(_06834_),
    .A2(_06826_));
 sg13g2_o21ai_1 _25829_ (.B1(_06834_),
    .Y(_06835_),
    .A1(_04990_),
    .A2(_06825_));
 sg13g2_nor2b_1 _25830_ (.A(_12144_),
    .B_N(net1027),
    .Y(_06836_));
 sg13g2_nor2_1 _25831_ (.A(net994),
    .B(_06836_),
    .Y(_06837_));
 sg13g2_a21oi_1 _25832_ (.A1(_05516_),
    .A2(_06837_),
    .Y(_06838_),
    .B1(_11939_));
 sg13g2_nand2_1 _25833_ (.Y(_06839_),
    .A(_06835_),
    .B(_06838_));
 sg13g2_buf_1 _25834_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06840_));
 sg13g2_nand2_1 _25835_ (.Y(_06841_),
    .A(net1150),
    .B(net1060));
 sg13g2_o21ai_1 _25836_ (.B1(_06841_),
    .Y(_06842_),
    .A1(net1060),
    .A2(_09824_));
 sg13g2_a22oi_1 _25837_ (.Y(_06843_),
    .B1(_06842_),
    .B2(_11965_),
    .A2(_06840_),
    .A1(_09888_));
 sg13g2_a21oi_1 _25838_ (.A1(_09861_),
    .A2(_06816_),
    .Y(_06844_),
    .B1(_11937_));
 sg13g2_nand4_1 _25839_ (.B(_06839_),
    .C(_06843_),
    .A(_06823_),
    .Y(_06845_),
    .D(_06844_));
 sg13g2_a21oi_1 _25840_ (.A1(_11968_),
    .A2(_06822_),
    .Y(_06846_),
    .B1(_06845_));
 sg13g2_buf_1 _25841_ (.A(net1060),
    .X(_06847_));
 sg13g2_buf_1 _25842_ (.A(net139),
    .X(_06848_));
 sg13g2_mux2_1 _25843_ (.A0(_09756_),
    .A1(_00237_),
    .S(net96),
    .X(_06849_));
 sg13g2_nand2_1 _25844_ (.Y(_06850_),
    .A(_09866_),
    .B(_03618_));
 sg13g2_o21ai_1 _25845_ (.B1(_06850_),
    .Y(_06851_),
    .A1(net828),
    .A2(_06849_));
 sg13g2_buf_1 _25846_ (.A(_09397_),
    .X(_06852_));
 sg13g2_mux2_1 _25847_ (.A0(_09664_),
    .A1(net385),
    .S(net139),
    .X(_06853_));
 sg13g2_nand2_1 _25848_ (.Y(_06854_),
    .A(net830),
    .B(_06853_));
 sg13g2_o21ai_1 _25849_ (.B1(_06854_),
    .Y(_06855_),
    .A1(net827),
    .A2(_08556_));
 sg13g2_a22oi_1 _25850_ (.Y(_06856_),
    .B1(_06855_),
    .B2(_11938_),
    .A2(_06851_),
    .A1(_11967_));
 sg13g2_nand2_1 _25851_ (.Y(_06857_),
    .A(_06723_),
    .B(_09843_));
 sg13g2_nand3_1 _25852_ (.B(_09842_),
    .C(_09841_),
    .A(net1137),
    .Y(_06858_));
 sg13g2_o21ai_1 _25853_ (.B1(_06858_),
    .Y(_06859_),
    .A1(_09841_),
    .A2(_06857_));
 sg13g2_nand2b_1 _25854_ (.Y(_06860_),
    .B(net172),
    .A_N(_09843_));
 sg13g2_a21oi_1 _25855_ (.A1(_06857_),
    .A2(_06860_),
    .Y(_06861_),
    .B1(net1137));
 sg13g2_o21ai_1 _25856_ (.B1(_06746_),
    .Y(_06862_),
    .A1(_06859_),
    .A2(_06861_));
 sg13g2_nand2_1 _25857_ (.Y(_06863_),
    .A(net1137),
    .B(_09841_));
 sg13g2_a21oi_1 _25858_ (.A1(_00178_),
    .A2(_06863_),
    .Y(_06864_),
    .B1(_09843_));
 sg13g2_nor2_1 _25859_ (.A(_06746_),
    .B(_06864_),
    .Y(_06865_));
 sg13g2_mux2_1 _25860_ (.A0(_06857_),
    .A1(_09843_),
    .S(net172),
    .X(_06866_));
 sg13g2_nand2_1 _25861_ (.Y(_06867_),
    .A(net1137),
    .B(_06865_));
 sg13g2_o21ai_1 _25862_ (.B1(_06867_),
    .Y(_06868_),
    .A1(_09858_),
    .A2(net1137));
 sg13g2_a21oi_1 _25863_ (.A1(_06865_),
    .A2(_06866_),
    .Y(_06869_),
    .B1(_06868_));
 sg13g2_nand2_1 _25864_ (.Y(_06870_),
    .A(_06862_),
    .B(_06869_));
 sg13g2_nand3_1 _25865_ (.B(_06856_),
    .C(_06870_),
    .A(_06846_),
    .Y(_06871_));
 sg13g2_o21ai_1 _25866_ (.B1(_06871_),
    .Y(_06872_),
    .A1(_06817_),
    .A2(_06818_));
 sg13g2_nand2_1 _25867_ (.Y(_06873_),
    .A(net11),
    .B(_06813_));
 sg13g2_o21ai_1 _25868_ (.B1(_06873_),
    .Y(_02545_),
    .A1(_06813_),
    .A2(_06872_));
 sg13g2_buf_1 _25869_ (.A(_12059_),
    .X(_06874_));
 sg13g2_a22oi_1 _25870_ (.Y(_06875_),
    .B1(_05322_),
    .B2(net994),
    .A2(_05315_),
    .A1(net1027));
 sg13g2_nor2_1 _25871_ (.A(net1026),
    .B(_03006_),
    .Y(_06876_));
 sg13g2_nor2b_1 _25872_ (.A(_05639_),
    .B_N(_06876_),
    .Y(_06877_));
 sg13g2_a21oi_1 _25873_ (.A1(net829),
    .A2(_06875_),
    .Y(_06878_),
    .B1(_06877_));
 sg13g2_nor2_1 _25874_ (.A(net829),
    .B(_05223_),
    .Y(_06879_));
 sg13g2_a21oi_1 _25875_ (.A1(net829),
    .A2(_05301_),
    .Y(_06880_),
    .B1(_06879_));
 sg13g2_nand3_1 _25876_ (.B(_05304_),
    .C(_05307_),
    .A(net1026),
    .Y(_06881_));
 sg13g2_o21ai_1 _25877_ (.B1(_06881_),
    .Y(_06882_),
    .A1(net829),
    .A2(_05229_));
 sg13g2_inv_1 _25878_ (.Y(_06883_),
    .A(_06882_));
 sg13g2_a22oi_1 _25879_ (.Y(_06884_),
    .B1(_06883_),
    .B2(net1027),
    .A2(_06880_),
    .A1(net994));
 sg13g2_nand2_1 _25880_ (.Y(_06885_),
    .A(net945),
    .B(_06884_));
 sg13g2_o21ai_1 _25881_ (.B1(_06885_),
    .Y(_06886_),
    .A1(net945),
    .A2(_06878_));
 sg13g2_inv_1 _25882_ (.Y(_06887_),
    .A(_06837_));
 sg13g2_o21ai_1 _25883_ (.B1(_09851_),
    .Y(_06888_),
    .A1(_05633_),
    .A2(_06887_));
 sg13g2_a21oi_1 _25884_ (.A1(_06832_),
    .A2(_06886_),
    .Y(_06889_),
    .B1(_06888_));
 sg13g2_nor2_1 _25885_ (.A(_11937_),
    .B(_06889_),
    .Y(_06890_));
 sg13g2_mux2_1 _25886_ (.A0(_09527_),
    .A1(net434),
    .S(net139),
    .X(_06891_));
 sg13g2_nand2_1 _25887_ (.Y(_06892_),
    .A(_09397_),
    .B(_06891_));
 sg13g2_o21ai_1 _25888_ (.B1(_06892_),
    .Y(_06893_),
    .A1(_06819_),
    .A2(_08738_));
 sg13g2_nor2_1 _25889_ (.A(_09768_),
    .B(net139),
    .Y(_06894_));
 sg13g2_a21oi_1 _25890_ (.A1(_04849_),
    .A2(_06848_),
    .Y(_06895_),
    .B1(_06894_));
 sg13g2_mux2_1 _25891_ (.A0(_10531_),
    .A1(_06895_),
    .S(net830),
    .X(_06896_));
 sg13g2_a22oi_1 _25892_ (.Y(_06897_),
    .B1(_06896_),
    .B2(_11965_),
    .A2(_06893_),
    .A1(_11968_));
 sg13g2_mux2_1 _25893_ (.A0(_09746_),
    .A1(_00239_),
    .S(_09833_),
    .X(_06898_));
 sg13g2_nand2_1 _25894_ (.Y(_06899_),
    .A(net1060),
    .B(_10838_));
 sg13g2_o21ai_1 _25895_ (.B1(_06899_),
    .Y(_06900_),
    .A1(_09866_),
    .A2(_06898_));
 sg13g2_mux2_1 _25896_ (.A0(_09624_),
    .A1(net386),
    .S(net139),
    .X(_06901_));
 sg13g2_nand2_1 _25897_ (.Y(_06902_),
    .A(net830),
    .B(_06901_));
 sg13g2_o21ai_1 _25898_ (.B1(_06902_),
    .Y(_06903_),
    .A1(net830),
    .A2(_08587_));
 sg13g2_a22oi_1 _25899_ (.Y(_06904_),
    .B1(_06903_),
    .B2(_11938_),
    .A2(_06900_),
    .A1(_11967_));
 sg13g2_and2_1 _25900_ (.A(_06897_),
    .B(_06904_),
    .X(_06905_));
 sg13g2_or2_1 _25901_ (.X(_06906_),
    .B(_06817_),
    .A(_09881_));
 sg13g2_nand4_1 _25902_ (.B(_06890_),
    .C(_06905_),
    .A(_06823_),
    .Y(_06907_),
    .D(_06906_));
 sg13g2_mux2_1 _25903_ (.A0(_06907_),
    .A1(net12),
    .S(_06813_),
    .X(_02546_));
 sg13g2_mux2_1 _25904_ (.A0(_09792_),
    .A1(_00241_),
    .S(net96),
    .X(_06908_));
 sg13g2_nand2_1 _25905_ (.Y(_06909_),
    .A(net828),
    .B(_10881_));
 sg13g2_o21ai_1 _25906_ (.B1(_06909_),
    .Y(_06910_),
    .A1(net828),
    .A2(_06908_));
 sg13g2_nand2_1 _25907_ (.Y(_06911_),
    .A(net945),
    .B(_05034_));
 sg13g2_o21ai_1 _25908_ (.B1(_06911_),
    .Y(_06912_),
    .A1(net945),
    .A2(_05385_));
 sg13g2_nand3_1 _25909_ (.B(_12057_),
    .C(_06912_),
    .A(_06824_),
    .Y(_06913_));
 sg13g2_nand3_1 _25910_ (.B(_12057_),
    .C(_05258_),
    .A(net945),
    .Y(_06914_));
 sg13g2_a21o_1 _25911_ (.A2(_05665_),
    .A1(_03005_),
    .B1(_06874_),
    .X(_06915_));
 sg13g2_a21o_1 _25912_ (.A2(_06915_),
    .A1(_06914_),
    .B1(_06824_),
    .X(_06916_));
 sg13g2_nand2_1 _25913_ (.Y(_06917_),
    .A(_12062_),
    .B(_05041_));
 sg13g2_o21ai_1 _25914_ (.B1(_06917_),
    .Y(_06918_),
    .A1(_12062_),
    .A2(_05252_));
 sg13g2_nand2_1 _25915_ (.Y(_06919_),
    .A(_06874_),
    .B(_06918_));
 sg13g2_o21ai_1 _25916_ (.B1(_06919_),
    .Y(_06920_),
    .A1(_12063_),
    .A2(_05393_));
 sg13g2_nand2_1 _25917_ (.Y(_06921_),
    .A(_03005_),
    .B(_06920_));
 sg13g2_nand4_1 _25918_ (.B(_06913_),
    .C(_06916_),
    .A(_06832_),
    .Y(_06922_),
    .D(_06921_));
 sg13g2_a21oi_1 _25919_ (.A1(_05673_),
    .A2(_06837_),
    .Y(_06923_),
    .B1(_11939_));
 sg13g2_mux2_1 _25920_ (.A0(_09707_),
    .A1(net428),
    .S(net139),
    .X(_06924_));
 sg13g2_nand2_1 _25921_ (.Y(_06925_),
    .A(_06819_),
    .B(_06924_));
 sg13g2_o21ai_1 _25922_ (.B1(_06925_),
    .Y(_06926_),
    .A1(net830),
    .A2(_09046_));
 sg13g2_mux2_1 _25923_ (.A0(_08565_),
    .A1(net654),
    .S(_09397_),
    .X(_06927_));
 sg13g2_o21ai_1 _25924_ (.B1(_06844_),
    .Y(_06928_),
    .A1(_00180_),
    .A2(_06927_));
 sg13g2_a221oi_1 _25925_ (.B2(_11968_),
    .C1(_06928_),
    .B1(_06926_),
    .A1(_06922_),
    .Y(_06929_),
    .A2(_06923_));
 sg13g2_mux2_1 _25926_ (.A0(_09616_),
    .A1(_09610_),
    .S(net139),
    .X(_06930_));
 sg13g2_nand2_1 _25927_ (.Y(_06931_),
    .A(net830),
    .B(_06930_));
 sg13g2_o21ai_1 _25928_ (.B1(_06931_),
    .Y(_06932_),
    .A1(net827),
    .A2(_08691_));
 sg13g2_mux2_1 _25929_ (.A0(_09814_),
    .A1(_00233_),
    .S(net96),
    .X(_06933_));
 sg13g2_nand2b_1 _25930_ (.Y(_06934_),
    .B(net828),
    .A_N(_10612_));
 sg13g2_o21ai_1 _25931_ (.B1(_06934_),
    .Y(_06935_),
    .A1(net828),
    .A2(_06933_));
 sg13g2_a22oi_1 _25932_ (.Y(_06936_),
    .B1(_06935_),
    .B2(_11965_),
    .A2(_06932_),
    .A1(_11938_));
 sg13g2_nand2_1 _25933_ (.Y(_06937_),
    .A(_06929_),
    .B(_06936_));
 sg13g2_a21oi_1 _25934_ (.A1(_11967_),
    .A2(_06910_),
    .Y(_06938_),
    .B1(_06937_));
 sg13g2_nor2_1 _25935_ (.A(net172),
    .B(_09881_),
    .Y(_06939_));
 sg13g2_nor2_1 _25936_ (.A(_06817_),
    .B(_06939_),
    .Y(_06940_));
 sg13g2_or2_1 _25937_ (.X(_06941_),
    .B(_06940_),
    .A(_06813_));
 sg13g2_nand2_1 _25938_ (.Y(_06942_),
    .A(net13),
    .B(_06813_));
 sg13g2_o21ai_1 _25939_ (.B1(_06942_),
    .Y(_02547_),
    .A1(_06938_),
    .A2(_06941_));
 sg13g2_mux2_1 _25940_ (.A0(_09802_),
    .A1(_00235_),
    .S(net96),
    .X(_06943_));
 sg13g2_nand2b_1 _25941_ (.Y(_06944_),
    .B(net828),
    .A_N(_10714_));
 sg13g2_o21ai_1 _25942_ (.B1(_06944_),
    .Y(_06945_),
    .A1(net828),
    .A2(_06943_));
 sg13g2_nor2_1 _25943_ (.A(_09466_),
    .B(_06848_),
    .Y(_06946_));
 sg13g2_a21oi_1 _25944_ (.A1(_09867_),
    .A2(net96),
    .Y(_06947_),
    .B1(_06946_));
 sg13g2_nand2_1 _25945_ (.Y(_06948_),
    .A(net827),
    .B(_06947_));
 sg13g2_nand3b_1 _25946_ (.B(_11935_),
    .C(_09865_),
    .Y(_06949_),
    .A_N(_09864_));
 sg13g2_a21oi_1 _25947_ (.A1(_09868_),
    .A2(_06948_),
    .Y(_06950_),
    .B1(_06949_));
 sg13g2_a21oi_1 _25948_ (.A1(_11965_),
    .A2(_06945_),
    .Y(_06951_),
    .B1(_06950_));
 sg13g2_mux2_1 _25949_ (.A0(_09496_),
    .A1(net435),
    .S(net96),
    .X(_06952_));
 sg13g2_nand2_1 _25950_ (.Y(_06953_),
    .A(net827),
    .B(_06952_));
 sg13g2_o21ai_1 _25951_ (.B1(_06953_),
    .Y(_06954_),
    .A1(net827),
    .A2(_08715_));
 sg13g2_inv_1 _25952_ (.Y(_06955_),
    .A(_00180_));
 sg13g2_nand2_1 _25953_ (.Y(_06956_),
    .A(net698),
    .B(net1060));
 sg13g2_o21ai_1 _25954_ (.B1(_06956_),
    .Y(_06957_),
    .A1(net1060),
    .A2(_09314_));
 sg13g2_a21oi_1 _25955_ (.A1(_06955_),
    .A2(_06957_),
    .Y(_06958_),
    .B1(_09859_));
 sg13g2_nand2_1 _25956_ (.Y(_06959_),
    .A(net945),
    .B(net994));
 sg13g2_mux2_1 _25957_ (.A0(_05071_),
    .A1(_05160_),
    .S(net829),
    .X(_06960_));
 sg13g2_o21ai_1 _25958_ (.B1(_06832_),
    .Y(_06961_),
    .A1(_06959_),
    .A2(_06960_));
 sg13g2_a22oi_1 _25959_ (.Y(_06962_),
    .B1(_05457_),
    .B2(net994),
    .A2(_05450_),
    .A1(net1027));
 sg13g2_a221oi_1 _25960_ (.B2(net829),
    .C1(net945),
    .B1(_06962_),
    .A1(_05053_),
    .Y(_06963_),
    .A2(_06876_));
 sg13g2_mux2_1 _25961_ (.A0(_05077_),
    .A1(_05166_),
    .S(net829),
    .X(_06964_));
 sg13g2_nand3_1 _25962_ (.B(net1027),
    .C(_06964_),
    .A(net945),
    .Y(_06965_));
 sg13g2_nand2b_1 _25963_ (.Y(_06966_),
    .B(_06965_),
    .A_N(_06963_));
 sg13g2_a21oi_1 _25964_ (.A1(_05061_),
    .A2(_06837_),
    .Y(_06967_),
    .B1(_11939_));
 sg13g2_o21ai_1 _25965_ (.B1(_06967_),
    .Y(_06968_),
    .A1(_06961_),
    .A2(_06966_));
 sg13g2_nand3_1 _25966_ (.B(_06958_),
    .C(_06968_),
    .A(_06844_),
    .Y(_06969_));
 sg13g2_a21oi_1 _25967_ (.A1(_11968_),
    .A2(_06954_),
    .Y(_06970_),
    .B1(_06969_));
 sg13g2_mux2_1 _25968_ (.A0(_09780_),
    .A1(_00243_),
    .S(net96),
    .X(_06971_));
 sg13g2_nand2_1 _25969_ (.Y(_06972_),
    .A(net828),
    .B(_03652_));
 sg13g2_o21ai_1 _25970_ (.B1(_06972_),
    .Y(_06973_),
    .A1(_06847_),
    .A2(_06971_));
 sg13g2_mux2_1 _25971_ (.A0(_09557_),
    .A1(_09574_),
    .S(net96),
    .X(_06974_));
 sg13g2_nand2_1 _25972_ (.Y(_06975_),
    .A(net827),
    .B(_06974_));
 sg13g2_o21ai_1 _25973_ (.B1(_06975_),
    .Y(_06976_),
    .A1(net827),
    .A2(_08784_));
 sg13g2_a22oi_1 _25974_ (.Y(_06977_),
    .B1(_06976_),
    .B2(_11938_),
    .A2(_06973_),
    .A1(_11967_));
 sg13g2_and3_1 _25975_ (.X(_06978_),
    .A(_06951_),
    .B(_06970_),
    .C(_06977_));
 sg13g2_nand2_1 _25976_ (.Y(_06979_),
    .A(net14),
    .B(_06813_));
 sg13g2_o21ai_1 _25977_ (.B1(_06979_),
    .Y(_02548_),
    .A1(_06941_),
    .A2(_06978_));
 sg13g2_mux4_1 _25978_ (.S0(_05547_),
    .A0(_09262_),
    .A1(_09248_),
    .A2(_09246_),
    .A3(_09252_),
    .S1(_06379_),
    .X(_06980_));
 sg13g2_mux4_1 _25979_ (.S0(_05547_),
    .A0(_09255_),
    .A1(_09264_),
    .A2(_09260_),
    .A3(_09245_),
    .S1(_06379_),
    .X(_06981_));
 sg13g2_nor2b_1 _25980_ (.A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B_N(_06981_),
    .Y(_06982_));
 sg13g2_a21oi_1 _25981_ (.A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .A2(_06980_),
    .Y(_06983_),
    .B1(_06982_));
 sg13g2_mux4_1 _25982_ (.S0(_05547_),
    .A0(_09253_),
    .A1(_09266_),
    .A2(_09249_),
    .A3(_09257_),
    .S1(_06379_),
    .X(_06984_));
 sg13g2_nand3b_1 _25983_ (.B(\cpu.gpio.r_spi_miso_src[1][3] ),
    .C(_06984_),
    .Y(_06985_),
    .A_N(_00150_));
 sg13g2_o21ai_1 _25984_ (.B1(_06985_),
    .Y(_06986_),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .A2(_06983_));
 sg13g2_mux4_1 _25985_ (.S0(_04873_),
    .A0(_09262_),
    .A1(_09248_),
    .A2(_09246_),
    .A3(_09252_),
    .S1(_06378_),
    .X(_06987_));
 sg13g2_mux4_1 _25986_ (.S0(_04873_),
    .A0(_09255_),
    .A1(_09264_),
    .A2(_09260_),
    .A3(_09245_),
    .S1(_06378_),
    .X(_06988_));
 sg13g2_nor2b_1 _25987_ (.A(\cpu.gpio.r_spi_miso_src[0][2] ),
    .B_N(_06988_),
    .Y(_06989_));
 sg13g2_a21oi_1 _25988_ (.A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .A2(_06987_),
    .Y(_06990_),
    .B1(_06989_));
 sg13g2_mux4_1 _25989_ (.S0(_04873_),
    .A0(_09253_),
    .A1(_09266_),
    .A2(_09249_),
    .A3(_09257_),
    .S1(_06378_),
    .X(_06991_));
 sg13g2_nand3b_1 _25990_ (.B(\cpu.gpio.r_spi_miso_src[0][3] ),
    .C(_06991_),
    .Y(_06992_),
    .A_N(_00110_));
 sg13g2_o21ai_1 _25991_ (.B1(_06992_),
    .Y(_06993_),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .A2(_06990_));
 sg13g2_mux2_1 _25992_ (.A0(_06986_),
    .A1(_06993_),
    .S(_11988_),
    .X(_06994_));
 sg13g2_nor2_1 _25993_ (.A(net1143),
    .B(_12036_),
    .Y(_06995_));
 sg13g2_nor2b_1 _25994_ (.A(_09318_),
    .B_N(_09356_),
    .Y(_06996_));
 sg13g2_a22oi_1 _25995_ (.Y(_06997_),
    .B1(_06996_),
    .B2(net595),
    .A2(_06995_),
    .A1(_09318_));
 sg13g2_nand3b_1 _25996_ (.B(_09321_),
    .C(net916),
    .Y(_06998_),
    .A_N(_06997_));
 sg13g2_buf_4 _25997_ (.X(_06999_),
    .A(_06998_));
 sg13g2_mux2_1 _25998_ (.A0(_06994_),
    .A1(_09343_),
    .S(_06999_),
    .X(_02588_));
 sg13g2_mux2_1 _25999_ (.A0(_09343_),
    .A1(_09342_),
    .S(_06999_),
    .X(_02589_));
 sg13g2_mux2_1 _26000_ (.A0(_09342_),
    .A1(_09346_),
    .S(_06999_),
    .X(_02590_));
 sg13g2_mux2_1 _26001_ (.A0(_09346_),
    .A1(_09340_),
    .S(_06999_),
    .X(_02591_));
 sg13g2_mux2_1 _26002_ (.A0(_09340_),
    .A1(_09348_),
    .S(_06999_),
    .X(_02592_));
 sg13g2_mux2_1 _26003_ (.A0(_09348_),
    .A1(_09347_),
    .S(_06999_),
    .X(_02593_));
 sg13g2_mux2_1 _26004_ (.A0(_09347_),
    .A1(_09341_),
    .S(_06999_),
    .X(_02594_));
 sg13g2_mux2_1 _26005_ (.A0(_09341_),
    .A1(\cpu.spi.r_in[7] ),
    .S(_06999_),
    .X(_02595_));
 sg13g2_nand2_1 _26006_ (.Y(_07000_),
    .A(net1144),
    .B(_09301_));
 sg13g2_nor2_1 _26007_ (.A(net1145),
    .B(_11999_),
    .Y(_07001_));
 sg13g2_buf_2 _26008_ (.A(_07001_),
    .X(_07002_));
 sg13g2_inv_1 _26009_ (.Y(_07003_),
    .A(net1144));
 sg13g2_a22oi_1 _26010_ (.Y(_07004_),
    .B1(_07002_),
    .B2(_07003_),
    .A2(_12037_),
    .A1(_09357_));
 sg13g2_nand4_1 _26011_ (.B(_12032_),
    .C(_12041_),
    .A(_07000_),
    .Y(_07005_),
    .D(_07004_));
 sg13g2_buf_1 _26012_ (.A(_07005_),
    .X(_07006_));
 sg13g2_buf_1 _26013_ (.A(_09290_),
    .X(_07007_));
 sg13g2_nand2b_1 _26014_ (.Y(_07008_),
    .B(_00225_),
    .A_N(_12044_));
 sg13g2_buf_1 _26015_ (.A(_00227_),
    .X(_07009_));
 sg13g2_buf_1 _26016_ (.A(_07009_),
    .X(_07010_));
 sg13g2_nor2_1 _26017_ (.A(_09290_),
    .B(net944),
    .Y(_07011_));
 sg13g2_a221oi_1 _26018_ (.B2(_07011_),
    .C1(net746),
    .B1(_07008_),
    .A1(net826),
    .Y(_07012_),
    .A2(net1057));
 sg13g2_nand2_1 _26019_ (.Y(_07013_),
    .A(\cpu.spi.r_out[0] ),
    .B(net58));
 sg13g2_o21ai_1 _26020_ (.B1(_07013_),
    .Y(_02603_),
    .A1(net58),
    .A2(_07012_));
 sg13g2_mux2_1 _26021_ (.A0(_00183_),
    .A1(_00225_),
    .S(net595),
    .X(_07014_));
 sg13g2_a22oi_1 _26022_ (.Y(_07015_),
    .B1(_07002_),
    .B2(_10087_),
    .A2(net746),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26023_ (.B1(_07015_),
    .Y(_07016_),
    .A1(net826),
    .A2(_07014_));
 sg13g2_mux2_1 _26024_ (.A0(_07016_),
    .A1(\cpu.spi.r_out[1] ),
    .S(net58),
    .X(_02604_));
 sg13g2_mux2_1 _26025_ (.A0(_00184_),
    .A1(_00183_),
    .S(net595),
    .X(_07017_));
 sg13g2_a22oi_1 _26026_ (.Y(_07018_),
    .B1(_07002_),
    .B2(net1048),
    .A2(net746),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26027_ (.B1(_07018_),
    .Y(_07019_),
    .A1(net826),
    .A2(_07017_));
 sg13g2_mux2_1 _26028_ (.A0(_07019_),
    .A1(\cpu.spi.r_out[2] ),
    .S(_07006_),
    .X(_02605_));
 sg13g2_mux2_1 _26029_ (.A0(_00289_),
    .A1(_00184_),
    .S(net595),
    .X(_07020_));
 sg13g2_a22oi_1 _26030_ (.Y(_07021_),
    .B1(_07002_),
    .B2(net1133),
    .A2(net746),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26031_ (.B1(_07021_),
    .Y(_07022_),
    .A1(net826),
    .A2(_07020_));
 sg13g2_mux2_1 _26032_ (.A0(_07022_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net58),
    .X(_02606_));
 sg13g2_mux2_1 _26033_ (.A0(_00185_),
    .A1(_00289_),
    .S(net595),
    .X(_07023_));
 sg13g2_a22oi_1 _26034_ (.Y(_07024_),
    .B1(_07002_),
    .B2(_10116_),
    .A2(net746),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26035_ (.B1(_07024_),
    .Y(_07025_),
    .A1(net826),
    .A2(_07023_));
 sg13g2_mux2_1 _26036_ (.A0(_07025_),
    .A1(\cpu.spi.r_out[4] ),
    .S(net58),
    .X(_02607_));
 sg13g2_mux2_1 _26037_ (.A0(_00186_),
    .A1(_00185_),
    .S(net595),
    .X(_07026_));
 sg13g2_a22oi_1 _26038_ (.Y(_07027_),
    .B1(_07002_),
    .B2(_10122_),
    .A2(net746),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26039_ (.B1(_07027_),
    .Y(_07028_),
    .A1(_07007_),
    .A2(_07026_));
 sg13g2_mux2_1 _26040_ (.A0(_07028_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net58),
    .X(_02608_));
 sg13g2_buf_1 _26041_ (.A(_00187_),
    .X(_07029_));
 sg13g2_mux2_1 _26042_ (.A0(_07029_),
    .A1(_00186_),
    .S(net595),
    .X(_07030_));
 sg13g2_a22oi_1 _26043_ (.Y(_07031_),
    .B1(_07002_),
    .B2(_10128_),
    .A2(_12024_),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26044_ (.B1(_07031_),
    .Y(_07032_),
    .A1(_07007_),
    .A2(_07030_));
 sg13g2_mux2_1 _26045_ (.A0(_07032_),
    .A1(\cpu.spi.r_out[6] ),
    .S(net58),
    .X(_02609_));
 sg13g2_buf_1 _26046_ (.A(_00283_),
    .X(_07033_));
 sg13g2_mux2_1 _26047_ (.A0(_07033_),
    .A1(_07029_),
    .S(_12044_),
    .X(_07034_));
 sg13g2_a22oi_1 _26048_ (.Y(_07035_),
    .B1(_07002_),
    .B2(_10131_),
    .A2(_12024_),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26049_ (.B1(_07035_),
    .Y(_07036_),
    .A1(net826),
    .A2(_07034_));
 sg13g2_mux2_1 _26050_ (.A0(_07036_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net58),
    .X(_02610_));
 sg13g2_or2_1 _26051_ (.X(_07037_),
    .B(_09366_),
    .A(net917));
 sg13g2_buf_1 _26052_ (.A(_07037_),
    .X(_07038_));
 sg13g2_nand2_1 _26053_ (.Y(_07039_),
    .A(net873),
    .B(_07038_));
 sg13g2_o21ai_1 _26054_ (.B1(_07039_),
    .Y(_02613_),
    .A1(net653),
    .A2(_07038_));
 sg13g2_buf_1 _26055_ (.A(_11975_),
    .X(_07040_));
 sg13g2_buf_1 _26056_ (.A(net943),
    .X(_07041_));
 sg13g2_nand2_1 _26057_ (.Y(_07042_),
    .A(net825),
    .B(_07038_));
 sg13g2_o21ai_1 _26058_ (.B1(_07042_),
    .Y(_02614_),
    .A1(_03019_),
    .A2(_07038_));
 sg13g2_nor2b_1 _26059_ (.A(_09294_),
    .B_N(_05112_),
    .Y(_07043_));
 sg13g2_buf_4 _26060_ (.X(_07044_),
    .A(_07043_));
 sg13g2_mux2_1 _26061_ (.A0(\cpu.spi.r_timeout[0] ),
    .A1(net868),
    .S(_07044_),
    .X(_02618_));
 sg13g2_mux2_1 _26062_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(net867),
    .S(_07044_),
    .X(_02619_));
 sg13g2_mux2_1 _26063_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(net866),
    .S(_07044_),
    .X(_02620_));
 sg13g2_mux2_1 _26064_ (.A0(\cpu.spi.r_timeout[3] ),
    .A1(net1016),
    .S(_07044_),
    .X(_02621_));
 sg13g2_mux2_1 _26065_ (.A0(\cpu.spi.r_timeout[4] ),
    .A1(net1015),
    .S(_07044_),
    .X(_02622_));
 sg13g2_mux2_1 _26066_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(net1014),
    .S(_07044_),
    .X(_02623_));
 sg13g2_mux2_1 _26067_ (.A0(\cpu.spi.r_timeout[6] ),
    .A1(_12279_),
    .S(_07044_),
    .X(_02624_));
 sg13g2_mux2_1 _26068_ (.A0(\cpu.spi.r_timeout[7] ),
    .A1(net1012),
    .S(_07044_),
    .X(_02625_));
 sg13g2_or2_1 _26069_ (.X(_07045_),
    .B(_09317_),
    .A(net1145));
 sg13g2_nand3_1 _26070_ (.B(_09339_),
    .C(_09351_),
    .A(_09320_),
    .Y(_07046_));
 sg13g2_or3_1 _26071_ (.A(_11973_),
    .B(_09324_),
    .C(_07046_),
    .X(_07047_));
 sg13g2_nand2_1 _26072_ (.Y(_07048_),
    .A(_09317_),
    .B(_07046_));
 sg13g2_nand4_1 _26073_ (.B(_07045_),
    .C(_07047_),
    .A(_12032_),
    .Y(_07049_),
    .D(_07048_));
 sg13g2_buf_2 _26074_ (.A(_07049_),
    .X(_07050_));
 sg13g2_buf_1 _26075_ (.A(_07050_),
    .X(_07051_));
 sg13g2_and2_1 _26076_ (.A(net870),
    .B(\cpu.spi.r_timeout[0] ),
    .X(_07052_));
 sg13g2_a21oi_1 _26077_ (.A1(net826),
    .A2(_00286_),
    .Y(_07053_),
    .B1(_07052_));
 sg13g2_nand2_1 _26078_ (.Y(_07054_),
    .A(_09326_),
    .B(net32));
 sg13g2_o21ai_1 _26079_ (.B1(_07054_),
    .Y(_02626_),
    .A1(net32),
    .A2(_07053_));
 sg13g2_nor3_1 _26080_ (.A(_09326_),
    .B(_09327_),
    .C(_07050_),
    .Y(_07055_));
 sg13g2_a21oi_1 _26081_ (.A1(_09326_),
    .A2(_09327_),
    .Y(_07056_),
    .B1(_07055_));
 sg13g2_nor2_1 _26082_ (.A(_09290_),
    .B(_07050_),
    .Y(_07057_));
 sg13g2_buf_2 _26083_ (.A(_07057_),
    .X(_07058_));
 sg13g2_a22oi_1 _26084_ (.Y(_07059_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[1] ),
    .A2(net32),
    .A1(_09327_));
 sg13g2_o21ai_1 _26085_ (.B1(_07059_),
    .Y(_02627_),
    .A1(net870),
    .A2(_07056_));
 sg13g2_a22oi_1 _26086_ (.Y(_07060_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[2] ),
    .A2(net32),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_o21ai_1 _26087_ (.B1(\cpu.spi.r_timeout_count[2] ),
    .Y(_07061_),
    .A1(_09326_),
    .A2(_09327_));
 sg13g2_o21ai_1 _26088_ (.B1(_07061_),
    .Y(_07062_),
    .A1(_09329_),
    .A2(net32));
 sg13g2_nand2_1 _26089_ (.Y(_07063_),
    .A(net826),
    .B(_07062_));
 sg13g2_nand2_1 _26090_ (.Y(_02628_),
    .A(_07060_),
    .B(_07063_));
 sg13g2_nor2_1 _26091_ (.A(_09331_),
    .B(_07050_),
    .Y(_07064_));
 sg13g2_a21oi_1 _26092_ (.A1(\cpu.spi.r_timeout_count[3] ),
    .A2(_09329_),
    .Y(_07065_),
    .B1(_07064_));
 sg13g2_a22oi_1 _26093_ (.Y(_07066_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[3] ),
    .A2(_07051_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_o21ai_1 _26094_ (.B1(_07066_),
    .Y(_02629_),
    .A1(net870),
    .A2(_07065_));
 sg13g2_nor2_1 _26095_ (.A(_09333_),
    .B(_07050_),
    .Y(_07067_));
 sg13g2_a21oi_1 _26096_ (.A1(\cpu.spi.r_timeout_count[4] ),
    .A2(_09331_),
    .Y(_07068_),
    .B1(_07067_));
 sg13g2_a22oi_1 _26097_ (.Y(_07069_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[4] ),
    .A2(_07051_),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_o21ai_1 _26098_ (.B1(_07069_),
    .Y(_02630_),
    .A1(net870),
    .A2(_07068_));
 sg13g2_nor2_1 _26099_ (.A(_09335_),
    .B(_07050_),
    .Y(_07070_));
 sg13g2_a21oi_1 _26100_ (.A1(\cpu.spi.r_timeout_count[5] ),
    .A2(_09333_),
    .Y(_07071_),
    .B1(_07070_));
 sg13g2_a22oi_1 _26101_ (.Y(_07072_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[5] ),
    .A2(net32),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_o21ai_1 _26102_ (.B1(_07072_),
    .Y(_02631_),
    .A1(net870),
    .A2(_07071_));
 sg13g2_nor2_1 _26103_ (.A(_09337_),
    .B(_07050_),
    .Y(_07073_));
 sg13g2_a21oi_1 _26104_ (.A1(\cpu.spi.r_timeout_count[6] ),
    .A2(_09335_),
    .Y(_07074_),
    .B1(_07073_));
 sg13g2_a22oi_1 _26105_ (.Y(_07075_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[6] ),
    .A2(net32),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_o21ai_1 _26106_ (.B1(_07075_),
    .Y(_02632_),
    .A1(net870),
    .A2(_07074_));
 sg13g2_nor3_1 _26107_ (.A(_09325_),
    .B(_09337_),
    .C(_07050_),
    .Y(_07076_));
 sg13g2_a21oi_1 _26108_ (.A1(_09325_),
    .A2(_09337_),
    .Y(_07077_),
    .B1(_07076_));
 sg13g2_a22oi_1 _26109_ (.Y(_07078_),
    .B1(_07058_),
    .B2(\cpu.spi.r_timeout[7] ),
    .A2(net32),
    .A1(_09325_));
 sg13g2_o21ai_1 _26110_ (.B1(_07078_),
    .Y(_02633_),
    .A1(net870),
    .A2(_07077_));
 sg13g2_buf_1 _26111_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07079_));
 sg13g2_nor2_1 _26112_ (.A(_07079_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07080_));
 sg13g2_nand2_1 _26113_ (.Y(_07081_),
    .A(_09954_),
    .B(_07080_));
 sg13g2_nor2_1 _26114_ (.A(net917),
    .B(_07081_),
    .Y(_07082_));
 sg13g2_buf_1 _26115_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07083_));
 sg13g2_buf_1 _26116_ (.A(net1106),
    .X(_07084_));
 sg13g2_buf_1 _26117_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07085_));
 sg13g2_buf_1 _26118_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07086_));
 sg13g2_buf_1 _26119_ (.A(_07086_),
    .X(_07087_));
 sg13g2_nor2_2 _26120_ (.A(_07085_),
    .B(net941),
    .Y(_07088_));
 sg13g2_buf_2 _26121_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07089_));
 sg13g2_inv_1 _26122_ (.Y(_07090_),
    .A(_07089_));
 sg13g2_nand3_1 _26123_ (.B(net942),
    .C(_07088_),
    .A(_07090_),
    .Y(_07091_));
 sg13g2_o21ai_1 _26124_ (.B1(_07091_),
    .Y(_07092_),
    .A1(net942),
    .A2(_07088_));
 sg13g2_and2_1 _26125_ (.A(_07082_),
    .B(_07092_),
    .X(_07093_));
 sg13g2_buf_2 _26126_ (.A(_07093_),
    .X(_07094_));
 sg13g2_mux2_1 _26127_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07094_),
    .X(_02646_));
 sg13g2_mux2_1 _26128_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07094_),
    .X(_02647_));
 sg13g2_mux2_1 _26129_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07094_),
    .X(_02648_));
 sg13g2_mux2_1 _26130_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07094_),
    .X(_02649_));
 sg13g2_mux2_1 _26131_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07094_),
    .X(_02650_));
 sg13g2_mux2_1 _26132_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07094_),
    .X(_02651_));
 sg13g2_xor2_1 _26133_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07095_));
 sg13g2_mux2_1 _26134_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07095_),
    .S(_07094_),
    .X(_02652_));
 sg13g2_and4_1 _26135_ (.A(_07089_),
    .B(_07084_),
    .C(_07082_),
    .D(_07088_),
    .X(_07096_));
 sg13g2_buf_1 _26136_ (.A(_07096_),
    .X(_07097_));
 sg13g2_mux2_1 _26137_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net175),
    .X(_02653_));
 sg13g2_mux2_1 _26138_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net175),
    .X(_02654_));
 sg13g2_mux2_1 _26139_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net175),
    .X(_02655_));
 sg13g2_mux2_1 _26140_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net175),
    .X(_02656_));
 sg13g2_mux2_1 _26141_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07097_),
    .X(_02657_));
 sg13g2_mux2_1 _26142_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net175),
    .X(_02658_));
 sg13g2_mux2_1 _26143_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net175),
    .X(_02659_));
 sg13g2_mux2_1 _26144_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07095_),
    .S(net175),
    .X(_02660_));
 sg13g2_buf_1 _26145_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07098_));
 sg13g2_buf_1 _26146_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07099_));
 sg13g2_buf_1 _26147_ (.A(_07099_),
    .X(_07100_));
 sg13g2_buf_1 _26148_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07101_));
 sg13g2_buf_1 _26149_ (.A(net1103),
    .X(_07102_));
 sg13g2_nor2_1 _26150_ (.A(net1070),
    .B(net1069),
    .Y(_07103_));
 sg13g2_and3_1 _26151_ (.X(_07104_),
    .A(_12008_),
    .B(_07103_),
    .C(_06367_));
 sg13g2_buf_2 _26152_ (.A(_07104_),
    .X(_07105_));
 sg13g2_nand2_2 _26153_ (.Y(_07106_),
    .A(net413),
    .B(_07105_));
 sg13g2_nand4_1 _26154_ (.B(net940),
    .C(net939),
    .A(net1104),
    .Y(_07107_),
    .D(_07106_));
 sg13g2_nor2_1 _26155_ (.A(net1104),
    .B(net1103),
    .Y(_07108_));
 sg13g2_o21ai_1 _26156_ (.B1(_07108_),
    .Y(_07109_),
    .A1(net940),
    .A2(_07106_));
 sg13g2_buf_1 _26157_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07110_));
 sg13g2_buf_1 _26158_ (.A(_07110_),
    .X(_07111_));
 sg13g2_a21o_1 _26159_ (.A2(_07109_),
    .A1(_07107_),
    .B1(_07111_),
    .X(_07112_));
 sg13g2_nand2_1 _26160_ (.Y(_07113_),
    .A(_07099_),
    .B(net1103));
 sg13g2_buf_1 _26161_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07114_));
 sg13g2_nor2_1 _26162_ (.A(_07114_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07115_));
 sg13g2_and2_1 _26163_ (.A(_09954_),
    .B(_07115_),
    .X(_07116_));
 sg13g2_buf_2 _26164_ (.A(_07116_),
    .X(_07117_));
 sg13g2_nor2b_1 _26165_ (.A(_07117_),
    .B_N(net1103),
    .Y(_07118_));
 sg13g2_inv_2 _26166_ (.Y(_07119_),
    .A(net1104));
 sg13g2_mux2_1 _26167_ (.A0(_07113_),
    .A1(_07118_),
    .S(_07119_),
    .X(_07120_));
 sg13g2_nand2b_1 _26168_ (.Y(_07121_),
    .B(_07117_),
    .A_N(net939));
 sg13g2_o21ai_1 _26169_ (.B1(_07121_),
    .Y(_07122_),
    .A1(net938),
    .A2(_07120_));
 sg13g2_nand3_1 _26170_ (.B(_07112_),
    .C(_07122_),
    .A(net1066),
    .Y(_07123_));
 sg13g2_buf_2 _26171_ (.A(_07123_),
    .X(_07124_));
 sg13g2_buf_1 _26172_ (.A(_07124_),
    .X(_07125_));
 sg13g2_nor2_1 _26173_ (.A(net1104),
    .B(_07110_),
    .Y(_07126_));
 sg13g2_xnor2_1 _26174_ (.Y(_07127_),
    .A(_07102_),
    .B(_07126_));
 sg13g2_buf_1 _26175_ (.A(_07127_),
    .X(_07128_));
 sg13g2_buf_1 _26176_ (.A(_07128_),
    .X(_07129_));
 sg13g2_nor2b_1 _26177_ (.A(net639),
    .B_N(_10080_),
    .Y(_07130_));
 sg13g2_a21oi_1 _26178_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net639),
    .Y(_07131_),
    .B1(_07130_));
 sg13g2_nand2_1 _26179_ (.Y(_07132_),
    .A(\cpu.uart.r_out[0] ),
    .B(net31));
 sg13g2_o21ai_1 _26180_ (.B1(_07132_),
    .Y(_02661_),
    .A1(net31),
    .A2(_07131_));
 sg13g2_nor2b_1 _26181_ (.A(net639),
    .B_N(_10087_),
    .Y(_07133_));
 sg13g2_a21oi_1 _26182_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net639),
    .Y(_07134_),
    .B1(_07133_));
 sg13g2_nand2_1 _26183_ (.Y(_07135_),
    .A(\cpu.uart.r_out[1] ),
    .B(net31));
 sg13g2_o21ai_1 _26184_ (.B1(_07135_),
    .Y(_02662_),
    .A1(net31),
    .A2(_07134_));
 sg13g2_nor2b_1 _26185_ (.A(_07128_),
    .B_N(_10164_),
    .Y(_07136_));
 sg13g2_a21oi_1 _26186_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net639),
    .Y(_07137_),
    .B1(_07136_));
 sg13g2_nand2_1 _26187_ (.Y(_07138_),
    .A(\cpu.uart.r_out[2] ),
    .B(_07124_));
 sg13g2_o21ai_1 _26188_ (.B1(_07138_),
    .Y(_02663_),
    .A1(net31),
    .A2(_07137_));
 sg13g2_nor2b_1 _26189_ (.A(_07128_),
    .B_N(net1133),
    .Y(_07139_));
 sg13g2_a21oi_1 _26190_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net639),
    .Y(_07140_),
    .B1(_07139_));
 sg13g2_nand2_1 _26191_ (.Y(_07141_),
    .A(\cpu.uart.r_out[3] ),
    .B(_07124_));
 sg13g2_o21ai_1 _26192_ (.B1(_07141_),
    .Y(_02664_),
    .A1(net31),
    .A2(_07140_));
 sg13g2_nor2b_1 _26193_ (.A(_07128_),
    .B_N(_10116_),
    .Y(_07142_));
 sg13g2_a21oi_1 _26194_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net639),
    .Y(_07143_),
    .B1(_07142_));
 sg13g2_nand2_1 _26195_ (.Y(_07144_),
    .A(\cpu.uart.r_out[4] ),
    .B(_07124_));
 sg13g2_o21ai_1 _26196_ (.B1(_07144_),
    .Y(_02665_),
    .A1(net31),
    .A2(_07143_));
 sg13g2_nor2b_1 _26197_ (.A(_07128_),
    .B_N(_10122_),
    .Y(_07145_));
 sg13g2_a21oi_1 _26198_ (.A1(\cpu.uart.r_out[6] ),
    .A2(_07129_),
    .Y(_07146_),
    .B1(_07145_));
 sg13g2_nand2_1 _26199_ (.Y(_07147_),
    .A(\cpu.uart.r_out[5] ),
    .B(_07124_));
 sg13g2_o21ai_1 _26200_ (.B1(_07147_),
    .Y(_02666_),
    .A1(net31),
    .A2(_07146_));
 sg13g2_nor2b_1 _26201_ (.A(_07128_),
    .B_N(_10128_),
    .Y(_07148_));
 sg13g2_a21oi_1 _26202_ (.A1(\cpu.uart.r_out[7] ),
    .A2(_07129_),
    .Y(_07149_),
    .B1(_07148_));
 sg13g2_nand2_1 _26203_ (.Y(_07150_),
    .A(\cpu.uart.r_out[6] ),
    .B(_07124_));
 sg13g2_o21ai_1 _26204_ (.B1(_07150_),
    .Y(_02667_),
    .A1(_07125_),
    .A2(_07149_));
 sg13g2_nor3_1 _26205_ (.A(_07033_),
    .B(_07124_),
    .C(net639),
    .Y(_07151_));
 sg13g2_a21o_1 _26206_ (.A2(_07125_),
    .A1(\cpu.uart.r_out[7] ),
    .B1(_07151_),
    .X(_02668_));
 sg13g2_nand2b_1 _26207_ (.Y(_07152_),
    .B(_09982_),
    .A_N(_09943_));
 sg13g2_nor3_1 _26208_ (.A(net1105),
    .B(_07086_),
    .C(net1106),
    .Y(_07153_));
 sg13g2_a22oi_1 _26209_ (.Y(_07154_),
    .B1(_07152_),
    .B2(_07153_),
    .A2(net1106),
    .A1(net1105));
 sg13g2_nor4_1 _26210_ (.A(_07089_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07086_),
    .D(net1106),
    .Y(_07155_));
 sg13g2_a21o_1 _26211_ (.A2(_07152_),
    .A1(net1105),
    .B1(_07086_),
    .X(_07156_));
 sg13g2_a22oi_1 _26212_ (.Y(_07157_),
    .B1(_07156_),
    .B2(net1106),
    .A2(_07155_),
    .A1(_07095_));
 sg13g2_o21ai_1 _26213_ (.B1(_07157_),
    .Y(_07158_),
    .A1(_07090_),
    .A2(_07154_));
 sg13g2_nor2_1 _26214_ (.A(_07090_),
    .B(_07085_),
    .Y(_07159_));
 sg13g2_nor2b_1 _26215_ (.A(net1106),
    .B_N(_07095_),
    .Y(_07160_));
 sg13g2_nand2_1 _26216_ (.Y(_07161_),
    .A(net1105),
    .B(net1106));
 sg13g2_nor2_1 _26217_ (.A(_07089_),
    .B(_07161_),
    .Y(_07162_));
 sg13g2_a21oi_1 _26218_ (.A1(_07159_),
    .A2(_07160_),
    .Y(_07163_),
    .B1(_07162_));
 sg13g2_nor3_1 _26219_ (.A(_07087_),
    .B(_07081_),
    .C(_07163_),
    .Y(_07164_));
 sg13g2_xor2_1 _26220_ (.B(_07088_),
    .A(_07084_),
    .X(_07165_));
 sg13g2_o21ai_1 _26221_ (.B1(net1066),
    .Y(_07166_),
    .A1(_09954_),
    .A2(_07165_));
 sg13g2_nor3_1 _26222_ (.A(_07158_),
    .B(_07164_),
    .C(_07166_),
    .Y(_07167_));
 sg13g2_and2_1 _26223_ (.A(_07089_),
    .B(net1105),
    .X(_07168_));
 sg13g2_buf_1 _26224_ (.A(_07168_),
    .X(_07169_));
 sg13g2_o21ai_1 _26225_ (.B1(net942),
    .Y(_07170_),
    .A1(net941),
    .A2(_07169_));
 sg13g2_nor2b_1 _26226_ (.A(_07155_),
    .B_N(_07170_),
    .Y(_07171_));
 sg13g2_and2_1 _26227_ (.A(_07167_),
    .B(_07171_),
    .X(_07172_));
 sg13g2_nor2_1 _26228_ (.A(_07079_),
    .B(_07167_),
    .Y(_07173_));
 sg13g2_a21oi_1 _26229_ (.A1(_07079_),
    .A2(_07172_),
    .Y(_02671_),
    .B1(_07173_));
 sg13g2_nand2_1 _26230_ (.Y(_07174_),
    .A(_07079_),
    .B(_07171_));
 sg13g2_inv_1 _26231_ (.Y(_07175_),
    .A(\cpu.uart.r_rcnt[1] ));
 sg13g2_a21oi_1 _26232_ (.A1(_07167_),
    .A2(_07174_),
    .Y(_07176_),
    .B1(_07175_));
 sg13g2_a21o_1 _26233_ (.A2(_07172_),
    .A1(_07080_),
    .B1(_07176_),
    .X(_02672_));
 sg13g2_buf_1 _26234_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07177_));
 sg13g2_nor2b_1 _26235_ (.A(_07110_),
    .B_N(net1103),
    .Y(_07178_));
 sg13g2_inv_1 _26236_ (.Y(_07179_),
    .A(_07110_));
 sg13g2_nor2_1 _26237_ (.A(net1103),
    .B(_07179_),
    .Y(_07180_));
 sg13g2_inv_1 _26238_ (.Y(_07181_),
    .A(_07099_));
 sg13g2_nand2_1 _26239_ (.Y(_07182_),
    .A(_07119_),
    .B(_07181_));
 sg13g2_nor3_1 _26240_ (.A(_07178_),
    .B(_07180_),
    .C(_07182_),
    .Y(_07183_));
 sg13g2_nand2_2 _26241_ (.Y(_07184_),
    .A(net1104),
    .B(_07178_));
 sg13g2_nand2_1 _26242_ (.Y(_07185_),
    .A(net1066),
    .B(_07184_));
 sg13g2_nor2_1 _26243_ (.A(_07183_),
    .B(_07185_),
    .Y(_07186_));
 sg13g2_nand2_1 _26244_ (.Y(_07187_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07128_));
 sg13g2_xor2_1 _26245_ (.B(_07187_),
    .A(\cpu.uart.r_x_invert ),
    .X(_07188_));
 sg13g2_nor2_1 _26246_ (.A(_00282_),
    .B(_07186_),
    .Y(_07189_));
 sg13g2_a21oi_1 _26247_ (.A1(_07186_),
    .A2(_07188_),
    .Y(_07190_),
    .B1(_07189_));
 sg13g2_nor3_2 _26248_ (.A(_07181_),
    .B(_07106_),
    .C(_07184_),
    .Y(_07191_));
 sg13g2_nand2_1 _26249_ (.Y(_07192_),
    .A(net1103),
    .B(net938));
 sg13g2_o21ai_1 _26250_ (.B1(_07192_),
    .Y(_07193_),
    .A1(net1103),
    .A2(_09954_));
 sg13g2_nand2b_1 _26251_ (.Y(_07194_),
    .B(_07126_),
    .A_N(_07117_));
 sg13g2_o21ai_1 _26252_ (.B1(_07194_),
    .Y(_07195_),
    .A1(_07119_),
    .A2(_07179_));
 sg13g2_a21oi_1 _26253_ (.A1(_07098_),
    .A2(_07113_),
    .Y(_07196_),
    .B1(_07180_));
 sg13g2_nor2_1 _26254_ (.A(_07117_),
    .B(_07196_),
    .Y(_07197_));
 sg13g2_a221oi_1 _26255_ (.B2(_07101_),
    .C1(_07197_),
    .B1(_07195_),
    .A1(_07100_),
    .Y(_07198_),
    .A2(_07193_));
 sg13g2_inv_1 _26256_ (.Y(_07199_),
    .A(_07198_));
 sg13g2_o21ai_1 _26257_ (.B1(net916),
    .Y(_07200_),
    .A1(_07191_),
    .A2(_07199_));
 sg13g2_mux2_1 _26258_ (.A0(_07177_),
    .A1(_07190_),
    .S(_07200_),
    .X(_02677_));
 sg13g2_nor4_2 _26259_ (.A(net1104),
    .B(_07100_),
    .C(_07102_),
    .Y(_07201_),
    .D(_07111_));
 sg13g2_a21oi_1 _26260_ (.A1(_07099_),
    .A2(_07115_),
    .Y(_07202_),
    .B1(net938));
 sg13g2_o21ai_1 _26261_ (.B1(net938),
    .Y(_07203_),
    .A1(_07099_),
    .A2(_07115_));
 sg13g2_o21ai_1 _26262_ (.B1(_07203_),
    .Y(_07204_),
    .A1(_07119_),
    .A2(_07202_));
 sg13g2_nand2_1 _26263_ (.Y(_07205_),
    .A(net939),
    .B(_07204_));
 sg13g2_nand3b_1 _26264_ (.B(net1066),
    .C(_07205_),
    .Y(_07206_),
    .A_N(_07201_));
 sg13g2_nor3_1 _26265_ (.A(_07152_),
    .B(_07191_),
    .C(_07206_),
    .Y(_07207_));
 sg13g2_and2_1 _26266_ (.A(net939),
    .B(net938),
    .X(_07208_));
 sg13g2_a22oi_1 _26267_ (.Y(_07209_),
    .B1(_07208_),
    .B2(_07182_),
    .A2(_07108_),
    .A1(_07179_));
 sg13g2_nand2_1 _26268_ (.Y(_07210_),
    .A(_07207_),
    .B(_07209_));
 sg13g2_nor2b_1 _26269_ (.A(_07114_),
    .B_N(_07207_),
    .Y(_07211_));
 sg13g2_a21oi_1 _26270_ (.A1(_07114_),
    .A2(_07210_),
    .Y(_07212_),
    .B1(_07211_));
 sg13g2_inv_1 _26271_ (.Y(_02680_),
    .A(_07212_));
 sg13g2_nand2_1 _26272_ (.Y(_07213_),
    .A(_07114_),
    .B(_07209_));
 sg13g2_nand2_1 _26273_ (.Y(_07214_),
    .A(_07207_),
    .B(_07213_));
 sg13g2_o21ai_1 _26274_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07215_),
    .A1(_07114_),
    .A2(_07210_));
 sg13g2_o21ai_1 _26275_ (.B1(_07215_),
    .Y(_02681_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07214_));
 sg13g2_nand2_1 _26276_ (.Y(_07216_),
    .A(net544),
    .B(net192));
 sg13g2_buf_1 _26277_ (.A(_07216_),
    .X(_07217_));
 sg13g2_buf_1 _26278_ (.A(net115),
    .X(_07218_));
 sg13g2_nand2_1 _26279_ (.Y(_07219_),
    .A(net193),
    .B(net384));
 sg13g2_buf_2 _26280_ (.A(_07219_),
    .X(_07220_));
 sg13g2_buf_1 _26281_ (.A(_07220_),
    .X(_07221_));
 sg13g2_buf_1 _26282_ (.A(_07220_),
    .X(_07222_));
 sg13g2_inv_1 _26283_ (.Y(_07223_),
    .A(_04885_));
 sg13g2_nand3_1 _26284_ (.B(_10241_),
    .C(_10236_),
    .A(_10234_),
    .Y(_07224_));
 sg13g2_buf_1 _26285_ (.A(_07224_),
    .X(_07225_));
 sg13g2_nor3_2 _26286_ (.A(_07223_),
    .B(_10200_),
    .C(_07225_),
    .Y(_07226_));
 sg13g2_nand2_1 _26287_ (.Y(_07227_),
    .A(net93),
    .B(_07226_));
 sg13g2_o21ai_1 _26288_ (.B1(_07227_),
    .Y(_07228_),
    .A1(_06794_),
    .A2(net94));
 sg13g2_nor2_1 _26289_ (.A(_10200_),
    .B(_07225_),
    .Y(_07229_));
 sg13g2_o21ai_1 _26290_ (.B1(net95),
    .Y(_07230_),
    .A1(net104),
    .A2(_07229_));
 sg13g2_a22oi_1 _26291_ (.Y(_02467_),
    .B1(_07230_),
    .B2(_07223_),
    .A2(_07228_),
    .A1(net95));
 sg13g2_and2_1 _26292_ (.A(_05361_),
    .B(_07226_),
    .X(_07231_));
 sg13g2_buf_1 _26293_ (.A(_07231_),
    .X(_07232_));
 sg13g2_nand2_1 _26294_ (.Y(_07233_),
    .A(net93),
    .B(_07232_));
 sg13g2_o21ai_1 _26295_ (.B1(_07233_),
    .Y(_07234_),
    .A1(net1049),
    .A2(net94));
 sg13g2_o21ai_1 _26296_ (.B1(net115),
    .Y(_07235_),
    .A1(net104),
    .A2(_07226_));
 sg13g2_inv_1 _26297_ (.Y(_07236_),
    .A(_05361_));
 sg13g2_a22oi_1 _26298_ (.Y(_02468_),
    .B1(_07235_),
    .B2(_07236_),
    .A2(_07234_),
    .A1(net95));
 sg13g2_nand3_1 _26299_ (.B(_07220_),
    .C(_07232_),
    .A(_05427_),
    .Y(_07237_));
 sg13g2_o21ai_1 _26300_ (.B1(_07237_),
    .Y(_07238_),
    .A1(net1048),
    .A2(net94));
 sg13g2_o21ai_1 _26301_ (.B1(net115),
    .Y(_07239_),
    .A1(net104),
    .A2(_07232_));
 sg13g2_inv_1 _26302_ (.Y(_07240_),
    .A(_05427_));
 sg13g2_a22oi_1 _26303_ (.Y(_02469_),
    .B1(_07239_),
    .B2(_07240_),
    .A2(_07238_),
    .A1(net95));
 sg13g2_inv_1 _26304_ (.Y(_07241_),
    .A(_05486_));
 sg13g2_nand4_1 _26305_ (.B(_05361_),
    .C(_05427_),
    .A(_04885_),
    .Y(_07242_),
    .D(_10185_));
 sg13g2_nor2_1 _26306_ (.A(_07225_),
    .B(_07242_),
    .Y(_07243_));
 sg13g2_o21ai_1 _26307_ (.B1(net115),
    .Y(_07244_),
    .A1(net103),
    .A2(_07243_));
 sg13g2_nor3_1 _26308_ (.A(_07241_),
    .B(_07225_),
    .C(_07242_),
    .Y(_07245_));
 sg13g2_nand2_1 _26309_ (.Y(_07246_),
    .A(net93),
    .B(_07245_));
 sg13g2_o21ai_1 _26310_ (.B1(_07246_),
    .Y(_07247_),
    .A1(net1054),
    .A2(net94));
 sg13g2_a22oi_1 _26311_ (.Y(_02470_),
    .B1(_07247_),
    .B2(net95),
    .A2(_07244_),
    .A1(_07241_));
 sg13g2_nand3_1 _26312_ (.B(_05486_),
    .C(_07232_),
    .A(_05427_),
    .Y(_07248_));
 sg13g2_nor3_1 _26313_ (.A(_05558_),
    .B(net134),
    .C(_07248_),
    .Y(_07249_));
 sg13g2_a21oi_1 _26314_ (.A1(_10117_),
    .A2(net103),
    .Y(_07250_),
    .B1(_07249_));
 sg13g2_a21oi_1 _26315_ (.A1(net93),
    .A2(_07248_),
    .Y(_07251_),
    .B1(net136));
 sg13g2_nand2b_1 _26316_ (.Y(_07252_),
    .B(_05558_),
    .A_N(_07251_));
 sg13g2_o21ai_1 _26317_ (.B1(_07252_),
    .Y(_02471_),
    .A1(net105),
    .A2(_07250_));
 sg13g2_nand2_1 _26318_ (.Y(_07253_),
    .A(_05558_),
    .B(_07245_));
 sg13g2_nor3_1 _26319_ (.A(_05606_),
    .B(net134),
    .C(_07253_),
    .Y(_07254_));
 sg13g2_a21oi_1 _26320_ (.A1(net1052),
    .A2(net103),
    .Y(_07255_),
    .B1(_07254_));
 sg13g2_and2_1 _26321_ (.A(_07220_),
    .B(_07253_),
    .X(_07256_));
 sg13g2_o21ai_1 _26322_ (.B1(_05606_),
    .Y(_07257_),
    .A1(net135),
    .A2(_07256_));
 sg13g2_o21ai_1 _26323_ (.B1(_07257_),
    .Y(_02472_),
    .A1(net105),
    .A2(_07255_));
 sg13g2_nand3_1 _26324_ (.B(_05427_),
    .C(_07226_),
    .A(_05361_),
    .Y(_07258_));
 sg13g2_nand3_1 _26325_ (.B(_05558_),
    .C(_05606_),
    .A(_05486_),
    .Y(_07259_));
 sg13g2_nor2_1 _26326_ (.A(_07258_),
    .B(_07259_),
    .Y(_07260_));
 sg13g2_nand3_1 _26327_ (.B(_07220_),
    .C(_07260_),
    .A(_05710_),
    .Y(_07261_));
 sg13g2_o21ai_1 _26328_ (.B1(_07261_),
    .Y(_07262_),
    .A1(_10129_),
    .A2(net94));
 sg13g2_o21ai_1 _26329_ (.B1(net115),
    .Y(_07263_),
    .A1(net104),
    .A2(_07260_));
 sg13g2_inv_1 _26330_ (.Y(_07264_),
    .A(_05710_));
 sg13g2_a22oi_1 _26331_ (.Y(_02473_),
    .B1(_07263_),
    .B2(_07264_),
    .A2(_07262_),
    .A1(net95));
 sg13g2_nand4_1 _26332_ (.B(_05606_),
    .C(_05710_),
    .A(_05558_),
    .Y(_07265_),
    .D(_07245_));
 sg13g2_buf_1 _26333_ (.A(_07265_),
    .X(_07266_));
 sg13g2_nor3_1 _26334_ (.A(_05122_),
    .B(net134),
    .C(_07266_),
    .Y(_07267_));
 sg13g2_a21oi_1 _26335_ (.A1(net1050),
    .A2(net103),
    .Y(_07268_),
    .B1(_07267_));
 sg13g2_a21oi_1 _26336_ (.A1(_07220_),
    .A2(_07266_),
    .Y(_07269_),
    .B1(_10148_));
 sg13g2_nand2b_1 _26337_ (.Y(_07270_),
    .B(_05122_),
    .A_N(_07269_));
 sg13g2_o21ai_1 _26338_ (.B1(_07270_),
    .Y(_02474_),
    .A1(net105),
    .A2(_07268_));
 sg13g2_nand3_1 _26339_ (.B(_05122_),
    .C(_07260_),
    .A(_05710_),
    .Y(_07271_));
 sg13g2_buf_1 _26340_ (.A(_07271_),
    .X(_07272_));
 sg13g2_nor2_1 _26341_ (.A(_05732_),
    .B(_07272_),
    .Y(_07273_));
 sg13g2_nand2_1 _26342_ (.Y(_07274_),
    .A(net93),
    .B(_07273_));
 sg13g2_o21ai_1 _26343_ (.B1(_07274_),
    .Y(_07275_),
    .A1(_10205_),
    .A2(net94));
 sg13g2_a21o_1 _26344_ (.A2(_07272_),
    .A1(net93),
    .B1(net135),
    .X(_07276_));
 sg13g2_a22oi_1 _26345_ (.Y(_02475_),
    .B1(_07276_),
    .B2(_05732_),
    .A2(_07275_),
    .A1(net95));
 sg13g2_inv_1 _26346_ (.Y(_07277_),
    .A(_05751_));
 sg13g2_nor3_1 _26347_ (.A(_05732_),
    .B(_07277_),
    .C(_07272_),
    .Y(_07278_));
 sg13g2_nand2_1 _26348_ (.Y(_07279_),
    .A(net93),
    .B(_07278_));
 sg13g2_o21ai_1 _26349_ (.B1(_07279_),
    .Y(_07280_),
    .A1(_10210_),
    .A2(net94));
 sg13g2_o21ai_1 _26350_ (.B1(net115),
    .Y(_07281_),
    .A1(_10159_),
    .A2(_07273_));
 sg13g2_a22oi_1 _26351_ (.Y(_02476_),
    .B1(_07281_),
    .B2(_07277_),
    .A2(_07280_),
    .A1(net95));
 sg13g2_nand2_1 _26352_ (.Y(_07282_),
    .A(_05020_),
    .B(_07278_));
 sg13g2_inv_1 _26353_ (.Y(_07283_),
    .A(_07282_));
 sg13g2_nand2_1 _26354_ (.Y(_07284_),
    .A(net93),
    .B(_07283_));
 sg13g2_o21ai_1 _26355_ (.B1(_07284_),
    .Y(_07285_),
    .A1(_10215_),
    .A2(net94));
 sg13g2_o21ai_1 _26356_ (.B1(net115),
    .Y(_07286_),
    .A1(_10159_),
    .A2(_07278_));
 sg13g2_a22oi_1 _26357_ (.Y(_02477_),
    .B1(_07286_),
    .B2(_05021_),
    .A2(_07285_),
    .A1(_07218_));
 sg13g2_nand4_1 _26358_ (.B(\cpu.intr.r_clock_count[24] ),
    .C(_05751_),
    .A(_05122_),
    .Y(_07287_),
    .D(_05020_));
 sg13g2_or2_1 _26359_ (.X(_07288_),
    .B(_07287_),
    .A(_07266_));
 sg13g2_buf_1 _26360_ (.A(_07288_),
    .X(_07289_));
 sg13g2_nor3_1 _26361_ (.A(_05171_),
    .B(net134),
    .C(_07289_),
    .Y(_07290_));
 sg13g2_a21oi_1 _26362_ (.A1(_10222_),
    .A2(net103),
    .Y(_07291_),
    .B1(_07290_));
 sg13g2_a21oi_1 _26363_ (.A1(_07220_),
    .A2(_07289_),
    .Y(_07292_),
    .B1(_10147_));
 sg13g2_nand2b_1 _26364_ (.Y(_07293_),
    .B(_05171_),
    .A_N(_07292_));
 sg13g2_o21ai_1 _26365_ (.B1(_07293_),
    .Y(_02478_),
    .A1(net105),
    .A2(_07291_));
 sg13g2_inv_1 _26366_ (.Y(_07294_),
    .A(_05171_));
 sg13g2_nor4_1 _26367_ (.A(_07294_),
    .B(_05186_),
    .C(net134),
    .D(_07282_),
    .Y(_07295_));
 sg13g2_a21oi_1 _26368_ (.A1(_10227_),
    .A2(_10142_),
    .Y(_07296_),
    .B1(_07295_));
 sg13g2_a21oi_1 _26369_ (.A1(_05171_),
    .A2(_07283_),
    .Y(_07297_),
    .B1(net134));
 sg13g2_o21ai_1 _26370_ (.B1(_05186_),
    .Y(_07298_),
    .A1(_10150_),
    .A2(_07297_));
 sg13g2_o21ai_1 _26371_ (.B1(_07298_),
    .Y(_02479_),
    .A1(net105),
    .A2(_07296_));
 sg13g2_nand3_1 _26372_ (.B(_05186_),
    .C(_05214_),
    .A(_05171_),
    .Y(_07299_));
 sg13g2_buf_1 _26373_ (.A(_07299_),
    .X(_07300_));
 sg13g2_nor2_1 _26374_ (.A(_07289_),
    .B(_07300_),
    .Y(_07301_));
 sg13g2_nand2_1 _26375_ (.Y(_07302_),
    .A(_07222_),
    .B(_07301_));
 sg13g2_o21ai_1 _26376_ (.B1(_07302_),
    .Y(_07303_),
    .A1(_10229_),
    .A2(_07221_));
 sg13g2_nand2_1 _26377_ (.Y(_07304_),
    .A(_05171_),
    .B(_05186_));
 sg13g2_o21ai_1 _26378_ (.B1(_07222_),
    .Y(_07305_),
    .A1(_07289_),
    .A2(_07304_));
 sg13g2_a21oi_1 _26379_ (.A1(net115),
    .A2(_07305_),
    .Y(_07306_),
    .B1(_05214_));
 sg13g2_a21oi_1 _26380_ (.A1(_07218_),
    .A2(_07303_),
    .Y(_02480_),
    .B1(_07306_));
 sg13g2_nor3_1 _26381_ (.A(_05262_),
    .B(_07282_),
    .C(_07300_),
    .Y(_07307_));
 sg13g2_a22oi_1 _26382_ (.Y(_07308_),
    .B1(_07221_),
    .B2(_07307_),
    .A2(_10142_),
    .A1(_10239_));
 sg13g2_o21ai_1 _26383_ (.B1(_07220_),
    .Y(_07309_),
    .A1(_07282_),
    .A2(_07300_));
 sg13g2_nand2_1 _26384_ (.Y(_07310_),
    .A(_07217_),
    .B(_07309_));
 sg13g2_nand2_1 _26385_ (.Y(_07311_),
    .A(_05262_),
    .B(_07310_));
 sg13g2_o21ai_1 _26386_ (.B1(_07311_),
    .Y(_02481_),
    .A1(_10149_),
    .A2(_07308_));
 sg13g2_nand2_1 _26387_ (.Y(_07312_),
    .A(_05262_),
    .B(_07301_));
 sg13g2_nor3_1 _26388_ (.A(_05276_),
    .B(_10158_),
    .C(_07312_),
    .Y(_07313_));
 sg13g2_a21oi_1 _26389_ (.A1(_10244_),
    .A2(_10182_),
    .Y(_07314_),
    .B1(_07313_));
 sg13g2_nor2b_1 _26390_ (.A(net192),
    .B_N(_07312_),
    .Y(_07315_));
 sg13g2_o21ai_1 _26391_ (.B1(_05276_),
    .Y(_07316_),
    .A1(_10150_),
    .A2(_07315_));
 sg13g2_o21ai_1 _26392_ (.B1(_07316_),
    .Y(_02482_),
    .A1(_10149_),
    .A2(_07314_));
 sg13g2_nor2_1 _26393_ (.A(\cpu.r_clk_invert ),
    .B(net691),
    .Y(_07317_));
 sg13g2_a21oi_1 _26394_ (.A1(_09252_),
    .A2(net682),
    .Y(_02549_),
    .B1(_07317_));
 sg13g2_nand2b_1 _26395_ (.Y(_07318_),
    .B(_09308_),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26396_ (.A(_07318_),
    .X(_07319_));
 sg13g2_nor2b_1 _26397_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net534),
    .Y(_07320_));
 sg13g2_nand3_1 _26398_ (.B(_03000_),
    .C(_03007_),
    .A(_09398_),
    .Y(_07321_));
 sg13g2_buf_2 _26399_ (.A(_07321_),
    .X(_07322_));
 sg13g2_nor2_1 _26400_ (.A(net659),
    .B(_07322_),
    .Y(_07323_));
 sg13g2_nor3_1 _26401_ (.A(_07319_),
    .B(_07320_),
    .C(_07323_),
    .Y(_00743_));
 sg13g2_nor2_1 _26402_ (.A(\cpu.dcache.r_valid[1] ),
    .B(_12293_),
    .Y(_07324_));
 sg13g2_nor2_1 _26403_ (.A(net658),
    .B(_07322_),
    .Y(_07325_));
 sg13g2_nor3_1 _26404_ (.A(_07319_),
    .B(_07324_),
    .C(_07325_),
    .Y(_00744_));
 sg13g2_nor2_1 _26405_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net421),
    .Y(_07326_));
 sg13g2_nor2_1 _26406_ (.A(net532),
    .B(_07322_),
    .Y(_07327_));
 sg13g2_nor3_1 _26407_ (.A(_07319_),
    .B(_07326_),
    .C(_07327_),
    .Y(_00745_));
 sg13g2_nor2_1 _26408_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net419),
    .Y(_07328_));
 sg13g2_nor2_1 _26409_ (.A(net531),
    .B(_07322_),
    .Y(_07329_));
 sg13g2_nor3_1 _26410_ (.A(_07319_),
    .B(_07328_),
    .C(_07329_),
    .Y(_00746_));
 sg13g2_inv_1 _26411_ (.Y(_07330_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _26412_ (.Y(_07331_),
    .A(_07322_));
 sg13g2_a221oi_1 _26413_ (.B2(net424),
    .C1(_07319_),
    .B1(_07331_),
    .A1(_07330_),
    .Y(_00747_),
    .A2(net259));
 sg13g2_nor2_1 _26414_ (.A(\cpu.dcache.r_valid[5] ),
    .B(net417),
    .Y(_07332_));
 sg13g2_nor2_1 _26415_ (.A(net528),
    .B(_07322_),
    .Y(_07333_));
 sg13g2_nor3_1 _26416_ (.A(_07319_),
    .B(_07332_),
    .C(_07333_),
    .Y(_00748_));
 sg13g2_nor2_1 _26417_ (.A(\cpu.dcache.r_valid[6] ),
    .B(net464),
    .Y(_07334_));
 sg13g2_nor2_1 _26418_ (.A(net593),
    .B(_07322_),
    .Y(_07335_));
 sg13g2_nor3_1 _26419_ (.A(_07319_),
    .B(_07334_),
    .C(_07335_),
    .Y(_00749_));
 sg13g2_nor2_1 _26420_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net382),
    .Y(_07336_));
 sg13g2_nor2_1 _26421_ (.A(net469),
    .B(_07322_),
    .Y(_07337_));
 sg13g2_nor3_1 _26422_ (.A(_07319_),
    .B(_07336_),
    .C(_07337_),
    .Y(_00750_));
 sg13g2_nor2_1 _26423_ (.A(net1131),
    .B(net1046),
    .Y(_07338_));
 sg13g2_nand3_1 _26424_ (.B(_07338_),
    .C(_04748_),
    .A(_10262_),
    .Y(_07339_));
 sg13g2_buf_1 _26425_ (.A(_07339_),
    .X(_07340_));
 sg13g2_nand2_1 _26426_ (.Y(_07341_),
    .A(_08311_),
    .B(net566));
 sg13g2_o21ai_1 _26427_ (.B1(_07341_),
    .Y(_07342_),
    .A1(_03788_),
    .A2(net566));
 sg13g2_and3_1 _26428_ (.X(_00799_),
    .A(net210),
    .B(_09309_),
    .C(_07342_));
 sg13g2_and4_1 _26429_ (.A(net734),
    .B(_11088_),
    .C(\cpu.dec.do_flush_all ),
    .D(_11580_),
    .X(_00932_));
 sg13g2_and4_1 _26430_ (.A(net734),
    .B(_11051_),
    .C(\cpu.dec.do_flush_all ),
    .D(net751),
    .X(_00950_));
 sg13g2_o21ai_1 _26431_ (.B1(net210),
    .Y(_07343_),
    .A1(_11943_),
    .A2(_10674_));
 sg13g2_nand2_1 _26432_ (.Y(_07344_),
    .A(net827),
    .B(_11943_));
 sg13g2_nand4_1 _26433_ (.B(_04091_),
    .C(net751),
    .A(net734),
    .Y(_07345_),
    .D(_10457_));
 sg13g2_mux2_1 _26434_ (.A0(_11022_),
    .A1(_09243_),
    .S(_07345_),
    .X(_07346_));
 sg13g2_o21ai_1 _26435_ (.B1(net797),
    .Y(_07347_),
    .A1(_03518_),
    .A2(net566));
 sg13g2_a221oi_1 _26436_ (.B2(net566),
    .C1(_07347_),
    .B1(_07346_),
    .A1(_07343_),
    .Y(_00951_),
    .A2(_07344_));
 sg13g2_or2_1 _26437_ (.X(_07348_),
    .B(_04792_),
    .A(_11594_));
 sg13g2_inv_1 _26438_ (.Y(_07349_),
    .A(_04816_));
 sg13g2_nor3_1 _26439_ (.A(_08352_),
    .B(_00300_),
    .C(_07349_),
    .Y(_07350_));
 sg13g2_nor4_2 _26440_ (.A(_08351_),
    .B(_08352_),
    .C(_00312_),
    .Y(_07351_),
    .D(_11943_));
 sg13g2_a22oi_1 _26441_ (.Y(_07352_),
    .B1(_12074_),
    .B2(_09307_),
    .A2(_09827_),
    .A1(_09398_));
 sg13g2_a21o_1 _26442_ (.A2(_07352_),
    .A1(_11614_),
    .B1(_08354_),
    .X(_07353_));
 sg13g2_and2_1 _26443_ (.A(_09307_),
    .B(_07353_),
    .X(_07354_));
 sg13g2_buf_1 _26444_ (.A(_07354_),
    .X(_07355_));
 sg13g2_o21ai_1 _26445_ (.B1(_07355_),
    .Y(_07356_),
    .A1(net1154),
    .A2(_07351_));
 sg13g2_a21oi_1 _26446_ (.A1(_07348_),
    .A2(_07350_),
    .Y(_01070_),
    .B1(_07356_));
 sg13g2_nand3_1 _26447_ (.B(_07355_),
    .C(_07351_),
    .A(_04816_),
    .Y(_07357_));
 sg13g2_a22oi_1 _26448_ (.Y(_07358_),
    .B1(_07351_),
    .B2(_11599_),
    .A2(_07355_),
    .A1(_08351_));
 sg13g2_o21ai_1 _26449_ (.B1(_07358_),
    .Y(_01071_),
    .A1(_04793_),
    .A2(_07357_));
 sg13g2_inv_1 _26450_ (.Y(_07359_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26451_ (.Y(_07360_),
    .B(_09308_),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26452_ (.A(_07360_),
    .X(_07361_));
 sg13g2_a21oi_1 _26453_ (.A1(_07359_),
    .A2(_06546_),
    .Y(_02426_),
    .B1(_07361_));
 sg13g2_nor2_1 _26454_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06457_),
    .Y(_07362_));
 sg13g2_nor2_1 _26455_ (.A(_07361_),
    .B(_07362_),
    .Y(_02427_));
 sg13g2_nor2_1 _26456_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06473_),
    .Y(_07363_));
 sg13g2_nor2_1 _26457_ (.A(_07361_),
    .B(_07363_),
    .Y(_02428_));
 sg13g2_inv_1 _26458_ (.Y(_07364_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26459_ (.A1(_07364_),
    .A2(_06608_),
    .Y(_02429_),
    .B1(_07361_));
 sg13g2_nor2_1 _26460_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06505_),
    .Y(_07365_));
 sg13g2_nor2_1 _26461_ (.A(_07361_),
    .B(_07365_),
    .Y(_02430_));
 sg13g2_inv_1 _26462_ (.Y(_07366_),
    .A(\cpu.icache.r_valid[5] ));
 sg13g2_a21oi_1 _26463_ (.A1(_07366_),
    .A2(_06518_),
    .Y(_02431_),
    .B1(_07361_));
 sg13g2_inv_1 _26464_ (.Y(_07367_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26465_ (.A1(_07367_),
    .A2(_06527_),
    .Y(_02432_),
    .B1(_07361_));
 sg13g2_nor2_1 _26466_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06541_),
    .Y(_07368_));
 sg13g2_nor2_1 _26467_ (.A(_07361_),
    .B(_07368_),
    .Y(_02433_));
 sg13g2_nand3_1 _26468_ (.B(_10032_),
    .C(net411),
    .A(net1133),
    .Y(_07369_));
 sg13g2_and2_1 _26469_ (.A(net193),
    .B(_04925_),
    .X(_07370_));
 sg13g2_buf_1 _26470_ (.A(_07370_),
    .X(_07371_));
 sg13g2_a22oi_1 _26471_ (.Y(_07372_),
    .B1(_07371_),
    .B2(net1000),
    .A2(_07369_),
    .A1(_09272_));
 sg13g2_nor2_1 _26472_ (.A(net614),
    .B(_07372_),
    .Y(_00319_));
 sg13g2_nor2_1 _26473_ (.A(_03000_),
    .B(_12055_),
    .Y(_07373_));
 sg13g2_nor2b_1 _26474_ (.A(_07373_),
    .B_N(_00317_),
    .Y(_00588_));
 sg13g2_a21oi_1 _26475_ (.A1(_12063_),
    .A2(_12109_),
    .Y(_00589_),
    .B1(_07373_));
 sg13g2_nand2b_1 _26476_ (.Y(_07374_),
    .B(_12070_),
    .A_N(net1027));
 sg13g2_a21oi_1 _26477_ (.A1(_06825_),
    .A2(_07374_),
    .Y(_00590_),
    .B1(_07373_));
 sg13g2_nor2_1 _26478_ (.A(_09314_),
    .B(net566),
    .Y(_07375_));
 sg13g2_a21oi_1 _26479_ (.A1(net1083),
    .A2(net566),
    .Y(_07376_),
    .B1(_07375_));
 sg13g2_nor2_1 _26480_ (.A(net614),
    .B(_07376_),
    .Y(_00800_));
 sg13g2_nand3_1 _26481_ (.B(net751),
    .C(_04216_),
    .A(net1152),
    .Y(_07377_));
 sg13g2_nand2_1 _26482_ (.Y(_07378_),
    .A(_11596_),
    .B(_07377_));
 sg13g2_nand2_1 _26483_ (.Y(_07379_),
    .A(net734),
    .B(_07378_));
 sg13g2_nor2_1 _26484_ (.A(_10649_),
    .B(_09376_),
    .Y(_07380_));
 sg13g2_nand3_1 _26485_ (.B(_10457_),
    .C(_07380_),
    .A(_04091_),
    .Y(_07381_));
 sg13g2_a21oi_1 _26486_ (.A1(net734),
    .A2(_07381_),
    .Y(_07382_),
    .B1(_09304_));
 sg13g2_nor2_1 _26487_ (.A(_03772_),
    .B(_07382_),
    .Y(_07383_));
 sg13g2_nor2_1 _26488_ (.A(_10649_),
    .B(_07383_),
    .Y(_07384_));
 sg13g2_a21oi_1 _26489_ (.A1(_10645_),
    .A2(_07383_),
    .Y(_07385_),
    .B1(_07384_));
 sg13g2_nand2b_1 _26490_ (.Y(_07386_),
    .B(_07385_),
    .A_N(_07378_));
 sg13g2_nand3_1 _26491_ (.B(_07379_),
    .C(_07386_),
    .A(_05808_),
    .Y(_00801_));
 sg13g2_mux2_1 _26492_ (.A0(net1069),
    .A1(_10721_),
    .S(net566),
    .X(_07387_));
 sg13g2_and2_1 _26493_ (.A(_09310_),
    .B(_07387_),
    .X(_00802_));
 sg13g2_nor3_1 _26494_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11595_),
    .C(_03476_),
    .Y(_07388_));
 sg13g2_nand3_1 _26495_ (.B(net751),
    .C(_07388_),
    .A(_08354_),
    .Y(_07389_));
 sg13g2_nand3_1 _26496_ (.B(_07353_),
    .C(_07389_),
    .A(_10252_),
    .Y(_07390_));
 sg13g2_nand3_1 _26497_ (.B(_11597_),
    .C(_07390_),
    .A(_08400_),
    .Y(_07391_));
 sg13g2_nand3_1 _26498_ (.B(_05292_),
    .C(_07391_),
    .A(_06852_),
    .Y(_07392_));
 sg13g2_o21ai_1 _26499_ (.B1(_07392_),
    .Y(_07393_),
    .A1(_06852_),
    .A2(net141));
 sg13g2_nand2_1 _26500_ (.Y(_00948_),
    .A(_05838_),
    .B(_07393_));
 sg13g2_nand2_1 _26501_ (.Y(_07394_),
    .A(_09398_),
    .B(_09376_));
 sg13g2_nand3_1 _26502_ (.B(\cpu.dec.do_flush_write ),
    .C(_11941_),
    .A(net734),
    .Y(_07395_));
 sg13g2_a21oi_1 _26503_ (.A1(_07394_),
    .A2(_07395_),
    .Y(_00949_),
    .B1(_06789_));
 sg13g2_nand2_1 _26504_ (.Y(_07396_),
    .A(\cpu.dec.io ),
    .B(_11941_));
 sg13g2_nand2_1 _26505_ (.Y(_07397_),
    .A(_04822_),
    .B(_09376_));
 sg13g2_a21oi_1 _26506_ (.A1(_07396_),
    .A2(_07397_),
    .Y(_00952_),
    .B1(_06789_));
 sg13g2_and2_1 _26507_ (.A(_09243_),
    .B(_07378_),
    .X(_07398_));
 sg13g2_nand2_1 _26508_ (.Y(_07399_),
    .A(\cpu.ex.r_prev_ie ),
    .B(net566));
 sg13g2_o21ai_1 _26509_ (.B1(_07399_),
    .Y(_07400_),
    .A1(_10094_),
    .A2(_07340_));
 sg13g2_nor2_1 _26510_ (.A(_07378_),
    .B(_07400_),
    .Y(_07401_));
 sg13g2_nor3_1 _26511_ (.A(_09365_),
    .B(_07398_),
    .C(_07401_),
    .Y(_00999_));
 sg13g2_a22oi_1 _26512_ (.Y(_07402_),
    .B1(_11615_),
    .B2(net1092),
    .A2(_11941_),
    .A1(_11595_));
 sg13g2_nor2_1 _26513_ (.A(net614),
    .B(_07402_),
    .Y(_01000_));
 sg13g2_and2_1 _26514_ (.A(_10645_),
    .B(_05818_),
    .X(_07403_));
 sg13g2_buf_1 _26515_ (.A(_07403_),
    .X(_07404_));
 sg13g2_mux2_1 _26516_ (.A0(_10503_),
    .A1(_09223_),
    .S(_07404_),
    .X(_07405_));
 sg13g2_nand2_1 _26517_ (.Y(_07406_),
    .A(net210),
    .B(_07405_));
 sg13g2_a21oi_1 _26518_ (.A1(_11596_),
    .A2(_07406_),
    .Y(_01076_),
    .B1(net567));
 sg13g2_nand2_1 _26519_ (.Y(_07407_),
    .A(_03532_),
    .B(_07404_));
 sg13g2_o21ai_1 _26520_ (.B1(_07407_),
    .Y(_07408_),
    .A1(_10420_),
    .A2(_07404_));
 sg13g2_nor2_1 _26521_ (.A(net687),
    .B(net210),
    .Y(_07409_));
 sg13g2_a21oi_1 _26522_ (.A1(_05809_),
    .A2(_07408_),
    .Y(_07410_),
    .B1(_07409_));
 sg13g2_nor2_1 _26523_ (.A(net614),
    .B(_07410_),
    .Y(_01077_));
 sg13g2_mux2_1 _26524_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_10137_),
    .S(_07404_),
    .X(_07411_));
 sg13g2_a21oi_1 _26525_ (.A1(_08359_),
    .A2(_07411_),
    .Y(_07412_),
    .B1(_08454_));
 sg13g2_nor2_1 _26526_ (.A(net614),
    .B(_07412_),
    .Y(_01078_));
 sg13g2_nor2b_1 _26527_ (.A(_00259_),
    .B_N(_05816_),
    .Y(_07413_));
 sg13g2_o21ai_1 _26528_ (.B1(_07413_),
    .Y(_07414_),
    .A1(_10645_),
    .A2(_00257_));
 sg13g2_a21o_1 _26529_ (.A2(_07414_),
    .A1(_05815_),
    .B1(_08457_),
    .X(_07415_));
 sg13g2_buf_1 _26530_ (.A(_07415_),
    .X(_07416_));
 sg13g2_nand2b_1 _26531_ (.Y(_07417_),
    .B(_05815_),
    .A_N(_07416_));
 sg13g2_buf_1 _26532_ (.A(_07417_),
    .X(_07418_));
 sg13g2_buf_1 _26533_ (.A(_07418_),
    .X(_07419_));
 sg13g2_nor2_2 _26534_ (.A(net1126),
    .B(_10872_),
    .Y(_07420_));
 sg13g2_nand2_1 _26535_ (.Y(_07421_),
    .A(_00290_),
    .B(_07420_));
 sg13g2_nor4_2 _26536_ (.A(net974),
    .B(net982),
    .C(net978),
    .Y(_07422_),
    .D(_07421_));
 sg13g2_a21oi_1 _26537_ (.A1(_03356_),
    .A2(_11088_),
    .Y(_07423_),
    .B1(_05815_));
 sg13g2_nor2_1 _26538_ (.A(_07416_),
    .B(_07423_),
    .Y(_07424_));
 sg13g2_buf_2 _26539_ (.A(_07424_),
    .X(_07425_));
 sg13g2_o21ai_1 _26540_ (.B1(_07425_),
    .Y(_07426_),
    .A1(net92),
    .A2(_07422_));
 sg13g2_and3_1 _26541_ (.X(_07427_),
    .A(_10137_),
    .B(net980),
    .C(_07422_));
 sg13g2_nor2_1 _26542_ (.A(_11051_),
    .B(_05813_),
    .Y(_07428_));
 sg13g2_nor2b_1 _26543_ (.A(_07428_),
    .B_N(_03356_),
    .Y(_07429_));
 sg13g2_buf_1 _26544_ (.A(_07429_),
    .X(_07430_));
 sg13g2_nor2_1 _26545_ (.A(_07430_),
    .B(_07416_),
    .Y(_07431_));
 sg13g2_a22oi_1 _26546_ (.Y(_07432_),
    .B1(_07427_),
    .B2(_07431_),
    .A2(_07426_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26547_ (.A(_09850_),
    .B(_07432_),
    .Y(_01079_));
 sg13g2_nor3_1 _26548_ (.A(net844),
    .B(_05293_),
    .C(net727),
    .Y(_07433_));
 sg13g2_buf_2 _26549_ (.A(_07433_),
    .X(_07434_));
 sg13g2_nor2_1 _26550_ (.A(_10308_),
    .B(_07421_),
    .Y(_07435_));
 sg13g2_a21oi_1 _26551_ (.A1(net1107),
    .A2(_07420_),
    .Y(_07436_),
    .B1(_05851_));
 sg13g2_a21o_1 _26552_ (.A2(_07435_),
    .A1(net982),
    .B1(_07436_),
    .X(_07437_));
 sg13g2_a22oi_1 _26553_ (.Y(_07438_),
    .B1(_07437_),
    .B2(_10420_),
    .A2(_07435_),
    .A1(_05926_));
 sg13g2_buf_2 _26554_ (.A(_07438_),
    .X(_07439_));
 sg13g2_nor2_2 _26555_ (.A(net92),
    .B(_07439_),
    .Y(_07440_));
 sg13g2_buf_1 _26556_ (.A(_07418_),
    .X(_07441_));
 sg13g2_buf_1 _26557_ (.A(_07425_),
    .X(_07442_));
 sg13g2_o21ai_1 _26558_ (.B1(net90),
    .Y(_07443_),
    .A1(_05881_),
    .A2(net91));
 sg13g2_a22oi_1 _26559_ (.Y(_07444_),
    .B1(_07443_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07440_),
    .A1(_07434_));
 sg13g2_nor2_1 _26560_ (.A(_09850_),
    .B(_07444_),
    .Y(_01080_));
 sg13g2_buf_1 _26561_ (.A(_09363_),
    .X(_07445_));
 sg13g2_buf_1 _26562_ (.A(_07445_),
    .X(_07446_));
 sg13g2_o21ai_1 _26563_ (.B1(_07425_),
    .Y(_07447_),
    .A1(_05889_),
    .A2(net92));
 sg13g2_nor2_1 _26564_ (.A(_10094_),
    .B(_07418_),
    .Y(_07448_));
 sg13g2_buf_2 _26565_ (.A(_07448_),
    .X(_07449_));
 sg13g2_buf_1 _26566_ (.A(_07449_),
    .X(_07450_));
 sg13g2_a22oi_1 _26567_ (.Y(_07451_),
    .B1(_07450_),
    .B2(_05889_),
    .A2(_07447_),
    .A1(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_nor2_1 _26568_ (.A(_07446_),
    .B(_07451_),
    .Y(_01081_));
 sg13g2_nand2_1 _26569_ (.Y(_07452_),
    .A(net981),
    .B(_04992_));
 sg13g2_nor3_1 _26570_ (.A(_05832_),
    .B(net1126),
    .C(_07452_),
    .Y(_07453_));
 sg13g2_buf_2 _26571_ (.A(_07453_),
    .X(_07454_));
 sg13g2_nor3_1 _26572_ (.A(_05832_),
    .B(net1126),
    .C(_05839_),
    .Y(_07455_));
 sg13g2_o21ai_1 _26573_ (.B1(_05819_),
    .Y(_07456_),
    .A1(_05844_),
    .A2(_07455_));
 sg13g2_buf_1 _26574_ (.A(_07456_),
    .X(_07457_));
 sg13g2_nor2_1 _26575_ (.A(_07439_),
    .B(_07457_),
    .Y(_07458_));
 sg13g2_o21ai_1 _26576_ (.B1(net90),
    .Y(_07459_),
    .A1(net91),
    .A2(_07458_));
 sg13g2_a22oi_1 _26577_ (.Y(_07460_),
    .B1(_07459_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07454_),
    .A1(_07440_));
 sg13g2_nor2_1 _26578_ (.A(net564),
    .B(_07460_),
    .Y(_01082_));
 sg13g2_nand3_1 _26579_ (.B(_05827_),
    .C(net981),
    .A(net982),
    .Y(_07461_));
 sg13g2_buf_1 _26580_ (.A(_07461_),
    .X(_07462_));
 sg13g2_nor2_2 _26581_ (.A(_07439_),
    .B(_07462_),
    .Y(_07463_));
 sg13g2_o21ai_1 _26582_ (.B1(net90),
    .Y(_07464_),
    .A1(net91),
    .A2(_07463_));
 sg13g2_a22oi_1 _26583_ (.Y(_07465_),
    .B1(_07464_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07463_),
    .A1(net69));
 sg13g2_nor2_1 _26584_ (.A(net564),
    .B(_07465_),
    .Y(_01083_));
 sg13g2_nor2_1 _26585_ (.A(net727),
    .B(_07452_),
    .Y(_07466_));
 sg13g2_buf_2 _26586_ (.A(_07466_),
    .X(_07467_));
 sg13g2_nor2_1 _26587_ (.A(_06022_),
    .B(_07439_),
    .Y(_07468_));
 sg13g2_o21ai_1 _26588_ (.B1(net90),
    .Y(_07469_),
    .A1(net91),
    .A2(_07468_));
 sg13g2_a22oi_1 _26589_ (.Y(_07470_),
    .B1(_07469_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07467_),
    .A1(_07440_));
 sg13g2_nor2_1 _26590_ (.A(net564),
    .B(_07470_),
    .Y(_01084_));
 sg13g2_nor2_2 _26591_ (.A(_05855_),
    .B(_07439_),
    .Y(_07471_));
 sg13g2_o21ai_1 _26592_ (.B1(net90),
    .Y(_07472_),
    .A1(net91),
    .A2(_07471_));
 sg13g2_a22oi_1 _26593_ (.Y(_07473_),
    .B1(_07472_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07471_),
    .A1(net69));
 sg13g2_nor2_1 _26594_ (.A(net564),
    .B(_07473_),
    .Y(_01085_));
 sg13g2_a21oi_1 _26595_ (.A1(net1107),
    .A2(_05863_),
    .Y(_07474_),
    .B1(_05293_));
 sg13g2_and2_1 _26596_ (.A(_06119_),
    .B(_07474_),
    .X(_07475_));
 sg13g2_buf_2 _26597_ (.A(_07475_),
    .X(_07476_));
 sg13g2_buf_1 _26598_ (.A(net565),
    .X(_07477_));
 sg13g2_o21ai_1 _26599_ (.B1(_05855_),
    .Y(_07478_),
    .A1(_05863_),
    .A2(_05917_));
 sg13g2_nand2_1 _26600_ (.Y(_07479_),
    .A(_05819_),
    .B(_07478_));
 sg13g2_nor2_1 _26601_ (.A(_07439_),
    .B(_07479_),
    .Y(_07480_));
 sg13g2_a21oi_1 _26602_ (.A1(_03356_),
    .A2(_11010_),
    .Y(_07481_),
    .B1(_05815_));
 sg13g2_nor2_1 _26603_ (.A(_07416_),
    .B(_07481_),
    .Y(_07482_));
 sg13g2_buf_2 _26604_ (.A(_07482_),
    .X(_07483_));
 sg13g2_buf_1 _26605_ (.A(_07483_),
    .X(_07484_));
 sg13g2_o21ai_1 _26606_ (.B1(net89),
    .Y(_07485_),
    .A1(net492),
    .A2(_07480_));
 sg13g2_a22oi_1 _26607_ (.Y(_07486_),
    .B1(_07485_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07476_),
    .A1(_07440_));
 sg13g2_nor2_1 _26608_ (.A(net564),
    .B(_07486_),
    .Y(_01086_));
 sg13g2_nor4_1 _26609_ (.A(_10419_),
    .B(net982),
    .C(net978),
    .D(net1107),
    .Y(_07487_));
 sg13g2_nand3_1 _26610_ (.B(net978),
    .C(net1107),
    .A(net974),
    .Y(_07488_));
 sg13g2_nand2b_1 _26611_ (.Y(_07489_),
    .B(_07488_),
    .A_N(_07487_));
 sg13g2_nand2b_1 _26612_ (.Y(_07490_),
    .B(net982),
    .A_N(net1107));
 sg13g2_a21oi_1 _26613_ (.A1(_07420_),
    .A2(_07490_),
    .Y(_07491_),
    .B1(_05925_));
 sg13g2_a22oi_1 _26614_ (.Y(_07492_),
    .B1(_07491_),
    .B2(_05964_),
    .A2(_07489_),
    .A1(_07420_));
 sg13g2_buf_2 _26615_ (.A(_07492_),
    .X(_07493_));
 sg13g2_nor3_2 _26616_ (.A(net844),
    .B(_05900_),
    .C(_07493_),
    .Y(_07494_));
 sg13g2_o21ai_1 _26617_ (.B1(net89),
    .Y(_07495_),
    .A1(net492),
    .A2(_07494_));
 sg13g2_a22oi_1 _26618_ (.Y(_07496_),
    .B1(_07495_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07494_),
    .A1(net69));
 sg13g2_nor2_1 _26619_ (.A(net564),
    .B(_07496_),
    .Y(_01087_));
 sg13g2_nor2_1 _26620_ (.A(net92),
    .B(_07493_),
    .Y(_07497_));
 sg13g2_o21ai_1 _26621_ (.B1(_07484_),
    .Y(_07498_),
    .A1(_07477_),
    .A2(_05928_));
 sg13g2_a22oi_1 _26622_ (.Y(_07499_),
    .B1(_07498_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07497_),
    .A1(_07434_));
 sg13g2_nor2_1 _26623_ (.A(net564),
    .B(_07499_),
    .Y(_01088_));
 sg13g2_o21ai_1 _26624_ (.B1(_07484_),
    .Y(_07500_),
    .A1(_07477_),
    .A2(_05935_));
 sg13g2_a22oi_1 _26625_ (.Y(_07501_),
    .B1(_07500_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07449_),
    .A1(_05935_));
 sg13g2_nor2_1 _26626_ (.A(net564),
    .B(_07501_),
    .Y(_01089_));
 sg13g2_nor2_1 _26627_ (.A(_05925_),
    .B(net1107),
    .Y(_07502_));
 sg13g2_a22oi_1 _26628_ (.Y(_07503_),
    .B1(_05926_),
    .B2(_07502_),
    .A2(_05893_),
    .A1(net1107));
 sg13g2_nor2b_1 _26629_ (.A(_07503_),
    .B_N(_07420_),
    .Y(_07504_));
 sg13g2_a21oi_1 _26630_ (.A1(_10420_),
    .A2(_07491_),
    .Y(_07505_),
    .B1(_07504_));
 sg13g2_buf_2 _26631_ (.A(_07505_),
    .X(_07506_));
 sg13g2_nor3_2 _26632_ (.A(net844),
    .B(_05900_),
    .C(_07506_),
    .Y(_07507_));
 sg13g2_o21ai_1 _26633_ (.B1(net90),
    .Y(_07508_),
    .A1(net91),
    .A2(_07507_));
 sg13g2_a22oi_1 _26634_ (.Y(_07509_),
    .B1(_07508_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07507_),
    .A1(net69));
 sg13g2_nor2_1 _26635_ (.A(_07446_),
    .B(_07509_),
    .Y(_01090_));
 sg13g2_buf_1 _26636_ (.A(_07445_),
    .X(_07510_));
 sg13g2_nor2_1 _26637_ (.A(_07457_),
    .B(_07493_),
    .Y(_07511_));
 sg13g2_o21ai_1 _26638_ (.B1(net89),
    .Y(_07512_),
    .A1(net492),
    .A2(_07511_));
 sg13g2_a22oi_1 _26639_ (.Y(_07513_),
    .B1(_07512_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07497_),
    .A1(_07454_));
 sg13g2_nor2_1 _26640_ (.A(net563),
    .B(_07513_),
    .Y(_01091_));
 sg13g2_nor2_2 _26641_ (.A(_07462_),
    .B(_07493_),
    .Y(_07514_));
 sg13g2_o21ai_1 _26642_ (.B1(net89),
    .Y(_07515_),
    .A1(net492),
    .A2(_07514_));
 sg13g2_a22oi_1 _26643_ (.Y(_07516_),
    .B1(_07515_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07514_),
    .A1(net69));
 sg13g2_nor2_1 _26644_ (.A(net563),
    .B(_07516_),
    .Y(_01092_));
 sg13g2_inv_1 _26645_ (.Y(_07517_),
    .A(_07493_));
 sg13g2_nor4_1 _26646_ (.A(_07430_),
    .B(net727),
    .C(_07416_),
    .D(_07452_),
    .Y(_07518_));
 sg13g2_nor2_1 _26647_ (.A(_06022_),
    .B(_07493_),
    .Y(_07519_));
 sg13g2_o21ai_1 _26648_ (.B1(net89),
    .Y(_07520_),
    .A1(net492),
    .A2(_07519_));
 sg13g2_a22oi_1 _26649_ (.Y(_07521_),
    .B1(_07520_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07518_),
    .A1(_07517_));
 sg13g2_nor2_1 _26650_ (.A(_07510_),
    .B(_07521_),
    .Y(_01093_));
 sg13g2_nor2_2 _26651_ (.A(_05855_),
    .B(_05916_),
    .Y(_07522_));
 sg13g2_o21ai_1 _26652_ (.B1(net89),
    .Y(_07523_),
    .A1(net492),
    .A2(_07522_));
 sg13g2_a22oi_1 _26653_ (.Y(_07524_),
    .B1(_07523_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07522_),
    .A1(net69));
 sg13g2_nor2_1 _26654_ (.A(net563),
    .B(_07524_),
    .Y(_01094_));
 sg13g2_nor2_1 _26655_ (.A(_07479_),
    .B(_07493_),
    .Y(_07525_));
 sg13g2_o21ai_1 _26656_ (.B1(net89),
    .Y(_07526_),
    .A1(net492),
    .A2(_07525_));
 sg13g2_a22oi_1 _26657_ (.Y(_07527_),
    .B1(_07526_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07497_),
    .A1(_07476_));
 sg13g2_nor2_1 _26658_ (.A(net563),
    .B(_07527_),
    .Y(_01095_));
 sg13g2_a21oi_1 _26659_ (.A1(_05964_),
    .A2(_07437_),
    .Y(_07528_),
    .B1(_07422_));
 sg13g2_buf_2 _26660_ (.A(_07528_),
    .X(_07529_));
 sg13g2_nor3_2 _26661_ (.A(net844),
    .B(_05900_),
    .C(_07529_),
    .Y(_07530_));
 sg13g2_o21ai_1 _26662_ (.B1(net89),
    .Y(_07531_),
    .A1(net492),
    .A2(_07530_));
 sg13g2_a22oi_1 _26663_ (.Y(_07532_),
    .B1(_07531_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07530_),
    .A1(net69));
 sg13g2_nor2_1 _26664_ (.A(net563),
    .B(_07532_),
    .Y(_01096_));
 sg13g2_nor2_1 _26665_ (.A(net92),
    .B(_07529_),
    .Y(_07533_));
 sg13g2_o21ai_1 _26666_ (.B1(_07483_),
    .Y(_07534_),
    .A1(net565),
    .A2(_05974_));
 sg13g2_a22oi_1 _26667_ (.Y(_07535_),
    .B1(_07534_),
    .B2(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A2(_07533_),
    .A1(_07434_));
 sg13g2_nor2_1 _26668_ (.A(_07510_),
    .B(_07535_),
    .Y(_01097_));
 sg13g2_o21ai_1 _26669_ (.B1(_07483_),
    .Y(_07536_),
    .A1(net565),
    .A2(_05979_));
 sg13g2_a22oi_1 _26670_ (.Y(_07537_),
    .B1(_07536_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07449_),
    .A1(_05979_));
 sg13g2_nor2_1 _26671_ (.A(net563),
    .B(_07537_),
    .Y(_01098_));
 sg13g2_nor2_1 _26672_ (.A(_07457_),
    .B(_07529_),
    .Y(_07538_));
 sg13g2_o21ai_1 _26673_ (.B1(_07483_),
    .Y(_07539_),
    .A1(net565),
    .A2(_07538_));
 sg13g2_a22oi_1 _26674_ (.Y(_07540_),
    .B1(_07539_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07533_),
    .A1(_07454_));
 sg13g2_nor2_1 _26675_ (.A(net563),
    .B(_07540_),
    .Y(_01099_));
 sg13g2_nor2_2 _26676_ (.A(_07462_),
    .B(_07529_),
    .Y(_07541_));
 sg13g2_o21ai_1 _26677_ (.B1(_07483_),
    .Y(_07542_),
    .A1(net565),
    .A2(_07541_));
 sg13g2_a22oi_1 _26678_ (.Y(_07543_),
    .B1(_07542_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07541_),
    .A1(net69));
 sg13g2_nor2_1 _26679_ (.A(net563),
    .B(_07543_),
    .Y(_01100_));
 sg13g2_buf_1 _26680_ (.A(_07445_),
    .X(_07544_));
 sg13g2_nor3_1 _26681_ (.A(net844),
    .B(net727),
    .C(_07506_),
    .Y(_07545_));
 sg13g2_o21ai_1 _26682_ (.B1(_07425_),
    .Y(_07546_),
    .A1(net92),
    .A2(_07545_));
 sg13g2_and2_1 _26683_ (.A(_04992_),
    .B(_07545_),
    .X(_07547_));
 sg13g2_a22oi_1 _26684_ (.Y(_07548_),
    .B1(_07547_),
    .B2(_07431_),
    .A2(_07546_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26685_ (.A(_07544_),
    .B(_07548_),
    .Y(_01101_));
 sg13g2_inv_1 _26686_ (.Y(_07549_),
    .A(_07529_));
 sg13g2_nor2_1 _26687_ (.A(_06022_),
    .B(_07529_),
    .Y(_07550_));
 sg13g2_o21ai_1 _26688_ (.B1(_07483_),
    .Y(_07551_),
    .A1(net565),
    .A2(_07550_));
 sg13g2_a22oi_1 _26689_ (.Y(_07552_),
    .B1(_07551_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07549_),
    .A1(_07518_));
 sg13g2_nor2_1 _26690_ (.A(net562),
    .B(_07552_),
    .Y(_01102_));
 sg13g2_nor2_2 _26691_ (.A(_05855_),
    .B(_07529_),
    .Y(_07553_));
 sg13g2_o21ai_1 _26692_ (.B1(_07483_),
    .Y(_07554_),
    .A1(net565),
    .A2(_07553_));
 sg13g2_a22oi_1 _26693_ (.Y(_07555_),
    .B1(_07554_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07553_),
    .A1(_07450_));
 sg13g2_nor2_1 _26694_ (.A(net562),
    .B(_07555_),
    .Y(_01103_));
 sg13g2_nor2b_2 _26695_ (.A(_07506_),
    .B_N(_05844_),
    .Y(_07556_));
 sg13g2_o21ai_1 _26696_ (.B1(net90),
    .Y(_07557_),
    .A1(net91),
    .A2(_07556_));
 sg13g2_a22oi_1 _26697_ (.Y(_07558_),
    .B1(_07557_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07556_),
    .A1(_07449_));
 sg13g2_nor2_1 _26698_ (.A(net562),
    .B(_07558_),
    .Y(_01104_));
 sg13g2_nor2_1 _26699_ (.A(net92),
    .B(_07506_),
    .Y(_07559_));
 sg13g2_nor2_1 _26700_ (.A(_07457_),
    .B(_07506_),
    .Y(_07560_));
 sg13g2_o21ai_1 _26701_ (.B1(net90),
    .Y(_07561_),
    .A1(net92),
    .A2(_07560_));
 sg13g2_a22oi_1 _26702_ (.Y(_07562_),
    .B1(_07561_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07559_),
    .A1(_07454_));
 sg13g2_nor2_1 _26703_ (.A(net562),
    .B(_07562_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26704_ (.B1(_07442_),
    .Y(_07563_),
    .A1(_06017_),
    .A2(_07441_));
 sg13g2_a22oi_1 _26705_ (.Y(_07564_),
    .B1(_07563_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07449_),
    .A1(_06017_));
 sg13g2_nor2_1 _26706_ (.A(net562),
    .B(_07564_),
    .Y(_01106_));
 sg13g2_o21ai_1 _26707_ (.B1(_07442_),
    .Y(_07565_),
    .A1(_06023_),
    .A2(net91));
 sg13g2_a22oi_1 _26708_ (.Y(_07566_),
    .B1(_07565_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07559_),
    .A1(_07467_));
 sg13g2_nor2_1 _26709_ (.A(net562),
    .B(_07566_),
    .Y(_01107_));
 sg13g2_o21ai_1 _26710_ (.B1(_07425_),
    .Y(_07567_),
    .A1(_06028_),
    .A2(_07441_));
 sg13g2_a22oi_1 _26711_ (.Y(_07568_),
    .B1(_07567_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07449_),
    .A1(_06028_));
 sg13g2_nor2_1 _26712_ (.A(net562),
    .B(_07568_),
    .Y(_01108_));
 sg13g2_nor2_1 _26713_ (.A(_07479_),
    .B(_07506_),
    .Y(_07569_));
 sg13g2_o21ai_1 _26714_ (.B1(_07425_),
    .Y(_07570_),
    .A1(_07419_),
    .A2(_07569_));
 sg13g2_a22oi_1 _26715_ (.Y(_07571_),
    .B1(_07570_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07559_),
    .A1(_07476_));
 sg13g2_nor2_1 _26716_ (.A(_07544_),
    .B(_07571_),
    .Y(_01109_));
 sg13g2_nor3_2 _26717_ (.A(net844),
    .B(_05900_),
    .C(_07439_),
    .Y(_07572_));
 sg13g2_o21ai_1 _26718_ (.B1(_07425_),
    .Y(_07573_),
    .A1(_07419_),
    .A2(_07572_));
 sg13g2_a22oi_1 _26719_ (.Y(_07574_),
    .B1(_07573_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07572_),
    .A1(_07449_));
 sg13g2_nor2_1 _26720_ (.A(net562),
    .B(_07574_),
    .Y(_01110_));
 sg13g2_buf_1 _26721_ (.A(_07445_),
    .X(_07575_));
 sg13g2_nand2_1 _26722_ (.Y(_07576_),
    .A(net1151),
    .B(_00257_));
 sg13g2_a21oi_1 _26723_ (.A1(_07413_),
    .A2(_07576_),
    .Y(_07577_),
    .B1(_07429_));
 sg13g2_nand2b_1 _26724_ (.Y(_07578_),
    .B(net275),
    .A_N(_07577_));
 sg13g2_buf_1 _26725_ (.A(_07578_),
    .X(_07579_));
 sg13g2_nor2_1 _26726_ (.A(net565),
    .B(_07579_),
    .Y(_07580_));
 sg13g2_nand2b_1 _26727_ (.Y(_07581_),
    .B(_05815_),
    .A_N(_07579_));
 sg13g2_buf_1 _26728_ (.A(_07581_),
    .X(_07582_));
 sg13g2_buf_1 _26729_ (.A(net144),
    .X(_07583_));
 sg13g2_nor2b_1 _26730_ (.A(_11051_),
    .B_N(_03356_),
    .Y(_07584_));
 sg13g2_a21oi_1 _26731_ (.A1(_05813_),
    .A2(_07584_),
    .Y(_07585_),
    .B1(_07579_));
 sg13g2_buf_2 _26732_ (.A(_07585_),
    .X(_07586_));
 sg13g2_buf_1 _26733_ (.A(_07586_),
    .X(_07587_));
 sg13g2_o21ai_1 _26734_ (.B1(net113),
    .Y(_07588_),
    .A1(_07422_),
    .A2(net114));
 sg13g2_a22oi_1 _26735_ (.Y(_07589_),
    .B1(_07588_),
    .B2(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A2(_07580_),
    .A1(_07427_));
 sg13g2_nor2_1 _26736_ (.A(net561),
    .B(_07589_),
    .Y(_01111_));
 sg13g2_nor2_1 _26737_ (.A(_07439_),
    .B(net144),
    .Y(_07590_));
 sg13g2_o21ai_1 _26738_ (.B1(net113),
    .Y(_07591_),
    .A1(_05881_),
    .A2(net114));
 sg13g2_a22oi_1 _26739_ (.Y(_07592_),
    .B1(_07591_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07590_),
    .A1(_07434_));
 sg13g2_nor2_1 _26740_ (.A(_07575_),
    .B(_07592_),
    .Y(_01112_));
 sg13g2_o21ai_1 _26741_ (.B1(_07586_),
    .Y(_07593_),
    .A1(_05889_),
    .A2(_07582_));
 sg13g2_nor2_1 _26742_ (.A(net544),
    .B(net144),
    .Y(_07594_));
 sg13g2_buf_2 _26743_ (.A(_07594_),
    .X(_07595_));
 sg13g2_buf_1 _26744_ (.A(_07595_),
    .X(_07596_));
 sg13g2_a22oi_1 _26745_ (.Y(_07597_),
    .B1(net79),
    .B2(_05889_),
    .A2(_07593_),
    .A1(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_nor2_1 _26746_ (.A(net561),
    .B(_07597_),
    .Y(_01113_));
 sg13g2_o21ai_1 _26747_ (.B1(net113),
    .Y(_07598_),
    .A1(_07458_),
    .A2(net114));
 sg13g2_a22oi_1 _26748_ (.Y(_07599_),
    .B1(_07598_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07590_),
    .A1(_07454_));
 sg13g2_nor2_1 _26749_ (.A(net561),
    .B(_07599_),
    .Y(_01114_));
 sg13g2_o21ai_1 _26750_ (.B1(net113),
    .Y(_07600_),
    .A1(_07463_),
    .A2(_07583_));
 sg13g2_a22oi_1 _26751_ (.Y(_07601_),
    .B1(_07600_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(_07596_),
    .A1(_07463_));
 sg13g2_nor2_1 _26752_ (.A(net561),
    .B(_07601_),
    .Y(_01115_));
 sg13g2_o21ai_1 _26753_ (.B1(net113),
    .Y(_07602_),
    .A1(_07468_),
    .A2(net114));
 sg13g2_a22oi_1 _26754_ (.Y(_07603_),
    .B1(_07602_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07590_),
    .A1(_07467_));
 sg13g2_nor2_1 _26755_ (.A(net561),
    .B(_07603_),
    .Y(_01116_));
 sg13g2_o21ai_1 _26756_ (.B1(net113),
    .Y(_07604_),
    .A1(_07471_),
    .A2(_07583_));
 sg13g2_a22oi_1 _26757_ (.Y(_07605_),
    .B1(_07604_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net79),
    .A1(_07471_));
 sg13g2_nor2_1 _26758_ (.A(_07575_),
    .B(_07605_),
    .Y(_01117_));
 sg13g2_a21oi_1 _26759_ (.A1(_03356_),
    .A2(\cpu.dec.imm[3] ),
    .Y(_07606_),
    .B1(_05815_));
 sg13g2_nor2_1 _26760_ (.A(_07579_),
    .B(_07606_),
    .Y(_07607_));
 sg13g2_buf_2 _26761_ (.A(_07607_),
    .X(_07608_));
 sg13g2_buf_1 _26762_ (.A(_07608_),
    .X(_07609_));
 sg13g2_o21ai_1 _26763_ (.B1(net112),
    .Y(_07610_),
    .A1(_07480_),
    .A2(net114));
 sg13g2_a22oi_1 _26764_ (.Y(_07611_),
    .B1(_07610_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07590_),
    .A1(_07476_));
 sg13g2_nor2_1 _26765_ (.A(net561),
    .B(_07611_),
    .Y(_01118_));
 sg13g2_o21ai_1 _26766_ (.B1(net112),
    .Y(_07612_),
    .A1(_07494_),
    .A2(net114));
 sg13g2_a22oi_1 _26767_ (.Y(_07613_),
    .B1(_07612_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net79),
    .A1(_07494_));
 sg13g2_nor2_1 _26768_ (.A(net561),
    .B(_07613_),
    .Y(_01119_));
 sg13g2_nor2_1 _26769_ (.A(_07493_),
    .B(net144),
    .Y(_07614_));
 sg13g2_o21ai_1 _26770_ (.B1(net112),
    .Y(_07615_),
    .A1(_05928_),
    .A2(net114));
 sg13g2_a22oi_1 _26771_ (.Y(_07616_),
    .B1(_07615_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07614_),
    .A1(_07434_));
 sg13g2_nor2_1 _26772_ (.A(net561),
    .B(_07616_),
    .Y(_01120_));
 sg13g2_buf_1 _26773_ (.A(_07445_),
    .X(_07617_));
 sg13g2_o21ai_1 _26774_ (.B1(_07609_),
    .Y(_07618_),
    .A1(_05935_),
    .A2(net114));
 sg13g2_a22oi_1 _26775_ (.Y(_07619_),
    .B1(_07618_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net79),
    .A1(_05935_));
 sg13g2_nor2_1 _26776_ (.A(_07617_),
    .B(_07619_),
    .Y(_01121_));
 sg13g2_buf_1 _26777_ (.A(net144),
    .X(_07620_));
 sg13g2_o21ai_1 _26778_ (.B1(net113),
    .Y(_07621_),
    .A1(_07507_),
    .A2(_07620_));
 sg13g2_a22oi_1 _26779_ (.Y(_07622_),
    .B1(_07621_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(_07596_),
    .A1(_07507_));
 sg13g2_nor2_1 _26780_ (.A(net560),
    .B(_07622_),
    .Y(_01122_));
 sg13g2_o21ai_1 _26781_ (.B1(net112),
    .Y(_07623_),
    .A1(_07511_),
    .A2(net111));
 sg13g2_a22oi_1 _26782_ (.Y(_07624_),
    .B1(_07623_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07614_),
    .A1(_07454_));
 sg13g2_nor2_1 _26783_ (.A(net560),
    .B(_07624_),
    .Y(_01123_));
 sg13g2_o21ai_1 _26784_ (.B1(net112),
    .Y(_07625_),
    .A1(_07514_),
    .A2(net111));
 sg13g2_a22oi_1 _26785_ (.Y(_07626_),
    .B1(_07625_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net79),
    .A1(_07514_));
 sg13g2_nor2_1 _26786_ (.A(net560),
    .B(_07626_),
    .Y(_01124_));
 sg13g2_o21ai_1 _26787_ (.B1(net112),
    .Y(_07627_),
    .A1(_07519_),
    .A2(net111));
 sg13g2_a22oi_1 _26788_ (.Y(_07628_),
    .B1(_07627_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07614_),
    .A1(_07467_));
 sg13g2_nor2_1 _26789_ (.A(net560),
    .B(_07628_),
    .Y(_01125_));
 sg13g2_o21ai_1 _26790_ (.B1(_07609_),
    .Y(_07629_),
    .A1(_07522_),
    .A2(_07620_));
 sg13g2_a22oi_1 _26791_ (.Y(_07630_),
    .B1(_07629_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net79),
    .A1(_07522_));
 sg13g2_nor2_1 _26792_ (.A(net560),
    .B(_07630_),
    .Y(_01126_));
 sg13g2_o21ai_1 _26793_ (.B1(net112),
    .Y(_07631_),
    .A1(_07525_),
    .A2(net111));
 sg13g2_a22oi_1 _26794_ (.Y(_07632_),
    .B1(_07631_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07614_),
    .A1(_07476_));
 sg13g2_nor2_1 _26795_ (.A(net560),
    .B(_07632_),
    .Y(_01127_));
 sg13g2_o21ai_1 _26796_ (.B1(net112),
    .Y(_07633_),
    .A1(_07530_),
    .A2(net111));
 sg13g2_a22oi_1 _26797_ (.Y(_07634_),
    .B1(_07633_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net79),
    .A1(_07530_));
 sg13g2_nor2_1 _26798_ (.A(_07617_),
    .B(_07634_),
    .Y(_01128_));
 sg13g2_nor2_1 _26799_ (.A(_07529_),
    .B(net144),
    .Y(_07635_));
 sg13g2_o21ai_1 _26800_ (.B1(_07608_),
    .Y(_07636_),
    .A1(_05974_),
    .A2(net111));
 sg13g2_a22oi_1 _26801_ (.Y(_07637_),
    .B1(_07636_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07635_),
    .A1(_07434_));
 sg13g2_nor2_1 _26802_ (.A(net560),
    .B(_07637_),
    .Y(_01129_));
 sg13g2_o21ai_1 _26803_ (.B1(_07608_),
    .Y(_07638_),
    .A1(_05979_),
    .A2(net111));
 sg13g2_a22oi_1 _26804_ (.Y(_07639_),
    .B1(_07638_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(net79),
    .A1(_05979_));
 sg13g2_nor2_1 _26805_ (.A(net560),
    .B(_07639_),
    .Y(_01130_));
 sg13g2_buf_1 _26806_ (.A(_07445_),
    .X(_07640_));
 sg13g2_o21ai_1 _26807_ (.B1(_07608_),
    .Y(_07641_),
    .A1(_07538_),
    .A2(net111));
 sg13g2_a22oi_1 _26808_ (.Y(_07642_),
    .B1(_07641_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07635_),
    .A1(_07454_));
 sg13g2_nor2_1 _26809_ (.A(net559),
    .B(_07642_),
    .Y(_01131_));
 sg13g2_buf_1 _26810_ (.A(net144),
    .X(_07643_));
 sg13g2_o21ai_1 _26811_ (.B1(_07608_),
    .Y(_07644_),
    .A1(_07541_),
    .A2(net110));
 sg13g2_a22oi_1 _26812_ (.Y(_07645_),
    .B1(_07644_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07595_),
    .A1(_07541_));
 sg13g2_nor2_1 _26813_ (.A(net559),
    .B(_07645_),
    .Y(_01132_));
 sg13g2_o21ai_1 _26814_ (.B1(net113),
    .Y(_07646_),
    .A1(_07545_),
    .A2(net110));
 sg13g2_a22oi_1 _26815_ (.Y(_07647_),
    .B1(_07646_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07580_),
    .A1(_07547_));
 sg13g2_nor2_1 _26816_ (.A(net559),
    .B(_07647_),
    .Y(_01133_));
 sg13g2_o21ai_1 _26817_ (.B1(_07608_),
    .Y(_07648_),
    .A1(_07550_),
    .A2(net110));
 sg13g2_a22oi_1 _26818_ (.Y(_07649_),
    .B1(_07648_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07635_),
    .A1(_07467_));
 sg13g2_nor2_1 _26819_ (.A(net559),
    .B(_07649_),
    .Y(_01134_));
 sg13g2_o21ai_1 _26820_ (.B1(_07608_),
    .Y(_07650_),
    .A1(_07553_),
    .A2(net110));
 sg13g2_a22oi_1 _26821_ (.Y(_07651_),
    .B1(_07650_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07595_),
    .A1(_07553_));
 sg13g2_nor2_1 _26822_ (.A(net559),
    .B(_07651_),
    .Y(_01135_));
 sg13g2_o21ai_1 _26823_ (.B1(_07587_),
    .Y(_07652_),
    .A1(_07556_),
    .A2(net110));
 sg13g2_a22oi_1 _26824_ (.Y(_07653_),
    .B1(_07652_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07595_),
    .A1(_07556_));
 sg13g2_nor2_1 _26825_ (.A(net559),
    .B(_07653_),
    .Y(_01136_));
 sg13g2_nor2_1 _26826_ (.A(_07506_),
    .B(net144),
    .Y(_07654_));
 sg13g2_o21ai_1 _26827_ (.B1(_07587_),
    .Y(_07655_),
    .A1(_07560_),
    .A2(_07643_));
 sg13g2_a22oi_1 _26828_ (.Y(_07656_),
    .B1(_07655_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07654_),
    .A1(_07454_));
 sg13g2_nor2_1 _26829_ (.A(net559),
    .B(_07656_),
    .Y(_01137_));
 sg13g2_o21ai_1 _26830_ (.B1(_07586_),
    .Y(_07657_),
    .A1(_06017_),
    .A2(net110));
 sg13g2_a22oi_1 _26831_ (.Y(_07658_),
    .B1(_07657_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07595_),
    .A1(_06017_));
 sg13g2_nor2_1 _26832_ (.A(_07640_),
    .B(_07658_),
    .Y(_01138_));
 sg13g2_o21ai_1 _26833_ (.B1(_07586_),
    .Y(_07659_),
    .A1(_06023_),
    .A2(net110));
 sg13g2_a22oi_1 _26834_ (.Y(_07660_),
    .B1(_07659_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07654_),
    .A1(_07467_));
 sg13g2_nor2_1 _26835_ (.A(net559),
    .B(_07660_),
    .Y(_01139_));
 sg13g2_o21ai_1 _26836_ (.B1(_07586_),
    .Y(_07661_),
    .A1(_06028_),
    .A2(_07643_));
 sg13g2_a22oi_1 _26837_ (.Y(_07662_),
    .B1(_07661_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07595_),
    .A1(_06028_));
 sg13g2_nor2_1 _26838_ (.A(_07640_),
    .B(_07662_),
    .Y(_01140_));
 sg13g2_buf_1 _26839_ (.A(_07445_),
    .X(_07663_));
 sg13g2_o21ai_1 _26840_ (.B1(_07586_),
    .Y(_07664_),
    .A1(_07569_),
    .A2(net110));
 sg13g2_a22oi_1 _26841_ (.Y(_07665_),
    .B1(_07664_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07654_),
    .A1(_07476_));
 sg13g2_nor2_1 _26842_ (.A(_07663_),
    .B(_07665_),
    .Y(_01141_));
 sg13g2_o21ai_1 _26843_ (.B1(_07586_),
    .Y(_07666_),
    .A1(_07572_),
    .A2(_07582_));
 sg13g2_a22oi_1 _26844_ (.Y(_07667_),
    .B1(_07666_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07595_),
    .A1(_07572_));
 sg13g2_nor2_1 _26845_ (.A(_07663_),
    .B(_07667_),
    .Y(_01142_));
 sg13g2_and2_1 _26846_ (.A(net455),
    .B(_06369_),
    .X(_07668_));
 sg13g2_buf_2 _26847_ (.A(_07668_),
    .X(_07669_));
 sg13g2_nand2_1 _26848_ (.Y(_07670_),
    .A(net946),
    .B(_07669_));
 sg13g2_nand2_1 _26849_ (.Y(_07671_),
    .A(net455),
    .B(_06369_));
 sg13g2_buf_2 _26850_ (.A(_07671_),
    .X(_07672_));
 sg13g2_nand2_1 _26851_ (.Y(_07673_),
    .A(\cpu.gpio.r_enable_in[0] ),
    .B(_07672_));
 sg13g2_a21oi_1 _26852_ (.A1(_07670_),
    .A2(_07673_),
    .Y(_01943_),
    .B1(net567));
 sg13g2_nand2_1 _26853_ (.Y(_07674_),
    .A(net999),
    .B(_07669_));
 sg13g2_nand2_1 _26854_ (.Y(_07675_),
    .A(\cpu.gpio.r_enable_in[1] ),
    .B(_07672_));
 sg13g2_a21oi_1 _26855_ (.A1(_07674_),
    .A2(_07675_),
    .Y(_01944_),
    .B1(net567));
 sg13g2_nand2_1 _26856_ (.Y(_07676_),
    .A(net864),
    .B(_07669_));
 sg13g2_nand2_1 _26857_ (.Y(_07677_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_07672_));
 sg13g2_buf_1 _26858_ (.A(_09368_),
    .X(_07678_));
 sg13g2_a21oi_1 _26859_ (.A1(_07676_),
    .A2(_07677_),
    .Y(_01945_),
    .B1(_07678_));
 sg13g2_nand2_1 _26860_ (.Y(_07679_),
    .A(net1054),
    .B(_07669_));
 sg13g2_nand2_1 _26861_ (.Y(_07680_),
    .A(\cpu.gpio.r_enable_in[3] ),
    .B(_07672_));
 sg13g2_a21oi_1 _26862_ (.A1(_07679_),
    .A2(_07680_),
    .Y(_01946_),
    .B1(net557));
 sg13g2_nand2_1 _26863_ (.Y(_07681_),
    .A(net1053),
    .B(_07669_));
 sg13g2_nand2_1 _26864_ (.Y(_07682_),
    .A(_09261_),
    .B(_07672_));
 sg13g2_a21oi_1 _26865_ (.A1(_07681_),
    .A2(_07682_),
    .Y(_01947_),
    .B1(net557));
 sg13g2_nand2_1 _26866_ (.Y(_07683_),
    .A(net1052),
    .B(_07669_));
 sg13g2_nand2_1 _26867_ (.Y(_07684_),
    .A(\cpu.gpio.r_enable_in[5] ),
    .B(_07672_));
 sg13g2_a21oi_1 _26868_ (.A1(_07683_),
    .A2(_07684_),
    .Y(_01948_),
    .B1(net557));
 sg13g2_nand2_1 _26869_ (.Y(_07685_),
    .A(net1051),
    .B(_07669_));
 sg13g2_nand2_1 _26870_ (.Y(_07686_),
    .A(\cpu.gpio.r_enable_in[6] ),
    .B(_07672_));
 sg13g2_a21oi_1 _26871_ (.A1(_07685_),
    .A2(_07686_),
    .Y(_01949_),
    .B1(_07678_));
 sg13g2_nand2_1 _26872_ (.Y(_07687_),
    .A(net1050),
    .B(_07669_));
 sg13g2_nand2_1 _26873_ (.Y(_07688_),
    .A(_09251_),
    .B(_07672_));
 sg13g2_a21oi_1 _26874_ (.A1(_07687_),
    .A2(_07688_),
    .Y(_01950_),
    .B1(net557));
 sg13g2_buf_1 _26875_ (.A(_06369_),
    .X(_07689_));
 sg13g2_nand3_1 _26876_ (.B(net407),
    .C(net109),
    .A(net1053),
    .Y(_07690_));
 sg13g2_nand2_1 _26877_ (.Y(_07691_),
    .A(net407),
    .B(_06369_));
 sg13g2_nand2_1 _26878_ (.Y(_07692_),
    .A(\cpu.gpio.r_enable_io[4] ),
    .B(_07691_));
 sg13g2_a21oi_1 _26879_ (.A1(_07690_),
    .A2(_07692_),
    .Y(_01951_),
    .B1(net557));
 sg13g2_nand3_1 _26880_ (.B(net407),
    .C(_07689_),
    .A(net1052),
    .Y(_07693_));
 sg13g2_nand2_1 _26881_ (.Y(_07694_),
    .A(_09265_),
    .B(_07691_));
 sg13g2_a21oi_1 _26882_ (.A1(_07693_),
    .A2(_07694_),
    .Y(_01952_),
    .B1(net557));
 sg13g2_nand3_1 _26883_ (.B(_05477_),
    .C(net109),
    .A(net1051),
    .Y(_07695_));
 sg13g2_nand2_1 _26884_ (.Y(_07696_),
    .A(\cpu.gpio.r_enable_io[6] ),
    .B(_07691_));
 sg13g2_a21oi_1 _26885_ (.A1(_07695_),
    .A2(_07696_),
    .Y(_01953_),
    .B1(net557));
 sg13g2_nand3_1 _26886_ (.B(_05477_),
    .C(_07689_),
    .A(net1050),
    .Y(_07697_));
 sg13g2_nand2_1 _26887_ (.Y(_07698_),
    .A(_09256_),
    .B(_07691_));
 sg13g2_a21oi_1 _26888_ (.A1(_07697_),
    .A2(_07698_),
    .Y(_01954_),
    .B1(net557));
 sg13g2_nand3_1 _26889_ (.B(_05184_),
    .C(_06369_),
    .A(net984),
    .Y(_07699_));
 sg13g2_buf_1 _26890_ (.A(_07699_),
    .X(_07700_));
 sg13g2_mux2_1 _26891_ (.A0(_10116_),
    .A1(net7),
    .S(_07700_),
    .X(_07701_));
 sg13g2_and2_1 _26892_ (.A(net693),
    .B(_07701_),
    .X(_01955_));
 sg13g2_mux2_1 _26893_ (.A0(net1052),
    .A1(net8),
    .S(_07700_),
    .X(_07702_));
 sg13g2_and2_1 _26894_ (.A(net693),
    .B(_07702_),
    .X(_01956_));
 sg13g2_mux2_1 _26895_ (.A0(net1051),
    .A1(net9),
    .S(_07700_),
    .X(_07703_));
 sg13g2_and2_1 _26896_ (.A(net693),
    .B(_07703_),
    .X(_01957_));
 sg13g2_mux2_1 _26897_ (.A0(_10131_),
    .A1(net10),
    .S(_07700_),
    .X(_07704_));
 sg13g2_and2_1 _26898_ (.A(net693),
    .B(_07704_),
    .X(_01958_));
 sg13g2_nand3_1 _26899_ (.B(_04864_),
    .C(net109),
    .A(net946),
    .Y(_07705_));
 sg13g2_nand2_1 _26900_ (.Y(_07706_),
    .A(_04864_),
    .B(_06369_));
 sg13g2_nand2_1 _26901_ (.Y(_07707_),
    .A(_04865_),
    .B(_07706_));
 sg13g2_nand3_1 _26902_ (.B(_07705_),
    .C(_07707_),
    .A(net728),
    .Y(_02004_));
 sg13g2_nand3_1 _26903_ (.B(_04864_),
    .C(net109),
    .A(net1056),
    .Y(_07708_));
 sg13g2_buf_1 _26904_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07709_));
 sg13g2_nand2_1 _26905_ (.Y(_07710_),
    .A(_07709_),
    .B(_07706_));
 sg13g2_buf_1 _26906_ (.A(_09368_),
    .X(_07711_));
 sg13g2_a21oi_1 _26907_ (.A1(_07708_),
    .A2(_07710_),
    .Y(_02005_),
    .B1(net556));
 sg13g2_nand3_1 _26908_ (.B(_04864_),
    .C(net109),
    .A(net1055),
    .Y(_07712_));
 sg13g2_nand2_1 _26909_ (.Y(_07713_),
    .A(\cpu.gpio.r_src_o[6][2] ),
    .B(_07706_));
 sg13g2_a21oi_1 _26910_ (.A1(_07712_),
    .A2(_07713_),
    .Y(_02006_),
    .B1(net556));
 sg13g2_nand3_1 _26911_ (.B(_04864_),
    .C(net109),
    .A(net1054),
    .Y(_07714_));
 sg13g2_nand2_1 _26912_ (.Y(_07715_),
    .A(\cpu.gpio.r_src_o[6][3] ),
    .B(_07706_));
 sg13g2_a21oi_1 _26913_ (.A1(_07714_),
    .A2(_07715_),
    .Y(_02007_),
    .B1(net556));
 sg13g2_nand2_1 _26914_ (.Y(_07716_),
    .A(_04868_),
    .B(_06369_));
 sg13g2_mux2_1 _26915_ (.A0(net1057),
    .A1(_04867_),
    .S(_07716_),
    .X(_07717_));
 sg13g2_and2_1 _26916_ (.A(_09310_),
    .B(_07717_),
    .X(_02012_));
 sg13g2_nand3_1 _26917_ (.B(_04868_),
    .C(net109),
    .A(net1056),
    .Y(_07718_));
 sg13g2_nand2_1 _26918_ (.Y(_07719_),
    .A(\cpu.gpio.r_uart_rx_src[1] ),
    .B(_07716_));
 sg13g2_a21oi_1 _26919_ (.A1(_07718_),
    .A2(_07719_),
    .Y(_02013_),
    .B1(_07711_));
 sg13g2_nand3_1 _26920_ (.B(_04868_),
    .C(net109),
    .A(net1055),
    .Y(_07720_));
 sg13g2_nand2_1 _26921_ (.Y(_07721_),
    .A(\cpu.gpio.r_uart_rx_src[2] ),
    .B(_07716_));
 sg13g2_a21oi_1 _26922_ (.A1(_07720_),
    .A2(_07721_),
    .Y(_02014_),
    .B1(_07711_));
 sg13g2_and2_1 _26923_ (.A(\cpu.i_wstrobe_d ),
    .B(_00318_),
    .X(_02271_));
 sg13g2_a21oi_1 _26924_ (.A1(_06402_),
    .A2(_06414_),
    .Y(_02272_),
    .B1(_06425_));
 sg13g2_xor2_1 _26925_ (.B(_06409_),
    .A(_06398_),
    .X(_07722_));
 sg13g2_nor2_1 _26926_ (.A(_06425_),
    .B(_07722_),
    .Y(_02273_));
 sg13g2_xnor2_1 _26927_ (.Y(_07723_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05276_));
 sg13g2_xnor2_1 _26928_ (.Y(_07724_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10207_));
 sg13g2_xnor2_1 _26929_ (.Y(_07725_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10224_));
 sg13g2_xnor2_1 _26930_ (.Y(_07726_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10161_));
 sg13g2_nand4_1 _26931_ (.B(_07724_),
    .C(_07725_),
    .A(_07723_),
    .Y(_07727_),
    .D(_07726_));
 sg13g2_xnor2_1 _26932_ (.Y(_07728_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05214_));
 sg13g2_xnor2_1 _26933_ (.Y(_07729_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05710_));
 sg13g2_xnor2_1 _26934_ (.Y(_07730_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05122_));
 sg13g2_xnor2_1 _26935_ (.Y(_07731_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04885_));
 sg13g2_nand4_1 _26936_ (.B(_07729_),
    .C(_07730_),
    .A(_07728_),
    .Y(_07732_),
    .D(_07731_));
 sg13g2_xnor2_1 _26937_ (.Y(_07733_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10230_));
 sg13g2_xnor2_1 _26938_ (.Y(_07734_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05751_));
 sg13g2_xnor2_1 _26939_ (.Y(_07735_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10189_));
 sg13g2_xnor2_1 _26940_ (.Y(_07736_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05171_));
 sg13g2_nand4_1 _26941_ (.B(_07734_),
    .C(_07735_),
    .A(_07733_),
    .Y(_07737_),
    .D(_07736_));
 sg13g2_xnor2_1 _26942_ (.Y(_07738_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05427_));
 sg13g2_xnor2_1 _26943_ (.Y(_07739_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05606_));
 sg13g2_xnor2_1 _26944_ (.Y(_07740_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10217_));
 sg13g2_xnor2_1 _26945_ (.Y(_07741_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10195_));
 sg13g2_nand4_1 _26946_ (.B(_07739_),
    .C(_07740_),
    .A(_07738_),
    .Y(_07742_),
    .D(_07741_));
 sg13g2_nor4_1 _26947_ (.A(_07727_),
    .B(_07732_),
    .C(_07737_),
    .D(_07742_),
    .Y(_07743_));
 sg13g2_xnor2_1 _26948_ (.Y(_07744_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05361_));
 sg13g2_xnor2_1 _26949_ (.Y(_07745_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05486_));
 sg13g2_xnor2_1 _26950_ (.Y(_07746_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10183_));
 sg13g2_xnor2_1 _26951_ (.Y(_07747_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10160_));
 sg13g2_nand4_1 _26952_ (.B(_07745_),
    .C(_07746_),
    .A(_07744_),
    .Y(_07748_),
    .D(_07747_));
 sg13g2_xnor2_1 _26953_ (.Y(_07749_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10199_));
 sg13g2_xnor2_1 _26954_ (.Y(_07750_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10177_));
 sg13g2_xnor2_1 _26955_ (.Y(_07751_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05558_));
 sg13g2_xnor2_1 _26956_ (.Y(_07752_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05262_));
 sg13g2_nand4_1 _26957_ (.B(_07750_),
    .C(_07751_),
    .A(_07749_),
    .Y(_07753_),
    .D(_07752_));
 sg13g2_xnor2_1 _26958_ (.Y(_07754_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05020_));
 sg13g2_xnor2_1 _26959_ (.Y(_07755_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05186_));
 sg13g2_xnor2_1 _26960_ (.Y(_07756_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10212_));
 sg13g2_xnor2_1 _26961_ (.Y(_07757_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10171_));
 sg13g2_nand4_1 _26962_ (.B(_07755_),
    .C(_07756_),
    .A(_07754_),
    .Y(_07758_),
    .D(_07757_));
 sg13g2_xnor2_1 _26963_ (.Y(_07759_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10234_));
 sg13g2_xnor2_1 _26964_ (.Y(_07760_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10166_));
 sg13g2_xnor2_1 _26965_ (.Y(_07761_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10241_));
 sg13g2_xnor2_1 _26966_ (.Y(_07762_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(\cpu.intr.r_clock_count[24] ));
 sg13g2_nand4_1 _26967_ (.B(_07760_),
    .C(_07761_),
    .A(_07759_),
    .Y(_07763_),
    .D(_07762_));
 sg13g2_nor4_1 _26968_ (.A(_07748_),
    .B(_07753_),
    .C(_07758_),
    .D(_07763_),
    .Y(_07764_));
 sg13g2_a22oi_1 _26969_ (.Y(_07765_),
    .B1(_07743_),
    .B2(_07764_),
    .A2(_07371_),
    .A1(net1049));
 sg13g2_nand3_1 _26970_ (.B(net193),
    .C(net411),
    .A(net1049),
    .Y(_07766_));
 sg13g2_nand2_1 _26971_ (.Y(_07767_),
    .A(_09274_),
    .B(_07766_));
 sg13g2_a21oi_1 _26972_ (.A1(_07765_),
    .A2(_07767_),
    .Y(_02434_),
    .B1(net556));
 sg13g2_and2_1 _26973_ (.A(net193),
    .B(_04888_),
    .X(_07768_));
 sg13g2_buf_1 _26974_ (.A(_07768_),
    .X(_07769_));
 sg13g2_nand2_1 _26975_ (.Y(_07770_),
    .A(net946),
    .B(_07769_));
 sg13g2_nand2_1 _26976_ (.Y(_07771_),
    .A(net193),
    .B(_04888_));
 sg13g2_buf_1 _26977_ (.A(_07771_),
    .X(_07772_));
 sg13g2_nand2_1 _26978_ (.Y(_07773_),
    .A(_09280_),
    .B(_07772_));
 sg13g2_a21oi_1 _26979_ (.A1(_07770_),
    .A2(_07773_),
    .Y(_02483_),
    .B1(net556));
 sg13g2_nand2_1 _26980_ (.Y(_07774_),
    .A(net1056),
    .B(_07769_));
 sg13g2_nand2_1 _26981_ (.Y(_07775_),
    .A(\cpu.intr.r_enable[1] ),
    .B(_07772_));
 sg13g2_a21oi_1 _26982_ (.A1(_07774_),
    .A2(_07775_),
    .Y(_02484_),
    .B1(net556));
 sg13g2_nand2_1 _26983_ (.Y(_07776_),
    .A(net1055),
    .B(_07769_));
 sg13g2_nand2_1 _26984_ (.Y(_07777_),
    .A(_09271_),
    .B(_07772_));
 sg13g2_a21oi_1 _26985_ (.A1(_07776_),
    .A2(_07777_),
    .Y(_02485_),
    .B1(net556));
 sg13g2_nand2_1 _26986_ (.Y(_07778_),
    .A(net1054),
    .B(_07769_));
 sg13g2_nand2_1 _26987_ (.Y(_07779_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07772_));
 sg13g2_a21oi_1 _26988_ (.A1(_07778_),
    .A2(_07779_),
    .Y(_02486_),
    .B1(net556));
 sg13g2_nand2_1 _26989_ (.Y(_07780_),
    .A(net1053),
    .B(_07769_));
 sg13g2_nand2_1 _26990_ (.Y(_07781_),
    .A(_09244_),
    .B(_07772_));
 sg13g2_buf_1 _26991_ (.A(_09368_),
    .X(_07782_));
 sg13g2_a21oi_1 _26992_ (.A1(_07780_),
    .A2(_07781_),
    .Y(_02487_),
    .B1(net555));
 sg13g2_nand2_1 _26993_ (.Y(_07783_),
    .A(net1052),
    .B(_07769_));
 sg13g2_nand2_1 _26994_ (.Y(_07784_),
    .A(_09276_),
    .B(_07772_));
 sg13g2_a21oi_1 _26995_ (.A1(_07783_),
    .A2(_07784_),
    .Y(_02488_),
    .B1(net555));
 sg13g2_nand3_1 _26996_ (.B(net193),
    .C(_04945_),
    .A(net1048),
    .Y(_07785_));
 sg13g2_inv_1 _26997_ (.Y(_07786_),
    .A(_10017_));
 sg13g2_a221oi_1 _26998_ (.B2(_09270_),
    .C1(_07786_),
    .B1(_07785_),
    .A1(net1055),
    .Y(_07787_),
    .A2(_07371_));
 sg13g2_nor2_1 _26999_ (.A(net558),
    .B(_07787_),
    .Y(_02489_));
 sg13g2_nand3b_1 _27000_ (.B(_06816_),
    .C(_09885_),
    .Y(_07788_),
    .A_N(_06807_));
 sg13g2_buf_1 _27001_ (.A(_07788_),
    .X(_07789_));
 sg13g2_o21ai_1 _27002_ (.B1(net916),
    .Y(_07790_),
    .A1(_06811_),
    .A2(_07789_));
 sg13g2_nor2b_1 _27003_ (.A(_09878_),
    .B_N(_09861_),
    .Y(_07791_));
 sg13g2_o21ai_1 _27004_ (.B1(net19),
    .Y(_07792_),
    .A1(_07789_),
    .A2(_07791_));
 sg13g2_nand2b_1 _27005_ (.Y(_02519_),
    .B(_07792_),
    .A_N(_07790_));
 sg13g2_nand3b_1 _27006_ (.B(_06840_),
    .C(_09841_),
    .Y(_07793_),
    .A_N(_09861_));
 sg13g2_a21o_1 _27007_ (.A2(_07793_),
    .A1(_06811_),
    .B1(_07789_),
    .X(_07794_));
 sg13g2_nand2_1 _27008_ (.Y(_07795_),
    .A(_09861_),
    .B(_06811_));
 sg13g2_nor2_1 _27009_ (.A(_09873_),
    .B(_07795_),
    .Y(_07796_));
 sg13g2_o21ai_1 _27010_ (.B1(net20),
    .Y(_07797_),
    .A1(_07789_),
    .A2(_07796_));
 sg13g2_nand3_1 _27011_ (.B(_07794_),
    .C(_07797_),
    .A(net728),
    .Y(_02520_));
 sg13g2_nor2b_1 _27012_ (.A(_09876_),
    .B_N(_09861_),
    .Y(_07798_));
 sg13g2_buf_1 _27013_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07799_));
 sg13g2_o21ai_1 _27014_ (.B1(_07799_),
    .Y(_07800_),
    .A1(_07789_),
    .A2(_07798_));
 sg13g2_nand2b_1 _27015_ (.Y(_02521_),
    .B(_07800_),
    .A_N(_07790_));
 sg13g2_nor3_1 _27016_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09848_),
    .C(_06840_),
    .Y(_07801_));
 sg13g2_nand3_1 _27017_ (.B(_06749_),
    .C(_07801_),
    .A(_06726_),
    .Y(_07802_));
 sg13g2_or4_1 _27018_ (.A(_09933_),
    .B(net1138),
    .C(_09886_),
    .D(_07802_),
    .X(_07803_));
 sg13g2_a21oi_1 _27019_ (.A1(_09888_),
    .A2(_07803_),
    .Y(_02522_),
    .B1(_07782_));
 sg13g2_nand2_1 _27020_ (.Y(_07804_),
    .A(_10132_),
    .B(_06768_));
 sg13g2_nand2_1 _27021_ (.Y(_07805_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06773_));
 sg13g2_a21oi_1 _27022_ (.A1(_07804_),
    .A2(_07805_),
    .Y(_02523_),
    .B1(_07782_));
 sg13g2_a21oi_1 _27023_ (.A1(_10153_),
    .A2(net582),
    .Y(_07806_),
    .B1(net983));
 sg13g2_nand2_1 _27024_ (.Y(_07807_),
    .A(_06771_),
    .B(_07806_));
 sg13g2_o21ai_1 _27025_ (.B1(net797),
    .Y(_07808_),
    .A1(_07033_),
    .A2(_07807_));
 sg13g2_a21o_1 _27026_ (.A2(_06785_),
    .A1(\cpu.qspi.r_mask[1] ),
    .B1(_07808_),
    .X(_02524_));
 sg13g2_nor2_1 _27027_ (.A(_07033_),
    .B(_06799_),
    .Y(_07809_));
 sg13g2_a21oi_1 _27028_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06799_),
    .Y(_07810_),
    .B1(_07809_));
 sg13g2_nor2_1 _27029_ (.A(net558),
    .B(_07810_),
    .Y(_02525_));
 sg13g2_nand2_1 _27030_ (.Y(_07811_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06773_));
 sg13g2_nand2_1 _27031_ (.Y(_07812_),
    .A(_10129_),
    .B(_06768_));
 sg13g2_nand3_1 _27032_ (.B(_07811_),
    .C(_07812_),
    .A(net728),
    .Y(_02526_));
 sg13g2_nor2_1 _27033_ (.A(_07029_),
    .B(_07807_),
    .Y(_07813_));
 sg13g2_a21oi_1 _27034_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06785_),
    .Y(_07814_),
    .B1(_07813_));
 sg13g2_nor2_1 _27035_ (.A(net558),
    .B(_07814_),
    .Y(_02527_));
 sg13g2_nand2_1 _27036_ (.Y(_07815_),
    .A(_07029_),
    .B(_06796_));
 sg13g2_o21ai_1 _27037_ (.B1(_07815_),
    .Y(_07816_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06796_));
 sg13g2_nand2_1 _27038_ (.Y(_02528_),
    .A(net647),
    .B(_07816_));
 sg13g2_nand3_1 _27039_ (.B(net543),
    .C(_06771_),
    .A(_03532_),
    .Y(_07817_));
 sg13g2_buf_1 _27040_ (.A(_07817_),
    .X(_07818_));
 sg13g2_nor2_1 _27041_ (.A(net946),
    .B(_07818_),
    .Y(_07819_));
 sg13g2_nor2b_1 _27042_ (.A(_09865_),
    .B_N(_07818_),
    .Y(_07820_));
 sg13g2_o21ai_1 _27043_ (.B1(net647),
    .Y(_02541_),
    .A1(_07819_),
    .A2(_07820_));
 sg13g2_nor2_1 _27044_ (.A(_10088_),
    .B(_07818_),
    .Y(_07821_));
 sg13g2_nor2b_1 _27045_ (.A(_09864_),
    .B_N(_07818_),
    .Y(_07822_));
 sg13g2_o21ai_1 _27046_ (.B1(net647),
    .Y(_02542_),
    .A1(_07821_),
    .A2(_07822_));
 sg13g2_nand2b_1 _27047_ (.Y(_07823_),
    .B(_11937_),
    .A_N(_06809_));
 sg13g2_nor4_1 _27048_ (.A(_09933_),
    .B(net1138),
    .C(_06725_),
    .D(_06734_),
    .Y(_07824_));
 sg13g2_nand3_1 _27049_ (.B(_07823_),
    .C(_07824_),
    .A(_09839_),
    .Y(_07825_));
 sg13g2_buf_1 _27050_ (.A(_07825_),
    .X(_07826_));
 sg13g2_nor2b_1 _27051_ (.A(net3),
    .B_N(_07826_),
    .Y(_07827_));
 sg13g2_or4_1 _27052_ (.A(_09848_),
    .B(_09840_),
    .C(_11935_),
    .D(_06840_),
    .X(_07828_));
 sg13g2_nor3_1 _27053_ (.A(_11937_),
    .B(net1136),
    .C(_07828_),
    .Y(_07829_));
 sg13g2_nor4_1 _27054_ (.A(_11935_),
    .B(_06840_),
    .C(_07826_),
    .D(_07829_),
    .Y(_07830_));
 sg13g2_nor3_1 _27055_ (.A(net691),
    .B(_07827_),
    .C(_07830_),
    .Y(_02543_));
 sg13g2_nor2b_1 _27056_ (.A(net6),
    .B_N(_07826_),
    .Y(_07831_));
 sg13g2_nor4_1 _27057_ (.A(_11937_),
    .B(net1136),
    .C(_09881_),
    .D(_07828_),
    .Y(_07832_));
 sg13g2_nor3_1 _27058_ (.A(_11935_),
    .B(_07826_),
    .C(_07832_),
    .Y(_07833_));
 sg13g2_nor3_1 _27059_ (.A(net691),
    .B(_07831_),
    .C(_07833_),
    .Y(_02544_));
 sg13g2_nor2_1 _27060_ (.A(net1144),
    .B(_07045_),
    .Y(_07834_));
 sg13g2_a221oi_1 _27061_ (.B2(_09317_),
    .C1(_07834_),
    .B1(_09216_),
    .A1(net1145),
    .Y(_07835_),
    .A2(_09315_));
 sg13g2_buf_2 _27062_ (.A(_07835_),
    .X(_07836_));
 sg13g2_nand3_1 _27063_ (.B(net1064),
    .C(_07836_),
    .A(_09322_),
    .Y(_07837_));
 sg13g2_o21ai_1 _27064_ (.B1(_07837_),
    .Y(_07838_),
    .A1(_09322_),
    .A2(_07836_));
 sg13g2_nand2_1 _27065_ (.Y(_02550_),
    .A(net647),
    .B(_07838_));
 sg13g2_inv_1 _27066_ (.Y(_07839_),
    .A(_11973_));
 sg13g2_nand2_1 _27067_ (.Y(_07840_),
    .A(_09322_),
    .B(_07839_));
 sg13g2_a21oi_1 _27068_ (.A1(_07836_),
    .A2(_07840_),
    .Y(_07841_),
    .B1(_09323_));
 sg13g2_inv_1 _27069_ (.Y(_07842_),
    .A(_09322_));
 sg13g2_and4_1 _27070_ (.A(_07842_),
    .B(_09323_),
    .C(_07839_),
    .D(_07836_),
    .X(_07843_));
 sg13g2_o21ai_1 _27071_ (.B1(net647),
    .Y(_02551_),
    .A1(_07841_),
    .A2(_07843_));
 sg13g2_nor2_1 _27072_ (.A(_09322_),
    .B(_09323_),
    .Y(_07844_));
 sg13g2_or2_1 _27073_ (.X(_07845_),
    .B(_07844_),
    .A(_11973_));
 sg13g2_a21oi_1 _27074_ (.A1(_07836_),
    .A2(_07845_),
    .Y(_07846_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27075_ (.A(\cpu.spi.r_bits[2] ),
    .B(_07839_),
    .C(_07844_),
    .D(_07836_),
    .X(_07847_));
 sg13g2_o21ai_1 _27076_ (.B1(net647),
    .Y(_02552_),
    .A1(_07846_),
    .A2(_07847_));
 sg13g2_nor4_2 _27077_ (.A(_12009_),
    .B(_04910_),
    .C(_09294_),
    .Y(_07848_),
    .D(net542));
 sg13g2_nand2_1 _27078_ (.Y(_07849_),
    .A(net774),
    .B(_07848_));
 sg13g2_buf_4 _27079_ (.X(_07850_),
    .A(_07849_));
 sg13g2_mux2_1 _27080_ (.A0(net1057),
    .A1(\cpu.spi.r_clk_count[0][0] ),
    .S(_07850_),
    .X(_07851_));
 sg13g2_and2_1 _27081_ (.A(net693),
    .B(_07851_),
    .X(_02553_));
 sg13g2_mux2_1 _27082_ (.A0(net1049),
    .A1(\cpu.spi.r_clk_count[0][1] ),
    .S(_07850_),
    .X(_07852_));
 sg13g2_and2_1 _27083_ (.A(net693),
    .B(_07852_),
    .X(_02554_));
 sg13g2_mux2_1 _27084_ (.A0(net1048),
    .A1(\cpu.spi.r_clk_count[0][2] ),
    .S(_07850_),
    .X(_07853_));
 sg13g2_and2_1 _27085_ (.A(net693),
    .B(_07853_),
    .X(_02555_));
 sg13g2_buf_1 _27086_ (.A(net797),
    .X(_07854_));
 sg13g2_mux2_1 _27087_ (.A0(net1133),
    .A1(\cpu.spi.r_clk_count[0][3] ),
    .S(_07850_),
    .X(_07855_));
 sg13g2_and2_1 _27088_ (.A(net638),
    .B(_07855_),
    .X(_02556_));
 sg13g2_mux2_1 _27089_ (.A0(_10116_),
    .A1(\cpu.spi.r_clk_count[0][4] ),
    .S(_07850_),
    .X(_07856_));
 sg13g2_and2_1 _27090_ (.A(net638),
    .B(_07856_),
    .X(_02557_));
 sg13g2_mux2_1 _27091_ (.A0(_10122_),
    .A1(\cpu.spi.r_clk_count[0][5] ),
    .S(_07850_),
    .X(_07857_));
 sg13g2_and2_1 _27092_ (.A(net638),
    .B(_07857_),
    .X(_02558_));
 sg13g2_mux2_1 _27093_ (.A0(_10128_),
    .A1(\cpu.spi.r_clk_count[0][6] ),
    .S(_07850_),
    .X(_07858_));
 sg13g2_and2_1 _27094_ (.A(net638),
    .B(_07858_),
    .X(_02559_));
 sg13g2_mux2_1 _27095_ (.A0(_10131_),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(_07850_),
    .X(_07859_));
 sg13g2_and2_1 _27096_ (.A(net638),
    .B(_07859_),
    .X(_02560_));
 sg13g2_nand2_1 _27097_ (.Y(_07860_),
    .A(net517),
    .B(_07848_));
 sg13g2_buf_2 _27098_ (.A(_07860_),
    .X(_07861_));
 sg13g2_nand2_1 _27099_ (.Y(_07862_),
    .A(\cpu.spi.r_clk_count[1][0] ),
    .B(_07861_));
 sg13g2_and2_1 _27100_ (.A(_12011_),
    .B(_07848_),
    .X(_07863_));
 sg13g2_buf_2 _27101_ (.A(_07863_),
    .X(_07864_));
 sg13g2_nand2_1 _27102_ (.Y(_07865_),
    .A(net946),
    .B(_07864_));
 sg13g2_a21oi_1 _27103_ (.A1(_07862_),
    .A2(_07865_),
    .Y(_02561_),
    .B1(net555));
 sg13g2_nand2_1 _27104_ (.Y(_07866_),
    .A(\cpu.spi.r_clk_count[1][1] ),
    .B(_07861_));
 sg13g2_nand2_1 _27105_ (.Y(_07867_),
    .A(net1056),
    .B(_07864_));
 sg13g2_a21oi_1 _27106_ (.A1(_07866_),
    .A2(_07867_),
    .Y(_02562_),
    .B1(net555));
 sg13g2_nand2_1 _27107_ (.Y(_07868_),
    .A(\cpu.spi.r_clk_count[1][2] ),
    .B(_07861_));
 sg13g2_nand2_1 _27108_ (.Y(_07869_),
    .A(net1055),
    .B(_07864_));
 sg13g2_a21oi_1 _27109_ (.A1(_07868_),
    .A2(_07869_),
    .Y(_02563_),
    .B1(net555));
 sg13g2_nand2_1 _27110_ (.Y(_07870_),
    .A(\cpu.spi.r_clk_count[1][3] ),
    .B(_07861_));
 sg13g2_nand2_1 _27111_ (.Y(_07871_),
    .A(net1054),
    .B(_07864_));
 sg13g2_a21oi_1 _27112_ (.A1(_07870_),
    .A2(_07871_),
    .Y(_02564_),
    .B1(net555));
 sg13g2_nand2_1 _27113_ (.Y(_07872_),
    .A(\cpu.spi.r_clk_count[1][4] ),
    .B(_07861_));
 sg13g2_nand2_1 _27114_ (.Y(_07873_),
    .A(net1053),
    .B(_07864_));
 sg13g2_a21oi_1 _27115_ (.A1(_07872_),
    .A2(_07873_),
    .Y(_02565_),
    .B1(net555));
 sg13g2_nand2_1 _27116_ (.Y(_07874_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(_07861_));
 sg13g2_nand2_1 _27117_ (.Y(_07875_),
    .A(net1052),
    .B(_07864_));
 sg13g2_a21oi_1 _27118_ (.A1(_07874_),
    .A2(_07875_),
    .Y(_02566_),
    .B1(net555));
 sg13g2_nand2_1 _27119_ (.Y(_07876_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_07861_));
 sg13g2_nand2_1 _27120_ (.Y(_07877_),
    .A(net1051),
    .B(_07864_));
 sg13g2_buf_1 _27121_ (.A(_09368_),
    .X(_07878_));
 sg13g2_a21oi_1 _27122_ (.A1(_07876_),
    .A2(_07877_),
    .Y(_02567_),
    .B1(net554));
 sg13g2_nand2_1 _27123_ (.Y(_07879_),
    .A(\cpu.spi.r_clk_count[1][7] ),
    .B(_07861_));
 sg13g2_nand2_1 _27124_ (.Y(_07880_),
    .A(net1050),
    .B(_07864_));
 sg13g2_a21oi_1 _27125_ (.A1(_07879_),
    .A2(_07880_),
    .Y(_02568_),
    .B1(_07878_));
 sg13g2_or4_1 _27126_ (.A(net872),
    .B(net663),
    .C(_04910_),
    .D(_09294_),
    .X(_07881_));
 sg13g2_buf_1 _27127_ (.A(_07881_),
    .X(_07882_));
 sg13g2_nor2_1 _27128_ (.A(net542),
    .B(_07882_),
    .Y(_07883_));
 sg13g2_buf_2 _27129_ (.A(_07883_),
    .X(_07884_));
 sg13g2_nand2_1 _27130_ (.Y(_07885_),
    .A(net946),
    .B(_07884_));
 sg13g2_buf_1 _27131_ (.A(_07882_),
    .X(_07886_));
 sg13g2_o21ai_1 _27132_ (.B1(_04932_),
    .Y(_07887_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27133_ (.A1(_07885_),
    .A2(_07887_),
    .Y(_02569_),
    .B1(net554));
 sg13g2_nand2_1 _27134_ (.Y(_07888_),
    .A(net1056),
    .B(_07884_));
 sg13g2_o21ai_1 _27135_ (.B1(_05345_),
    .Y(_07889_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27136_ (.A1(_07888_),
    .A2(_07889_),
    .Y(_02570_),
    .B1(net554));
 sg13g2_nand2_1 _27137_ (.Y(_07890_),
    .A(net1055),
    .B(_07884_));
 sg13g2_o21ai_1 _27138_ (.B1(_05413_),
    .Y(_07891_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27139_ (.A1(_07890_),
    .A2(_07891_),
    .Y(_02571_),
    .B1(net554));
 sg13g2_nand2_1 _27140_ (.Y(_07892_),
    .A(net1054),
    .B(_07884_));
 sg13g2_o21ai_1 _27141_ (.B1(_05478_),
    .Y(_07893_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27142_ (.A1(_07892_),
    .A2(_07893_),
    .Y(_02572_),
    .B1(net554));
 sg13g2_nand2_1 _27143_ (.Y(_07894_),
    .A(net1053),
    .B(_07884_));
 sg13g2_o21ai_1 _27144_ (.B1(_05569_),
    .Y(_07895_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27145_ (.A1(_07894_),
    .A2(_07895_),
    .Y(_02573_),
    .B1(net554));
 sg13g2_nand2_1 _27146_ (.Y(_07896_),
    .A(net1052),
    .B(_07884_));
 sg13g2_o21ai_1 _27147_ (.B1(_05617_),
    .Y(_07897_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27148_ (.A1(_07896_),
    .A2(_07897_),
    .Y(_02574_),
    .B1(net554));
 sg13g2_nand2_1 _27149_ (.Y(_07898_),
    .A(net1051),
    .B(_07884_));
 sg13g2_o21ai_1 _27150_ (.B1(_05714_),
    .Y(_07899_),
    .A1(net438),
    .A2(net88));
 sg13g2_a21oi_1 _27151_ (.A1(_07898_),
    .A2(_07899_),
    .Y(_02575_),
    .B1(net554));
 sg13g2_nand2_1 _27152_ (.Y(_07900_),
    .A(net1050),
    .B(_07884_));
 sg13g2_o21ai_1 _27153_ (.B1(_05109_),
    .Y(_07901_),
    .A1(net438),
    .A2(_07882_));
 sg13g2_a21oi_1 _27154_ (.A1(_07900_),
    .A2(_07901_),
    .Y(_02576_),
    .B1(_07878_));
 sg13g2_o21ai_1 _27155_ (.B1(_09297_),
    .Y(_07902_),
    .A1(_09320_),
    .A2(_09288_));
 sg13g2_nor2_1 _27156_ (.A(_07010_),
    .B(_09320_),
    .Y(_07903_));
 sg13g2_nor3_1 _27157_ (.A(_09298_),
    .B(\cpu.spi.r_state[5] ),
    .C(_12043_),
    .Y(_07904_));
 sg13g2_buf_1 _27158_ (.A(_07904_),
    .X(_07905_));
 sg13g2_nand2_1 _27159_ (.Y(_07906_),
    .A(_07009_),
    .B(_07905_));
 sg13g2_nor2_1 _27160_ (.A(net1144),
    .B(_07906_),
    .Y(_07907_));
 sg13g2_a21oi_1 _27161_ (.A1(_09296_),
    .A2(_07903_),
    .Y(_07908_),
    .B1(_07907_));
 sg13g2_nand3_1 _27162_ (.B(_07902_),
    .C(_07908_),
    .A(_07000_),
    .Y(_07909_));
 sg13g2_buf_2 _27163_ (.A(_07909_),
    .X(_07910_));
 sg13g2_buf_1 _27164_ (.A(_07910_),
    .X(_07911_));
 sg13g2_buf_1 _27165_ (.A(_07906_),
    .X(_07912_));
 sg13g2_nand2b_1 _27166_ (.Y(_07913_),
    .B(net660),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _27167_ (.B1(_07913_),
    .Y(_07914_),
    .A1(net596),
    .A2(_04932_));
 sg13g2_mux2_1 _27168_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net660),
    .X(_07915_));
 sg13g2_nor2_1 _27169_ (.A(net661),
    .B(_07915_),
    .Y(_07916_));
 sg13g2_a21oi_1 _27170_ (.A1(net662),
    .A2(_07914_),
    .Y(_07917_),
    .B1(_07916_));
 sg13g2_nor2_1 _27171_ (.A(net491),
    .B(_07917_),
    .Y(_07918_));
 sg13g2_buf_1 _27172_ (.A(_07905_),
    .X(_07919_));
 sg13g2_mux2_1 _27173_ (.A0(_00316_),
    .A1(_00315_),
    .S(net1028),
    .X(_07920_));
 sg13g2_nor2_1 _27174_ (.A(net1028),
    .B(_04932_),
    .Y(_07921_));
 sg13g2_a21oi_1 _27175_ (.A1(net874),
    .A2(_00316_),
    .Y(_07922_),
    .B1(_07921_));
 sg13g2_nand2_1 _27176_ (.Y(_07923_),
    .A(net825),
    .B(_07922_));
 sg13g2_o21ai_1 _27177_ (.B1(_07923_),
    .Y(_07924_),
    .A1(net825),
    .A2(_07920_));
 sg13g2_nand2_1 _27178_ (.Y(_07925_),
    .A(net106),
    .B(_07924_));
 sg13g2_o21ai_1 _27179_ (.B1(_07925_),
    .Y(_07926_),
    .A1(_09207_),
    .A2(net87));
 sg13g2_nor2_1 _27180_ (.A(net388),
    .B(_07924_),
    .Y(_07927_));
 sg13g2_nor3_1 _27181_ (.A(_09207_),
    .B(_07919_),
    .C(_07927_),
    .Y(_07928_));
 sg13g2_a221oi_1 _27182_ (.B2(net1065),
    .C1(_07928_),
    .B1(_07926_),
    .A1(net944),
    .Y(_07929_),
    .A2(_07919_));
 sg13g2_nor3_1 _27183_ (.A(_07910_),
    .B(_07918_),
    .C(_07929_),
    .Y(_07930_));
 sg13g2_a21oi_1 _27184_ (.A1(_09207_),
    .A2(net30),
    .Y(_07931_),
    .B1(_07930_));
 sg13g2_nor2_1 _27185_ (.A(net558),
    .B(_07931_),
    .Y(_02577_));
 sg13g2_nand2b_1 _27186_ (.Y(_07932_),
    .B(net663),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _27187_ (.B1(_07932_),
    .Y(_07933_),
    .A1(net660),
    .A2(_05345_));
 sg13g2_mux2_1 _27188_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net748),
    .X(_07934_));
 sg13g2_nor2_1 _27189_ (.A(net747),
    .B(_07934_),
    .Y(_07935_));
 sg13g2_a21oi_1 _27190_ (.A1(net747),
    .A2(_07933_),
    .Y(_07936_),
    .B1(_07935_));
 sg13g2_o21ai_1 _27191_ (.B1(_09207_),
    .Y(_07937_),
    .A1(net491),
    .A2(_07936_));
 sg13g2_nor2_1 _27192_ (.A(_09316_),
    .B(_07937_),
    .Y(_07938_));
 sg13g2_o21ai_1 _27193_ (.B1(_09208_),
    .Y(_07939_),
    .A1(_07911_),
    .A2(_07938_));
 sg13g2_nor2_1 _27194_ (.A(net874),
    .B(_05345_),
    .Y(_07940_));
 sg13g2_a21oi_1 _27195_ (.A1(_11993_),
    .A2(_00095_),
    .Y(_07941_),
    .B1(_07940_));
 sg13g2_nand2_1 _27196_ (.Y(_07942_),
    .A(net1028),
    .B(_00094_));
 sg13g2_o21ai_1 _27197_ (.B1(_07942_),
    .Y(_07943_),
    .A1(net874),
    .A2(_05344_));
 sg13g2_nor2_1 _27198_ (.A(_07041_),
    .B(_07943_),
    .Y(_07944_));
 sg13g2_a21oi_1 _27199_ (.A1(_07041_),
    .A2(_07941_),
    .Y(_07945_),
    .B1(_07944_));
 sg13g2_nor2_1 _27200_ (.A(net106),
    .B(_09209_),
    .Y(_07946_));
 sg13g2_a21oi_1 _27201_ (.A1(net87),
    .A2(_07945_),
    .Y(_07947_),
    .B1(_07946_));
 sg13g2_nand2_1 _27202_ (.Y(_07948_),
    .A(_09207_),
    .B(_09208_));
 sg13g2_or2_1 _27203_ (.X(_07949_),
    .B(_09208_),
    .A(_09207_));
 sg13g2_a221oi_1 _27204_ (.B2(_07949_),
    .C1(_07905_),
    .B1(_07948_),
    .A1(net387),
    .Y(_07950_),
    .A2(_07945_));
 sg13g2_a221oi_1 _27205_ (.B2(net1065),
    .C1(_07950_),
    .B1(_07947_),
    .A1(net944),
    .Y(_07951_),
    .A2(net553));
 sg13g2_nor2_1 _27206_ (.A(_07910_),
    .B(_07951_),
    .Y(_07952_));
 sg13g2_o21ai_1 _27207_ (.B1(_07952_),
    .Y(_07953_),
    .A1(net491),
    .A2(_07936_));
 sg13g2_buf_1 _27208_ (.A(_09368_),
    .X(_07954_));
 sg13g2_a21oi_1 _27209_ (.A1(_07939_),
    .A2(_07953_),
    .Y(_02578_),
    .B1(net552));
 sg13g2_nand2b_1 _27210_ (.Y(_07955_),
    .B(net660),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _27211_ (.B1(_07955_),
    .Y(_07956_),
    .A1(net596),
    .A2(_05413_));
 sg13g2_mux2_1 _27212_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net663),
    .X(_07957_));
 sg13g2_nor2_1 _27213_ (.A(net661),
    .B(_07957_),
    .Y(_07958_));
 sg13g2_a21oi_1 _27214_ (.A1(net662),
    .A2(_07956_),
    .Y(_07959_),
    .B1(_07958_));
 sg13g2_nor2_1 _27215_ (.A(net491),
    .B(_07959_),
    .Y(_07960_));
 sg13g2_xnor2_1 _27216_ (.Y(_07961_),
    .A(\cpu.spi.r_count[2] ),
    .B(_09209_));
 sg13g2_nand2_1 _27217_ (.Y(_07962_),
    .A(net1028),
    .B(_00104_));
 sg13g2_o21ai_1 _27218_ (.B1(_07962_),
    .Y(_07963_),
    .A1(net873),
    .A2(_05412_));
 sg13g2_nor2_1 _27219_ (.A(net1029),
    .B(_05413_),
    .Y(_07964_));
 sg13g2_a21oi_1 _27220_ (.A1(_11979_),
    .A2(_00105_),
    .Y(_07965_),
    .B1(_07964_));
 sg13g2_nand2_1 _27221_ (.Y(_07966_),
    .A(_07040_),
    .B(_07965_));
 sg13g2_o21ai_1 _27222_ (.B1(_07966_),
    .Y(_07967_),
    .A1(net825),
    .A2(_07963_));
 sg13g2_nand2_1 _27223_ (.Y(_07968_),
    .A(net106),
    .B(_07967_));
 sg13g2_o21ai_1 _27224_ (.B1(_07968_),
    .Y(_07969_),
    .A1(net87),
    .A2(_07961_));
 sg13g2_nor2_1 _27225_ (.A(net388),
    .B(_07967_),
    .Y(_07970_));
 sg13g2_nor3_1 _27226_ (.A(net553),
    .B(_07970_),
    .C(_07961_),
    .Y(_07971_));
 sg13g2_a221oi_1 _27227_ (.B2(net1065),
    .C1(_07971_),
    .B1(_07969_),
    .A1(net944),
    .Y(_07972_),
    .A2(net553));
 sg13g2_nor3_1 _27228_ (.A(_07910_),
    .B(_07960_),
    .C(_07972_),
    .Y(_07973_));
 sg13g2_a21oi_1 _27229_ (.A1(\cpu.spi.r_count[2] ),
    .A2(net30),
    .Y(_07974_),
    .B1(_07973_));
 sg13g2_nor2_1 _27230_ (.A(net558),
    .B(_07974_),
    .Y(_02579_));
 sg13g2_nand2b_1 _27231_ (.Y(_07975_),
    .B(net660),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _27232_ (.B1(_07975_),
    .Y(_07976_),
    .A1(net596),
    .A2(_05478_));
 sg13g2_mux2_1 _27233_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net663),
    .X(_07977_));
 sg13g2_nor2_1 _27234_ (.A(net661),
    .B(_07977_),
    .Y(_07978_));
 sg13g2_a21oi_1 _27235_ (.A1(net662),
    .A2(_07976_),
    .Y(_07979_),
    .B1(_07978_));
 sg13g2_nor2_1 _27236_ (.A(net491),
    .B(_07979_),
    .Y(_07980_));
 sg13g2_xor2_1 _27237_ (.B(_09210_),
    .A(_09206_),
    .X(_07981_));
 sg13g2_nand2_1 _27238_ (.Y(_07982_),
    .A(net1028),
    .B(_00114_));
 sg13g2_o21ai_1 _27239_ (.B1(_07982_),
    .Y(_07983_),
    .A1(net873),
    .A2(_05476_));
 sg13g2_nor2_1 _27240_ (.A(net1029),
    .B(_05478_),
    .Y(_07984_));
 sg13g2_a21oi_1 _27241_ (.A1(net874),
    .A2(_00115_),
    .Y(_07985_),
    .B1(_07984_));
 sg13g2_nand2_1 _27242_ (.Y(_07986_),
    .A(net943),
    .B(_07985_));
 sg13g2_o21ai_1 _27243_ (.B1(_07986_),
    .Y(_07987_),
    .A1(net825),
    .A2(_07983_));
 sg13g2_nand2_1 _27244_ (.Y(_07988_),
    .A(net106),
    .B(_07987_));
 sg13g2_o21ai_1 _27245_ (.B1(_07988_),
    .Y(_07989_),
    .A1(net87),
    .A2(_07981_));
 sg13g2_nor2_1 _27246_ (.A(net388),
    .B(_07987_),
    .Y(_07990_));
 sg13g2_nor3_1 _27247_ (.A(net553),
    .B(_07981_),
    .C(_07990_),
    .Y(_07991_));
 sg13g2_a221oi_1 _27248_ (.B2(net1065),
    .C1(_07991_),
    .B1(_07989_),
    .A1(net944),
    .Y(_07992_),
    .A2(net553));
 sg13g2_nor3_1 _27249_ (.A(_07910_),
    .B(_07980_),
    .C(_07992_),
    .Y(_07993_));
 sg13g2_a21oi_1 _27250_ (.A1(_09206_),
    .A2(net30),
    .Y(_07994_),
    .B1(_07993_));
 sg13g2_nor2_1 _27251_ (.A(net558),
    .B(_07994_),
    .Y(_02580_));
 sg13g2_nand2b_1 _27252_ (.Y(_07995_),
    .B(net660),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _27253_ (.B1(_07995_),
    .Y(_07996_),
    .A1(net596),
    .A2(_05569_));
 sg13g2_mux2_1 _27254_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net663),
    .X(_07997_));
 sg13g2_nor2_1 _27255_ (.A(net661),
    .B(_07997_),
    .Y(_07998_));
 sg13g2_a21oi_1 _27256_ (.A1(net661),
    .A2(_07996_),
    .Y(_07999_),
    .B1(_07998_));
 sg13g2_nor2_1 _27257_ (.A(net491),
    .B(_07999_),
    .Y(_08000_));
 sg13g2_nor2_1 _27258_ (.A(_09206_),
    .B(_09210_),
    .Y(_08001_));
 sg13g2_xnor2_1 _27259_ (.Y(_08002_),
    .A(\cpu.spi.r_count[4] ),
    .B(_08001_));
 sg13g2_nand2_1 _27260_ (.Y(_08003_),
    .A(net1028),
    .B(_00125_));
 sg13g2_o21ai_1 _27261_ (.B1(_08003_),
    .Y(_08004_),
    .A1(net873),
    .A2(_05568_));
 sg13g2_nor2_1 _27262_ (.A(net1029),
    .B(_05569_),
    .Y(_08005_));
 sg13g2_a21oi_1 _27263_ (.A1(net874),
    .A2(_00126_),
    .Y(_08006_),
    .B1(_08005_));
 sg13g2_nand2_1 _27264_ (.Y(_08007_),
    .A(net943),
    .B(_08006_));
 sg13g2_o21ai_1 _27265_ (.B1(_08007_),
    .Y(_08008_),
    .A1(net825),
    .A2(_08004_));
 sg13g2_nand2_1 _27266_ (.Y(_08009_),
    .A(net106),
    .B(_08008_));
 sg13g2_o21ai_1 _27267_ (.B1(_08009_),
    .Y(_08010_),
    .A1(net87),
    .A2(_08002_));
 sg13g2_nor2_1 _27268_ (.A(net388),
    .B(_08008_),
    .Y(_08011_));
 sg13g2_nor3_1 _27269_ (.A(_07905_),
    .B(_08002_),
    .C(_08011_),
    .Y(_08012_));
 sg13g2_a221oi_1 _27270_ (.B2(net1065),
    .C1(_08012_),
    .B1(_08010_),
    .A1(net944),
    .Y(_08013_),
    .A2(net553));
 sg13g2_nor3_1 _27271_ (.A(_07910_),
    .B(_08000_),
    .C(_08013_),
    .Y(_08014_));
 sg13g2_a21oi_1 _27272_ (.A1(\cpu.spi.r_count[4] ),
    .A2(net30),
    .Y(_08015_),
    .B1(_08014_));
 sg13g2_nor2_1 _27273_ (.A(net558),
    .B(_08015_),
    .Y(_02581_));
 sg13g2_nand2b_1 _27274_ (.Y(_08016_),
    .B(_12015_),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _27275_ (.B1(_08016_),
    .Y(_08017_),
    .A1(_12011_),
    .A2(_05617_));
 sg13g2_mux2_1 _27276_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(_12004_),
    .X(_08018_));
 sg13g2_nor2_1 _27277_ (.A(_12014_),
    .B(_08018_),
    .Y(_08019_));
 sg13g2_a21oi_1 _27278_ (.A1(net661),
    .A2(_08017_),
    .Y(_08020_),
    .B1(_08019_));
 sg13g2_nand2_1 _27279_ (.Y(_08021_),
    .A(_11977_),
    .B(_00132_));
 sg13g2_o21ai_1 _27280_ (.B1(_08021_),
    .Y(_08022_),
    .A1(_11978_),
    .A2(_05616_));
 sg13g2_nor2_1 _27281_ (.A(_11977_),
    .B(_05617_),
    .Y(_08023_));
 sg13g2_a21oi_1 _27282_ (.A1(net1029),
    .A2(_00133_),
    .Y(_08024_),
    .B1(_08023_));
 sg13g2_nand2_1 _27283_ (.Y(_08025_),
    .A(net943),
    .B(_08024_));
 sg13g2_o21ai_1 _27284_ (.B1(_08025_),
    .Y(_08026_),
    .A1(net943),
    .A2(_08022_));
 sg13g2_xnor2_1 _27285_ (.Y(_08027_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09211_));
 sg13g2_nor2_1 _27286_ (.A(_07905_),
    .B(_08027_),
    .Y(_08028_));
 sg13g2_o21ai_1 _27287_ (.B1(_08028_),
    .Y(_08029_),
    .A1(net388),
    .A2(_08026_));
 sg13g2_nand2_1 _27288_ (.Y(_08030_),
    .A(net106),
    .B(_08026_));
 sg13g2_o21ai_1 _27289_ (.B1(_08030_),
    .Y(_08031_),
    .A1(net106),
    .A2(_08027_));
 sg13g2_nand2_1 _27290_ (.Y(_08032_),
    .A(net1145),
    .B(_08031_));
 sg13g2_nand3_1 _27291_ (.B(_08029_),
    .C(_08032_),
    .A(_07912_),
    .Y(_08033_));
 sg13g2_o21ai_1 _27292_ (.B1(_08033_),
    .Y(_08034_),
    .A1(_07912_),
    .A2(_08020_));
 sg13g2_nor2_1 _27293_ (.A(net30),
    .B(_08034_),
    .Y(_08035_));
 sg13g2_a21oi_1 _27294_ (.A1(\cpu.spi.r_count[5] ),
    .A2(net30),
    .Y(_08036_),
    .B1(_08035_));
 sg13g2_nor2_1 _27295_ (.A(net558),
    .B(_08036_),
    .Y(_02582_));
 sg13g2_nand2b_1 _27296_ (.Y(_08037_),
    .B(net660),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _27297_ (.B1(_08037_),
    .Y(_08038_),
    .A1(net596),
    .A2(_05714_));
 sg13g2_mux2_1 _27298_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net663),
    .X(_08039_));
 sg13g2_nor2_1 _27299_ (.A(net661),
    .B(_08039_),
    .Y(_08040_));
 sg13g2_a21oi_1 _27300_ (.A1(net661),
    .A2(_08038_),
    .Y(_08041_),
    .B1(_08040_));
 sg13g2_nor2_1 _27301_ (.A(net491),
    .B(_08041_),
    .Y(_08042_));
 sg13g2_xnor2_1 _27302_ (.Y(_08043_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09212_));
 sg13g2_nand2_1 _27303_ (.Y(_08044_),
    .A(net1028),
    .B(_00144_));
 sg13g2_o21ai_1 _27304_ (.B1(_08044_),
    .Y(_08045_),
    .A1(net874),
    .A2(_05713_));
 sg13g2_nor2_1 _27305_ (.A(net1029),
    .B(_05714_),
    .Y(_08046_));
 sg13g2_a21oi_1 _27306_ (.A1(net874),
    .A2(_00145_),
    .Y(_08047_),
    .B1(_08046_));
 sg13g2_nand2_1 _27307_ (.Y(_08048_),
    .A(net943),
    .B(_08047_));
 sg13g2_o21ai_1 _27308_ (.B1(_08048_),
    .Y(_08049_),
    .A1(net825),
    .A2(_08045_));
 sg13g2_nand2_1 _27309_ (.Y(_08050_),
    .A(net106),
    .B(_08049_));
 sg13g2_o21ai_1 _27310_ (.B1(_08050_),
    .Y(_08051_),
    .A1(net87),
    .A2(_08043_));
 sg13g2_nor2_1 _27311_ (.A(net388),
    .B(_08049_),
    .Y(_08052_));
 sg13g2_nor3_1 _27312_ (.A(_07905_),
    .B(_08052_),
    .C(_08043_),
    .Y(_08053_));
 sg13g2_a221oi_1 _27313_ (.B2(net1065),
    .C1(_08053_),
    .B1(_08051_),
    .A1(net944),
    .Y(_08054_),
    .A2(net553));
 sg13g2_nor3_1 _27314_ (.A(_07910_),
    .B(_08042_),
    .C(_08054_),
    .Y(_08055_));
 sg13g2_a21oi_1 _27315_ (.A1(\cpu.spi.r_count[6] ),
    .A2(net30),
    .Y(_08056_),
    .B1(_08055_));
 sg13g2_nor2_1 _27316_ (.A(net692),
    .B(_08056_),
    .Y(_02583_));
 sg13g2_nand2b_1 _27317_ (.Y(_08057_),
    .B(_12004_),
    .A_N(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_o21ai_1 _27318_ (.B1(_08057_),
    .Y(_08058_),
    .A1(net660),
    .A2(_05109_));
 sg13g2_mux2_1 _27319_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(net748),
    .X(_08059_));
 sg13g2_nor2_1 _27320_ (.A(net747),
    .B(_08059_),
    .Y(_08060_));
 sg13g2_a21oi_1 _27321_ (.A1(net747),
    .A2(_08058_),
    .Y(_08061_),
    .B1(_08060_));
 sg13g2_nor2_1 _27322_ (.A(_07906_),
    .B(_08061_),
    .Y(_08062_));
 sg13g2_nor3_1 _27323_ (.A(_09214_),
    .B(_09316_),
    .C(_08062_),
    .Y(_08063_));
 sg13g2_o21ai_1 _27324_ (.B1(_09205_),
    .Y(_08064_),
    .A1(net30),
    .A2(_08063_));
 sg13g2_nor2_1 _27325_ (.A(net1029),
    .B(_05109_),
    .Y(_08065_));
 sg13g2_a21oi_1 _27326_ (.A1(_11979_),
    .A2(_00157_),
    .Y(_08066_),
    .B1(_08065_));
 sg13g2_nand2_1 _27327_ (.Y(_08067_),
    .A(_11977_),
    .B(_00156_));
 sg13g2_o21ai_1 _27328_ (.B1(_08067_),
    .Y(_08068_),
    .A1(net1029),
    .A2(_05108_));
 sg13g2_nor2_1 _27329_ (.A(_07040_),
    .B(_08068_),
    .Y(_08069_));
 sg13g2_a21oi_1 _27330_ (.A1(net943),
    .A2(_08066_),
    .Y(_08070_),
    .B1(_08069_));
 sg13g2_nor2_1 _27331_ (.A(_09359_),
    .B(net387),
    .Y(_08071_));
 sg13g2_a21oi_1 _27332_ (.A1(_09359_),
    .A2(_08070_),
    .Y(_08072_),
    .B1(_08071_));
 sg13g2_nor2_1 _27333_ (.A(_09205_),
    .B(_08070_),
    .Y(_08073_));
 sg13g2_nor2b_1 _27334_ (.A(_09214_),
    .B_N(_09205_),
    .Y(_08074_));
 sg13g2_a21oi_1 _27335_ (.A1(_09214_),
    .A2(_08073_),
    .Y(_08075_),
    .B1(_08074_));
 sg13g2_o21ai_1 _27336_ (.B1(net491),
    .Y(_08076_),
    .A1(net553),
    .A2(_08075_));
 sg13g2_a21oi_1 _27337_ (.A1(net1065),
    .A2(_08072_),
    .Y(_08077_),
    .B1(_08076_));
 sg13g2_or3_1 _27338_ (.A(_07911_),
    .B(_08062_),
    .C(_08077_),
    .X(_08078_));
 sg13g2_a21oi_1 _27339_ (.A1(_08064_),
    .A2(_08078_),
    .Y(_02584_),
    .B1(net552));
 sg13g2_buf_1 _27340_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08079_));
 sg13g2_inv_1 _27341_ (.Y(_08080_),
    .A(_08079_));
 sg13g2_a21oi_1 _27342_ (.A1(_09315_),
    .A2(_09288_),
    .Y(_08081_),
    .B1(net944));
 sg13g2_or2_1 _27343_ (.X(_08082_),
    .B(net1145),
    .A(_09298_));
 sg13g2_buf_1 _27344_ (.A(_08082_),
    .X(_08083_));
 sg13g2_nand2_1 _27345_ (.Y(_08084_),
    .A(_09320_),
    .B(_08083_));
 sg13g2_nor3_1 _27346_ (.A(_09357_),
    .B(_09320_),
    .C(_08083_),
    .Y(_08085_));
 sg13g2_a21oi_1 _27347_ (.A1(net943),
    .A2(net873),
    .Y(_08086_),
    .B1(_09216_));
 sg13g2_nor3_1 _27348_ (.A(_00280_),
    .B(_08085_),
    .C(_08086_),
    .Y(_08087_));
 sg13g2_a21oi_1 _27349_ (.A1(_00280_),
    .A2(_08084_),
    .Y(_08088_),
    .B1(_08087_));
 sg13g2_nand2b_1 _27350_ (.Y(_08089_),
    .B(_08088_),
    .A_N(_08081_));
 sg13g2_buf_1 _27351_ (.A(_08089_),
    .X(_08090_));
 sg13g2_nor3_1 _27352_ (.A(net825),
    .B(net873),
    .C(_08090_),
    .Y(_08091_));
 sg13g2_inv_1 _27353_ (.Y(_08092_),
    .A(_08090_));
 sg13g2_a21oi_1 _27354_ (.A1(_08083_),
    .A2(_08092_),
    .Y(_08093_),
    .B1(net795));
 sg13g2_o21ai_1 _27355_ (.B1(_08093_),
    .Y(_02585_),
    .A1(_08080_),
    .A2(_08091_));
 sg13g2_nand2_1 _27356_ (.Y(_08094_),
    .A(_11976_),
    .B(net873));
 sg13g2_buf_1 _27357_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08095_));
 sg13g2_o21ai_1 _27358_ (.B1(_08095_),
    .Y(_08096_),
    .A1(_08090_),
    .A2(_08094_));
 sg13g2_nand2_1 _27359_ (.Y(_02586_),
    .A(_08093_),
    .B(_08096_));
 sg13g2_buf_1 _27360_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08097_));
 sg13g2_inv_1 _27361_ (.Y(_08098_),
    .A(_08097_));
 sg13g2_nor3_1 _27362_ (.A(_11976_),
    .B(net873),
    .C(_08090_),
    .Y(_08099_));
 sg13g2_o21ai_1 _27363_ (.B1(_08093_),
    .Y(_02587_),
    .A1(_08098_),
    .A2(_08099_));
 sg13g2_nand2_1 _27364_ (.Y(_08100_),
    .A(_09320_),
    .B(_09352_));
 sg13g2_nor3_1 _27365_ (.A(_07010_),
    .B(_09296_),
    .C(_09288_),
    .Y(_08101_));
 sg13g2_a221oi_1 _27366_ (.B2(_09317_),
    .C1(_08101_),
    .B1(_08100_),
    .A1(_09300_),
    .Y(_08102_),
    .A2(_09301_));
 sg13g2_buf_1 _27367_ (.A(_08102_),
    .X(_08103_));
 sg13g2_o21ai_1 _27368_ (.B1(_08103_),
    .Y(_08104_),
    .A1(net1144),
    .A2(net870));
 sg13g2_a22oi_1 _27369_ (.Y(_08105_),
    .B1(_08104_),
    .B2(_09275_),
    .A2(_08103_),
    .A1(net1064));
 sg13g2_nor2_1 _27370_ (.A(net692),
    .B(_08105_),
    .Y(_02596_));
 sg13g2_nor4_2 _27371_ (.A(_12009_),
    .B(_04910_),
    .C(net581),
    .Y(_08106_),
    .D(_09294_));
 sg13g2_and2_1 _27372_ (.A(net774),
    .B(_08106_),
    .X(_08107_));
 sg13g2_buf_1 _27373_ (.A(_08107_),
    .X(_08108_));
 sg13g2_nor2b_1 _27374_ (.A(_08108_),
    .B_N(\cpu.spi.r_mode[0][0] ),
    .Y(_08109_));
 sg13g2_a21oi_1 _27375_ (.A1(net946),
    .A2(_08108_),
    .Y(_08110_),
    .B1(_08109_));
 sg13g2_nor2_1 _27376_ (.A(net692),
    .B(_08110_),
    .Y(_02597_));
 sg13g2_nor2b_1 _27377_ (.A(_08108_),
    .B_N(_11991_),
    .Y(_08111_));
 sg13g2_a21oi_1 _27378_ (.A1(net1056),
    .A2(_08108_),
    .Y(_08112_),
    .B1(_08111_));
 sg13g2_nor2_1 _27379_ (.A(net692),
    .B(_08112_),
    .Y(_02598_));
 sg13g2_nand2_2 _27380_ (.Y(_08113_),
    .A(net517),
    .B(_08106_));
 sg13g2_mux2_1 _27381_ (.A0(net1057),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_08113_),
    .X(_08114_));
 sg13g2_and2_1 _27382_ (.A(net638),
    .B(_08114_),
    .X(_02599_));
 sg13g2_mux2_1 _27383_ (.A0(net1049),
    .A1(_11992_),
    .S(_08113_),
    .X(_08115_));
 sg13g2_and2_1 _27384_ (.A(net638),
    .B(_08115_),
    .X(_02600_));
 sg13g2_o21ai_1 _27385_ (.B1(\cpu.spi.r_mode[2][0] ),
    .Y(_08116_),
    .A1(net581),
    .A2(_07886_));
 sg13g2_nor2_1 _27386_ (.A(net581),
    .B(_07882_),
    .Y(_08117_));
 sg13g2_nand2_1 _27387_ (.Y(_08118_),
    .A(net946),
    .B(_08117_));
 sg13g2_a21oi_1 _27388_ (.A1(_08116_),
    .A2(_08118_),
    .Y(_02601_),
    .B1(net552));
 sg13g2_o21ai_1 _27389_ (.B1(_11996_),
    .Y(_08119_),
    .A1(net581),
    .A2(net88));
 sg13g2_nand2_1 _27390_ (.Y(_08120_),
    .A(net1056),
    .B(_08117_));
 sg13g2_a21oi_1 _27391_ (.A1(_08119_),
    .A2(_08120_),
    .Y(_02602_),
    .B1(net552));
 sg13g2_nand2b_1 _27392_ (.Y(_08121_),
    .B(_09217_),
    .A_N(\cpu.spi.r_ready ));
 sg13g2_nor2b_1 _27393_ (.A(_09298_),
    .B_N(_07834_),
    .Y(_08122_));
 sg13g2_nor2b_1 _27394_ (.A(_08122_),
    .B_N(_08103_),
    .Y(_08123_));
 sg13g2_nand3b_1 _27395_ (.B(_09316_),
    .C(_08123_),
    .Y(_08124_),
    .A_N(_09298_));
 sg13g2_a21oi_1 _27396_ (.A1(_08121_),
    .A2(_08124_),
    .Y(_08125_),
    .B1(net1064));
 sg13g2_nor2_1 _27397_ (.A(\cpu.spi.r_ready ),
    .B(_08123_),
    .Y(_08126_));
 sg13g2_o21ai_1 _27398_ (.B1(net647),
    .Y(_02611_),
    .A1(_08125_),
    .A2(_08126_));
 sg13g2_nand2_1 _27399_ (.Y(_08127_),
    .A(_09355_),
    .B(_07836_));
 sg13g2_nand2_1 _27400_ (.Y(_08128_),
    .A(\cpu.spi.r_searching ),
    .B(_08127_));
 sg13g2_o21ai_1 _27401_ (.B1(_12030_),
    .Y(_08129_),
    .A1(net624),
    .A2(net581));
 sg13g2_or2_1 _27402_ (.X(_08130_),
    .B(_08129_),
    .A(_08127_));
 sg13g2_a21oi_1 _27403_ (.A1(_08128_),
    .A2(_08130_),
    .Y(_02612_),
    .B1(net552));
 sg13g2_nor2b_1 _27404_ (.A(_08108_),
    .B_N(\cpu.spi.r_src[0] ),
    .Y(_08131_));
 sg13g2_a21oi_1 _27405_ (.A1(net1055),
    .A2(_08108_),
    .Y(_08132_),
    .B1(_08131_));
 sg13g2_nor2_1 _27406_ (.A(net692),
    .B(_08132_),
    .Y(_02615_));
 sg13g2_mux2_1 _27407_ (.A0(_10164_),
    .A1(\cpu.spi.r_src[1] ),
    .S(_08113_),
    .X(_08133_));
 sg13g2_and2_1 _27408_ (.A(net638),
    .B(_08133_),
    .X(_02616_));
 sg13g2_o21ai_1 _27409_ (.B1(_11985_),
    .Y(_08134_),
    .A1(net581),
    .A2(_07886_));
 sg13g2_nand2_1 _27410_ (.Y(_08135_),
    .A(net1055),
    .B(_08117_));
 sg13g2_a21oi_1 _27411_ (.A1(_08134_),
    .A2(_08135_),
    .Y(_02617_),
    .B1(net552));
 sg13g2_and2_1 _27412_ (.A(net412),
    .B(_07105_),
    .X(_08136_));
 sg13g2_buf_2 _27413_ (.A(_08136_),
    .X(_08137_));
 sg13g2_nand2_1 _27414_ (.Y(_08138_),
    .A(net901),
    .B(_08137_));
 sg13g2_nand2_1 _27415_ (.Y(_08139_),
    .A(net412),
    .B(_07105_));
 sg13g2_buf_2 _27416_ (.A(_08139_),
    .X(_08140_));
 sg13g2_nand2_1 _27417_ (.Y(_08141_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08140_));
 sg13g2_nand3_1 _27418_ (.B(_08138_),
    .C(_08141_),
    .A(net728),
    .Y(_02634_));
 sg13g2_nand2_2 _27419_ (.Y(_08142_),
    .A(net411),
    .B(_07105_));
 sg13g2_mux2_1 _27420_ (.A0(net1048),
    .A1(_09976_),
    .S(_08142_),
    .X(_08143_));
 sg13g2_and2_1 _27421_ (.A(_07854_),
    .B(_08143_),
    .X(_02635_));
 sg13g2_mux2_1 _27422_ (.A0(net1133),
    .A1(\cpu.uart.r_div_value[11] ),
    .S(_08142_),
    .X(_08144_));
 sg13g2_and2_1 _27423_ (.A(_07854_),
    .B(_08144_),
    .X(_02636_));
 sg13g2_nand2_1 _27424_ (.Y(_08145_),
    .A(_10088_),
    .B(_08137_));
 sg13g2_nand2_1 _27425_ (.Y(_08146_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27426_ (.A1(_08145_),
    .A2(_08146_),
    .Y(_02637_),
    .B1(net552));
 sg13g2_nand2_1 _27427_ (.Y(_08147_),
    .A(_10106_),
    .B(_08137_));
 sg13g2_nand2_1 _27428_ (.Y(_08148_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27429_ (.A1(_08147_),
    .A2(_08148_),
    .Y(_02638_),
    .B1(net552));
 sg13g2_nand2_1 _27430_ (.Y(_08149_),
    .A(_10111_),
    .B(_08137_));
 sg13g2_nand2_1 _27431_ (.Y(_08150_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27432_ (.A1(_08149_),
    .A2(_08150_),
    .Y(_02639_),
    .B1(_07954_));
 sg13g2_nand2_1 _27433_ (.Y(_08151_),
    .A(net1053),
    .B(_08137_));
 sg13g2_nand2_1 _27434_ (.Y(_08152_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27435_ (.A1(_08151_),
    .A2(_08152_),
    .Y(_02640_),
    .B1(_07954_));
 sg13g2_nand2_1 _27436_ (.Y(_08153_),
    .A(_10123_),
    .B(_08137_));
 sg13g2_nand2_1 _27437_ (.Y(_08154_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27438_ (.A1(_08153_),
    .A2(_08154_),
    .Y(_02641_),
    .B1(net682));
 sg13g2_nand2_1 _27439_ (.Y(_08155_),
    .A(net1051),
    .B(_08137_));
 sg13g2_nand2_1 _27440_ (.Y(_08156_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27441_ (.A1(_08155_),
    .A2(_08156_),
    .Y(_02642_),
    .B1(net682));
 sg13g2_nand2_1 _27442_ (.Y(_08157_),
    .A(net1050),
    .B(_08137_));
 sg13g2_nand2_1 _27443_ (.Y(_08158_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08140_));
 sg13g2_a21oi_1 _27444_ (.A1(_08157_),
    .A2(_08158_),
    .Y(_02643_),
    .B1(net682));
 sg13g2_mux2_1 _27445_ (.A0(_10081_),
    .A1(\cpu.uart.r_div_value[8] ),
    .S(_08142_),
    .X(_08159_));
 sg13g2_and2_1 _27446_ (.A(net750),
    .B(_08159_),
    .X(_02644_));
 sg13g2_mux2_1 _27447_ (.A0(net1049),
    .A1(\cpu.uart.r_div_value[9] ),
    .S(_08142_),
    .X(_08160_));
 sg13g2_and2_1 _27448_ (.A(net750),
    .B(_08160_),
    .X(_02645_));
 sg13g2_nand3_1 _27449_ (.B(net415),
    .C(_07105_),
    .A(_10144_),
    .Y(_08161_));
 sg13g2_nor2_1 _27450_ (.A(net1071),
    .B(_04851_),
    .Y(_08162_));
 sg13g2_nand4_1 _27451_ (.B(_07103_),
    .C(_05045_),
    .A(net662),
    .Y(_08163_),
    .D(_08162_));
 sg13g2_or2_1 _27452_ (.X(_08164_),
    .B(_08163_),
    .A(_09287_));
 sg13g2_nand4_1 _27453_ (.B(net797),
    .C(_08161_),
    .A(_09279_),
    .Y(_08165_),
    .D(_08164_));
 sg13g2_nand2b_1 _27454_ (.Y(_02669_),
    .B(_08165_),
    .A_N(net175));
 sg13g2_nand2_1 _27455_ (.Y(_08166_),
    .A(net504),
    .B(_07105_));
 sg13g2_mux2_1 _27456_ (.A0(_10144_),
    .A1(\cpu.uart.r_r_invert ),
    .S(_08166_),
    .X(_08167_));
 sg13g2_and2_1 _27457_ (.A(net750),
    .B(_08167_),
    .X(_02670_));
 sg13g2_a21oi_1 _27458_ (.A1(_07089_),
    .A2(_09954_),
    .Y(_08168_),
    .B1(net1106));
 sg13g2_a21oi_1 _27459_ (.A1(_07090_),
    .A2(_09954_),
    .Y(_08169_),
    .B1(_07161_));
 sg13g2_a221oi_1 _27460_ (.B2(_08168_),
    .C1(_08169_),
    .B1(_07088_),
    .A1(_07087_),
    .Y(_08170_),
    .A2(_07083_));
 sg13g2_a21oi_1 _27461_ (.A1(_07081_),
    .A2(_08170_),
    .Y(_08171_),
    .B1(_07158_));
 sg13g2_buf_2 _27462_ (.A(_08171_),
    .X(_08172_));
 sg13g2_o21ai_1 _27463_ (.B1(_08172_),
    .Y(_08173_),
    .A1(net941),
    .A2(_07161_));
 sg13g2_xnor2_1 _27464_ (.Y(_08174_),
    .A(_07090_),
    .B(_08173_));
 sg13g2_nor2_1 _27465_ (.A(_09364_),
    .B(_08174_),
    .Y(_02673_));
 sg13g2_o21ai_1 _27466_ (.B1(_08172_),
    .Y(_08175_),
    .A1(_07089_),
    .A2(net942));
 sg13g2_nand2_1 _27467_ (.Y(_08176_),
    .A(net1105),
    .B(_08175_));
 sg13g2_nand2b_1 _27468_ (.Y(_08177_),
    .B(net941),
    .A_N(net942));
 sg13g2_o21ai_1 _27469_ (.B1(_08177_),
    .Y(_08178_),
    .A1(net941),
    .A2(_07160_));
 sg13g2_nand3_1 _27470_ (.B(_08172_),
    .C(_08178_),
    .A(_07159_),
    .Y(_08179_));
 sg13g2_a21oi_1 _27471_ (.A1(_08176_),
    .A2(_08179_),
    .Y(_02674_),
    .B1(net682));
 sg13g2_nand2_1 _27472_ (.Y(_08180_),
    .A(_07089_),
    .B(net1105));
 sg13g2_nor3_1 _27473_ (.A(net941),
    .B(net942),
    .C(_08180_),
    .Y(_08181_));
 sg13g2_o21ai_1 _27474_ (.B1(_08172_),
    .Y(_08182_),
    .A1(net942),
    .A2(_07169_));
 sg13g2_a22oi_1 _27475_ (.Y(_08183_),
    .B1(_08182_),
    .B2(net941),
    .A2(_08181_),
    .A1(_08172_));
 sg13g2_nor2_1 _27476_ (.A(_09364_),
    .B(_08183_),
    .Y(_02675_));
 sg13g2_a21oi_1 _27477_ (.A1(_07169_),
    .A2(_08172_),
    .Y(_08184_),
    .B1(net942));
 sg13g2_nor2b_1 _27478_ (.A(net941),
    .B_N(net1105),
    .Y(_08185_));
 sg13g2_a21oi_1 _27479_ (.A1(_08172_),
    .A2(_08185_),
    .Y(_08186_),
    .B1(_09368_));
 sg13g2_nor2b_1 _27480_ (.A(_08184_),
    .B_N(_08186_),
    .Y(_02676_));
 sg13g2_nor2_1 _27481_ (.A(net940),
    .B(_07184_),
    .Y(_08187_));
 sg13g2_o21ai_1 _27482_ (.B1(_08187_),
    .Y(_08188_),
    .A1(_09278_),
    .A2(_07117_));
 sg13g2_a21oi_1 _27483_ (.A1(_10080_),
    .A2(net415),
    .Y(_08189_),
    .B1(net413));
 sg13g2_o21ai_1 _27484_ (.B1(net542),
    .Y(_08190_),
    .A1(_00225_),
    .A2(net582));
 sg13g2_nand3_1 _27485_ (.B(_07201_),
    .C(_08190_),
    .A(net912),
    .Y(_08191_));
 sg13g2_o21ai_1 _27486_ (.B1(_08191_),
    .Y(_08192_),
    .A1(_07184_),
    .A2(_08189_));
 sg13g2_nand2_1 _27487_ (.Y(_08193_),
    .A(_07105_),
    .B(_08192_));
 sg13g2_nand2_1 _27488_ (.Y(_08194_),
    .A(_09278_),
    .B(_08193_));
 sg13g2_a21oi_1 _27489_ (.A1(_08188_),
    .A2(_08194_),
    .Y(_02678_),
    .B1(net682));
 sg13g2_mux2_1 _27490_ (.A0(_10081_),
    .A1(\cpu.uart.r_x_invert ),
    .S(_08166_),
    .X(_08195_));
 sg13g2_and2_1 _27491_ (.A(net750),
    .B(_08195_),
    .X(_02679_));
 sg13g2_nand4_1 _27492_ (.B(net940),
    .C(_07179_),
    .A(_07098_),
    .Y(_08196_),
    .D(_07106_));
 sg13g2_o21ai_1 _27493_ (.B1(_08196_),
    .Y(_08197_),
    .A1(_07179_),
    .A2(_07182_));
 sg13g2_a221oi_1 _27494_ (.B2(_07118_),
    .C1(_07199_),
    .B1(_08197_),
    .A1(_07106_),
    .Y(_08198_),
    .A2(_07201_));
 sg13g2_buf_2 _27495_ (.A(_08198_),
    .X(_08199_));
 sg13g2_a21oi_1 _27496_ (.A1(_07117_),
    .A2(_07191_),
    .Y(_08200_),
    .B1(_07181_));
 sg13g2_nand3_1 _27497_ (.B(_08199_),
    .C(_08200_),
    .A(_07192_),
    .Y(_08201_));
 sg13g2_o21ai_1 _27498_ (.B1(_08201_),
    .Y(_08202_),
    .A1(net940),
    .A2(_08199_));
 sg13g2_nor2_1 _27499_ (.A(net692),
    .B(_08202_),
    .Y(_02682_));
 sg13g2_o21ai_1 _27500_ (.B1(_08199_),
    .Y(_08203_),
    .A1(net940),
    .A2(_07208_));
 sg13g2_nand2_1 _27501_ (.Y(_08204_),
    .A(net1104),
    .B(_08203_));
 sg13g2_nand4_1 _27502_ (.B(net940),
    .C(_07192_),
    .A(_07119_),
    .Y(_08205_),
    .D(_08199_));
 sg13g2_a21oi_1 _27503_ (.A1(_08204_),
    .A2(_08205_),
    .Y(_02683_),
    .B1(net682));
 sg13g2_nand2_1 _27504_ (.Y(_08206_),
    .A(net1104),
    .B(net940));
 sg13g2_nand2b_1 _27505_ (.Y(_08207_),
    .B(_07191_),
    .A_N(_07117_));
 sg13g2_o21ai_1 _27506_ (.B1(_08207_),
    .Y(_08208_),
    .A1(net939),
    .A2(_08206_));
 sg13g2_a21oi_1 _27507_ (.A1(_08199_),
    .A2(_08208_),
    .Y(_08209_),
    .B1(net938));
 sg13g2_nor2b_1 _27508_ (.A(_08206_),
    .B_N(_08207_),
    .Y(_08210_));
 sg13g2_or2_1 _27509_ (.X(_08211_),
    .B(_08210_),
    .A(net939));
 sg13g2_and3_1 _27510_ (.X(_08212_),
    .A(net938),
    .B(_08199_),
    .C(_08211_));
 sg13g2_nor3_1 _27511_ (.A(net691),
    .B(_08209_),
    .C(_08212_),
    .Y(_02684_));
 sg13g2_o21ai_1 _27512_ (.B1(_08199_),
    .Y(_08213_),
    .A1(net938),
    .A2(_08210_));
 sg13g2_nor4_1 _27513_ (.A(_07119_),
    .B(_07181_),
    .C(net939),
    .D(_07179_),
    .Y(_08214_));
 sg13g2_a22oi_1 _27514_ (.Y(_08215_),
    .B1(_08214_),
    .B2(_08199_),
    .A2(_08213_),
    .A1(net939));
 sg13g2_nor2_1 _27515_ (.A(net692),
    .B(_08215_),
    .Y(_02685_));
 sg13g2_nand2_1 _27516_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(net622),
    .B(_10715_));
 sg13g2_nand2b_1 _27517_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07382_),
    .A_N(_07378_));
 sg13g2_nor3_1 _27518_ (.A(_09933_),
    .B(_09840_),
    .C(_07802_),
    .Y(_08216_));
 sg13g2_nor2b_1 _27519_ (.A(_09886_),
    .B_N(_08216_),
    .Y(_08217_));
 sg13g2_a22oi_1 _27520_ (.Y(_08218_),
    .B1(_09855_),
    .B2(_08217_),
    .A2(net773),
    .A1(_09851_));
 sg13g2_inv_1 _27521_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08218_));
 sg13g2_nor2_1 _27522_ (.A(net1138),
    .B(net773),
    .Y(_08219_));
 sg13g2_a22oi_1 _27523_ (.Y(_08220_),
    .B1(_08216_),
    .B2(_08219_),
    .A2(_09853_),
    .A1(_09847_));
 sg13g2_nor2_1 _27524_ (.A(_06847_),
    .B(_08220_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27525_ (.A(_00189_),
    .B(_08220_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27526_ (.S0(_04867_),
    .A0(_09255_),
    .A1(_09264_),
    .A2(_09260_),
    .A3(_09245_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08221_));
 sg13g2_mux4_1 _27527_ (.S0(_04867_),
    .A0(_09262_),
    .A1(_09248_),
    .A2(_09246_),
    .A3(_09252_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08222_));
 sg13g2_mux2_1 _27528_ (.A0(_08221_),
    .A1(_08222_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27529_ (.S0(_04858_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_05333_),
    .X(_08223_));
 sg13g2_mux4_1 _27530_ (.S0(_04858_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_05333_),
    .X(_08224_));
 sg13g2_nor2b_1 _27531_ (.A(_05401_),
    .B_N(_08224_),
    .Y(_08225_));
 sg13g2_a21oi_1 _27532_ (.A1(_05401_),
    .A2(_08223_),
    .Y(_08226_),
    .B1(_08225_));
 sg13g2_nand2b_1 _27533_ (.Y(_08227_),
    .B(net1098),
    .A_N(_04858_));
 sg13g2_nand3_1 _27534_ (.B(_05333_),
    .C(net1101),
    .A(_04858_),
    .Y(_08228_));
 sg13g2_o21ai_1 _27535_ (.B1(_08228_),
    .Y(_08229_),
    .A1(_05333_),
    .A2(_08227_));
 sg13g2_nand3_1 _27536_ (.B(_00182_),
    .C(_08229_),
    .A(_05469_),
    .Y(_08230_));
 sg13g2_o21ai_1 _27537_ (.B1(_08230_),
    .Y(net15),
    .A1(_05469_),
    .A2(_08226_));
 sg13g2_mux4_1 _27538_ (.S0(_05540_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_05597_),
    .X(_08231_));
 sg13g2_mux4_1 _27539_ (.S0(_05540_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_05597_),
    .X(_08232_));
 sg13g2_nor2b_1 _27540_ (.A(_05687_),
    .B_N(_08232_),
    .Y(_08233_));
 sg13g2_a21oi_1 _27541_ (.A1(_05687_),
    .A2(_08231_),
    .Y(_08234_),
    .B1(_08233_));
 sg13g2_nand2b_1 _27542_ (.Y(_08235_),
    .B(net1098),
    .A_N(_05540_));
 sg13g2_nand3_1 _27543_ (.B(_05597_),
    .C(net1101),
    .A(_05540_),
    .Y(_08236_));
 sg13g2_o21ai_1 _27544_ (.B1(_08236_),
    .Y(_08237_),
    .A1(_05597_),
    .A2(_08235_));
 sg13g2_nand3_1 _27545_ (.B(_00181_),
    .C(_08237_),
    .A(_05101_),
    .Y(_08238_));
 sg13g2_o21ai_1 _27546_ (.B1(_08238_),
    .Y(net16),
    .A1(_05101_),
    .A2(_08234_));
 sg13g2_mux4_1 _27547_ (.S0(_04859_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_06384_),
    .X(_08239_));
 sg13g2_mux4_1 _27548_ (.S0(_04859_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_06384_),
    .X(_08240_));
 sg13g2_nor2b_1 _27549_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08240_),
    .Y(_08241_));
 sg13g2_a21oi_1 _27550_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08239_),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_nand2b_1 _27551_ (.Y(_08243_),
    .B(net1098),
    .A_N(_04859_));
 sg13g2_nand3_1 _27552_ (.B(net1101),
    .C(_06384_),
    .A(_04859_),
    .Y(_08244_));
 sg13g2_o21ai_1 _27553_ (.B1(_08244_),
    .Y(_08245_),
    .A1(_06384_),
    .A2(_08243_));
 sg13g2_nand3_1 _27554_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08245_),
    .A(_00106_),
    .Y(_08246_));
 sg13g2_o21ai_1 _27555_ (.B1(_08246_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08242_));
 sg13g2_mux4_1 _27556_ (.S0(_05541_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_06385_),
    .X(_08247_));
 sg13g2_mux4_1 _27557_ (.S0(_05541_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_06385_),
    .X(_08248_));
 sg13g2_nor2b_1 _27558_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08248_),
    .Y(_08249_));
 sg13g2_a21oi_1 _27559_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08247_),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_nand2b_1 _27560_ (.Y(_08251_),
    .B(net1098),
    .A_N(_05541_));
 sg13g2_nand3_1 _27561_ (.B(net1101),
    .C(_06385_),
    .A(_05541_),
    .Y(_08252_));
 sg13g2_o21ai_1 _27562_ (.B1(_08252_),
    .Y(_08253_),
    .A1(_06385_),
    .A2(_08251_));
 sg13g2_nand3_1 _27563_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08253_),
    .A(_00146_),
    .Y(_08254_));
 sg13g2_o21ai_1 _27564_ (.B1(_08254_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08250_));
 sg13g2_xor2_1 _27565_ (.B(clknet_leaf_83_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27566_ (.S0(_05549_),
    .A0(net1123),
    .A1(net1124),
    .A2(_08079_),
    .A3(_08095_),
    .S1(_06388_),
    .X(_08255_));
 sg13g2_mux4_1 _27567_ (.S0(_05549_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_06388_),
    .X(_08256_));
 sg13g2_nor2b_1 _27568_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08256_),
    .Y(_08257_));
 sg13g2_a21oi_1 _27569_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08255_),
    .Y(_08258_),
    .B1(_08257_));
 sg13g2_nand2b_1 _27570_ (.Y(_08259_),
    .B(_08097_),
    .A_N(_05549_));
 sg13g2_nand3_1 _27571_ (.B(net1101),
    .C(_06388_),
    .A(_05549_),
    .Y(_08260_));
 sg13g2_o21ai_1 _27572_ (.B1(_08260_),
    .Y(_08261_),
    .A1(_06388_),
    .A2(_08259_));
 sg13g2_nand3_1 _27573_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08261_),
    .A(_00149_),
    .Y(_08262_));
 sg13g2_o21ai_1 _27574_ (.B1(_08262_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08258_));
 sg13g2_mux4_1 _27575_ (.S0(_04848_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_06391_),
    .X(_08263_));
 sg13g2_mux4_1 _27576_ (.S0(_04848_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_06391_),
    .X(_08264_));
 sg13g2_nor2b_1 _27577_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08264_),
    .Y(_08265_));
 sg13g2_a21oi_1 _27578_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08263_),
    .Y(_08266_),
    .B1(_08265_));
 sg13g2_nand2b_1 _27579_ (.Y(_08267_),
    .B(net1098),
    .A_N(_04848_));
 sg13g2_nand3_1 _27580_ (.B(net1101),
    .C(_06391_),
    .A(_04848_),
    .Y(_08268_));
 sg13g2_o21ai_1 _27581_ (.B1(_08268_),
    .Y(_08269_),
    .A1(_06391_),
    .A2(_08267_));
 sg13g2_nand3_1 _27582_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08269_),
    .A(_00108_),
    .Y(_08270_));
 sg13g2_o21ai_1 _27583_ (.B1(_08270_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08266_));
 sg13g2_mux4_1 _27584_ (.S0(_05545_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_06392_),
    .X(_08271_));
 sg13g2_mux4_1 _27585_ (.S0(_05545_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(net1122),
    .S1(_06392_),
    .X(_08272_));
 sg13g2_nor2b_1 _27586_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08272_),
    .Y(_08273_));
 sg13g2_a21oi_1 _27587_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08271_),
    .Y(_08274_),
    .B1(_08273_));
 sg13g2_nand2b_1 _27588_ (.Y(_08275_),
    .B(net1098),
    .A_N(_05545_));
 sg13g2_nand3_1 _27589_ (.B(net1101),
    .C(_06392_),
    .A(_05545_),
    .Y(_08276_));
 sg13g2_o21ai_1 _27590_ (.B1(_08276_),
    .Y(_08277_),
    .A1(_06392_),
    .A2(_08275_));
 sg13g2_nand3_1 _27591_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08277_),
    .A(_00148_),
    .Y(_08278_));
 sg13g2_o21ai_1 _27592_ (.B1(_08278_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08274_));
 sg13g2_mux4_1 _27593_ (.S0(_04865_),
    .A0(net1123),
    .A1(net1124),
    .A2(net1100),
    .A3(net1099),
    .S1(_07709_),
    .X(_08279_));
 sg13g2_mux4_1 _27594_ (.S0(_04865_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(_07177_),
    .A2(_12048_),
    .A3(net1122),
    .S1(_07709_),
    .X(_08280_));
 sg13g2_nor2b_1 _27595_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08280_),
    .Y(_08281_));
 sg13g2_a21oi_1 _27596_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08279_),
    .Y(_08282_),
    .B1(_08281_));
 sg13g2_nand2b_1 _27597_ (.Y(_08283_),
    .B(net1098),
    .A_N(_04865_));
 sg13g2_nand3_1 _27598_ (.B(net1101),
    .C(_07709_),
    .A(_04865_),
    .Y(_08284_));
 sg13g2_o21ai_1 _27599_ (.B1(_08284_),
    .Y(_08285_),
    .A1(_07709_),
    .A2(_08283_));
 sg13g2_nand3_1 _27600_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08285_),
    .A(_00107_),
    .Y(_08286_));
 sg13g2_o21ai_1 _27601_ (.B1(_08286_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08282_));
 sg13g2_mux4_1 _27602_ (.S0(_05548_),
    .A0(_12027_),
    .A1(_12021_),
    .A2(net1100),
    .A3(net1099),
    .S1(_06394_),
    .X(_08287_));
 sg13g2_mux4_1 _27603_ (.S0(_05548_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1102),
    .A2(net1121),
    .A3(_12029_),
    .S1(_06394_),
    .X(_08288_));
 sg13g2_nor2b_1 _27604_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08288_),
    .Y(_08289_));
 sg13g2_a21oi_1 _27605_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08287_),
    .Y(_08290_),
    .B1(_08289_));
 sg13g2_nand2b_1 _27606_ (.Y(_08291_),
    .B(net1098),
    .A_N(_05548_));
 sg13g2_nand3_1 _27607_ (.B(_07799_),
    .C(_06394_),
    .A(_05548_),
    .Y(_08292_));
 sg13g2_o21ai_1 _27608_ (.B1(_08292_),
    .Y(_08293_),
    .A1(_06394_),
    .A2(_08291_));
 sg13g2_nand3_1 _27609_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08293_),
    .A(_00147_),
    .Y(_08294_));
 sg13g2_o21ai_1 _27610_ (.B1(_08294_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08290_));
 sg13g2_dfrbp_1 _27611_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1157),
    .D(_00319_),
    .Q_N(_14930_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27612_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1158),
    .D(_00320_),
    .Q_N(_14929_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27613_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1159),
    .D(_00321_),
    .Q_N(_14928_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27614_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1160),
    .D(_00322_),
    .Q_N(_14927_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27615_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1161),
    .D(_00323_),
    .Q_N(_14926_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27617_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27618_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1162),
    .D(_00324_),
    .Q_N(_14925_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1163),
    .D(_00325_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1164),
    .D(_00326_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1165),
    .D(_00327_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1166),
    .D(_00328_),
    .Q_N(_00131_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1167),
    .D(_00329_),
    .Q_N(_00143_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1168),
    .D(_00330_),
    .Q_N(_00155_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1169),
    .D(_00331_),
    .Q_N(_14924_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1170),
    .D(_00332_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1171),
    .D(_00333_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1172),
    .D(_00334_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1173),
    .D(_00335_),
    .Q_N(_14923_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1174),
    .D(_00336_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1175),
    .D(_00337_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1176),
    .D(_00338_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1177),
    .D(_00339_),
    .Q_N(_00153_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1178),
    .D(_00340_),
    .Q_N(_00313_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1179),
    .D(_00341_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1180),
    .D(_00342_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1181),
    .D(_00343_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1182),
    .D(_00344_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1183),
    .D(_00345_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1184),
    .D(_00346_),
    .Q_N(_14922_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1185),
    .D(_00347_),
    .Q_N(_00142_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1186),
    .D(_00348_),
    .Q_N(_00154_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1187),
    .D(_00349_),
    .Q_N(_14921_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1188),
    .D(_00350_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1189),
    .D(_00351_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1190),
    .D(_00352_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1191),
    .D(_00353_),
    .Q_N(_00152_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1192),
    .D(_00354_),
    .Q_N(_00314_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1193),
    .D(_00355_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1194),
    .D(_00356_),
    .Q_N(_14920_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1195),
    .D(_00357_),
    .Q_N(_14919_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1196),
    .D(_00358_),
    .Q_N(_14918_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1197),
    .D(_00359_),
    .Q_N(_14917_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1198),
    .D(_00360_),
    .Q_N(_14916_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1199),
    .D(_00361_),
    .Q_N(_14915_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1200),
    .D(_00362_),
    .Q_N(_14914_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1201),
    .D(_00363_),
    .Q_N(_14913_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1202),
    .D(_00364_),
    .Q_N(_14912_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1203),
    .D(_00365_),
    .Q_N(_14911_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1204),
    .D(_00366_),
    .Q_N(_14910_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1205),
    .D(_00367_),
    .Q_N(_14909_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1206),
    .D(_00368_),
    .Q_N(_14908_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1207),
    .D(_00369_),
    .Q_N(_14907_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1208),
    .D(_00370_),
    .Q_N(_14906_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1209),
    .D(_00371_),
    .Q_N(_14905_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1210),
    .D(_00372_),
    .Q_N(_14904_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1211),
    .D(_00373_),
    .Q_N(_14903_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1212),
    .D(_00374_),
    .Q_N(_14902_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1213),
    .D(_00375_),
    .Q_N(_14901_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1214),
    .D(_00376_),
    .Q_N(_14900_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1215),
    .D(_00377_),
    .Q_N(_14899_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1216),
    .D(_00378_),
    .Q_N(_14898_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1217),
    .D(_00379_),
    .Q_N(_14897_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1218),
    .D(_00380_),
    .Q_N(_14896_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1219),
    .D(_00381_),
    .Q_N(_14895_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1220),
    .D(_00382_),
    .Q_N(_14894_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1221),
    .D(_00383_),
    .Q_N(_14893_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1222),
    .D(_00384_),
    .Q_N(_14892_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1223),
    .D(_00385_),
    .Q_N(_14891_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1224),
    .D(_00386_),
    .Q_N(_14890_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1225),
    .D(_00387_),
    .Q_N(_14889_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1226),
    .D(_00388_),
    .Q_N(_14888_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1227),
    .D(_00389_),
    .Q_N(_14887_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1228),
    .D(_00390_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1229),
    .D(_00391_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1230),
    .D(_00392_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1231),
    .D(_00393_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_00394_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1233),
    .D(_00395_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1234),
    .D(_00396_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1235),
    .D(_00397_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1236),
    .D(_00398_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1237),
    .D(_00399_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1238),
    .D(_00400_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1239),
    .D(_00401_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1240),
    .D(_00402_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1241),
    .D(_00403_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1242),
    .D(_00404_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1243),
    .D(_00405_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1244),
    .D(_00406_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1245),
    .D(_00407_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1246),
    .D(_00408_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1247),
    .D(_00409_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1248),
    .D(_00410_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1249),
    .D(_00411_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1250),
    .D(_00412_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1251),
    .D(_00413_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1252),
    .D(_00414_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1253),
    .D(_00415_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1254),
    .D(_00416_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1255),
    .D(_00417_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1256),
    .D(_00418_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1257),
    .D(_00419_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1258),
    .D(_00420_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1259),
    .D(_00421_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1260),
    .D(_00422_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1261),
    .D(_00423_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1262),
    .D(_00424_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1263),
    .D(_00425_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1264),
    .D(_00426_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1265),
    .D(_00427_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1266),
    .D(_00428_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1267),
    .D(_00429_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1268),
    .D(_00430_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1269),
    .D(_00431_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1270),
    .D(_00432_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1271),
    .D(_00433_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1272),
    .D(_00434_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1273),
    .D(_00435_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1274),
    .D(_00436_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1275),
    .D(_00437_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1276),
    .D(_00438_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1277),
    .D(_00439_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1278),
    .D(_00440_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1279),
    .D(_00441_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1280),
    .D(_00442_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1281),
    .D(_00443_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1282),
    .D(_00444_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1283),
    .D(_00445_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1284),
    .D(_00446_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1285),
    .D(_00447_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1286),
    .D(_00448_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1287),
    .D(_00449_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1288),
    .D(_00450_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1289),
    .D(_00451_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1290),
    .D(_00452_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1291),
    .D(_00453_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1292),
    .D(_00454_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1293),
    .D(_00455_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1294),
    .D(_00456_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1295),
    .D(_00457_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1296),
    .D(_00458_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1297),
    .D(_00459_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1298),
    .D(_00460_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1299),
    .D(_00461_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1300),
    .D(_00462_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1301),
    .D(_00463_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1302),
    .D(_00464_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1303),
    .D(_00465_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1304),
    .D(_00466_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1305),
    .D(_00467_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1306),
    .D(_00468_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1307),
    .D(_00469_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1308),
    .D(_00470_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1309),
    .D(_00471_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1310),
    .D(_00472_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1311),
    .D(_00473_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1312),
    .D(_00474_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1313),
    .D(_00475_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1314),
    .D(_00476_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1315),
    .D(_00477_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1316),
    .D(_00478_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1317),
    .D(_00479_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1318),
    .D(_00480_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1319),
    .D(_00481_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1320),
    .D(_00482_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1321),
    .D(_00483_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1322),
    .D(_00484_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1323),
    .D(_00485_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1324),
    .D(_00486_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1325),
    .D(_00487_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1326),
    .D(_00488_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1327),
    .D(_00489_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1328),
    .D(_00490_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1329),
    .D(_00491_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1330),
    .D(_00492_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1331),
    .D(_00493_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1332),
    .D(_00494_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1333),
    .D(_00495_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1334),
    .D(_00496_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1335),
    .D(_00497_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1336),
    .D(_00498_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1337),
    .D(_00499_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1338),
    .D(_00500_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1339),
    .D(_00501_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1340),
    .D(_00502_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1341),
    .D(_00503_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1342),
    .D(_00504_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1343),
    .D(_00505_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1344),
    .D(_00506_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1345),
    .D(_00507_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1346),
    .D(_00508_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1347),
    .D(_00509_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1348),
    .D(_00510_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1349),
    .D(_00511_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1350),
    .D(_00512_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1351),
    .D(_00513_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1352),
    .D(_00514_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1353),
    .D(_00515_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1354),
    .D(_00516_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1355),
    .D(_00517_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1356),
    .D(_00518_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1357),
    .D(_00519_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1358),
    .D(_00520_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1359),
    .D(_00521_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1360),
    .D(_00522_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1361),
    .D(_00523_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1362),
    .D(_00524_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1363),
    .D(_00525_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1364),
    .D(_00526_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1365),
    .D(_00527_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1366),
    .D(_00528_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1367),
    .D(_00529_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1368),
    .D(_00530_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1369),
    .D(_00531_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1370),
    .D(_00532_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1371),
    .D(_00533_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1372),
    .D(_00534_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1373),
    .D(_00535_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1374),
    .D(_00536_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1375),
    .D(_00537_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1376),
    .D(_00538_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1377),
    .D(_00539_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1378),
    .D(_00540_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1379),
    .D(_00541_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1380),
    .D(_00542_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1381),
    .D(_00543_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1382),
    .D(_00544_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1383),
    .D(_00545_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1384),
    .D(_00546_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1385),
    .D(_00547_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1386),
    .D(_00548_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1387),
    .D(_00549_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1388),
    .D(_00550_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1389),
    .D(_00551_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1390),
    .D(_00552_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1391),
    .D(_00553_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1392),
    .D(_00554_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1393),
    .D(_00555_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1394),
    .D(_00556_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1395),
    .D(_00557_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1396),
    .D(_00558_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1397),
    .D(_00559_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1398),
    .D(_00560_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1399),
    .D(_00561_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1400),
    .D(_00562_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1401),
    .D(_00563_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1402),
    .D(_00564_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1403),
    .D(_00565_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1404),
    .D(_00566_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1405),
    .D(_00567_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1406),
    .D(_00568_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1407),
    .D(_00569_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1408),
    .D(_00570_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1409),
    .D(_00571_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1410),
    .D(_00572_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1411),
    .D(_00573_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1412),
    .D(_00574_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1413),
    .D(_00575_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1414),
    .D(_00576_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1415),
    .D(_00577_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1416),
    .D(_00578_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1417),
    .D(_00579_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1418),
    .D(_00580_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1419),
    .D(_00581_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1420),
    .D(_00582_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1421),
    .D(_00583_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1422),
    .D(_00584_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1423),
    .D(_00585_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1424),
    .D(_00586_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1425),
    .D(_00587_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1426),
    .D(_00588_),
    .Q_N(_00317_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1427),
    .D(_00589_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1428),
    .D(_00590_),
    .Q_N(_00278_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1429),
    .D(_00591_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1430),
    .D(_00592_),
    .Q_N(_00248_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1431),
    .D(_00593_),
    .Q_N(_00249_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1432),
    .D(_00594_),
    .Q_N(_00250_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1433),
    .D(_00595_),
    .Q_N(_00251_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1434),
    .D(_00596_),
    .Q_N(_00252_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1435),
    .D(_00597_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1436),
    .D(_00598_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1437),
    .D(_00599_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1438),
    .D(_00600_),
    .Q_N(_00253_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1439),
    .D(_00601_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1440),
    .D(_00602_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1441),
    .D(_00603_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1442),
    .D(_00604_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1443),
    .D(_00605_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1444),
    .D(_00606_),
    .Q_N(_00244_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1445),
    .D(_00607_),
    .Q_N(_00245_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1446),
    .D(_00608_),
    .Q_N(_00246_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1447),
    .D(_00609_),
    .Q_N(_00247_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1448),
    .D(_00610_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1449),
    .D(_00611_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1450),
    .D(_00612_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1451),
    .D(_00613_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1452),
    .D(_00614_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1453),
    .D(_00615_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1454),
    .D(_00616_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1455),
    .D(_00617_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1456),
    .D(_00618_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1457),
    .D(_00619_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1458),
    .D(_00620_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1459),
    .D(_00621_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1460),
    .D(_00622_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1461),
    .D(_00623_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1462),
    .D(_00624_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1463),
    .D(_00625_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1464),
    .D(_00626_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1465),
    .D(_00627_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1466),
    .D(_00628_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1467),
    .D(_00629_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1468),
    .D(_00630_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1469),
    .D(_00631_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1470),
    .D(_00632_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1471),
    .D(_00633_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1472),
    .D(_00634_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1473),
    .D(_00635_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1474),
    .D(_00636_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1475),
    .D(_00637_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1476),
    .D(_00638_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1477),
    .D(_00639_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1478),
    .D(_00640_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1479),
    .D(_00641_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1480),
    .D(_00642_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1481),
    .D(_00643_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1482),
    .D(_00644_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1483),
    .D(_00645_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1484),
    .D(_00646_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1485),
    .D(_00647_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1486),
    .D(_00648_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1487),
    .D(_00649_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1488),
    .D(_00650_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1489),
    .D(_00651_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1490),
    .D(_00652_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1491),
    .D(_00653_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1492),
    .D(_00654_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1493),
    .D(_00655_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1494),
    .D(_00656_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1495),
    .D(_00657_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1496),
    .D(_00658_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1497),
    .D(_00659_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1498),
    .D(_00660_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1499),
    .D(_00661_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1500),
    .D(_00662_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1501),
    .D(_00663_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1502),
    .D(_00664_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1503),
    .D(_00665_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1504),
    .D(_00666_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1505),
    .D(_00667_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1506),
    .D(_00668_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1507),
    .D(_00669_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1508),
    .D(_00670_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1509),
    .D(_00671_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1510),
    .D(_00672_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1511),
    .D(_00673_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1512),
    .D(_00674_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1513),
    .D(_00675_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1514),
    .D(_00676_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1515),
    .D(_00677_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1516),
    .D(_00678_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1517),
    .D(_00679_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1518),
    .D(_00680_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1519),
    .D(_00681_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1520),
    .D(_00682_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1521),
    .D(_00683_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1522),
    .D(_00684_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1523),
    .D(_00685_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1524),
    .D(_00686_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1525),
    .D(_00687_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1526),
    .D(_00688_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1527),
    .D(_00689_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1528),
    .D(_00690_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1529),
    .D(_00691_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1530),
    .D(_00692_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1531),
    .D(_00693_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1532),
    .D(_00694_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1533),
    .D(_00695_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1534),
    .D(_00696_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1535),
    .D(_00697_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1536),
    .D(_00698_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1537),
    .D(_00699_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1538),
    .D(_00700_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1539),
    .D(_00701_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1540),
    .D(_00702_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1541),
    .D(_00703_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1542),
    .D(_00704_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1543),
    .D(_00705_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1544),
    .D(_00706_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1545),
    .D(_00707_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1546),
    .D(_00708_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1547),
    .D(_00709_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1548),
    .D(_00710_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1549),
    .D(_00711_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1550),
    .D(_00712_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1551),
    .D(_00713_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1552),
    .D(_00714_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1553),
    .D(_00715_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1554),
    .D(_00716_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1555),
    .D(_00717_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1556),
    .D(_00718_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1557),
    .D(_00719_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1558),
    .D(_00720_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1559),
    .D(_00721_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1560),
    .D(_00722_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1561),
    .D(_00723_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1562),
    .D(_00724_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1563),
    .D(_00725_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1564),
    .D(_00726_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1565),
    .D(_00727_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1566),
    .D(_00728_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1567),
    .D(_00729_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1568),
    .D(_00730_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1569),
    .D(_00731_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1570),
    .D(_00732_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1571),
    .D(_00733_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1572),
    .D(_00734_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1573),
    .D(_00735_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1574),
    .D(_00736_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1575),
    .D(_00737_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1576),
    .D(_00738_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1577),
    .D(_00739_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1578),
    .D(_00740_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1579),
    .D(_00741_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1580),
    .D(_00742_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1581),
    .D(_00743_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1582),
    .D(_00744_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1583),
    .D(_00745_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1584),
    .D(_00746_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1585),
    .D(_00747_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1586),
    .D(_00748_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1587),
    .D(_00749_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1588),
    .D(_00750_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1589),
    .D(_00751_),
    .Q_N(_14543_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1590),
    .D(_00752_),
    .Q_N(_00300_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1591),
    .D(_00753_),
    .Q_N(_14542_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1592),
    .D(_00754_),
    .Q_N(_00275_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1593),
    .D(_00755_),
    .Q_N(_14541_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1594),
    .D(_00756_),
    .Q_N(_14540_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1595),
    .D(_00757_),
    .Q_N(_14539_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1596),
    .D(_00758_),
    .Q_N(_14538_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1597),
    .D(_00759_),
    .Q_N(_14537_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1598),
    .D(_00760_),
    .Q_N(_14536_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1599),
    .D(_00761_),
    .Q_N(_14535_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1600),
    .D(_00762_),
    .Q_N(_14534_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1601),
    .D(_00763_),
    .Q_N(_14533_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1602),
    .D(_00764_),
    .Q_N(_14532_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1603),
    .D(_00765_),
    .Q_N(_14531_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1604),
    .D(_00766_),
    .Q_N(_14530_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1605),
    .D(_00767_),
    .Q_N(_14529_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1606),
    .D(_00768_),
    .Q_N(_14528_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1607),
    .D(_00769_),
    .Q_N(_14527_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1608),
    .D(_00770_),
    .Q_N(_14526_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1609),
    .D(_00771_),
    .Q_N(_14525_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1610),
    .D(_00772_),
    .Q_N(_14524_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1611),
    .D(_00773_),
    .Q_N(_14523_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1612),
    .D(_00774_),
    .Q_N(_14522_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1613),
    .D(_00775_),
    .Q_N(_14521_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1614),
    .D(_00776_),
    .Q_N(_00260_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1615),
    .D(_00777_),
    .Q_N(_14520_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1616),
    .D(_00778_),
    .Q_N(_14519_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1617),
    .D(_00779_),
    .Q_N(_14931_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1618),
    .D(_00011_),
    .Q_N(_14932_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1619),
    .D(_00012_),
    .Q_N(_14933_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1620),
    .D(_00013_),
    .Q_N(_14934_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1621),
    .D(_00014_),
    .Q_N(_14935_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1622),
    .D(_00015_),
    .Q_N(_14936_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1623),
    .D(_00016_),
    .Q_N(_14937_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1624),
    .D(_00017_),
    .Q_N(_14938_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1625),
    .D(_00018_),
    .Q_N(_14939_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1626),
    .D(_00019_),
    .Q_N(_14940_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1627),
    .D(_00020_),
    .Q_N(_14518_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1628),
    .D(_00780_),
    .Q_N(_14517_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1629),
    .D(_00781_),
    .Q_N(_14516_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1630),
    .D(_00782_),
    .Q_N(_14515_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1631),
    .D(_00783_),
    .Q_N(_14941_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1632),
    .D(_00052_),
    .Q_N(_14514_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1633),
    .D(_00784_),
    .Q_N(_14513_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1634),
    .D(_00785_),
    .Q_N(_14512_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1635),
    .D(_00786_),
    .Q_N(_14511_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1636),
    .D(_00787_),
    .Q_N(_14510_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1637),
    .D(_00788_),
    .Q_N(_14509_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1638),
    .D(_00789_),
    .Q_N(_14508_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1639),
    .D(_00790_),
    .Q_N(_14507_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1640),
    .D(_00791_),
    .Q_N(_14506_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_inv$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1641),
    .D(_00792_),
    .Q_N(_14505_),
    .Q(\cpu.dec.r_rs2_inv ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1642),
    .D(_00793_),
    .Q_N(_14504_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1643),
    .D(_00794_),
    .Q_N(_14503_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1644),
    .D(_00795_),
    .Q_N(_00312_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1645),
    .D(_00796_),
    .Q_N(_14502_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1646),
    .D(_00797_),
    .Q_N(_00276_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1647),
    .D(_00798_),
    .Q_N(_14501_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1648),
    .D(_00799_),
    .Q_N(_14500_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1649),
    .D(_00800_),
    .Q_N(_00192_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1650),
    .D(_00801_),
    .Q_N(_14942_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1651),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00193_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1652),
    .D(_00802_),
    .Q_N(_14499_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1653),
    .D(_00803_),
    .Q_N(_14498_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1654),
    .D(_00804_),
    .Q_N(_14497_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1655),
    .D(_00805_),
    .Q_N(_14496_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1656),
    .D(_00806_),
    .Q_N(_14495_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1657),
    .D(_00807_),
    .Q_N(_14494_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1658),
    .D(_00808_),
    .Q_N(_14493_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1659),
    .D(_00809_),
    .Q_N(_14492_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1660),
    .D(_00810_),
    .Q_N(_14491_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1661),
    .D(_00811_),
    .Q_N(_14490_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1662),
    .D(_00812_),
    .Q_N(_14489_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1663),
    .D(_00813_),
    .Q_N(_14488_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1664),
    .D(_00814_),
    .Q_N(_14487_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1665),
    .D(_00815_),
    .Q_N(_14486_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1666),
    .D(_00816_),
    .Q_N(_14485_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1667),
    .D(_00817_),
    .Q_N(_14484_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1668),
    .D(_00818_),
    .Q_N(_14483_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1669),
    .D(_00819_),
    .Q_N(_14482_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1670),
    .D(_00820_),
    .Q_N(_14481_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1671),
    .D(_00821_),
    .Q_N(_14480_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1672),
    .D(_00822_),
    .Q_N(_14479_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1673),
    .D(_00823_),
    .Q_N(_14478_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1674),
    .D(_00824_),
    .Q_N(_14477_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1675),
    .D(_00825_),
    .Q_N(_14476_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1676),
    .D(_00826_),
    .Q_N(_14475_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1677),
    .D(_00827_),
    .Q_N(_14474_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1678),
    .D(_00828_),
    .Q_N(_14473_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1679),
    .D(_00829_),
    .Q_N(_14472_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1680),
    .D(_00830_),
    .Q_N(_14471_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1681),
    .D(_00831_),
    .Q_N(_14470_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1682),
    .D(_00832_),
    .Q_N(_14469_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1683),
    .D(_00833_),
    .Q_N(_14468_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1684),
    .D(_00834_),
    .Q_N(_14467_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1685),
    .D(_00835_),
    .Q_N(_14466_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1686),
    .D(_00836_),
    .Q_N(_14465_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1687),
    .D(_00837_),
    .Q_N(_14464_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1688),
    .D(_00838_),
    .Q_N(_14463_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1689),
    .D(_00839_),
    .Q_N(_14462_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1690),
    .D(_00840_),
    .Q_N(_14461_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1691),
    .D(_00841_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1692),
    .D(_00842_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1693),
    .D(_00843_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1694),
    .D(_00844_),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1695),
    .D(_00845_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1696),
    .D(_00846_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1697),
    .D(_00847_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1698),
    .D(_00848_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1699),
    .D(_00849_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1700),
    .D(_00850_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1701),
    .D(_00851_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1702),
    .D(_00852_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1703),
    .D(_00853_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1704),
    .D(_00854_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1705),
    .D(_00855_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1706),
    .D(_00856_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1707),
    .D(_00857_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1708),
    .D(_00858_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1709),
    .D(_00859_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1710),
    .D(_00860_),
    .Q_N(_14441_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1711),
    .D(_00861_),
    .Q_N(_14440_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1712),
    .D(_00862_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1713),
    .D(_00863_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1714),
    .D(_00864_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1715),
    .D(_00865_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1716),
    .D(_00866_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1717),
    .D(_00867_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1718),
    .D(_00868_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1719),
    .D(_00869_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1720),
    .D(_00870_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1721),
    .D(_00871_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1722),
    .D(_00872_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1723),
    .D(_00873_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1724),
    .D(_00874_),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1725),
    .D(_00875_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1726),
    .D(_00876_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1727),
    .D(_00877_),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1728),
    .D(_00878_),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1729),
    .D(_00879_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1730),
    .D(_00880_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1731),
    .D(_00881_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1732),
    .D(_00882_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1733),
    .D(_00883_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1734),
    .D(_00884_),
    .Q_N(_00270_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1735),
    .D(_00885_),
    .Q_N(_00271_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1736),
    .D(_00886_),
    .Q_N(_00272_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1737),
    .D(_00887_),
    .Q_N(_00273_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1738),
    .D(_00888_),
    .Q_N(_00274_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1739),
    .D(_00889_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1740),
    .D(_00890_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1741),
    .D(_00891_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1742),
    .D(_00892_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1743),
    .D(_00893_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1744),
    .D(_00894_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1745),
    .D(_00895_),
    .Q_N(_00266_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1746),
    .D(_00896_),
    .Q_N(_00267_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1747),
    .D(_00897_),
    .Q_N(_00268_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1748),
    .D(_00898_),
    .Q_N(_00269_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1749),
    .D(_00899_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1750),
    .D(_00900_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1751),
    .D(_00901_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1752),
    .D(_00902_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1753),
    .D(_00903_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1754),
    .D(_00904_),
    .Q_N(_14411_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1755),
    .D(_00905_),
    .Q_N(_14410_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1756),
    .D(_00906_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1757),
    .D(_00907_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1758),
    .D(_00908_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1759),
    .D(_00909_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1760),
    .D(_00910_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1761),
    .D(_00911_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1762),
    .D(_00912_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1763),
    .D(_00913_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1764),
    .D(_00914_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1765),
    .D(_00915_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1766),
    .D(_00916_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1767),
    .D(_00917_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1768),
    .D(_00918_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1769),
    .D(_00919_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1770),
    .D(_00920_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1771),
    .D(_00921_),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1772),
    .D(_00922_),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1773),
    .D(_00923_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1774),
    .D(_00924_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1775),
    .D(_00925_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1776),
    .D(_00926_),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1777),
    .D(_00927_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1778),
    .D(_00928_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1779),
    .D(_00929_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1780),
    .D(_00930_),
    .Q_N(_14943_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1781),
    .D(_00053_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1782),
    .D(_00931_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1783),
    .D(_00932_),
    .Q_N(_14944_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1784),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1785),
    .D(_00933_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1786),
    .D(_00934_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1787),
    .D(_00935_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1788),
    .D(_00936_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1789),
    .D(_00937_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1790),
    .D(_00938_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1791),
    .D(_00939_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1792),
    .D(_00940_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1793),
    .D(_00941_),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1794),
    .D(_00942_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1795),
    .D(_00943_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1796),
    .D(_00944_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1797),
    .D(_00945_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1798),
    .D(_00946_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1799),
    .D(_00947_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1800),
    .D(_00948_),
    .Q_N(_00189_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1801),
    .D(_00949_),
    .Q_N(_14367_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1802),
    .D(_00950_),
    .Q_N(_14366_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1803),
    .D(_00951_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1804),
    .D(_00952_),
    .Q_N(_00197_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1805),
    .D(_00953_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1806),
    .D(_00954_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1807),
    .D(_00955_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1808),
    .D(_00956_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1809),
    .D(_00957_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1810),
    .D(_00958_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1811),
    .D(_00959_),
    .Q_N(_14358_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1812),
    .D(_00960_),
    .Q_N(_14357_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1813),
    .D(_00961_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1814),
    .D(_00962_),
    .Q_N(_14355_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1815),
    .D(_00963_),
    .Q_N(_14354_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1816),
    .D(_00964_),
    .Q_N(_14353_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1817),
    .D(_00965_),
    .Q_N(_14352_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1818),
    .D(_00966_),
    .Q_N(_14351_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1819),
    .D(_00967_),
    .Q_N(_14945_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1820),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14946_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1821),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00167_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1822),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00168_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1823),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00169_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1824),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00170_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1825),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00171_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1826),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1827),
    .D(_00968_),
    .Q_N(_00311_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1828),
    .D(_00969_),
    .Q_N(_00310_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1829),
    .D(_00970_),
    .Q_N(_00309_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1830),
    .D(_00971_),
    .Q_N(_00308_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1831),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1832),
    .D(_00972_),
    .Q_N(_00307_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1833),
    .D(_00973_),
    .Q_N(_00306_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1834),
    .D(_00974_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1835),
    .D(_00975_),
    .Q_N(_00305_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1836),
    .D(_00976_),
    .Q_N(_00304_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1837),
    .D(_00977_),
    .Q_N(_00303_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1838),
    .D(_00978_),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1839),
    .D(_00979_),
    .Q_N(_00302_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1840),
    .D(_00980_),
    .Q_N(_14346_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1841),
    .D(_00981_),
    .Q_N(_14947_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1842),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1843),
    .D(_00982_),
    .Q_N(_00301_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1844),
    .D(_00983_),
    .Q_N(_14948_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1845),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00127_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1846),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00139_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1847),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00151_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1848),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1849),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00164_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1850),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00165_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1851),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00166_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1852),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14949_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1853),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14950_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1854),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14951_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1855),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14952_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1856),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00199_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1857),
    .D(_00984_),
    .Q_N(_00200_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1858),
    .D(_00985_),
    .Q_N(_00292_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1859),
    .D(_00986_),
    .Q_N(_00291_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1860),
    .D(_00987_),
    .Q_N(_00196_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1861),
    .D(_00988_),
    .Q_N(_00195_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1862),
    .D(_00989_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1863),
    .D(_00990_),
    .Q_N(_00299_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1864),
    .D(_00991_),
    .Q_N(_00191_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1865),
    .D(_00992_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1866),
    .D(_00993_),
    .Q_N(_00298_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1867),
    .D(_00994_),
    .Q_N(_00297_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1868),
    .D(_00995_),
    .Q_N(_00296_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1869),
    .D(_00996_),
    .Q_N(_00295_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1870),
    .D(_00997_),
    .Q_N(_00294_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1871),
    .D(_00998_),
    .Q_N(_00293_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1872),
    .D(_00999_),
    .Q_N(_14345_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1873),
    .D(_01000_),
    .Q_N(_00198_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1874),
    .D(_01001_),
    .Q_N(_14344_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1875),
    .D(_01002_),
    .Q_N(_14343_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1876),
    .D(_01003_),
    .Q_N(_14342_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1877),
    .D(_01004_),
    .Q_N(_14341_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1878),
    .D(_01005_),
    .Q_N(_14340_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1879),
    .D(_01006_),
    .Q_N(_14339_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1880),
    .D(_01007_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1881),
    .D(_01008_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1882),
    .D(_01009_),
    .Q_N(_14336_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1883),
    .D(_01010_),
    .Q_N(_14335_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1884),
    .D(_01011_),
    .Q_N(_14334_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1885),
    .D(_01012_),
    .Q_N(_14333_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1886),
    .D(_01013_),
    .Q_N(_14332_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1887),
    .D(_01014_),
    .Q_N(_14331_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1888),
    .D(_01015_),
    .Q_N(_14330_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1889),
    .D(_01016_),
    .Q_N(_14329_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1890),
    .D(_01017_),
    .Q_N(_14328_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1891),
    .D(_01018_),
    .Q_N(_14327_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1892),
    .D(_01019_),
    .Q_N(_14326_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1893),
    .D(_01020_),
    .Q_N(_14325_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1894),
    .D(_01021_),
    .Q_N(_14324_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1895),
    .D(_01022_),
    .Q_N(_14323_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1896),
    .D(_01023_),
    .Q_N(_14322_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1897),
    .D(_01024_),
    .Q_N(_14321_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1898),
    .D(_01025_),
    .Q_N(_14320_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1899),
    .D(_01026_),
    .Q_N(_14319_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1900),
    .D(_01027_),
    .Q_N(_14318_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1901),
    .D(_01028_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1902),
    .D(_01029_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1903),
    .D(_01030_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1904),
    .D(_01031_),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1905),
    .D(_01032_),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1906),
    .D(_01033_),
    .Q_N(_00259_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1907),
    .D(_01034_),
    .Q_N(_00241_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1908),
    .D(_01035_),
    .Q_N(_00243_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1909),
    .D(_01036_),
    .Q_N(_14312_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1910),
    .D(_01037_),
    .Q_N(_14311_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1911),
    .D(_01038_),
    .Q_N(_14310_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1912),
    .D(_01039_),
    .Q_N(_14309_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1913),
    .D(_01040_),
    .Q_N(_00277_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1914),
    .D(_01041_),
    .Q_N(_14308_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1915),
    .D(_01042_),
    .Q_N(_00230_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1916),
    .D(_01043_),
    .Q_N(_00229_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1917),
    .D(_01044_),
    .Q_N(_00231_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1918),
    .D(_01045_),
    .Q_N(_00233_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1919),
    .D(_01046_),
    .Q_N(_00235_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1920),
    .D(_01047_),
    .Q_N(_00237_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1921),
    .D(_01048_),
    .Q_N(_00239_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1922),
    .D(_01049_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1923),
    .D(_01050_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1924),
    .D(_01051_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1925),
    .D(_01052_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1926),
    .D(_01053_),
    .Q_N(_14953_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1927),
    .D(_00054_),
    .Q_N(_00258_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1928),
    .D(_01054_),
    .Q_N(_00225_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1929),
    .D(_01055_),
    .Q_N(_14303_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1930),
    .D(_01056_),
    .Q_N(_14302_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1931),
    .D(_01057_),
    .Q_N(_14301_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1932),
    .D(_01058_),
    .Q_N(_14300_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1933),
    .D(_01059_),
    .Q_N(_14299_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1934),
    .D(_01060_),
    .Q_N(_14298_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1935),
    .D(_01061_),
    .Q_N(_00183_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1936),
    .D(_01062_),
    .Q_N(_00184_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1937),
    .D(_01063_),
    .Q_N(_00289_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1938),
    .D(_01064_),
    .Q_N(_00185_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1939),
    .D(_01065_),
    .Q_N(_00186_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1940),
    .D(_01066_),
    .Q_N(_00187_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1941),
    .D(_01067_),
    .Q_N(_00283_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1942),
    .D(_01068_),
    .Q_N(_14297_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1943),
    .D(_01069_),
    .Q_N(_14296_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1944),
    .D(_01070_),
    .Q_N(_14295_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1945),
    .D(_01071_),
    .Q_N(_14294_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1946),
    .D(_01072_),
    .Q_N(_00290_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1947),
    .D(_01073_),
    .Q_N(_14293_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1948),
    .D(_01074_),
    .Q_N(_00188_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1949),
    .D(_01075_),
    .Q_N(_14292_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1950),
    .D(_01076_),
    .Q_N(_00257_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1951),
    .D(_01077_),
    .Q_N(_14291_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1952),
    .D(_01078_),
    .Q_N(_14290_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1953),
    .D(_01079_),
    .Q_N(_14289_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1954),
    .D(_01080_),
    .Q_N(_14288_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1955),
    .D(_01081_),
    .Q_N(_14287_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1956),
    .D(_01082_),
    .Q_N(_14286_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1957),
    .D(_01083_),
    .Q_N(_14285_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1958),
    .D(_01084_),
    .Q_N(_14284_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1959),
    .D(_01085_),
    .Q_N(_14283_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1960),
    .D(_01086_),
    .Q_N(_14282_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1961),
    .D(_01087_),
    .Q_N(_14281_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1962),
    .D(_01088_),
    .Q_N(_14280_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1963),
    .D(_01089_),
    .Q_N(_14279_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1964),
    .D(_01090_),
    .Q_N(_14278_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1965),
    .D(_01091_),
    .Q_N(_14277_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1966),
    .D(_01092_),
    .Q_N(_14276_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1967),
    .D(_01093_),
    .Q_N(_14275_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1968),
    .D(_01094_),
    .Q_N(_14274_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1969),
    .D(_01095_),
    .Q_N(_14273_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1970),
    .D(_01096_),
    .Q_N(_14272_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1971),
    .D(_01097_),
    .Q_N(_14271_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1972),
    .D(_01098_),
    .Q_N(_14270_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1973),
    .D(_01099_),
    .Q_N(_14269_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1974),
    .D(_01100_),
    .Q_N(_14268_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1975),
    .D(_01101_),
    .Q_N(_14267_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1976),
    .D(_01102_),
    .Q_N(_14266_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1977),
    .D(_01103_),
    .Q_N(_14265_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1978),
    .D(_01104_),
    .Q_N(_14264_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1979),
    .D(_01105_),
    .Q_N(_14263_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1980),
    .D(_01106_),
    .Q_N(_14262_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1981),
    .D(_01107_),
    .Q_N(_14261_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1982),
    .D(_01108_),
    .Q_N(_14260_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1983),
    .D(_01109_),
    .Q_N(_14259_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1984),
    .D(_01110_),
    .Q_N(_14258_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1985),
    .D(_01111_),
    .Q_N(_14257_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1986),
    .D(_01112_),
    .Q_N(_14256_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1987),
    .D(_01113_),
    .Q_N(_14255_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1988),
    .D(_01114_),
    .Q_N(_14254_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1989),
    .D(_01115_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1990),
    .D(_01116_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1991),
    .D(_01117_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1992),
    .D(_01118_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1993),
    .D(_01119_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1994),
    .D(_01120_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1995),
    .D(_01121_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1996),
    .D(_01122_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1997),
    .D(_01123_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1998),
    .D(_01124_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1999),
    .D(_01125_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2000),
    .D(_01126_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2001),
    .D(_01127_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2002),
    .D(_01128_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2003),
    .D(_01129_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2004),
    .D(_01130_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2005),
    .D(_01131_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2006),
    .D(_01132_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2007),
    .D(_01133_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2008),
    .D(_01134_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2009),
    .D(_01135_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2010),
    .D(_01136_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2011),
    .D(_01137_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2012),
    .D(_01138_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2013),
    .D(_01139_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2014),
    .D(_01140_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2015),
    .D(_01141_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2016),
    .D(_01142_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2017),
    .D(_01143_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2018),
    .D(_01144_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2019),
    .D(_01145_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2020),
    .D(_01146_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2021),
    .D(_01147_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2022),
    .D(_01148_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2023),
    .D(_01149_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2024),
    .D(_01150_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2025),
    .D(_01151_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2026),
    .D(_01152_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2027),
    .D(_01153_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2028),
    .D(_01154_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2029),
    .D(_01155_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2030),
    .D(_01156_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2031),
    .D(_01157_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2032),
    .D(_01158_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2033),
    .D(_01159_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2034),
    .D(_01160_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2035),
    .D(_01161_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2036),
    .D(_01162_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2037),
    .D(_01163_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2038),
    .D(_01164_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2039),
    .D(_01165_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2040),
    .D(_01166_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2041),
    .D(_01167_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2042),
    .D(_01168_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2043),
    .D(_01169_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2044),
    .D(_01170_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2045),
    .D(_01171_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2046),
    .D(_01172_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2047),
    .D(_01173_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2048),
    .D(_01174_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2049),
    .D(_01175_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2050),
    .D(_01176_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2051),
    .D(_01177_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2052),
    .D(_01178_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2053),
    .D(_01179_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2054),
    .D(_01180_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2055),
    .D(_01181_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2056),
    .D(_01182_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2057),
    .D(_01183_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2058),
    .D(_01184_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2059),
    .D(_01185_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2060),
    .D(_01186_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2061),
    .D(_01187_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2062),
    .D(_01188_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2063),
    .D(_01189_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2064),
    .D(_01190_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2065),
    .D(_01191_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2066),
    .D(_01192_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2067),
    .D(_01193_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2068),
    .D(_01194_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2069),
    .D(_01195_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2070),
    .D(_01196_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2071),
    .D(_01197_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2072),
    .D(_01198_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2073),
    .D(_01199_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2074),
    .D(_01200_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2075),
    .D(_01201_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2076),
    .D(_01202_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2077),
    .D(_01203_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2078),
    .D(_01204_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2079),
    .D(_01205_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2080),
    .D(_01206_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2081),
    .D(_01207_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2082),
    .D(_01208_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2083),
    .D(_01209_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2084),
    .D(_01210_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2085),
    .D(_01211_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2086),
    .D(_01212_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2087),
    .D(_01213_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2088),
    .D(_01214_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2089),
    .D(_01215_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2090),
    .D(_01216_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2091),
    .D(_01217_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2092),
    .D(_01218_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2093),
    .D(_01219_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2094),
    .D(_01220_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2095),
    .D(_01221_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2096),
    .D(_01222_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2097),
    .D(_01223_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2098),
    .D(_01224_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2099),
    .D(_01225_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2100),
    .D(_01226_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2101),
    .D(_01227_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2102),
    .D(_01228_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2103),
    .D(_01229_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2104),
    .D(_01230_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2105),
    .D(_01231_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2106),
    .D(_01232_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2107),
    .D(_01233_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2108),
    .D(_01234_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2109),
    .D(_01235_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2110),
    .D(_01236_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2111),
    .D(_01237_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2112),
    .D(_01238_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2113),
    .D(_01239_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2114),
    .D(_01240_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2115),
    .D(_01241_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2116),
    .D(_01242_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2117),
    .D(_01243_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2118),
    .D(_01244_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2119),
    .D(_01245_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2120),
    .D(_01246_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2121),
    .D(_01247_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2122),
    .D(_01248_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2123),
    .D(_01249_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2124),
    .D(_01250_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2125),
    .D(_01251_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2126),
    .D(_01252_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2127),
    .D(_01253_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2128),
    .D(_01254_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2129),
    .D(_01255_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2130),
    .D(_01256_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2131),
    .D(_01257_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2132),
    .D(_01258_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2133),
    .D(_01259_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2134),
    .D(_01260_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2135),
    .D(_01261_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2136),
    .D(_01262_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2137),
    .D(_01263_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2138),
    .D(_01264_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2139),
    .D(_01265_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2140),
    .D(_01266_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2141),
    .D(_01267_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2142),
    .D(_01268_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2143),
    .D(_01269_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2144),
    .D(_01270_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2145),
    .D(_01271_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2146),
    .D(_01272_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2147),
    .D(_01273_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2148),
    .D(_01274_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2149),
    .D(_01275_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2150),
    .D(_01276_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2151),
    .D(_01277_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2152),
    .D(_01278_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2153),
    .D(_01279_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2154),
    .D(_01280_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2155),
    .D(_01281_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2156),
    .D(_01282_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2157),
    .D(_01283_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2158),
    .D(_01284_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2159),
    .D(_01285_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2160),
    .D(_01286_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2161),
    .D(_01287_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2162),
    .D(_01288_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2163),
    .D(_01289_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2164),
    .D(_01290_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2165),
    .D(_01291_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2166),
    .D(_01292_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2167),
    .D(_01293_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2168),
    .D(_01294_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2169),
    .D(_01295_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2170),
    .D(_01296_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2171),
    .D(_01297_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2172),
    .D(_01298_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2173),
    .D(_01299_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2174),
    .D(_01300_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2175),
    .D(_01301_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2176),
    .D(_01302_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2177),
    .D(_01303_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2178),
    .D(_01304_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2179),
    .D(_01305_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2180),
    .D(_01306_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2181),
    .D(_01307_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2182),
    .D(_01308_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2183),
    .D(_01309_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2184),
    .D(_01310_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2185),
    .D(_01311_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2186),
    .D(_01312_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2187),
    .D(_01313_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2188),
    .D(_01314_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2189),
    .D(_01315_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2190),
    .D(_01316_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2191),
    .D(_01317_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2192),
    .D(_01318_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2193),
    .D(_01319_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2194),
    .D(_01320_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2195),
    .D(_01321_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2196),
    .D(_01322_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2197),
    .D(_01323_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2198),
    .D(_01324_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2199),
    .D(_01325_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2200),
    .D(_01326_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2201),
    .D(_01327_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2202),
    .D(_01328_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2203),
    .D(_01329_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2204),
    .D(_01330_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2205),
    .D(_01331_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2206),
    .D(_01332_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2207),
    .D(_01333_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2208),
    .D(_01334_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2209),
    .D(_01335_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2210),
    .D(_01336_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2211),
    .D(_01337_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2212),
    .D(_01338_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2213),
    .D(_01339_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2214),
    .D(_01340_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2215),
    .D(_01341_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2216),
    .D(_01342_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2217),
    .D(_01343_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2218),
    .D(_01344_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2219),
    .D(_01345_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2220),
    .D(_01346_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2221),
    .D(_01347_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2222),
    .D(_01348_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2223),
    .D(_01349_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2224),
    .D(_01350_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2225),
    .D(_01351_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2226),
    .D(_01352_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2227),
    .D(_01353_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2228),
    .D(_01354_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2229),
    .D(_01355_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2230),
    .D(_01356_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2231),
    .D(_01357_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2232),
    .D(_01358_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2233),
    .D(_01359_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2234),
    .D(_01360_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2235),
    .D(_01361_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2236),
    .D(_01362_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2237),
    .D(_01363_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2238),
    .D(_01364_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2239),
    .D(_01365_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2240),
    .D(_01366_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2241),
    .D(_01367_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2242),
    .D(_01368_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2243),
    .D(_01369_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2244),
    .D(_01370_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2245),
    .D(_01371_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2246),
    .D(_01372_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2247),
    .D(_01373_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2248),
    .D(_01374_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2249),
    .D(_01375_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2250),
    .D(_01376_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2251),
    .D(_01377_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2252),
    .D(_01378_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2253),
    .D(_01379_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2254),
    .D(_01380_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2255),
    .D(_01381_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2256),
    .D(_01382_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2257),
    .D(_01383_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2258),
    .D(_01384_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2259),
    .D(_01385_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2260),
    .D(_01386_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2261),
    .D(_01387_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2262),
    .D(_01388_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2263),
    .D(_01389_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2264),
    .D(_01390_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2265),
    .D(_01391_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2266),
    .D(_01392_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2267),
    .D(_01393_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2268),
    .D(_01394_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2269),
    .D(_01395_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2270),
    .D(_01396_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2271),
    .D(_01397_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2272),
    .D(_01398_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2273),
    .D(_01399_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2274),
    .D(_01400_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2275),
    .D(_01401_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2276),
    .D(_01402_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2277),
    .D(_01403_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2278),
    .D(_01404_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2279),
    .D(_01405_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2280),
    .D(_01406_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2281),
    .D(_01407_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2282),
    .D(_01408_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2283),
    .D(_01409_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2284),
    .D(_01410_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2285),
    .D(_01411_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2286),
    .D(_01412_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2287),
    .D(_01413_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2288),
    .D(_01414_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2289),
    .D(_01415_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2290),
    .D(_01416_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2291),
    .D(_01417_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2292),
    .D(_01418_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2293),
    .D(_01419_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2294),
    .D(_01420_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2295),
    .D(_01421_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2296),
    .D(_01422_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2297),
    .D(_01423_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2298),
    .D(_01424_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2299),
    .D(_01425_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2300),
    .D(_01426_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2301),
    .D(_01427_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2302),
    .D(_01428_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2303),
    .D(_01429_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2304),
    .D(_01430_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2305),
    .D(_01431_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2306),
    .D(_01432_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2307),
    .D(_01433_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2308),
    .D(_01434_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2309),
    .D(_01435_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2310),
    .D(_01436_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2311),
    .D(_01437_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2312),
    .D(_01438_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2313),
    .D(_01439_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2314),
    .D(_01440_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2315),
    .D(_01441_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2316),
    .D(_01442_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2317),
    .D(_01443_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2318),
    .D(_01444_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2319),
    .D(_01445_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2320),
    .D(_01446_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2321),
    .D(_01447_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2322),
    .D(_01448_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2323),
    .D(_01449_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2324),
    .D(_01450_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2325),
    .D(_01451_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2326),
    .D(_01452_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2327),
    .D(_01453_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2328),
    .D(_01454_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2329),
    .D(_01455_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2330),
    .D(_01456_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2331),
    .D(_01457_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2332),
    .D(_01458_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2333),
    .D(_01459_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2334),
    .D(_01460_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2335),
    .D(_01461_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2336),
    .D(_01462_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2337),
    .D(_01463_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2338),
    .D(_01464_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2339),
    .D(_01465_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2340),
    .D(_01466_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2341),
    .D(_01467_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2342),
    .D(_01468_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2343),
    .D(_01469_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2344),
    .D(_01470_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2345),
    .D(_01471_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2346),
    .D(_01472_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2347),
    .D(_01473_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2348),
    .D(_01474_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2349),
    .D(_01475_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2350),
    .D(_01476_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2351),
    .D(_01477_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2352),
    .D(_01478_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2353),
    .D(_01479_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2354),
    .D(_01480_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2355),
    .D(_01481_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2356),
    .D(_01482_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2357),
    .D(_01483_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2358),
    .D(_01484_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2359),
    .D(_01485_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2360),
    .D(_01486_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2361),
    .D(_01487_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2362),
    .D(_01488_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2363),
    .D(_01489_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2364),
    .D(_01490_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2365),
    .D(_01491_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2366),
    .D(_01492_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2367),
    .D(_01493_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2368),
    .D(_01494_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2369),
    .D(_01495_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2370),
    .D(_01496_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2371),
    .D(_01497_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2372),
    .D(_01498_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2373),
    .D(_01499_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2374),
    .D(_01500_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2375),
    .D(_01501_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2376),
    .D(_01502_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2377),
    .D(_01503_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2378),
    .D(_01504_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2379),
    .D(_01505_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2380),
    .D(_01506_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2381),
    .D(_01507_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2382),
    .D(_01508_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2383),
    .D(_01509_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2384),
    .D(_01510_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2385),
    .D(_01511_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2386),
    .D(_01512_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2387),
    .D(_01513_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2388),
    .D(_01514_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2389),
    .D(_01515_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2390),
    .D(_01516_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2391),
    .D(_01517_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2392),
    .D(_01518_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2393),
    .D(_01519_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2394),
    .D(_01520_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2395),
    .D(_01521_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2396),
    .D(_01522_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2397),
    .D(_01523_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2398),
    .D(_01524_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2399),
    .D(_01525_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2400),
    .D(_01526_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2401),
    .D(_01527_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2402),
    .D(_01528_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2403),
    .D(_01529_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2404),
    .D(_01530_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2405),
    .D(_01531_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2406),
    .D(_01532_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2407),
    .D(_01533_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2408),
    .D(_01534_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2409),
    .D(_01535_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2410),
    .D(_01536_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2411),
    .D(_01537_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2412),
    .D(_01538_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2413),
    .D(_01539_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2414),
    .D(_01540_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2415),
    .D(_01541_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2416),
    .D(_01542_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2417),
    .D(_01543_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2418),
    .D(_01544_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2419),
    .D(_01545_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2420),
    .D(_01546_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2421),
    .D(_01547_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2422),
    .D(_01548_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2423),
    .D(_01549_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2424),
    .D(_01550_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2425),
    .D(_01551_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2426),
    .D(_01552_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2427),
    .D(_01553_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2428),
    .D(_01554_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2429),
    .D(_01555_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2430),
    .D(_01556_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2431),
    .D(_01557_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2432),
    .D(_01558_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2433),
    .D(_01559_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2434),
    .D(_01560_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2435),
    .D(_01561_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2436),
    .D(_01562_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2437),
    .D(_01563_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2438),
    .D(_01564_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2439),
    .D(_01565_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2440),
    .D(_01566_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2441),
    .D(_01567_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2442),
    .D(_01568_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2443),
    .D(_01569_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2444),
    .D(_01570_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2445),
    .D(_01571_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2446),
    .D(_01572_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2447),
    .D(_01573_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2448),
    .D(_01574_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2449),
    .D(_01575_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2450),
    .D(_01576_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2451),
    .D(_01577_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2452),
    .D(_01578_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2453),
    .D(_01579_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2454),
    .D(_01580_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2455),
    .D(_01581_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2456),
    .D(_01582_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2457),
    .D(_01583_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2458),
    .D(_01584_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2459),
    .D(_01585_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2460),
    .D(_01586_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2461),
    .D(_01587_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2462),
    .D(_01588_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2463),
    .D(_01589_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2464),
    .D(_01590_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2465),
    .D(_01591_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2466),
    .D(_01592_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2467),
    .D(_01593_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2468),
    .D(_01594_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2469),
    .D(_01595_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2470),
    .D(_01596_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2471),
    .D(_01597_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2472),
    .D(_01598_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2473),
    .D(_01599_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2474),
    .D(_01600_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2475),
    .D(_01601_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2476),
    .D(_01602_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2477),
    .D(_01603_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2478),
    .D(_01604_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2479),
    .D(_01605_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2480),
    .D(_01606_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2481),
    .D(_01607_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2482),
    .D(_01608_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2483),
    .D(_01609_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2484),
    .D(_01610_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2485),
    .D(_01611_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2486),
    .D(_01612_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2487),
    .D(_01613_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2488),
    .D(_01614_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2489),
    .D(_01615_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2490),
    .D(_01616_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2491),
    .D(_01617_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2492),
    .D(_01618_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2493),
    .D(_01619_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2494),
    .D(_01620_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2495),
    .D(_01621_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2496),
    .D(_01622_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2497),
    .D(_01623_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2498),
    .D(_01624_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2499),
    .D(_01625_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2500),
    .D(_01626_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2501),
    .D(_01627_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2502),
    .D(_01628_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2503),
    .D(_01629_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2504),
    .D(_01630_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2505),
    .D(_01631_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2506),
    .D(_01632_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2507),
    .D(_01633_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2508),
    .D(_01634_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2509),
    .D(_01635_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2510),
    .D(_01636_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2511),
    .D(_01637_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2512),
    .D(_01638_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2513),
    .D(_01639_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2514),
    .D(_01640_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2515),
    .D(_01641_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2516),
    .D(_01642_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2517),
    .D(_01643_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2518),
    .D(_01644_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2519),
    .D(_01645_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2520),
    .D(_01646_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2521),
    .D(_01647_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2522),
    .D(_01648_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2523),
    .D(_01649_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2524),
    .D(_01650_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2525),
    .D(_01651_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2526),
    .D(_01652_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2527),
    .D(_01653_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2528),
    .D(_01654_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2529),
    .D(_01655_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2530),
    .D(_01656_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2531),
    .D(_01657_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2532),
    .D(_01658_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2533),
    .D(_01659_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2534),
    .D(_01660_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2535),
    .D(_01661_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2536),
    .D(_01662_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2537),
    .D(_01663_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2538),
    .D(_01664_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2539),
    .D(_01665_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2540),
    .D(_01666_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2541),
    .D(_01667_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2542),
    .D(_01668_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2543),
    .D(_01669_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2544),
    .D(_01670_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2545),
    .D(_01671_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2546),
    .D(_01672_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2547),
    .D(_01673_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2548),
    .D(_01674_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2549),
    .D(_01675_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2550),
    .D(_01676_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net2551),
    .D(_01677_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2552),
    .D(_01678_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2553),
    .D(_01679_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2554),
    .D(_01680_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2555),
    .D(_01681_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2556),
    .D(_01682_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2557),
    .D(_01683_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2558),
    .D(_01684_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2559),
    .D(_01685_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2560),
    .D(_01686_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2561),
    .D(_01687_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2562),
    .D(_01688_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2563),
    .D(_01689_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2564),
    .D(_01690_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2565),
    .D(_01691_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2566),
    .D(_01692_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2567),
    .D(_01693_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2568),
    .D(_01694_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2569),
    .D(_01695_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2570),
    .D(_01696_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2571),
    .D(_01697_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2572),
    .D(_01698_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2573),
    .D(_01699_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2574),
    .D(_01700_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2575),
    .D(_01701_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2576),
    .D(_01702_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2577),
    .D(_01703_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2578),
    .D(_01704_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2579),
    .D(_01705_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2580),
    .D(_01706_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2581),
    .D(_01707_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2582),
    .D(_01708_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2583),
    .D(_01709_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2584),
    .D(_01710_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2585),
    .D(_01711_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2586),
    .D(_01712_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2587),
    .D(_01713_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2588),
    .D(_01714_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2589),
    .D(_01715_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2590),
    .D(_01716_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2591),
    .D(_01717_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2592),
    .D(_01718_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2593),
    .D(_01719_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2594),
    .D(_01720_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2595),
    .D(_01721_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2596),
    .D(_01722_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2597),
    .D(_01723_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2598),
    .D(_01724_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2599),
    .D(_01725_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2600),
    .D(_01726_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2601),
    .D(_01727_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2602),
    .D(_01728_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2603),
    .D(_01729_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2604),
    .D(_01730_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2605),
    .D(_01731_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2606),
    .D(_01732_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2607),
    .D(_01733_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2608),
    .D(_01734_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2609),
    .D(_01735_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2610),
    .D(_01736_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2611),
    .D(_01737_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2612),
    .D(_01738_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2613),
    .D(_01739_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2614),
    .D(_01740_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2615),
    .D(_01741_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2616),
    .D(_01742_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2617),
    .D(_01743_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2618),
    .D(_01744_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2619),
    .D(_01745_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2620),
    .D(_01746_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2621),
    .D(_01747_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2622),
    .D(_01748_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2623),
    .D(_01749_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2624),
    .D(_01750_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2625),
    .D(_01751_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2626),
    .D(_01752_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2627),
    .D(_01753_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2628),
    .D(_01754_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2629),
    .D(_01755_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2630),
    .D(_01756_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2631),
    .D(_01757_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2632),
    .D(_01758_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2633),
    .D(_01759_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2634),
    .D(_01760_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2635),
    .D(_01761_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2636),
    .D(_01762_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2637),
    .D(_01763_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2638),
    .D(_01764_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2639),
    .D(_01765_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2640),
    .D(_01766_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2641),
    .D(_01767_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2642),
    .D(_01768_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2643),
    .D(_01769_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2644),
    .D(_01770_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2645),
    .D(_01771_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2646),
    .D(_01772_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2647),
    .D(_01773_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2648),
    .D(_01774_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2649),
    .D(_01775_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2650),
    .D(_01776_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2651),
    .D(_01777_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2652),
    .D(_01778_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2653),
    .D(_01779_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2654),
    .D(_01780_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2655),
    .D(_01781_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2656),
    .D(_01782_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2657),
    .D(_01783_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2658),
    .D(_01784_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2659),
    .D(_01785_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2660),
    .D(_01786_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2661),
    .D(_01787_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2662),
    .D(_01788_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2663),
    .D(_01789_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2664),
    .D(_01790_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2665),
    .D(_01791_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2666),
    .D(_01792_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2667),
    .D(_01793_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2668),
    .D(_01794_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2669),
    .D(_01795_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2670),
    .D(_01796_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2671),
    .D(_01797_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2672),
    .D(_01798_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2673),
    .D(_01799_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2674),
    .D(_01800_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2675),
    .D(_01801_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2676),
    .D(_01802_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2677),
    .D(_01803_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2678),
    .D(_01804_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2679),
    .D(_01805_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2680),
    .D(_01806_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2681),
    .D(_01807_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2682),
    .D(_01808_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2683),
    .D(_01809_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2684),
    .D(_01810_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2685),
    .D(_01811_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2686),
    .D(_01812_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2687),
    .D(_01813_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2688),
    .D(_01814_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2689),
    .D(_01815_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2690),
    .D(_01816_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2691),
    .D(_01817_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2692),
    .D(_01818_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2693),
    .D(_01819_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2694),
    .D(_01820_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2695),
    .D(_01821_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2696),
    .D(_01822_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2697),
    .D(_01823_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2698),
    .D(_01824_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2699),
    .D(_01825_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2700),
    .D(_01826_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2701),
    .D(_01827_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2702),
    .D(_01828_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2703),
    .D(_01829_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2704),
    .D(_01830_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2705),
    .D(_01831_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2706),
    .D(_01832_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2707),
    .D(_01833_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2708),
    .D(_01834_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2709),
    .D(_01835_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2710),
    .D(_01836_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2711),
    .D(_01837_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2712),
    .D(_01838_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2713),
    .D(_01839_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2714),
    .D(_01840_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2715),
    .D(_01841_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2716),
    .D(_01842_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2717),
    .D(_01843_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2718),
    .D(_01844_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2719),
    .D(_01845_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2720),
    .D(_01846_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2721),
    .D(_01847_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2722),
    .D(_01848_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2723),
    .D(_01849_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2724),
    .D(_01850_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2725),
    .D(_01851_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2726),
    .D(_01852_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2727),
    .D(_01853_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2728),
    .D(_01854_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2729),
    .D(_01855_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2730),
    .D(_01856_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2731),
    .D(_01857_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2732),
    .D(_01858_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2733),
    .D(_01859_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2734),
    .D(_01860_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2735),
    .D(_01861_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2736),
    .D(_01862_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2737),
    .D(_01863_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2738),
    .D(_01864_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2739),
    .D(_01865_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2740),
    .D(_01866_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2741),
    .D(_01867_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2742),
    .D(_01868_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2743),
    .D(_01869_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2744),
    .D(_01870_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2745),
    .D(_01871_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2746),
    .D(_01872_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2747),
    .D(_01873_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2748),
    .D(_01874_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2749),
    .D(_01875_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2750),
    .D(_01876_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2751),
    .D(_01877_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2752),
    .D(_01878_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2753),
    .D(_01879_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2754),
    .D(_01880_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2755),
    .D(_01881_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2756),
    .D(_01882_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2757),
    .D(_01883_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2758),
    .D(_01884_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2759),
    .D(_01885_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2760),
    .D(_01886_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2761),
    .D(_01887_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2762),
    .D(_01888_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2763),
    .D(_01889_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2764),
    .D(_01890_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2765),
    .D(_01891_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2766),
    .D(_01892_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2767),
    .D(_01893_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2768),
    .D(_01894_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2769),
    .D(_01895_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2770),
    .D(_01896_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2771),
    .D(_01897_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2772),
    .D(_01898_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2773),
    .D(_01899_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2774),
    .D(_01900_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2775),
    .D(_01901_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2776),
    .D(_01902_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2777),
    .D(_01903_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2778),
    .D(_01904_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2779),
    .D(_01905_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2780),
    .D(_01906_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2781),
    .D(_01907_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2782),
    .D(_01908_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2783),
    .D(_01909_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2784),
    .D(_01910_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2785),
    .D(_01911_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2786),
    .D(_01912_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2787),
    .D(_01913_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2788),
    .D(_01914_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2789),
    .D(_01915_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2790),
    .D(_01916_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2791),
    .D(_01917_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2792),
    .D(_01918_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2793),
    .D(_01919_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2794),
    .D(_01920_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2795),
    .D(_01921_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2796),
    .D(_01922_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2797),
    .D(_01923_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2798),
    .D(_01924_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2799),
    .D(_01925_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2800),
    .D(_01926_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2801),
    .D(_01927_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2802),
    .D(_01928_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2803),
    .D(_01929_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2804),
    .D(_01930_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2805),
    .D(_01931_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2806),
    .D(_01932_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2807),
    .D(_01933_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2808),
    .D(_01934_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2809),
    .D(_01935_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2810),
    .D(_01936_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2811),
    .D(_01937_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2812),
    .D(_01938_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2813),
    .D(_01939_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2814),
    .D(_01940_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2815),
    .D(_01941_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2816),
    .D(_01942_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2817),
    .D(_01943_),
    .Q_N(_13425_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2818),
    .D(_01944_),
    .Q_N(_13424_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2819),
    .D(_01945_),
    .Q_N(_13423_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2820),
    .D(_01946_),
    .Q_N(_13422_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2821),
    .D(_01947_),
    .Q_N(_13421_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2822),
    .D(_01948_),
    .Q_N(_13420_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net2823),
    .D(_01949_),
    .Q_N(_13419_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2824),
    .D(_01950_),
    .Q_N(_13418_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2825),
    .D(_01951_),
    .Q_N(_13417_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2826),
    .D(_01952_),
    .Q_N(_13416_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2827),
    .D(_01953_),
    .Q_N(_13415_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2828),
    .D(_01954_),
    .Q_N(_13414_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2829),
    .D(_01955_),
    .Q_N(_13413_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2830),
    .D(_01956_),
    .Q_N(_13412_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2831),
    .D(_01957_),
    .Q_N(_13411_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2832),
    .D(_01958_),
    .Q_N(_13410_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2833),
    .D(_01959_),
    .Q_N(_13409_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2834),
    .D(_01960_),
    .Q_N(_13408_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2835),
    .D(_01961_),
    .Q_N(_13407_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2836),
    .D(_01962_),
    .Q_N(_13406_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2837),
    .D(_01963_),
    .Q_N(_13405_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2838),
    .D(_01964_),
    .Q_N(_13404_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2839),
    .D(_01965_),
    .Q_N(_13403_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2840),
    .D(_01966_),
    .Q_N(_13402_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2841),
    .D(_01967_),
    .Q_N(_13401_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2842),
    .D(_01968_),
    .Q_N(_13400_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2843),
    .D(_01969_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net2844),
    .D(_01970_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2845),
    .D(_01971_),
    .Q_N(_00119_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2846),
    .D(_01972_),
    .Q_N(_13399_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2847),
    .D(_01973_),
    .Q_N(_00138_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2848),
    .D(_01974_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2849),
    .D(_01975_),
    .Q_N(_00162_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2850),
    .D(_01976_),
    .Q_N(_13398_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2851),
    .D(_01977_),
    .Q_N(_13397_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2852),
    .D(_01978_),
    .Q_N(_00182_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2853),
    .D(_01979_),
    .Q_N(_13396_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2854),
    .D(_01980_),
    .Q_N(_13395_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2855),
    .D(_01981_),
    .Q_N(_13394_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2856),
    .D(_01982_),
    .Q_N(_00181_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2857),
    .D(_01983_),
    .Q_N(_13393_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2858),
    .D(_01984_),
    .Q_N(_13392_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2859),
    .D(_01985_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2860),
    .D(_01986_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2861),
    .D(_01987_),
    .Q_N(_00116_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2862),
    .D(_01988_),
    .Q_N(_13391_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2863),
    .D(_01989_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2864),
    .D(_01990_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2865),
    .D(_01991_),
    .Q_N(_00158_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2866),
    .D(_01992_),
    .Q_N(_13390_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2867),
    .D(_01993_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2868),
    .D(_01994_),
    .Q_N(_00149_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2869),
    .D(_01995_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2870),
    .D(_01996_),
    .Q_N(_13389_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2871),
    .D(_01997_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2872),
    .D(_01998_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2873),
    .D(_01999_),
    .Q_N(_00118_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2874),
    .D(_02000_),
    .Q_N(_13388_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2875),
    .D(_02001_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2876),
    .D(_02002_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2877),
    .D(_02003_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2878),
    .D(_02004_),
    .Q_N(_13387_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2879),
    .D(_02005_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2880),
    .D(_02006_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2881),
    .D(_02007_),
    .Q_N(_00117_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2882),
    .D(_02008_),
    .Q_N(_13386_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2883),
    .D(_02009_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2884),
    .D(_02010_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2885),
    .D(_02011_),
    .Q_N(_00159_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2886),
    .D(_02012_),
    .Q_N(_13385_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2887),
    .D(_02013_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2888),
    .D(_02014_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2889),
    .D(_02015_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2890),
    .D(_02016_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2891),
    .D(_02017_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2892),
    .D(_02018_),
    .Q_N(_00215_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2893),
    .D(_02019_),
    .Q_N(_13384_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2894),
    .D(_02020_),
    .Q_N(_13383_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2895),
    .D(_02021_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2896),
    .D(_02022_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2897),
    .D(_02023_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2898),
    .D(_02024_),
    .Q_N(_00218_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2899),
    .D(_02025_),
    .Q_N(_00220_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2900),
    .D(_02026_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2901),
    .D(_02027_),
    .Q_N(_00222_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2902),
    .D(_02028_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2903),
    .D(_02029_),
    .Q_N(_00214_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2904),
    .D(_02030_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2905),
    .D(_02031_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2906),
    .D(_02032_),
    .Q_N(_00177_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2907),
    .D(_02033_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2908),
    .D(_02034_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2909),
    .D(_02035_),
    .Q_N(_00216_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2910),
    .D(_02036_),
    .Q_N(_13382_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2911),
    .D(_02037_),
    .Q_N(_00217_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2912),
    .D(_02038_),
    .Q_N(_13381_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2913),
    .D(_02039_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2914),
    .D(_02040_),
    .Q_N(_00219_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2915),
    .D(_02041_),
    .Q_N(_00221_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2916),
    .D(_02042_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2917),
    .D(_02043_),
    .Q_N(_00213_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2918),
    .D(_02044_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2919),
    .D(_02045_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2920),
    .D(_02046_),
    .Q_N(_00176_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2921),
    .D(_02047_),
    .Q_N(_13380_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2922),
    .D(_02048_),
    .Q_N(_13379_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2923),
    .D(_02049_),
    .Q_N(_13378_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2924),
    .D(_02050_),
    .Q_N(_13377_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2925),
    .D(_02051_),
    .Q_N(_13376_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2926),
    .D(_02052_),
    .Q_N(_13375_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2927),
    .D(_02053_),
    .Q_N(_13374_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2928),
    .D(_02054_),
    .Q_N(_13373_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2929),
    .D(_02055_),
    .Q_N(_13372_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2930),
    .D(_02056_),
    .Q_N(_13371_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2931),
    .D(_02057_),
    .Q_N(_13370_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2932),
    .D(_02058_),
    .Q_N(_13369_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2933),
    .D(_02059_),
    .Q_N(_13368_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2934),
    .D(_02060_),
    .Q_N(_13367_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2935),
    .D(_02061_),
    .Q_N(_13366_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2936),
    .D(_02062_),
    .Q_N(_13365_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2937),
    .D(_02063_),
    .Q_N(_13364_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2938),
    .D(_02064_),
    .Q_N(_13363_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2939),
    .D(_02065_),
    .Q_N(_13362_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2940),
    .D(_02066_),
    .Q_N(_13361_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2941),
    .D(_02067_),
    .Q_N(_13360_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2942),
    .D(_02068_),
    .Q_N(_13359_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2943),
    .D(_02069_),
    .Q_N(_13358_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2944),
    .D(_02070_),
    .Q_N(_13357_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2945),
    .D(_02071_),
    .Q_N(_13356_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2946),
    .D(_02072_),
    .Q_N(_13355_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2947),
    .D(_02073_),
    .Q_N(_13354_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2948),
    .D(_02074_),
    .Q_N(_13353_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2949),
    .D(_02075_),
    .Q_N(_13352_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2950),
    .D(_02076_),
    .Q_N(_13351_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2951),
    .D(_02077_),
    .Q_N(_13350_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2952),
    .D(_02078_),
    .Q_N(_13349_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2953),
    .D(_02079_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2954),
    .D(_02080_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2955),
    .D(_02081_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2956),
    .D(_02082_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2957),
    .D(_02083_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2958),
    .D(_02084_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2959),
    .D(_02085_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2960),
    .D(_02086_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2961),
    .D(_02087_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2962),
    .D(_02088_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2963),
    .D(_02089_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2964),
    .D(_02090_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2965),
    .D(_02091_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2966),
    .D(_02092_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2967),
    .D(_02093_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2968),
    .D(_02094_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2969),
    .D(_02095_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2970),
    .D(_02096_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2971),
    .D(_02097_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2972),
    .D(_02098_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2973),
    .D(_02099_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2974),
    .D(_02100_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2975),
    .D(_02101_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2976),
    .D(_02102_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2977),
    .D(_02103_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2978),
    .D(_02104_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2979),
    .D(_02105_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2980),
    .D(_02106_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2981),
    .D(_02107_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2982),
    .D(_02108_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2983),
    .D(_02109_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2984),
    .D(_02110_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2985),
    .D(_02111_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2986),
    .D(_02112_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2987),
    .D(_02113_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2988),
    .D(_02114_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2989),
    .D(_02115_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2990),
    .D(_02116_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2991),
    .D(_02117_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2992),
    .D(_02118_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2993),
    .D(_02119_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2994),
    .D(_02120_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2995),
    .D(_02121_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2996),
    .D(_02122_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2997),
    .D(_02123_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2998),
    .D(_02124_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2999),
    .D(_02125_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3000),
    .D(_02126_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3001),
    .D(_02127_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3002),
    .D(_02128_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3003),
    .D(_02129_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3004),
    .D(_02130_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3005),
    .D(_02131_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3006),
    .D(_02132_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3007),
    .D(_02133_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3008),
    .D(_02134_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3009),
    .D(_02135_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3010),
    .D(_02136_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3011),
    .D(_02137_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3012),
    .D(_02138_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3013),
    .D(_02139_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3014),
    .D(_02140_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3015),
    .D(_02141_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3016),
    .D(_02142_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3017),
    .D(_02143_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3018),
    .D(_02144_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3019),
    .D(_02145_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3020),
    .D(_02146_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3021),
    .D(_02147_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3022),
    .D(_02148_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3023),
    .D(_02149_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3024),
    .D(_02150_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3025),
    .D(_02151_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3026),
    .D(_02152_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3027),
    .D(_02153_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3028),
    .D(_02154_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3029),
    .D(_02155_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3030),
    .D(_02156_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3031),
    .D(_02157_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3032),
    .D(_02158_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3033),
    .D(_02159_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3034),
    .D(_02160_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3035),
    .D(_02161_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3036),
    .D(_02162_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3037),
    .D(_02163_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3038),
    .D(_02164_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3039),
    .D(_02165_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3040),
    .D(_02166_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3041),
    .D(_02167_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3042),
    .D(_02168_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3043),
    .D(_02169_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3044),
    .D(_02170_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3045),
    .D(_02171_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3046),
    .D(_02172_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3047),
    .D(_02173_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3048),
    .D(_02174_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3049),
    .D(_02175_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3050),
    .D(_02176_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3051),
    .D(_02177_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3052),
    .D(_02178_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3053),
    .D(_02179_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3054),
    .D(_02180_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3055),
    .D(_02181_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3056),
    .D(_02182_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3057),
    .D(_02183_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3058),
    .D(_02184_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3059),
    .D(_02185_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3060),
    .D(_02186_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3061),
    .D(_02187_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3062),
    .D(_02188_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3063),
    .D(_02189_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3064),
    .D(_02190_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3065),
    .D(_02191_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3066),
    .D(_02192_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3067),
    .D(_02193_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3068),
    .D(_02194_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3069),
    .D(_02195_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3070),
    .D(_02196_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3071),
    .D(_02197_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3072),
    .D(_02198_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3073),
    .D(_02199_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3074),
    .D(_02200_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3075),
    .D(_02201_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3076),
    .D(_02202_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3077),
    .D(_02203_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3078),
    .D(_02204_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3079),
    .D(_02205_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3080),
    .D(_02206_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3081),
    .D(_02207_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3082),
    .D(_02208_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3083),
    .D(_02209_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3084),
    .D(_02210_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3085),
    .D(_02211_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3086),
    .D(_02212_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3087),
    .D(_02213_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3088),
    .D(_02214_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3089),
    .D(_02215_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3090),
    .D(_02216_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3091),
    .D(_02217_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3092),
    .D(_02218_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3093),
    .D(_02219_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3094),
    .D(_02220_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3095),
    .D(_02221_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3096),
    .D(_02222_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3097),
    .D(_02223_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3098),
    .D(_02224_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3099),
    .D(_02225_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3100),
    .D(_02226_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3101),
    .D(_02227_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3102),
    .D(_02228_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3103),
    .D(_02229_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3104),
    .D(_02230_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3105),
    .D(_02231_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3106),
    .D(_02232_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3107),
    .D(_02233_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3108),
    .D(_02234_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3109),
    .D(_02235_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3110),
    .D(_02236_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3111),
    .D(_02237_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3112),
    .D(_02238_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3113),
    .D(_02239_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3114),
    .D(_02240_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3115),
    .D(_02241_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3116),
    .D(_02242_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3117),
    .D(_02243_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3118),
    .D(_02244_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3119),
    .D(_02245_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3120),
    .D(_02246_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3121),
    .D(_02247_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3122),
    .D(_02248_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3123),
    .D(_02249_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3124),
    .D(_02250_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3125),
    .D(_02251_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3126),
    .D(_02252_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3127),
    .D(_02253_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3128),
    .D(_02254_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3129),
    .D(_02255_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3130),
    .D(_02256_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3131),
    .D(_02257_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3132),
    .D(_02258_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3133),
    .D(_02259_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3134),
    .D(_02260_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3135),
    .D(_02261_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3136),
    .D(_02262_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3137),
    .D(_02263_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3138),
    .D(_02264_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3139),
    .D(_02265_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3140),
    .D(_02266_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3141),
    .D(_02267_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3142),
    .D(_02268_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3143),
    .D(_02269_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3144),
    .D(_02270_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3145),
    .D(_02271_),
    .Q_N(_00318_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3146),
    .D(_02272_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3147),
    .D(_02273_),
    .Q_N(_00256_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3148),
    .D(_02274_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3149),
    .D(_02275_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3150),
    .D(_02276_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3151),
    .D(_02277_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3152),
    .D(_02278_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3153),
    .D(_02279_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3154),
    .D(_02280_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3155),
    .D(_02281_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3156),
    .D(_02282_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3157),
    .D(_02283_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3158),
    .D(_02284_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3159),
    .D(_02285_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3160),
    .D(_02286_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3161),
    .D(_02287_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3162),
    .D(_02288_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3163),
    .D(_02289_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3164),
    .D(_02290_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3165),
    .D(_02291_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3166),
    .D(_02292_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3167),
    .D(_02293_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3168),
    .D(_02294_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3169),
    .D(_02295_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3170),
    .D(_02296_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3171),
    .D(_02297_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3172),
    .D(_02298_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3173),
    .D(_02299_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3174),
    .D(_02300_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3175),
    .D(_02301_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3176),
    .D(_02302_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3177),
    .D(_02303_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3178),
    .D(_02304_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3179),
    .D(_02305_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3180),
    .D(_02306_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3181),
    .D(_02307_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3182),
    .D(_02308_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3183),
    .D(_02309_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3184),
    .D(_02310_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3185),
    .D(_02311_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3186),
    .D(_02312_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3187),
    .D(_02313_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3188),
    .D(_02314_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3189),
    .D(_02315_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3190),
    .D(_02316_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3191),
    .D(_02317_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3192),
    .D(_02318_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3193),
    .D(_02319_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3194),
    .D(_02320_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3195),
    .D(_02321_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3196),
    .D(_02322_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3197),
    .D(_02323_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3198),
    .D(_02324_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3199),
    .D(_02325_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3200),
    .D(_02326_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3201),
    .D(_02327_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3202),
    .D(_02328_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3203),
    .D(_02329_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3204),
    .D(_02330_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3205),
    .D(_02331_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3206),
    .D(_02332_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3207),
    .D(_02333_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3208),
    .D(_02334_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3209),
    .D(_02335_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3210),
    .D(_02336_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3211),
    .D(_02337_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3212),
    .D(_02338_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3213),
    .D(_02339_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3214),
    .D(_02340_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3215),
    .D(_02341_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3216),
    .D(_02342_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3217),
    .D(_02343_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3218),
    .D(_02344_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3219),
    .D(_02345_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3220),
    .D(_02346_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3221),
    .D(_02347_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3222),
    .D(_02348_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3223),
    .D(_02349_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3224),
    .D(_02350_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3225),
    .D(_02351_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3226),
    .D(_02352_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3227),
    .D(_02353_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3228),
    .D(_02354_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3229),
    .D(_02355_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net3230),
    .D(_02356_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3231),
    .D(_02357_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3232),
    .D(_02358_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3233),
    .D(_02359_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3234),
    .D(_02360_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3235),
    .D(_02361_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3236),
    .D(_02362_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3237),
    .D(_02363_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3238),
    .D(_02364_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3239),
    .D(_02365_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3240),
    .D(_02366_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3241),
    .D(_02367_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3242),
    .D(_02368_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3243),
    .D(_02369_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3244),
    .D(_02370_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3245),
    .D(_02371_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3246),
    .D(_02372_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3247),
    .D(_02373_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3248),
    .D(_02374_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3249),
    .D(_02375_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3250),
    .D(_02376_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3251),
    .D(_02377_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3252),
    .D(_02378_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3253),
    .D(_02379_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3254),
    .D(_02380_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3255),
    .D(_02381_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3256),
    .D(_02382_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3257),
    .D(_02383_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3258),
    .D(_02384_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3259),
    .D(_02385_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3260),
    .D(_02386_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3261),
    .D(_02387_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3262),
    .D(_02388_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3263),
    .D(_02389_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3264),
    .D(_02390_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3265),
    .D(_02391_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3266),
    .D(_02392_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3267),
    .D(_02393_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3268),
    .D(_02394_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3269),
    .D(_02395_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3270),
    .D(_02396_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3271),
    .D(_02397_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3272),
    .D(_02398_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3273),
    .D(_02399_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3274),
    .D(_02400_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3275),
    .D(_02401_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3276),
    .D(_02402_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3277),
    .D(_02403_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3278),
    .D(_02404_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3279),
    .D(_02405_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3280),
    .D(_02406_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3281),
    .D(_02407_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3282),
    .D(_02408_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3283),
    .D(_02409_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3284),
    .D(_02410_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3285),
    .D(_02411_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3286),
    .D(_02412_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3287),
    .D(_02413_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3288),
    .D(_02414_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3289),
    .D(_02415_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3290),
    .D(_02416_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3291),
    .D(_02417_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3292),
    .D(_02418_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3293),
    .D(_02419_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3294),
    .D(_02420_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3295),
    .D(_02421_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3296),
    .D(_02422_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3297),
    .D(_02423_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3298),
    .D(_02424_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3299),
    .D(_02425_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3300),
    .D(_02426_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3301),
    .D(_02427_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3302),
    .D(_02428_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3303),
    .D(_02429_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3304),
    .D(_02430_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3305),
    .D(_02431_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3306),
    .D(_02432_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3307),
    .D(_02433_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3308),
    .D(_02434_),
    .Q_N(_12995_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3309),
    .D(_02435_),
    .Q_N(_12994_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3310),
    .D(_02436_),
    .Q_N(_12993_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3311),
    .D(_02437_),
    .Q_N(_12992_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3312),
    .D(_02438_),
    .Q_N(_12991_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3313),
    .D(_02439_),
    .Q_N(_12990_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3314),
    .D(_02440_),
    .Q_N(_12989_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3315),
    .D(_02441_),
    .Q_N(_12988_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3316),
    .D(_02442_),
    .Q_N(_12987_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3317),
    .D(_02443_),
    .Q_N(_12986_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3318),
    .D(_02444_),
    .Q_N(_12985_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3319),
    .D(_02445_),
    .Q_N(_12984_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3320),
    .D(_02446_),
    .Q_N(_12983_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3321),
    .D(_02447_),
    .Q_N(_12982_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3322),
    .D(_02448_),
    .Q_N(_12981_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3323),
    .D(_02449_),
    .Q_N(_12980_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3324),
    .D(_02450_),
    .Q_N(_12979_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3325),
    .D(_02451_),
    .Q_N(_12978_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3326),
    .D(_02452_),
    .Q_N(_12977_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3327),
    .D(_02453_),
    .Q_N(_12976_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3328),
    .D(_02454_),
    .Q_N(_12975_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3329),
    .D(_02455_),
    .Q_N(_12974_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3330),
    .D(_02456_),
    .Q_N(_12973_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3331),
    .D(_02457_),
    .Q_N(_12972_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3332),
    .D(_02458_),
    .Q_N(_12971_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3333),
    .D(_02459_),
    .Q_N(_12970_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3334),
    .D(_02460_),
    .Q_N(_12969_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3335),
    .D(_02461_),
    .Q_N(_12968_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3336),
    .D(_02462_),
    .Q_N(_12967_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3337),
    .D(_02463_),
    .Q_N(_12966_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3338),
    .D(_02464_),
    .Q_N(_12965_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3339),
    .D(_02465_),
    .Q_N(_12964_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3340),
    .D(_02466_),
    .Q_N(_14954_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3341),
    .D(_00036_),
    .Q_N(_00288_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3342),
    .D(_00037_),
    .Q_N(_14955_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3343),
    .D(_00038_),
    .Q_N(_14956_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3344),
    .D(_00039_),
    .Q_N(_14957_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3345),
    .D(_00040_),
    .Q_N(_14958_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3346),
    .D(_00041_),
    .Q_N(_14959_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3347),
    .D(_00042_),
    .Q_N(_12963_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3348),
    .D(_02467_),
    .Q_N(_12962_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3349),
    .D(_02468_),
    .Q_N(_12961_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3350),
    .D(_02469_),
    .Q_N(_12960_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3351),
    .D(_02470_),
    .Q_N(_14960_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3352),
    .D(_00043_),
    .Q_N(_12959_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3353),
    .D(_02471_),
    .Q_N(_12958_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3354),
    .D(_02472_),
    .Q_N(_12957_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3355),
    .D(_02473_),
    .Q_N(_12956_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3356),
    .D(_02474_),
    .Q_N(_12955_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3357),
    .D(_02475_),
    .Q_N(_12954_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3358),
    .D(_02476_),
    .Q_N(_12953_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3359),
    .D(_02477_),
    .Q_N(_12952_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3360),
    .D(_02478_),
    .Q_N(_12951_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3361),
    .D(_02479_),
    .Q_N(_12950_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3362),
    .D(_02480_),
    .Q_N(_14961_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3363),
    .D(_00044_),
    .Q_N(_12949_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3364),
    .D(_02481_),
    .Q_N(_12948_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3365),
    .D(_02482_),
    .Q_N(_14962_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3366),
    .D(_00045_),
    .Q_N(_14963_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3367),
    .D(_00046_),
    .Q_N(_14964_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3368),
    .D(_00047_),
    .Q_N(_14965_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3369),
    .D(_00048_),
    .Q_N(_14966_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3370),
    .D(_00049_),
    .Q_N(_14967_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3371),
    .D(_00050_),
    .Q_N(_14968_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3372),
    .D(_00051_),
    .Q_N(_12947_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3373),
    .D(_02483_),
    .Q_N(_12946_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3374),
    .D(_02484_),
    .Q_N(_12945_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3375),
    .D(_02485_),
    .Q_N(_12944_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3376),
    .D(_02486_),
    .Q_N(_12943_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3377),
    .D(_02487_),
    .Q_N(_12942_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3378),
    .D(_02488_),
    .Q_N(_12941_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3379),
    .D(_02489_),
    .Q_N(_14969_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3380),
    .D(_00055_),
    .Q_N(_00287_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3381),
    .D(_00056_),
    .Q_N(_14970_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3382),
    .D(_00057_),
    .Q_N(_14971_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3383),
    .D(_00058_),
    .Q_N(_14972_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3384),
    .D(_00059_),
    .Q_N(_14973_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3385),
    .D(_00060_),
    .Q_N(_14974_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3386),
    .D(_00061_),
    .Q_N(_14975_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3387),
    .D(_00062_),
    .Q_N(_14976_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3388),
    .D(_00063_),
    .Q_N(_14977_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3389),
    .D(_00064_),
    .Q_N(_14978_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3390),
    .D(_00065_),
    .Q_N(_14979_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3391),
    .D(_00066_),
    .Q_N(_14980_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3392),
    .D(_00067_),
    .Q_N(_14981_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3393),
    .D(_00068_),
    .Q_N(_14982_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3394),
    .D(_00069_),
    .Q_N(_14983_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3395),
    .D(_00070_),
    .Q_N(_14984_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3396),
    .D(_00071_),
    .Q_N(_14985_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3397),
    .D(_00072_),
    .Q_N(_14986_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3398),
    .D(_00073_),
    .Q_N(_14987_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3399),
    .D(_00074_),
    .Q_N(_14988_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3400),
    .D(_00075_),
    .Q_N(_14989_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3401),
    .D(_00076_),
    .Q_N(_14990_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3402),
    .D(_00077_),
    .Q_N(_14991_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3403),
    .D(_00078_),
    .Q_N(_12940_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3404),
    .D(_02490_),
    .Q_N(_12939_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3405),
    .D(_02491_),
    .Q_N(_12938_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3406),
    .D(_02492_),
    .Q_N(_12937_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3407),
    .D(_02493_),
    .Q_N(_12936_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3408),
    .D(_02494_),
    .Q_N(_12935_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3409),
    .D(_02495_),
    .Q_N(_12934_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3410),
    .D(_02496_),
    .Q_N(_12933_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3411),
    .D(_02497_),
    .Q_N(_12932_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3412),
    .D(_02498_),
    .Q_N(_12931_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3413),
    .D(_02499_),
    .Q_N(_12930_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3414),
    .D(_02500_),
    .Q_N(_12929_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3415),
    .D(_02501_),
    .Q_N(_12928_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3416),
    .D(_02502_),
    .Q_N(_12927_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3417),
    .D(_02503_),
    .Q_N(_12926_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3418),
    .D(_02504_),
    .Q_N(_12925_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3419),
    .D(_02505_),
    .Q_N(_12924_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3420),
    .D(_02506_),
    .Q_N(_12923_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3421),
    .D(_02507_),
    .Q_N(_12922_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3422),
    .D(_02508_),
    .Q_N(_12921_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3423),
    .D(_02509_),
    .Q_N(_12920_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3424),
    .D(_02510_),
    .Q_N(_12919_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3425),
    .D(_02511_),
    .Q_N(_12918_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3426),
    .D(_02512_),
    .Q_N(_12917_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3427),
    .D(_02513_),
    .Q_N(_12916_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3428),
    .D(_02514_),
    .Q_N(_00178_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3429),
    .D(_02515_),
    .Q_N(_12915_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3430),
    .D(_02516_),
    .Q_N(_00179_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net3431),
    .D(_02517_),
    .Q_N(_12914_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3432),
    .D(_02518_),
    .Q_N(_00254_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3433),
    .D(_02519_),
    .Q_N(_12913_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3434),
    .D(_02520_),
    .Q_N(_12912_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3435),
    .D(_02521_),
    .Q_N(_12911_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3436),
    .D(_02522_),
    .Q_N(_12910_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3437),
    .D(_02523_),
    .Q_N(_12909_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3438),
    .D(_02524_),
    .Q_N(_12908_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3439),
    .D(_02525_),
    .Q_N(_12907_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3440),
    .D(_02526_),
    .Q_N(_12906_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3441),
    .D(_02527_),
    .Q_N(_12905_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3442),
    .D(_02528_),
    .Q_N(_12904_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3443),
    .D(_02529_),
    .Q_N(_12903_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3444),
    .D(_02530_),
    .Q_N(_12902_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3445),
    .D(_02531_),
    .Q_N(_12901_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3446),
    .D(_02532_),
    .Q_N(_12900_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3447),
    .D(_02533_),
    .Q_N(_12899_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3448),
    .D(_02534_),
    .Q_N(_12898_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3449),
    .D(_02535_),
    .Q_N(_12897_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3450),
    .D(_02536_),
    .Q_N(_12896_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3451),
    .D(_02537_),
    .Q_N(_12895_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3452),
    .D(_02538_),
    .Q_N(_12894_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3453),
    .D(_02539_),
    .Q_N(_12893_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3454),
    .D(_02540_),
    .Q_N(_12892_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3455),
    .D(_02541_),
    .Q_N(_12891_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3456),
    .D(_02542_),
    .Q_N(_14992_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3457),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14993_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3458),
    .D(_00021_),
    .Q_N(_00279_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3459),
    .D(_00008_),
    .Q_N(_14994_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3460),
    .D(_00022_),
    .Q_N(_14995_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3461),
    .D(_00023_),
    .Q_N(_14996_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3462),
    .D(_00009_),
    .Q_N(_14997_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3463),
    .D(_00024_),
    .Q_N(_14998_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3464),
    .D(_00010_),
    .Q_N(_14999_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3465),
    .D(_00025_),
    .Q_N(_15000_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3466),
    .D(_00026_),
    .Q_N(_15001_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3467),
    .D(_00001_),
    .Q_N(_15002_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3468),
    .D(_00027_),
    .Q_N(_15003_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3469),
    .D(_00002_),
    .Q_N(_15004_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3470),
    .D(_00028_),
    .Q_N(_15005_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3471),
    .D(_00003_),
    .Q_N(_15006_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3472),
    .D(_00004_),
    .Q_N(_15007_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3473),
    .D(_00005_),
    .Q_N(_15008_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3474),
    .D(_00006_),
    .Q_N(_00180_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3475),
    .D(_00007_),
    .Q_N(_12890_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3476),
    .D(_02543_),
    .Q_N(_12889_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3477),
    .D(_02544_),
    .Q_N(_12888_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3478),
    .D(_02545_),
    .Q_N(_12887_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3479),
    .D(_02546_),
    .Q_N(_12886_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3480),
    .D(_02547_),
    .Q_N(_12885_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3481),
    .D(_02548_),
    .Q_N(_15009_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3482),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_15010_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3483),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00255_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3484),
    .D(_02549_),
    .Q_N(_12884_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3485),
    .D(_02550_),
    .Q_N(_12883_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3486),
    .D(_02551_),
    .Q_N(_12882_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3487),
    .D(_02552_),
    .Q_N(_12881_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3488),
    .D(_02553_),
    .Q_N(_00316_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3489),
    .D(_02554_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3490),
    .D(_02555_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3491),
    .D(_02556_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3492),
    .D(_02557_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3493),
    .D(_02558_),
    .Q_N(_00133_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3494),
    .D(_02559_),
    .Q_N(_00145_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3495),
    .D(_02560_),
    .Q_N(_00157_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3496),
    .D(_02561_),
    .Q_N(_00315_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3497),
    .D(_02562_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3498),
    .D(_02563_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3499),
    .D(_02564_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3500),
    .D(_02565_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3501),
    .D(_02566_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3502),
    .D(_02567_),
    .Q_N(_00144_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3503),
    .D(_02568_),
    .Q_N(_00156_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3504),
    .D(_02569_),
    .Q_N(_12880_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3505),
    .D(_02570_),
    .Q_N(_12879_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3506),
    .D(_02571_),
    .Q_N(_12878_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3507),
    .D(_02572_),
    .Q_N(_12877_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3508),
    .D(_02573_),
    .Q_N(_12876_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3509),
    .D(_02574_),
    .Q_N(_12875_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3510),
    .D(_02575_),
    .Q_N(_12874_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3511),
    .D(_02576_),
    .Q_N(_12873_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3512),
    .D(_02577_),
    .Q_N(_12872_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3513),
    .D(_02578_),
    .Q_N(_12871_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3514),
    .D(_02579_),
    .Q_N(_12870_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3515),
    .D(_02580_),
    .Q_N(_12869_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3516),
    .D(_02581_),
    .Q_N(_12868_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3517),
    .D(_02582_),
    .Q_N(_12867_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3518),
    .D(_02583_),
    .Q_N(_12866_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3519),
    .D(_02584_),
    .Q_N(_12865_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3520),
    .D(_02585_),
    .Q_N(_12864_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3521),
    .D(_02586_),
    .Q_N(_12863_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3522),
    .D(_02587_),
    .Q_N(_12862_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3523),
    .D(_02588_),
    .Q_N(_12861_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3524),
    .D(_02589_),
    .Q_N(_12860_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3525),
    .D(_02590_),
    .Q_N(_12859_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3526),
    .D(_02591_),
    .Q_N(_12858_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3527),
    .D(_02592_),
    .Q_N(_12857_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3528),
    .D(_02593_),
    .Q_N(_12856_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3529),
    .D(_02594_),
    .Q_N(_12855_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3530),
    .D(_02595_),
    .Q_N(_00224_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3531),
    .D(_02596_),
    .Q_N(_12854_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3532),
    .D(_02597_),
    .Q_N(_00226_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3533),
    .D(_02598_),
    .Q_N(_12853_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3534),
    .D(_02599_),
    .Q_N(_12852_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3535),
    .D(_02600_),
    .Q_N(_12851_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3536),
    .D(_02601_),
    .Q_N(_12850_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3537),
    .D(_02602_),
    .Q_N(_12849_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3538),
    .D(_02603_),
    .Q_N(_12848_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3539),
    .D(_02604_),
    .Q_N(_12847_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3540),
    .D(_02605_),
    .Q_N(_12846_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3541),
    .D(_02606_),
    .Q_N(_12845_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3542),
    .D(_02607_),
    .Q_N(_12844_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3543),
    .D(_02608_),
    .Q_N(_12843_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3544),
    .D(_02609_),
    .Q_N(_12842_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3545),
    .D(_02610_),
    .Q_N(_12841_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3546),
    .D(_02611_),
    .Q_N(_12840_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3547),
    .D(_02612_),
    .Q_N(_00223_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3548),
    .D(_02613_),
    .Q_N(_12839_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3549),
    .D(_02614_),
    .Q_N(_12838_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3550),
    .D(_02615_),
    .Q_N(_00284_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3551),
    .D(_02616_),
    .Q_N(_00285_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3552),
    .D(_02617_),
    .Q_N(_15011_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3553),
    .D(_00029_),
    .Q_N(_15012_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3554),
    .D(_00030_),
    .Q_N(_00227_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3555),
    .D(_00031_),
    .Q_N(_15013_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3556),
    .D(_00032_),
    .Q_N(_15014_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3557),
    .D(_00033_),
    .Q_N(_00280_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3558),
    .D(_00034_),
    .Q_N(_15015_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3559),
    .D(_00035_),
    .Q_N(_00228_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3560),
    .D(_02618_),
    .Q_N(_12837_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3561),
    .D(_02619_),
    .Q_N(_12836_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3562),
    .D(_02620_),
    .Q_N(_12835_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3563),
    .D(_02621_),
    .Q_N(_12834_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3564),
    .D(_02622_),
    .Q_N(_12833_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3565),
    .D(_02623_),
    .Q_N(_12832_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3566),
    .D(_02624_),
    .Q_N(_12831_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3567),
    .D(_02625_),
    .Q_N(_12830_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3568),
    .D(_02626_),
    .Q_N(_00286_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3569),
    .D(_02627_),
    .Q_N(_12829_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3570),
    .D(_02628_),
    .Q_N(_12828_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3571),
    .D(_02629_),
    .Q_N(_12827_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3572),
    .D(_02630_),
    .Q_N(_12826_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3573),
    .D(_02631_),
    .Q_N(_12825_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3574),
    .D(_02632_),
    .Q_N(_12824_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3575),
    .D(_02633_),
    .Q_N(_15016_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3576),
    .D(_00079_),
    .Q_N(_00281_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3577),
    .D(_00080_),
    .Q_N(_15017_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3578),
    .D(_00081_),
    .Q_N(_15018_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3579),
    .D(_00082_),
    .Q_N(_15019_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3580),
    .D(_00083_),
    .Q_N(_15020_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3581),
    .D(_00084_),
    .Q_N(_15021_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3582),
    .D(_00085_),
    .Q_N(_15022_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3583),
    .D(_00086_),
    .Q_N(_15023_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3584),
    .D(_00087_),
    .Q_N(_15024_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3585),
    .D(_00088_),
    .Q_N(_15025_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3586),
    .D(_00089_),
    .Q_N(_15026_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3587),
    .D(_00090_),
    .Q_N(_12823_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3588),
    .D(_02634_),
    .Q_N(_12822_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3589),
    .D(_02635_),
    .Q_N(_12821_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3590),
    .D(_02636_),
    .Q_N(_12820_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3591),
    .D(_02637_),
    .Q_N(_12819_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3592),
    .D(_02638_),
    .Q_N(_12818_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3593),
    .D(_02639_),
    .Q_N(_12817_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3594),
    .D(_02640_),
    .Q_N(_12816_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3595),
    .D(_02641_),
    .Q_N(_12815_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3596),
    .D(_02642_),
    .Q_N(_12814_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3597),
    .D(_02643_),
    .Q_N(_12813_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3598),
    .D(_02644_),
    .Q_N(_12812_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3599),
    .D(_02645_),
    .Q_N(_12811_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3600),
    .D(_02646_),
    .Q_N(_12810_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3601),
    .D(_02647_),
    .Q_N(_12809_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3602),
    .D(_02648_),
    .Q_N(_12808_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3603),
    .D(_02649_),
    .Q_N(_12807_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3604),
    .D(_02650_),
    .Q_N(_12806_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3605),
    .D(_02651_),
    .Q_N(_12805_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3606),
    .D(_02652_),
    .Q_N(_12804_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3607),
    .D(_02653_),
    .Q_N(_12803_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3608),
    .D(_02654_),
    .Q_N(_12802_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3609),
    .D(_02655_),
    .Q_N(_12801_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3610),
    .D(_02656_),
    .Q_N(_12800_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3611),
    .D(_02657_),
    .Q_N(_12799_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3612),
    .D(_02658_),
    .Q_N(_12798_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3613),
    .D(_02659_),
    .Q_N(_12797_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3614),
    .D(_02660_),
    .Q_N(_12796_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3615),
    .D(_02661_),
    .Q_N(_12795_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3616),
    .D(_02662_),
    .Q_N(_12794_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3617),
    .D(_02663_),
    .Q_N(_12793_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3618),
    .D(_02664_),
    .Q_N(_12792_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3619),
    .D(_02665_),
    .Q_N(_12791_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3620),
    .D(_02666_),
    .Q_N(_12790_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3621),
    .D(_02667_),
    .Q_N(_12789_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3622),
    .D(_02668_),
    .Q_N(_15027_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3623),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12788_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3624),
    .D(_02669_),
    .Q_N(_12787_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3625),
    .D(_02670_),
    .Q_N(_12786_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3626),
    .D(_02671_),
    .Q_N(_12785_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3627),
    .D(_02672_),
    .Q_N(_12784_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3628),
    .D(_02673_),
    .Q_N(_12783_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3629),
    .D(_02674_),
    .Q_N(_12782_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3630),
    .D(_02675_),
    .Q_N(_12781_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3631),
    .D(_02676_),
    .Q_N(_12780_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3632),
    .D(_02677_),
    .Q_N(_12779_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3633),
    .D(_02678_),
    .Q_N(_12778_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3634),
    .D(_02679_),
    .Q_N(_00282_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3635),
    .D(_02680_),
    .Q_N(_12777_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3636),
    .D(_02681_),
    .Q_N(_12776_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3637),
    .D(_02682_),
    .Q_N(_12775_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3638),
    .D(_02683_),
    .Q_N(_12774_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3639),
    .D(_02684_),
    .Q_N(_12773_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3640),
    .D(_02685_),
    .Q_N(_15028_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3641),
    .D(_00000_),
    .Q_N(_12772_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_03839_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_03838_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_06730_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07911_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_07125_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_07051_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_04227_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02953_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02900_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02835_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02801_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02776_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02768_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02704_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_12754_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12729_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12721_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12671_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12627_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12602_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12594_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12544_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12492_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12422_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12388_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12363_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12355_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12289_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12241_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12207_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12194_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_07006_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_02927_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_02892_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12516_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_12484_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_11762_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_11728_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_11705_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_10049_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_10038_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_10037_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_07450_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_05377_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_05292_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_05291_));
 sg13g2_buf_2 fanout73 (.A(_05182_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_05178_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04238_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_04098_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_11624_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_11588_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_07596_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_05009_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_05006_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04821_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04820_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_04214_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_11612_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_11583_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_09359_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_07886_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_07484_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_07442_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_07441_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_07419_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_07222_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_07221_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_07218_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_06848_),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(_06712_));
 sg13g2_buf_2 fanout98 (.A(_04328_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04313_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04132_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_03288_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_03190_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_10182_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_10159_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_10149_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_09358_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09121_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_09052_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_07689_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_07643_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_07620_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_07609_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_07587_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_07583_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_07217_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_04390_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04318_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04276_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_04200_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_04195_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_04183_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_04165_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_04162_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04131_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_03767_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_03705_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_03699_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_03685_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_03205_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_03195_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_03085_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_11770_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_11458_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_10158_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_10150_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_10148_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_10034_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_09941_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_09833_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_09132_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_09120_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_09051_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_08897_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_07582_),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_06718_));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_06715_));
 sg13g2_buf_2 fanout147 (.A(_04207_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_04205_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_04186_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_04180_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_04178_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_04176_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_04166_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04153_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04151_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04149_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04139_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04130_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04102_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04099_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_03754_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03743_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03681_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03672_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03621_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03576_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_11832_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_11547_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_11356_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_10143_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_10100_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_09855_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_08997_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_08896_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_07097_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_05243_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_05137_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_04297_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_04148_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_04138_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_04101_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03725_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03634_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_03231_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03200_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03074_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_11744_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_11607_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_11570_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_11491_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_11460_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_10142_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_10032_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_09113_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_04320_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_04095_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03573_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_03259_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_03185_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_03095_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_03090_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_03087_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_03086_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_03071_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_11745_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_11673_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_11507_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_11383_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_09957_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_05809_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_04201_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_03706_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03266_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03131_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03089_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_03079_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_03077_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03076_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_03072_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03070_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_11638_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_11255_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_11229_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_11190_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_11126_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_11093_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_11064_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_10533_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_09956_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_09127_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_09111_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_06357_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_06312_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_06267_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_06258_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_06225_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_06182_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_06173_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_06163_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_06132_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_06086_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_06075_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_06046_),
    .X(net243));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(_06037_));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_06015_));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_05996_));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_05989_));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(_05972_));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(_05956_));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_05953_));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_05945_));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(_05924_));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(_05905_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_05898_));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_05871_));
 sg13g2_buf_2 fanout256 (.A(_03078_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_03075_),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_03056_));
 sg13g2_buf_2 fanout259 (.A(_03054_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_11249_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_11246_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_11242_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_11219_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_11161_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_11155_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_11015_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_10980_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_10799_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_10478_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_09930_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_09912_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_09907_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_09158_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_09071_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_08456_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_06592_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_06590_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_06589_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_06356_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_06348_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_06339_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_06330_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_06321_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_06311_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_06303_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_06294_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_06285_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_06276_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_06266_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_06257_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_06248_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_06235_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_06224_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_06209_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_06200_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_06191_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06181_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06172_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06162_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_06154_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_06145_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_06131_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_06122_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06105_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06095_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06085_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06074_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06065_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06056_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06045_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_06034_));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_06031_));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_06026_));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_06020_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_06011_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_06008_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_06005_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_06002_));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_05982_));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_05977_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_05968_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05962_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_05959_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_05938_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_05931_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05920_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_05913_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_05909_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_05892_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_05884_));
 sg13g2_buf_2 fanout331 (.A(_03856_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_03832_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_03162_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_03092_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_12667_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_11574_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_11222_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_10798_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_10477_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_10272_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_09895_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_09175_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_09125_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_09046_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_09015_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_08993_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_08918_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_06673_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_06671_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_06670_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_06631_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06629_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06628_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_06615_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_06608_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_06571_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_06569_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_06568_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_06495_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_06494_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_06347_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_06338_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_06329_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_06320_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_06302_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_06293_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_06284_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_06275_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_06247_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_06234_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_06208_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_06199_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_06190_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_06153_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_06144_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_06121_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_06104_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_06094_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_06064_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_06055_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_04894_),
    .X(net381));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_03068_));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_03067_));
 sg13g2_buf_2 fanout384 (.A(_10156_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_09657_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_09642_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_09321_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_09217_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_09124_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_09069_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_08805_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_08784_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_08762_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_08738_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_08715_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_08487_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_06694_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_06692_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_06691_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_06652_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_06650_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_06649_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_06553_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_06546_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_06431_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_06430_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_05477_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_05032_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_05031_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_05026_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_04945_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_04925_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_04903_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_04892_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_04888_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_04883_),
    .X(net416));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(_03060_));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_03059_));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(_03053_));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_03052_));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_03050_));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_03049_));
 sg13g2_buf_2 fanout423 (.A(_02955_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_12665_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_11593_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_10155_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_09724_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_09701_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_09680_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_09610_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_09589_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_09574_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_09543_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_09513_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_09485_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_08670_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_08587_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_06781_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_06237_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_06134_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_06102_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_06053_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_05993_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_05942_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_05906_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_05876_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_05875_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_05184_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_05183_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_05030_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_04961_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_04957_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_04891_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_04882_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_04846_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_04758_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_04754_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_03811_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_03782_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_03536_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_03531_),
    .X(net461));
 sg13g2_buf_1 fanout462 (.A(_03529_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_03115_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_03062_));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_03061_));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(_03040_));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_03022_));
 sg13g2_buf_2 fanout468 (.A(_03021_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_02890_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_02706_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_12664_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_12546_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_12535_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_12424_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_12166_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_12157_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_12131_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_12127_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_12123_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_12117_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_12108_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_12098_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_10269_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_10204_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_10025_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_08691_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_08615_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_08556_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_08500_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_08398_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_07912_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_07477_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_06366_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_06365_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_06364_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_05973_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_05921_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_04963_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_04960_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_04959_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_04956_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_04890_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_04881_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_04862_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_04857_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_04756_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_04747_),
    .X(net507));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(_04740_));
 sg13g2_buf_2 fanout509 (.A(_04115_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_03810_),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_03566_));
 sg13g2_buf_2 fanout512 (.A(_03563_),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_03562_));
 sg13g2_buf_2 fanout514 (.A(_03555_),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_03554_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(_03539_));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(_03535_));
 sg13g2_buf_2 fanout518 (.A(_03534_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_03533_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_03528_),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_03525_));
 sg13g2_buf_2 fanout522 (.A(_03118_),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_03117_));
 sg13g2_buf_2 fanout524 (.A(_03114_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(_03041_));
 sg13g2_buf_2 fanout526 (.A(_03039_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_02837_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_12718_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_12663_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_12534_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_12482_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_12352_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_12293_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_12153_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_11630_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_11622_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_11516_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_10538_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_10481_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_10358_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_10292_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_10153_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_10137_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_10094_));
 sg13g2_buf_2 fanout545 (.A(_10024_),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(_09021_));
 sg13g2_buf_2 fanout547 (.A(_08931_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_08616_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_08522_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_08506_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_08499_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_07954_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_07919_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_07878_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_07782_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_07711_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_07678_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_07663_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_07640_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_07617_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_07575_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_07544_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_07510_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_07446_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_07430_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_07340_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_06789_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_06238_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_06232_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_06135_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_06129_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_05998_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_05963_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_05947_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_05910_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_05886_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_05153_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_05146_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_05140_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_04869_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_04842_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_04835_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_03789_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_03783_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_03776_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_03775_),
    .X(net586));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(_03559_));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(_03550_));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_03544_));
 sg13g2_buf_2 fanout590 (.A(_03532_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_03526_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_03038_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_02765_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_12591_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_12044_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_12011_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_11621_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_11523_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_11257_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_11100_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_10937_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_10334_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_10326_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_10318_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_10314_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_10302_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_10297_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_10291_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_10248_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_10247_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_10093_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_10023_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_10021_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_09850_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_09547_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_09516_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_09493_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_09457_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_09454_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_09447_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_09438_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_09382_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_09369_),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(_09223_));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(_09002_));
 sg13g2_buf_2 fanout626 (.A(_08956_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_08930_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_08925_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_08739_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_08716_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_08588_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_08557_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_08521_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_08516_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_08511_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_08505_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_08498_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_07854_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_07129_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_06242_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_06212_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_06139_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_06108_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_05999_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_05948_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_05887_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_05838_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_05042_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_04982_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_04979_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_03796_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_03795_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_03788_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_03785_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_03778_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_03527_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_03020_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_12189_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_12054_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_12015_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_12014_),
    .X(net661));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(_12010_));
 sg13g2_buf_2 fanout663 (.A(_12004_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_11413_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10989_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_10749_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_10662_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_10624_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_10540_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_10507_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_10499_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_10350_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_10337_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_10317_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_10313_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_10301_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_10296_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_10092_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_10030_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_10022_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_10020_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_09889_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_09489_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_09446_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_09442_),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(_09422_));
 sg13g2_buf_2 fanout687 (.A(_09416_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_09413_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_09394_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_09390_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_09365_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_09364_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_09310_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_09237_),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(_09222_));
 sg13g2_buf_2 fanout696 (.A(_09122_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_08819_),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(_08810_));
 sg13g2_buf_2 fanout699 (.A(_08766_),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_08704_));
 sg13g2_buf_2 fanout701 (.A(_08649_),
    .X(net701));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_08642_));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(_08634_));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_08629_));
 sg13g2_buf_2 fanout705 (.A(_08620_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_08593_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_08561_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_08520_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_08515_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_08510_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_08504_),
    .X(net711));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_08474_));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_08470_));
 sg13g2_buf_2 fanout714 (.A(_08466_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_06244_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_06217_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_06216_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_06214_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_06141_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_06113_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_06112_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_06110_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_05997_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_05946_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_05914_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_05885_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_05878_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_05808_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_04743_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_04742_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_03780_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_03556_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_03530_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_03483_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_03099_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_03064_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_03063_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_03045_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_03044_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_03043_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_03031_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_03029_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_03026_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_03019_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_12188_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_12024_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_12009_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_12001_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_11946_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_11936_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_11580_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_11144_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_10966_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_10955_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_10733_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_10558_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_10509_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_10506_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_10502_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_10484_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_10432_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10431_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10346_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_10339_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_10336_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_10332_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_10316_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_10307_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_10300_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_10295_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_10091_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_10019_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_09853_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_09824_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_09728_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_09710_),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(_09628_),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(_09625_),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(_09566_));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_09565_));
 sg13g2_buf_8 fanout781 (.A(_09509_),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(_09506_),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(_09473_),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(_09470_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_09460_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_09430_),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_09419_));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(_09412_));
 sg13g2_buf_8 fanout789 (.A(_09410_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_09408_));
 sg13g2_buf_8 fanout791 (.A(_09407_),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_09403_));
 sg13g2_buf_8 fanout793 (.A(_09401_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_09393_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_09363_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_09314_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_09309_),
    .X(net797));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_09236_));
 sg13g2_buf_2 fanout799 (.A(_09221_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_08920_),
    .X(net800));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_08743_));
 sg13g2_buf_2 fanout802 (.A(_08719_),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(_08703_),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(_08641_),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_08637_));
 sg13g2_buf_8 fanout806 (.A(_08633_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_08628_),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(_08627_),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_08617_));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_08597_));
 sg13g2_buf_2 fanout811 (.A(_08560_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_08534_),
    .X(net812));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_08531_));
 sg13g2_buf_2 fanout814 (.A(_08528_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_08525_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_08509_),
    .X(net816));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_08476_));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_08473_));
 sg13g2_buf_8 fanout819 (.A(_08469_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_08465_),
    .X(net820));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(_08463_));
 sg13g2_buf_2 fanout822 (.A(_08443_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_08411_),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_08314_));
 sg13g2_buf_2 fanout825 (.A(_07041_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_07007_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_06852_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_06847_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_06824_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_06819_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_06220_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_06219_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_06218_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_06116_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_06115_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_06114_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_05984_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_05983_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_05969_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_05933_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_05932_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_05874_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_05873_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_05845_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_05843_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_04822_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_04109_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_03692_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_03518_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_03098_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_03069_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_03066_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_03065_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_03051_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_03048_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_03046_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_03042_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_03037_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_03035_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_03033_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_03030_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_03028_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_03025_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_12766_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_12581_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_12255_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_12250_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_12201_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_12069_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_12030_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_12008_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_12000_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_11993_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_11979_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_11444_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_11122_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_11095_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_11068_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_10653_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_10633_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_10557_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_10446_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_10435_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_10430_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_10425_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_10417_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_10415_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_10403_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_10323_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_10315_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_10311_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_10299_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_10294_),
    .X(net893));
 sg13g2_buf_1 fanout894 (.A(_10188_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_10181_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_10170_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_10165_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_10145_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_10133_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_10090_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_10082_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_10018_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_09926_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_09742_),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_09635_));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(_09629_));
 sg13g2_buf_2 fanout907 (.A(_09558_),
    .X(net907));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(_09537_));
 sg13g2_buf_2 fanout909 (.A(_09524_),
    .X(net909));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(_09479_));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(_09471_));
 sg13g2_buf_2 fanout912 (.A(_09435_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_09402_),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(_09400_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_09313_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_09308_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_09304_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09235_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_09220_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_08919_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_08875_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_08852_),
    .X(net922));
 sg13g2_buf_4 fanout923 (.X(net923),
    .A(_08632_));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_08595_));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_08580_));
 sg13g2_buf_2 fanout926 (.A(_08565_),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_08542_));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(_08533_));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(_08530_));
 sg13g2_buf_2 fanout930 (.A(_08524_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_08508_),
    .X(net931));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_08484_));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(_08475_));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_08464_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_08462_));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_08377_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_08303_));
 sg13g2_buf_2 fanout938 (.A(_07111_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_07102_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_07100_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_07087_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_07084_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_07040_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_07010_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_06874_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_06794_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_06511_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_06510_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_06509_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_06507_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_06491_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_06490_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_06488_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_06486_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_06479_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_06478_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_06477_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_06474_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_06455_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_06454_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_06453_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_06450_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_06447_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_06444_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_06441_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_06438_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_06418_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_06413_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_06406_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_06395_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_05992_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_05991_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_05990_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_05964_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05941_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05940_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_05939_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_05925_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_05872_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_05851_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_05841_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_05832_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_05293_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_04849_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_04733_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_04614_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_04581_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_04229_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_03900_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_03517_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_03036_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_03034_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_03032_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_03005_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_02759_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_02755_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_02751_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_02747_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_12762_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_12694_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_12659_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_12655_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_12643_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_12628_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_12541_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_12454_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_12447_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_12443_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_12437_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_12339_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_12335_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_12283_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_12279_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_12275_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_12271_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_12260_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_12257_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_12252_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_12247_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_12227_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_12220_),
    .X(net1021));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(_12216_));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(_12209_));
 sg13g2_buf_2 fanout1024 (.A(_12196_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_12080_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_12062_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_12057_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_11980_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_11978_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_11945_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_11120_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_10945_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_10942_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_10416_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_10414_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_10410_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_10404_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_10402_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_10373_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_10364_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_10362_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_10310_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_10303_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_10298_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_10293_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_10257_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_10176_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_10164_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_10144_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_10132_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_10129_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_10123_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_10117_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_10111_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_10106_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_10088_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_10081_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_10027_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_09922_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_09866_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_09737_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_09523_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_09449_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_09318_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_09311_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_09307_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_09239_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_09234_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_09229_),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(_09227_));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(_09225_));
 sg13g2_buf_2 fanout1072 (.A(_09219_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_09203_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_09196_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_09131_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_09038_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_09006_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_08899_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_08883_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_08825_),
    .X(net1080));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(_08579_));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(_08541_));
 sg13g2_buf_2 fanout1083 (.A(_08540_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_08529_),
    .X(net1084));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(_08526_));
 sg13g2_buf_2 fanout1086 (.A(_08489_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_08483_),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(_08461_));
 sg13g2_buf_1 fanout1089 (.A(_08460_),
    .X(net1089));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(_08369_));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(_08367_));
 sg13g2_buf_2 fanout1092 (.A(_08362_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_08334_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_08316_),
    .X(net1094));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(_08302_));
 sg13g2_buf_4 fanout1096 (.X(net1096),
    .A(_08300_));
 sg13g2_buf_2 fanout1097 (.A(_08296_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_08097_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_08095_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_08079_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_07799_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_07177_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_07101_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_07098_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_07085_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_07083_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_05819_),
    .X(net1107));
 sg13g2_buf_4 fanout1108 (.X(net1108),
    .A(_02933_));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(_02922_));
 sg13g2_buf_4 fanout1110 (.X(net1110),
    .A(_02918_));
 sg13g2_buf_2 fanout1111 (.A(_02909_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_12226_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_12215_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_12208_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_12195_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_12119_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_12104_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_12087_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_12082_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_12052_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_12048_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_12029_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_12027_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_12021_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_11838_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_11433_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_11218_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_10375_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_10374_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_10259_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_10255_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_10253_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_10110_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_09921_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_09890_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_09886_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_09862_),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_09856_),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(_09758_),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(_09431_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_09392_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_09372_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_09356_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_09300_),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_09289_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(_09218_),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(_09130_),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(_09037_),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(_08492_),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(_08491_),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(_08403_),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(_08400_),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(_08372_));
 sg13g2_buf_2 fanout1154 (.A(_08352_),
    .X(net1154));
 sg13g2_buf_2 fanout1155 (.A(_08349_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(_08297_),
    .X(net1156));
 sg13g2_tiehi _27611__1157 (.L_HI(net1157));
 sg13g2_tiehi _27612__1158 (.L_HI(net1158));
 sg13g2_tiehi _27613__1159 (.L_HI(net1159));
 sg13g2_tiehi _27614__1160 (.L_HI(net1160));
 sg13g2_tiehi _27615__1161 (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.dec.r_rs2_inv$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_count[0]$_SDFFE_PN0P__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_count[1]$_SDFFE_PN0P__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_count[2]$_SDFFE_PN0P__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_count[3]$_SDFFE_PN0P__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_count[4]$_SDFFE_PN0P__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_count[5]$_SDFFE_PN0P__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_count[6]$_SDFFE_PN0P__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_count[7]$_SDFFE_PN0P__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_SDFFE_PN0P__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_SDFFE_PN0P__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_SDFFE_PN0P__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_SDFFE_PN0P__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_SDFFE_PN0P__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_SDFFE_PN0P__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.spi.r_src[0]$_SDFFE_PN0P__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.spi.r_src[1]$_SDFFE_PN0P__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.spi.r_src[2]$_SDFFE_PN0P__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3614  (.L_HI(net3614));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3615  (.L_HI(net3615));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3616  (.L_HI(net3616));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3617  (.L_HI(net3617));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3618  (.L_HI(net3618));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3619  (.L_HI(net3619));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3620  (.L_HI(net3620));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3621  (.L_HI(net3621));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3622  (.L_HI(net3622));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3623  (.L_HI(net3623));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3624  (.L_HI(net3624));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3625  (.L_HI(net3625));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3626  (.L_HI(net3626));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3627  (.L_HI(net3627));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3628  (.L_HI(net3628));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3629  (.L_HI(net3629));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3630  (.L_HI(net3630));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3631  (.L_HI(net3631));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3632  (.L_HI(net3632));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3633  (.L_HI(net3633));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3634  (.L_HI(net3634));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3635  (.L_HI(net3635));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3636  (.L_HI(net3636));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3637  (.L_HI(net3637));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3638  (.L_HI(net3638));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3639  (.L_HI(net3639));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3640  (.L_HI(net3640));
 sg13g2_tiehi \r_reset$_DFF_P__3641  (.L_HI(net3641));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_310_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_131_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2 (.A(_00000_));
 sg13g2_antennanp ANTENNA_3 (.A(_00230_));
 sg13g2_antennanp ANTENNA_4 (.A(_00237_));
 sg13g2_antennanp ANTENNA_5 (.A(_00237_));
 sg13g2_antennanp ANTENNA_6 (.A(_00237_));
 sg13g2_antennanp ANTENNA_7 (.A(_00752_));
 sg13g2_antennanp ANTENNA_8 (.A(_00752_));
 sg13g2_antennanp ANTENNA_9 (.A(_00800_));
 sg13g2_antennanp ANTENNA_10 (.A(_00800_));
 sg13g2_antennanp ANTENNA_11 (.A(_01061_));
 sg13g2_antennanp ANTENNA_12 (.A(_01063_));
 sg13g2_antennanp ANTENNA_13 (.A(_02909_));
 sg13g2_antennanp ANTENNA_14 (.A(_02909_));
 sg13g2_antennanp ANTENNA_15 (.A(_02909_));
 sg13g2_antennanp ANTENNA_16 (.A(_02909_));
 sg13g2_antennanp ANTENNA_17 (.A(_02909_));
 sg13g2_antennanp ANTENNA_18 (.A(_02909_));
 sg13g2_antennanp ANTENNA_19 (.A(_02909_));
 sg13g2_antennanp ANTENNA_20 (.A(_02909_));
 sg13g2_antennanp ANTENNA_21 (.A(_02909_));
 sg13g2_antennanp ANTENNA_22 (.A(_02918_));
 sg13g2_antennanp ANTENNA_23 (.A(_02918_));
 sg13g2_antennanp ANTENNA_24 (.A(_02918_));
 sg13g2_antennanp ANTENNA_25 (.A(_02918_));
 sg13g2_antennanp ANTENNA_26 (.A(_02918_));
 sg13g2_antennanp ANTENNA_27 (.A(_02918_));
 sg13g2_antennanp ANTENNA_28 (.A(_02918_));
 sg13g2_antennanp ANTENNA_29 (.A(_02918_));
 sg13g2_antennanp ANTENNA_30 (.A(_02918_));
 sg13g2_antennanp ANTENNA_31 (.A(_02922_));
 sg13g2_antennanp ANTENNA_32 (.A(_02922_));
 sg13g2_antennanp ANTENNA_33 (.A(_02922_));
 sg13g2_antennanp ANTENNA_34 (.A(_02922_));
 sg13g2_antennanp ANTENNA_35 (.A(_02922_));
 sg13g2_antennanp ANTENNA_36 (.A(_02922_));
 sg13g2_antennanp ANTENNA_37 (.A(_02922_));
 sg13g2_antennanp ANTENNA_38 (.A(_02922_));
 sg13g2_antennanp ANTENNA_39 (.A(_02922_));
 sg13g2_antennanp ANTENNA_40 (.A(_02933_));
 sg13g2_antennanp ANTENNA_41 (.A(_02933_));
 sg13g2_antennanp ANTENNA_42 (.A(_02933_));
 sg13g2_antennanp ANTENNA_43 (.A(_02933_));
 sg13g2_antennanp ANTENNA_44 (.A(_02933_));
 sg13g2_antennanp ANTENNA_45 (.A(_02933_));
 sg13g2_antennanp ANTENNA_46 (.A(_02933_));
 sg13g2_antennanp ANTENNA_47 (.A(_02933_));
 sg13g2_antennanp ANTENNA_48 (.A(_02933_));
 sg13g2_antennanp ANTENNA_49 (.A(_03019_));
 sg13g2_antennanp ANTENNA_50 (.A(_03019_));
 sg13g2_antennanp ANTENNA_51 (.A(_03019_));
 sg13g2_antennanp ANTENNA_52 (.A(_03020_));
 sg13g2_antennanp ANTENNA_53 (.A(_03020_));
 sg13g2_antennanp ANTENNA_54 (.A(_03020_));
 sg13g2_antennanp ANTENNA_55 (.A(_03161_));
 sg13g2_antennanp ANTENNA_56 (.A(_03533_));
 sg13g2_antennanp ANTENNA_57 (.A(_03533_));
 sg13g2_antennanp ANTENNA_58 (.A(_03533_));
 sg13g2_antennanp ANTENNA_59 (.A(_03533_));
 sg13g2_antennanp ANTENNA_60 (.A(_03535_));
 sg13g2_antennanp ANTENNA_61 (.A(_03535_));
 sg13g2_antennanp ANTENNA_62 (.A(_03535_));
 sg13g2_antennanp ANTENNA_63 (.A(_03535_));
 sg13g2_antennanp ANTENNA_64 (.A(_03535_));
 sg13g2_antennanp ANTENNA_65 (.A(_03535_));
 sg13g2_antennanp ANTENNA_66 (.A(_03535_));
 sg13g2_antennanp ANTENNA_67 (.A(_03535_));
 sg13g2_antennanp ANTENNA_68 (.A(_04699_));
 sg13g2_antennanp ANTENNA_69 (.A(_04699_));
 sg13g2_antennanp ANTENNA_70 (.A(_04699_));
 sg13g2_antennanp ANTENNA_71 (.A(_04699_));
 sg13g2_antennanp ANTENNA_72 (.A(_04843_));
 sg13g2_antennanp ANTENNA_73 (.A(_04890_));
 sg13g2_antennanp ANTENNA_74 (.A(_04890_));
 sg13g2_antennanp ANTENNA_75 (.A(_04890_));
 sg13g2_antennanp ANTENNA_76 (.A(_04890_));
 sg13g2_antennanp ANTENNA_77 (.A(_04914_));
 sg13g2_antennanp ANTENNA_78 (.A(_04954_));
 sg13g2_antennanp ANTENNA_79 (.A(_05005_));
 sg13g2_antennanp ANTENNA_80 (.A(_05175_));
 sg13g2_antennanp ANTENNA_81 (.A(_05207_));
 sg13g2_antennanp ANTENNA_82 (.A(_05231_));
 sg13g2_antennanp ANTENNA_83 (.A(_05267_));
 sg13g2_antennanp ANTENNA_84 (.A(_05282_));
 sg13g2_antennanp ANTENNA_85 (.A(_05373_));
 sg13g2_antennanp ANTENNA_86 (.A(_05437_));
 sg13g2_antennanp ANTENNA_87 (.A(_05577_));
 sg13g2_antennanp ANTENNA_88 (.A(_05649_));
 sg13g2_antennanp ANTENNA_89 (.A(_05722_));
 sg13g2_antennanp ANTENNA_90 (.A(_05737_));
 sg13g2_antennanp ANTENNA_91 (.A(_05783_));
 sg13g2_antennanp ANTENNA_92 (.A(_05789_));
 sg13g2_antennanp ANTENNA_93 (.A(_05795_));
 sg13g2_antennanp ANTENNA_94 (.A(_05800_));
 sg13g2_antennanp ANTENNA_95 (.A(_05800_));
 sg13g2_antennanp ANTENNA_96 (.A(_05805_));
 sg13g2_antennanp ANTENNA_97 (.A(_05838_));
 sg13g2_antennanp ANTENNA_98 (.A(_05838_));
 sg13g2_antennanp ANTENNA_99 (.A(_05838_));
 sg13g2_antennanp ANTENNA_100 (.A(_06038_));
 sg13g2_antennanp ANTENNA_101 (.A(_06479_));
 sg13g2_antennanp ANTENNA_102 (.A(_06479_));
 sg13g2_antennanp ANTENNA_103 (.A(_06479_));
 sg13g2_antennanp ANTENNA_104 (.A(_06479_));
 sg13g2_antennanp ANTENNA_105 (.A(_06479_));
 sg13g2_antennanp ANTENNA_106 (.A(_06479_));
 sg13g2_antennanp ANTENNA_107 (.A(_06479_));
 sg13g2_antennanp ANTENNA_108 (.A(_06479_));
 sg13g2_antennanp ANTENNA_109 (.A(_06479_));
 sg13g2_antennanp ANTENNA_110 (.A(_06822_));
 sg13g2_antennanp ANTENNA_111 (.A(_06856_));
 sg13g2_antennanp ANTENNA_112 (.A(_06905_));
 sg13g2_antennanp ANTENNA_113 (.A(_06949_));
 sg13g2_antennanp ANTENNA_114 (.A(_06978_));
 sg13g2_antennanp ANTENNA_115 (.A(_07663_));
 sg13g2_antennanp ANTENNA_116 (.A(_07663_));
 sg13g2_antennanp ANTENNA_117 (.A(_07663_));
 sg13g2_antennanp ANTENNA_118 (.A(_07663_));
 sg13g2_antennanp ANTENNA_119 (.A(_08220_));
 sg13g2_antennanp ANTENNA_120 (.A(_08220_));
 sg13g2_antennanp ANTENNA_121 (.A(_08377_));
 sg13g2_antennanp ANTENNA_122 (.A(_08377_));
 sg13g2_antennanp ANTENNA_123 (.A(_08377_));
 sg13g2_antennanp ANTENNA_124 (.A(_08411_));
 sg13g2_antennanp ANTENNA_125 (.A(_08411_));
 sg13g2_antennanp ANTENNA_126 (.A(_08411_));
 sg13g2_antennanp ANTENNA_127 (.A(_08411_));
 sg13g2_antennanp ANTENNA_128 (.A(_08443_));
 sg13g2_antennanp ANTENNA_129 (.A(_08443_));
 sg13g2_antennanp ANTENNA_130 (.A(_08443_));
 sg13g2_antennanp ANTENNA_131 (.A(_08486_));
 sg13g2_antennanp ANTENNA_132 (.A(_08491_));
 sg13g2_antennanp ANTENNA_133 (.A(_08491_));
 sg13g2_antennanp ANTENNA_134 (.A(_08491_));
 sg13g2_antennanp ANTENNA_135 (.A(_08556_));
 sg13g2_antennanp ANTENNA_136 (.A(_08556_));
 sg13g2_antennanp ANTENNA_137 (.A(_08556_));
 sg13g2_antennanp ANTENNA_138 (.A(_08565_));
 sg13g2_antennanp ANTENNA_139 (.A(_08565_));
 sg13g2_antennanp ANTENNA_140 (.A(_08565_));
 sg13g2_antennanp ANTENNA_141 (.A(_08565_));
 sg13g2_antennanp ANTENNA_142 (.A(_08669_));
 sg13g2_antennanp ANTENNA_143 (.A(_08691_));
 sg13g2_antennanp ANTENNA_144 (.A(_08691_));
 sg13g2_antennanp ANTENNA_145 (.A(_08691_));
 sg13g2_antennanp ANTENNA_146 (.A(_08735_));
 sg13g2_antennanp ANTENNA_147 (.A(_08784_));
 sg13g2_antennanp ANTENNA_148 (.A(_08784_));
 sg13g2_antennanp ANTENNA_149 (.A(_08784_));
 sg13g2_antennanp ANTENNA_150 (.A(_08804_));
 sg13g2_antennanp ANTENNA_151 (.A(_08839_));
 sg13g2_antennanp ANTENNA_152 (.A(_08839_));
 sg13g2_antennanp ANTENNA_153 (.A(_08839_));
 sg13g2_antennanp ANTENNA_154 (.A(_08894_));
 sg13g2_antennanp ANTENNA_155 (.A(_08894_));
 sg13g2_antennanp ANTENNA_156 (.A(_08894_));
 sg13g2_antennanp ANTENNA_157 (.A(_08940_));
 sg13g2_antennanp ANTENNA_158 (.A(_08976_));
 sg13g2_antennanp ANTENNA_159 (.A(_09068_));
 sg13g2_antennanp ANTENNA_160 (.A(_09123_));
 sg13g2_antennanp ANTENNA_161 (.A(_09223_));
 sg13g2_antennanp ANTENNA_162 (.A(_09223_));
 sg13g2_antennanp ANTENNA_163 (.A(_09223_));
 sg13g2_antennanp ANTENNA_164 (.A(_09223_));
 sg13g2_antennanp ANTENNA_165 (.A(_09225_));
 sg13g2_antennanp ANTENNA_166 (.A(_09225_));
 sg13g2_antennanp ANTENNA_167 (.A(_09225_));
 sg13g2_antennanp ANTENNA_168 (.A(_09225_));
 sg13g2_antennanp ANTENNA_169 (.A(_09227_));
 sg13g2_antennanp ANTENNA_170 (.A(_09227_));
 sg13g2_antennanp ANTENNA_171 (.A(_09227_));
 sg13g2_antennanp ANTENNA_172 (.A(_09227_));
 sg13g2_antennanp ANTENNA_173 (.A(_09240_));
 sg13g2_antennanp ANTENNA_174 (.A(_09240_));
 sg13g2_antennanp ANTENNA_175 (.A(_09240_));
 sg13g2_antennanp ANTENNA_176 (.A(_09240_));
 sg13g2_antennanp ANTENNA_177 (.A(_09240_));
 sg13g2_antennanp ANTENNA_178 (.A(_09240_));
 sg13g2_antennanp ANTENNA_179 (.A(_09282_));
 sg13g2_antennanp ANTENNA_180 (.A(_09282_));
 sg13g2_antennanp ANTENNA_181 (.A(_09282_));
 sg13g2_antennanp ANTENNA_182 (.A(_09282_));
 sg13g2_antennanp ANTENNA_183 (.A(_09284_));
 sg13g2_antennanp ANTENNA_184 (.A(_09284_));
 sg13g2_antennanp ANTENNA_185 (.A(_09284_));
 sg13g2_antennanp ANTENNA_186 (.A(_09284_));
 sg13g2_antennanp ANTENNA_187 (.A(_09310_));
 sg13g2_antennanp ANTENNA_188 (.A(_09310_));
 sg13g2_antennanp ANTENNA_189 (.A(_09310_));
 sg13g2_antennanp ANTENNA_190 (.A(_09363_));
 sg13g2_antennanp ANTENNA_191 (.A(_09363_));
 sg13g2_antennanp ANTENNA_192 (.A(_09363_));
 sg13g2_antennanp ANTENNA_193 (.A(_09363_));
 sg13g2_antennanp ANTENNA_194 (.A(_09365_));
 sg13g2_antennanp ANTENNA_195 (.A(_09365_));
 sg13g2_antennanp ANTENNA_196 (.A(_09365_));
 sg13g2_antennanp ANTENNA_197 (.A(_09365_));
 sg13g2_antennanp ANTENNA_198 (.A(_09435_));
 sg13g2_antennanp ANTENNA_199 (.A(_09435_));
 sg13g2_antennanp ANTENNA_200 (.A(_09435_));
 sg13g2_antennanp ANTENNA_201 (.A(_09463_));
 sg13g2_antennanp ANTENNA_202 (.A(_09463_));
 sg13g2_antennanp ANTENNA_203 (.A(_09463_));
 sg13g2_antennanp ANTENNA_204 (.A(_09463_));
 sg13g2_antennanp ANTENNA_205 (.A(_09463_));
 sg13g2_antennanp ANTENNA_206 (.A(_09463_));
 sg13g2_antennanp ANTENNA_207 (.A(_09463_));
 sg13g2_antennanp ANTENNA_208 (.A(_09463_));
 sg13g2_antennanp ANTENNA_209 (.A(_09463_));
 sg13g2_antennanp ANTENNA_210 (.A(_09463_));
 sg13g2_antennanp ANTENNA_211 (.A(_09463_));
 sg13g2_antennanp ANTENNA_212 (.A(_09463_));
 sg13g2_antennanp ANTENNA_213 (.A(_09463_));
 sg13g2_antennanp ANTENNA_214 (.A(_09463_));
 sg13g2_antennanp ANTENNA_215 (.A(_09463_));
 sg13g2_antennanp ANTENNA_216 (.A(_09512_));
 sg13g2_antennanp ANTENNA_217 (.A(_09512_));
 sg13g2_antennanp ANTENNA_218 (.A(_09558_));
 sg13g2_antennanp ANTENNA_219 (.A(_09558_));
 sg13g2_antennanp ANTENNA_220 (.A(_09558_));
 sg13g2_antennanp ANTENNA_221 (.A(_09558_));
 sg13g2_antennanp ANTENNA_222 (.A(_09573_));
 sg13g2_antennanp ANTENNA_223 (.A(_09588_));
 sg13g2_antennanp ANTENNA_224 (.A(_09639_));
 sg13g2_antennanp ANTENNA_225 (.A(_09700_));
 sg13g2_antennanp ANTENNA_226 (.A(_09854_));
 sg13g2_antennanp ANTENNA_227 (.A(_09897_));
 sg13g2_antennanp ANTENNA_228 (.A(_09899_));
 sg13g2_antennanp ANTENNA_229 (.A(_10089_));
 sg13g2_antennanp ANTENNA_230 (.A(_10089_));
 sg13g2_antennanp ANTENNA_231 (.A(_10089_));
 sg13g2_antennanp ANTENNA_232 (.A(_10089_));
 sg13g2_antennanp ANTENNA_233 (.A(_10089_));
 sg13g2_antennanp ANTENNA_234 (.A(_10089_));
 sg13g2_antennanp ANTENNA_235 (.A(_10116_));
 sg13g2_antennanp ANTENNA_236 (.A(_10116_));
 sg13g2_antennanp ANTENNA_237 (.A(_10116_));
 sg13g2_antennanp ANTENNA_238 (.A(_10116_));
 sg13g2_antennanp ANTENNA_239 (.A(_10116_));
 sg13g2_antennanp ANTENNA_240 (.A(_10116_));
 sg13g2_antennanp ANTENNA_241 (.A(_10116_));
 sg13g2_antennanp ANTENNA_242 (.A(_10116_));
 sg13g2_antennanp ANTENNA_243 (.A(_10137_));
 sg13g2_antennanp ANTENNA_244 (.A(_10137_));
 sg13g2_antennanp ANTENNA_245 (.A(_10137_));
 sg13g2_antennanp ANTENNA_246 (.A(_10137_));
 sg13g2_antennanp ANTENNA_247 (.A(_10137_));
 sg13g2_antennanp ANTENNA_248 (.A(_10137_));
 sg13g2_antennanp ANTENNA_249 (.A(_10137_));
 sg13g2_antennanp ANTENNA_250 (.A(_10137_));
 sg13g2_antennanp ANTENNA_251 (.A(_10137_));
 sg13g2_antennanp ANTENNA_252 (.A(_10137_));
 sg13g2_antennanp ANTENNA_253 (.A(_10204_));
 sg13g2_antennanp ANTENNA_254 (.A(_10204_));
 sg13g2_antennanp ANTENNA_255 (.A(_10204_));
 sg13g2_antennanp ANTENNA_256 (.A(_10204_));
 sg13g2_antennanp ANTENNA_257 (.A(_10210_));
 sg13g2_antennanp ANTENNA_258 (.A(_10210_));
 sg13g2_antennanp ANTENNA_259 (.A(_10210_));
 sg13g2_antennanp ANTENNA_260 (.A(_10210_));
 sg13g2_antennanp ANTENNA_261 (.A(_10210_));
 sg13g2_antennanp ANTENNA_262 (.A(_10210_));
 sg13g2_antennanp ANTENNA_263 (.A(_10210_));
 sg13g2_antennanp ANTENNA_264 (.A(_10210_));
 sg13g2_antennanp ANTENNA_265 (.A(_10210_));
 sg13g2_antennanp ANTENNA_266 (.A(_10210_));
 sg13g2_antennanp ANTENNA_267 (.A(_10210_));
 sg13g2_antennanp ANTENNA_268 (.A(_10210_));
 sg13g2_antennanp ANTENNA_269 (.A(_10383_));
 sg13g2_antennanp ANTENNA_270 (.A(_10383_));
 sg13g2_antennanp ANTENNA_271 (.A(_10383_));
 sg13g2_antennanp ANTENNA_272 (.A(_10383_));
 sg13g2_antennanp ANTENNA_273 (.A(_10721_));
 sg13g2_antennanp ANTENNA_274 (.A(_10721_));
 sg13g2_antennanp ANTENNA_275 (.A(_10721_));
 sg13g2_antennanp ANTENNA_276 (.A(_10721_));
 sg13g2_antennanp ANTENNA_277 (.A(_10721_));
 sg13g2_antennanp ANTENNA_278 (.A(_10819_));
 sg13g2_antennanp ANTENNA_279 (.A(_10819_));
 sg13g2_antennanp ANTENNA_280 (.A(_10819_));
 sg13g2_antennanp ANTENNA_281 (.A(_10819_));
 sg13g2_antennanp ANTENNA_282 (.A(_10819_));
 sg13g2_antennanp ANTENNA_283 (.A(_10819_));
 sg13g2_antennanp ANTENNA_284 (.A(_10819_));
 sg13g2_antennanp ANTENNA_285 (.A(_10819_));
 sg13g2_antennanp ANTENNA_286 (.A(_10819_));
 sg13g2_antennanp ANTENNA_287 (.A(_12000_));
 sg13g2_antennanp ANTENNA_288 (.A(_12000_));
 sg13g2_antennanp ANTENNA_289 (.A(_12000_));
 sg13g2_antennanp ANTENNA_290 (.A(_12000_));
 sg13g2_antennanp ANTENNA_291 (.A(_12010_));
 sg13g2_antennanp ANTENNA_292 (.A(_12010_));
 sg13g2_antennanp ANTENNA_293 (.A(_12010_));
 sg13g2_antennanp ANTENNA_294 (.A(_12010_));
 sg13g2_antennanp ANTENNA_295 (.A(_12010_));
 sg13g2_antennanp ANTENNA_296 (.A(_12010_));
 sg13g2_antennanp ANTENNA_297 (.A(_12010_));
 sg13g2_antennanp ANTENNA_298 (.A(_12010_));
 sg13g2_antennanp ANTENNA_299 (.A(_12010_));
 sg13g2_antennanp ANTENNA_300 (.A(_12010_));
 sg13g2_antennanp ANTENNA_301 (.A(_12010_));
 sg13g2_antennanp ANTENNA_302 (.A(_12010_));
 sg13g2_antennanp ANTENNA_303 (.A(_12010_));
 sg13g2_antennanp ANTENNA_304 (.A(_12010_));
 sg13g2_antennanp ANTENNA_305 (.A(_12052_));
 sg13g2_antennanp ANTENNA_306 (.A(_12052_));
 sg13g2_antennanp ANTENNA_307 (.A(_12052_));
 sg13g2_antennanp ANTENNA_308 (.A(_12052_));
 sg13g2_antennanp ANTENNA_309 (.A(_12052_));
 sg13g2_antennanp ANTENNA_310 (.A(_12052_));
 sg13g2_antennanp ANTENNA_311 (.A(_12052_));
 sg13g2_antennanp ANTENNA_312 (.A(_12052_));
 sg13g2_antennanp ANTENNA_313 (.A(_12052_));
 sg13g2_antennanp ANTENNA_314 (.A(_12087_));
 sg13g2_antennanp ANTENNA_315 (.A(_12087_));
 sg13g2_antennanp ANTENNA_316 (.A(_12087_));
 sg13g2_antennanp ANTENNA_317 (.A(_12087_));
 sg13g2_antennanp ANTENNA_318 (.A(_12087_));
 sg13g2_antennanp ANTENNA_319 (.A(_12087_));
 sg13g2_antennanp ANTENNA_320 (.A(_12087_));
 sg13g2_antennanp ANTENNA_321 (.A(_12087_));
 sg13g2_antennanp ANTENNA_322 (.A(_12087_));
 sg13g2_antennanp ANTENNA_323 (.A(_12119_));
 sg13g2_antennanp ANTENNA_324 (.A(_12119_));
 sg13g2_antennanp ANTENNA_325 (.A(_12119_));
 sg13g2_antennanp ANTENNA_326 (.A(_12119_));
 sg13g2_antennanp ANTENNA_327 (.A(_12119_));
 sg13g2_antennanp ANTENNA_328 (.A(_12119_));
 sg13g2_antennanp ANTENNA_329 (.A(_12119_));
 sg13g2_antennanp ANTENNA_330 (.A(_12119_));
 sg13g2_antennanp ANTENNA_331 (.A(_12119_));
 sg13g2_antennanp ANTENNA_332 (.A(_12119_));
 sg13g2_antennanp ANTENNA_333 (.A(_12201_));
 sg13g2_antennanp ANTENNA_334 (.A(_12201_));
 sg13g2_antennanp ANTENNA_335 (.A(_12201_));
 sg13g2_antennanp ANTENNA_336 (.A(_12209_));
 sg13g2_antennanp ANTENNA_337 (.A(_12209_));
 sg13g2_antennanp ANTENNA_338 (.A(_12209_));
 sg13g2_antennanp ANTENNA_339 (.A(_12209_));
 sg13g2_antennanp ANTENNA_340 (.A(_12209_));
 sg13g2_antennanp ANTENNA_341 (.A(_12209_));
 sg13g2_antennanp ANTENNA_342 (.A(_12216_));
 sg13g2_antennanp ANTENNA_343 (.A(_12216_));
 sg13g2_antennanp ANTENNA_344 (.A(_12216_));
 sg13g2_antennanp ANTENNA_345 (.A(_12216_));
 sg13g2_antennanp ANTENNA_346 (.A(_12216_));
 sg13g2_antennanp ANTENNA_347 (.A(_12216_));
 sg13g2_antennanp ANTENNA_348 (.A(_12220_));
 sg13g2_antennanp ANTENNA_349 (.A(_12220_));
 sg13g2_antennanp ANTENNA_350 (.A(_12220_));
 sg13g2_antennanp ANTENNA_351 (.A(_12220_));
 sg13g2_antennanp ANTENNA_352 (.A(_12220_));
 sg13g2_antennanp ANTENNA_353 (.A(_12220_));
 sg13g2_antennanp ANTENNA_354 (.A(_12220_));
 sg13g2_antennanp ANTENNA_355 (.A(_12220_));
 sg13g2_antennanp ANTENNA_356 (.A(_12220_));
 sg13g2_antennanp ANTENNA_357 (.A(_12227_));
 sg13g2_antennanp ANTENNA_358 (.A(_12227_));
 sg13g2_antennanp ANTENNA_359 (.A(_12227_));
 sg13g2_antennanp ANTENNA_360 (.A(_12227_));
 sg13g2_antennanp ANTENNA_361 (.A(_12227_));
 sg13g2_antennanp ANTENNA_362 (.A(_12227_));
 sg13g2_antennanp ANTENNA_363 (.A(_12227_));
 sg13g2_antennanp ANTENNA_364 (.A(_12227_));
 sg13g2_antennanp ANTENNA_365 (.A(_12227_));
 sg13g2_antennanp ANTENNA_366 (.A(_12250_));
 sg13g2_antennanp ANTENNA_367 (.A(_12250_));
 sg13g2_antennanp ANTENNA_368 (.A(_12250_));
 sg13g2_antennanp ANTENNA_369 (.A(_12255_));
 sg13g2_antennanp ANTENNA_370 (.A(_12255_));
 sg13g2_antennanp ANTENNA_371 (.A(_12255_));
 sg13g2_antennanp ANTENNA_372 (.A(clk));
 sg13g2_antennanp ANTENNA_373 (.A(clk));
 sg13g2_antennanp ANTENNA_374 (.A(\cpu.d_flush_all ));
 sg13g2_antennanp ANTENNA_375 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_376 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_377 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_378 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_379 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_380 (.A(net1));
 sg13g2_antennanp ANTENNA_381 (.A(net1));
 sg13g2_antennanp ANTENNA_382 (.A(net1));
 sg13g2_antennanp ANTENNA_383 (.A(net1));
 sg13g2_antennanp ANTENNA_384 (.A(net1));
 sg13g2_antennanp ANTENNA_385 (.A(net1));
 sg13g2_antennanp ANTENNA_386 (.A(net1));
 sg13g2_antennanp ANTENNA_387 (.A(net1));
 sg13g2_antennanp ANTENNA_388 (.A(net3));
 sg13g2_antennanp ANTENNA_389 (.A(net3));
 sg13g2_antennanp ANTENNA_390 (.A(net12));
 sg13g2_antennanp ANTENNA_391 (.A(net12));
 sg13g2_antennanp ANTENNA_392 (.A(net13));
 sg13g2_antennanp ANTENNA_393 (.A(net13));
 sg13g2_antennanp ANTENNA_394 (.A(net14));
 sg13g2_antennanp ANTENNA_395 (.A(net14));
 sg13g2_antennanp ANTENNA_396 (.A(net517));
 sg13g2_antennanp ANTENNA_397 (.A(net517));
 sg13g2_antennanp ANTENNA_398 (.A(net517));
 sg13g2_antennanp ANTENNA_399 (.A(net517));
 sg13g2_antennanp ANTENNA_400 (.A(net517));
 sg13g2_antennanp ANTENNA_401 (.A(net517));
 sg13g2_antennanp ANTENNA_402 (.A(net517));
 sg13g2_antennanp ANTENNA_403 (.A(net517));
 sg13g2_antennanp ANTENNA_404 (.A(net517));
 sg13g2_antennanp ANTENNA_405 (.A(net517));
 sg13g2_antennanp ANTENNA_406 (.A(net517));
 sg13g2_antennanp ANTENNA_407 (.A(net517));
 sg13g2_antennanp ANTENNA_408 (.A(net520));
 sg13g2_antennanp ANTENNA_409 (.A(net520));
 sg13g2_antennanp ANTENNA_410 (.A(net520));
 sg13g2_antennanp ANTENNA_411 (.A(net520));
 sg13g2_antennanp ANTENNA_412 (.A(net520));
 sg13g2_antennanp ANTENNA_413 (.A(net520));
 sg13g2_antennanp ANTENNA_414 (.A(net520));
 sg13g2_antennanp ANTENNA_415 (.A(net520));
 sg13g2_antennanp ANTENNA_416 (.A(net544));
 sg13g2_antennanp ANTENNA_417 (.A(net544));
 sg13g2_antennanp ANTENNA_418 (.A(net544));
 sg13g2_antennanp ANTENNA_419 (.A(net544));
 sg13g2_antennanp ANTENNA_420 (.A(net544));
 sg13g2_antennanp ANTENNA_421 (.A(net544));
 sg13g2_antennanp ANTENNA_422 (.A(net544));
 sg13g2_antennanp ANTENNA_423 (.A(net544));
 sg13g2_antennanp ANTENNA_424 (.A(net544));
 sg13g2_antennanp ANTENNA_425 (.A(net544));
 sg13g2_antennanp ANTENNA_426 (.A(net544));
 sg13g2_antennanp ANTENNA_427 (.A(net544));
 sg13g2_antennanp ANTENNA_428 (.A(net544));
 sg13g2_antennanp ANTENNA_429 (.A(net544));
 sg13g2_antennanp ANTENNA_430 (.A(net653));
 sg13g2_antennanp ANTENNA_431 (.A(net653));
 sg13g2_antennanp ANTENNA_432 (.A(net653));
 sg13g2_antennanp ANTENNA_433 (.A(net653));
 sg13g2_antennanp ANTENNA_434 (.A(net653));
 sg13g2_antennanp ANTENNA_435 (.A(net653));
 sg13g2_antennanp ANTENNA_436 (.A(net653));
 sg13g2_antennanp ANTENNA_437 (.A(net653));
 sg13g2_antennanp ANTENNA_438 (.A(net653));
 sg13g2_antennanp ANTENNA_439 (.A(net728));
 sg13g2_antennanp ANTENNA_440 (.A(net728));
 sg13g2_antennanp ANTENNA_441 (.A(net728));
 sg13g2_antennanp ANTENNA_442 (.A(net728));
 sg13g2_antennanp ANTENNA_443 (.A(net728));
 sg13g2_antennanp ANTENNA_444 (.A(net728));
 sg13g2_antennanp ANTENNA_445 (.A(net728));
 sg13g2_antennanp ANTENNA_446 (.A(net728));
 sg13g2_antennanp ANTENNA_447 (.A(net795));
 sg13g2_antennanp ANTENNA_448 (.A(net795));
 sg13g2_antennanp ANTENNA_449 (.A(net795));
 sg13g2_antennanp ANTENNA_450 (.A(net795));
 sg13g2_antennanp ANTENNA_451 (.A(net795));
 sg13g2_antennanp ANTENNA_452 (.A(net795));
 sg13g2_antennanp ANTENNA_453 (.A(net795));
 sg13g2_antennanp ANTENNA_454 (.A(net795));
 sg13g2_antennanp ANTENNA_455 (.A(net795));
 sg13g2_antennanp ANTENNA_456 (.A(net795));
 sg13g2_antennanp ANTENNA_457 (.A(net795));
 sg13g2_antennanp ANTENNA_458 (.A(net795));
 sg13g2_antennanp ANTENNA_459 (.A(net795));
 sg13g2_antennanp ANTENNA_460 (.A(net795));
 sg13g2_antennanp ANTENNA_461 (.A(net795));
 sg13g2_antennanp ANTENNA_462 (.A(net795));
 sg13g2_antennanp ANTENNA_463 (.A(net797));
 sg13g2_antennanp ANTENNA_464 (.A(net797));
 sg13g2_antennanp ANTENNA_465 (.A(net797));
 sg13g2_antennanp ANTENNA_466 (.A(net797));
 sg13g2_antennanp ANTENNA_467 (.A(net797));
 sg13g2_antennanp ANTENNA_468 (.A(net797));
 sg13g2_antennanp ANTENNA_469 (.A(net797));
 sg13g2_antennanp ANTENNA_470 (.A(net797));
 sg13g2_antennanp ANTENNA_471 (.A(net797));
 sg13g2_antennanp ANTENNA_472 (.A(net797));
 sg13g2_antennanp ANTENNA_473 (.A(net797));
 sg13g2_antennanp ANTENNA_474 (.A(net797));
 sg13g2_antennanp ANTENNA_475 (.A(net797));
 sg13g2_antennanp ANTENNA_476 (.A(net797));
 sg13g2_antennanp ANTENNA_477 (.A(net797));
 sg13g2_antennanp ANTENNA_478 (.A(net797));
 sg13g2_antennanp ANTENNA_479 (.A(net797));
 sg13g2_antennanp ANTENNA_480 (.A(net797));
 sg13g2_antennanp ANTENNA_481 (.A(net809));
 sg13g2_antennanp ANTENNA_482 (.A(net809));
 sg13g2_antennanp ANTENNA_483 (.A(net809));
 sg13g2_antennanp ANTENNA_484 (.A(net809));
 sg13g2_antennanp ANTENNA_485 (.A(net809));
 sg13g2_antennanp ANTENNA_486 (.A(net809));
 sg13g2_antennanp ANTENNA_487 (.A(net809));
 sg13g2_antennanp ANTENNA_488 (.A(net809));
 sg13g2_antennanp ANTENNA_489 (.A(net809));
 sg13g2_antennanp ANTENNA_490 (.A(net809));
 sg13g2_antennanp ANTENNA_491 (.A(net809));
 sg13g2_antennanp ANTENNA_492 (.A(net809));
 sg13g2_antennanp ANTENNA_493 (.A(net809));
 sg13g2_antennanp ANTENNA_494 (.A(net809));
 sg13g2_antennanp ANTENNA_495 (.A(net809));
 sg13g2_antennanp ANTENNA_496 (.A(net810));
 sg13g2_antennanp ANTENNA_497 (.A(net810));
 sg13g2_antennanp ANTENNA_498 (.A(net810));
 sg13g2_antennanp ANTENNA_499 (.A(net810));
 sg13g2_antennanp ANTENNA_500 (.A(net810));
 sg13g2_antennanp ANTENNA_501 (.A(net810));
 sg13g2_antennanp ANTENNA_502 (.A(net810));
 sg13g2_antennanp ANTENNA_503 (.A(net810));
 sg13g2_antennanp ANTENNA_504 (.A(net810));
 sg13g2_antennanp ANTENNA_505 (.A(net810));
 sg13g2_antennanp ANTENNA_506 (.A(net810));
 sg13g2_antennanp ANTENNA_507 (.A(net810));
 sg13g2_antennanp ANTENNA_508 (.A(net810));
 sg13g2_antennanp ANTENNA_509 (.A(net810));
 sg13g2_antennanp ANTENNA_510 (.A(net810));
 sg13g2_antennanp ANTENNA_511 (.A(net810));
 sg13g2_antennanp ANTENNA_512 (.A(net812));
 sg13g2_antennanp ANTENNA_513 (.A(net812));
 sg13g2_antennanp ANTENNA_514 (.A(net812));
 sg13g2_antennanp ANTENNA_515 (.A(net812));
 sg13g2_antennanp ANTENNA_516 (.A(net812));
 sg13g2_antennanp ANTENNA_517 (.A(net812));
 sg13g2_antennanp ANTENNA_518 (.A(net812));
 sg13g2_antennanp ANTENNA_519 (.A(net812));
 sg13g2_antennanp ANTENNA_520 (.A(net812));
 sg13g2_antennanp ANTENNA_521 (.A(net812));
 sg13g2_antennanp ANTENNA_522 (.A(net812));
 sg13g2_antennanp ANTENNA_523 (.A(net812));
 sg13g2_antennanp ANTENNA_524 (.A(net812));
 sg13g2_antennanp ANTENNA_525 (.A(net812));
 sg13g2_antennanp ANTENNA_526 (.A(net812));
 sg13g2_antennanp ANTENNA_527 (.A(net812));
 sg13g2_antennanp ANTENNA_528 (.A(net812));
 sg13g2_antennanp ANTENNA_529 (.A(net812));
 sg13g2_antennanp ANTENNA_530 (.A(net812));
 sg13g2_antennanp ANTENNA_531 (.A(net812));
 sg13g2_antennanp ANTENNA_532 (.A(net812));
 sg13g2_antennanp ANTENNA_533 (.A(net812));
 sg13g2_antennanp ANTENNA_534 (.A(net812));
 sg13g2_antennanp ANTENNA_535 (.A(net861));
 sg13g2_antennanp ANTENNA_536 (.A(net861));
 sg13g2_antennanp ANTENNA_537 (.A(net861));
 sg13g2_antennanp ANTENNA_538 (.A(net861));
 sg13g2_antennanp ANTENNA_539 (.A(net861));
 sg13g2_antennanp ANTENNA_540 (.A(net861));
 sg13g2_antennanp ANTENNA_541 (.A(net861));
 sg13g2_antennanp ANTENNA_542 (.A(net861));
 sg13g2_antennanp ANTENNA_543 (.A(net861));
 sg13g2_antennanp ANTENNA_544 (.A(net861));
 sg13g2_antennanp ANTENNA_545 (.A(net861));
 sg13g2_antennanp ANTENNA_546 (.A(net861));
 sg13g2_antennanp ANTENNA_547 (.A(net861));
 sg13g2_antennanp ANTENNA_548 (.A(net861));
 sg13g2_antennanp ANTENNA_549 (.A(net861));
 sg13g2_antennanp ANTENNA_550 (.A(net861));
 sg13g2_antennanp ANTENNA_551 (.A(net862));
 sg13g2_antennanp ANTENNA_552 (.A(net862));
 sg13g2_antennanp ANTENNA_553 (.A(net862));
 sg13g2_antennanp ANTENNA_554 (.A(net862));
 sg13g2_antennanp ANTENNA_555 (.A(net862));
 sg13g2_antennanp ANTENNA_556 (.A(net862));
 sg13g2_antennanp ANTENNA_557 (.A(net862));
 sg13g2_antennanp ANTENNA_558 (.A(net862));
 sg13g2_antennanp ANTENNA_559 (.A(net862));
 sg13g2_antennanp ANTENNA_560 (.A(net862));
 sg13g2_antennanp ANTENNA_561 (.A(net862));
 sg13g2_antennanp ANTENNA_562 (.A(net862));
 sg13g2_antennanp ANTENNA_563 (.A(net862));
 sg13g2_antennanp ANTENNA_564 (.A(net862));
 sg13g2_antennanp ANTENNA_565 (.A(net901));
 sg13g2_antennanp ANTENNA_566 (.A(net901));
 sg13g2_antennanp ANTENNA_567 (.A(net901));
 sg13g2_antennanp ANTENNA_568 (.A(net901));
 sg13g2_antennanp ANTENNA_569 (.A(net901));
 sg13g2_antennanp ANTENNA_570 (.A(net901));
 sg13g2_antennanp ANTENNA_571 (.A(net901));
 sg13g2_antennanp ANTENNA_572 (.A(net901));
 sg13g2_antennanp ANTENNA_573 (.A(net907));
 sg13g2_antennanp ANTENNA_574 (.A(net907));
 sg13g2_antennanp ANTENNA_575 (.A(net907));
 sg13g2_antennanp ANTENNA_576 (.A(net907));
 sg13g2_antennanp ANTENNA_577 (.A(net907));
 sg13g2_antennanp ANTENNA_578 (.A(net907));
 sg13g2_antennanp ANTENNA_579 (.A(net907));
 sg13g2_antennanp ANTENNA_580 (.A(net907));
 sg13g2_antennanp ANTENNA_581 (.A(net907));
 sg13g2_antennanp ANTENNA_582 (.A(net907));
 sg13g2_antennanp ANTENNA_583 (.A(net907));
 sg13g2_antennanp ANTENNA_584 (.A(net907));
 sg13g2_antennanp ANTENNA_585 (.A(net907));
 sg13g2_antennanp ANTENNA_586 (.A(net907));
 sg13g2_antennanp ANTENNA_587 (.A(net916));
 sg13g2_antennanp ANTENNA_588 (.A(net916));
 sg13g2_antennanp ANTENNA_589 (.A(net916));
 sg13g2_antennanp ANTENNA_590 (.A(net916));
 sg13g2_antennanp ANTENNA_591 (.A(net916));
 sg13g2_antennanp ANTENNA_592 (.A(net916));
 sg13g2_antennanp ANTENNA_593 (.A(net916));
 sg13g2_antennanp ANTENNA_594 (.A(net916));
 sg13g2_antennanp ANTENNA_595 (.A(net916));
 sg13g2_antennanp ANTENNA_596 (.A(net916));
 sg13g2_antennanp ANTENNA_597 (.A(net916));
 sg13g2_antennanp ANTENNA_598 (.A(net916));
 sg13g2_antennanp ANTENNA_599 (.A(net916));
 sg13g2_antennanp ANTENNA_600 (.A(net916));
 sg13g2_antennanp ANTENNA_601 (.A(net916));
 sg13g2_antennanp ANTENNA_602 (.A(net916));
 sg13g2_antennanp ANTENNA_603 (.A(net917));
 sg13g2_antennanp ANTENNA_604 (.A(net917));
 sg13g2_antennanp ANTENNA_605 (.A(net917));
 sg13g2_antennanp ANTENNA_606 (.A(net917));
 sg13g2_antennanp ANTENNA_607 (.A(net917));
 sg13g2_antennanp ANTENNA_608 (.A(net917));
 sg13g2_antennanp ANTENNA_609 (.A(net917));
 sg13g2_antennanp ANTENNA_610 (.A(net917));
 sg13g2_antennanp ANTENNA_611 (.A(net917));
 sg13g2_antennanp ANTENNA_612 (.A(net917));
 sg13g2_antennanp ANTENNA_613 (.A(net917));
 sg13g2_antennanp ANTENNA_614 (.A(net917));
 sg13g2_antennanp ANTENNA_615 (.A(net917));
 sg13g2_antennanp ANTENNA_616 (.A(net917));
 sg13g2_antennanp ANTENNA_617 (.A(net917));
 sg13g2_antennanp ANTENNA_618 (.A(net917));
 sg13g2_antennanp ANTENNA_619 (.A(net917));
 sg13g2_antennanp ANTENNA_620 (.A(net917));
 sg13g2_antennanp ANTENNA_621 (.A(net917));
 sg13g2_antennanp ANTENNA_622 (.A(net917));
 sg13g2_antennanp ANTENNA_623 (.A(net917));
 sg13g2_antennanp ANTENNA_624 (.A(net917));
 sg13g2_antennanp ANTENNA_625 (.A(net917));
 sg13g2_antennanp ANTENNA_626 (.A(net917));
 sg13g2_antennanp ANTENNA_627 (.A(net917));
 sg13g2_antennanp ANTENNA_628 (.A(net917));
 sg13g2_antennanp ANTENNA_629 (.A(net917));
 sg13g2_antennanp ANTENNA_630 (.A(net917));
 sg13g2_antennanp ANTENNA_631 (.A(net917));
 sg13g2_antennanp ANTENNA_632 (.A(net917));
 sg13g2_antennanp ANTENNA_633 (.A(net917));
 sg13g2_antennanp ANTENNA_634 (.A(net917));
 sg13g2_antennanp ANTENNA_635 (.A(net917));
 sg13g2_antennanp ANTENNA_636 (.A(net917));
 sg13g2_antennanp ANTENNA_637 (.A(net993));
 sg13g2_antennanp ANTENNA_638 (.A(net993));
 sg13g2_antennanp ANTENNA_639 (.A(net993));
 sg13g2_antennanp ANTENNA_640 (.A(net993));
 sg13g2_antennanp ANTENNA_641 (.A(net993));
 sg13g2_antennanp ANTENNA_642 (.A(net993));
 sg13g2_antennanp ANTENNA_643 (.A(net993));
 sg13g2_antennanp ANTENNA_644 (.A(net993));
 sg13g2_antennanp ANTENNA_645 (.A(net993));
 sg13g2_antennanp ANTENNA_646 (.A(net993));
 sg13g2_antennanp ANTENNA_647 (.A(net993));
 sg13g2_antennanp ANTENNA_648 (.A(net993));
 sg13g2_antennanp ANTENNA_649 (.A(net993));
 sg13g2_antennanp ANTENNA_650 (.A(net993));
 sg13g2_antennanp ANTENNA_651 (.A(net993));
 sg13g2_antennanp ANTENNA_652 (.A(net993));
 sg13g2_antennanp ANTENNA_653 (.A(net1020));
 sg13g2_antennanp ANTENNA_654 (.A(net1020));
 sg13g2_antennanp ANTENNA_655 (.A(net1020));
 sg13g2_antennanp ANTENNA_656 (.A(net1020));
 sg13g2_antennanp ANTENNA_657 (.A(net1020));
 sg13g2_antennanp ANTENNA_658 (.A(net1020));
 sg13g2_antennanp ANTENNA_659 (.A(net1020));
 sg13g2_antennanp ANTENNA_660 (.A(net1020));
 sg13g2_antennanp ANTENNA_661 (.A(net1020));
 sg13g2_antennanp ANTENNA_662 (.A(net1020));
 sg13g2_antennanp ANTENNA_663 (.A(net1020));
 sg13g2_antennanp ANTENNA_664 (.A(net1020));
 sg13g2_antennanp ANTENNA_665 (.A(net1020));
 sg13g2_antennanp ANTENNA_666 (.A(net1020));
 sg13g2_antennanp ANTENNA_667 (.A(net1020));
 sg13g2_antennanp ANTENNA_668 (.A(net1020));
 sg13g2_antennanp ANTENNA_669 (.A(net1020));
 sg13g2_antennanp ANTENNA_670 (.A(net1020));
 sg13g2_antennanp ANTENNA_671 (.A(net1020));
 sg13g2_antennanp ANTENNA_672 (.A(net1020));
 sg13g2_antennanp ANTENNA_673 (.A(net1020));
 sg13g2_antennanp ANTENNA_674 (.A(net1020));
 sg13g2_antennanp ANTENNA_675 (.A(net1020));
 sg13g2_antennanp ANTENNA_676 (.A(net1020));
 sg13g2_antennanp ANTENNA_677 (.A(net1020));
 sg13g2_antennanp ANTENNA_678 (.A(net1020));
 sg13g2_antennanp ANTENNA_679 (.A(net1020));
 sg13g2_antennanp ANTENNA_680 (.A(net1020));
 sg13g2_antennanp ANTENNA_681 (.A(net1020));
 sg13g2_antennanp ANTENNA_682 (.A(net1020));
 sg13g2_antennanp ANTENNA_683 (.A(net1020));
 sg13g2_antennanp ANTENNA_684 (.A(net1020));
 sg13g2_antennanp ANTENNA_685 (.A(net1020));
 sg13g2_antennanp ANTENNA_686 (.A(net1020));
 sg13g2_antennanp ANTENNA_687 (.A(net1021));
 sg13g2_antennanp ANTENNA_688 (.A(net1021));
 sg13g2_antennanp ANTENNA_689 (.A(net1021));
 sg13g2_antennanp ANTENNA_690 (.A(net1021));
 sg13g2_antennanp ANTENNA_691 (.A(net1021));
 sg13g2_antennanp ANTENNA_692 (.A(net1021));
 sg13g2_antennanp ANTENNA_693 (.A(net1021));
 sg13g2_antennanp ANTENNA_694 (.A(net1021));
 sg13g2_antennanp ANTENNA_695 (.A(net1021));
 sg13g2_antennanp ANTENNA_696 (.A(net1021));
 sg13g2_antennanp ANTENNA_697 (.A(net1021));
 sg13g2_antennanp ANTENNA_698 (.A(net1021));
 sg13g2_antennanp ANTENNA_699 (.A(net1021));
 sg13g2_antennanp ANTENNA_700 (.A(net1021));
 sg13g2_antennanp ANTENNA_701 (.A(net1071));
 sg13g2_antennanp ANTENNA_702 (.A(net1071));
 sg13g2_antennanp ANTENNA_703 (.A(net1071));
 sg13g2_antennanp ANTENNA_704 (.A(net1071));
 sg13g2_antennanp ANTENNA_705 (.A(net1071));
 sg13g2_antennanp ANTENNA_706 (.A(net1071));
 sg13g2_antennanp ANTENNA_707 (.A(net1071));
 sg13g2_antennanp ANTENNA_708 (.A(net1071));
 sg13g2_antennanp ANTENNA_709 (.A(net1071));
 sg13g2_antennanp ANTENNA_710 (.A(net1108));
 sg13g2_antennanp ANTENNA_711 (.A(net1108));
 sg13g2_antennanp ANTENNA_712 (.A(net1108));
 sg13g2_antennanp ANTENNA_713 (.A(net1108));
 sg13g2_antennanp ANTENNA_714 (.A(net1108));
 sg13g2_antennanp ANTENNA_715 (.A(net1108));
 sg13g2_antennanp ANTENNA_716 (.A(net1108));
 sg13g2_antennanp ANTENNA_717 (.A(net1108));
 sg13g2_antennanp ANTENNA_718 (.A(net1108));
 sg13g2_antennanp ANTENNA_719 (.A(net1108));
 sg13g2_antennanp ANTENNA_720 (.A(net1108));
 sg13g2_antennanp ANTENNA_721 (.A(net1108));
 sg13g2_antennanp ANTENNA_722 (.A(net1108));
 sg13g2_antennanp ANTENNA_723 (.A(net1108));
 sg13g2_antennanp ANTENNA_724 (.A(net1108));
 sg13g2_antennanp ANTENNA_725 (.A(net1108));
 sg13g2_antennanp ANTENNA_726 (.A(net1108));
 sg13g2_antennanp ANTENNA_727 (.A(net1108));
 sg13g2_antennanp ANTENNA_728 (.A(net1108));
 sg13g2_antennanp ANTENNA_729 (.A(net1108));
 sg13g2_antennanp ANTENNA_730 (.A(net1109));
 sg13g2_antennanp ANTENNA_731 (.A(net1109));
 sg13g2_antennanp ANTENNA_732 (.A(net1109));
 sg13g2_antennanp ANTENNA_733 (.A(net1109));
 sg13g2_antennanp ANTENNA_734 (.A(net1109));
 sg13g2_antennanp ANTENNA_735 (.A(net1109));
 sg13g2_antennanp ANTENNA_736 (.A(net1109));
 sg13g2_antennanp ANTENNA_737 (.A(net1109));
 sg13g2_antennanp ANTENNA_738 (.A(net1109));
 sg13g2_antennanp ANTENNA_739 (.A(net1109));
 sg13g2_antennanp ANTENNA_740 (.A(net1109));
 sg13g2_antennanp ANTENNA_741 (.A(net1109));
 sg13g2_antennanp ANTENNA_742 (.A(net1109));
 sg13g2_antennanp ANTENNA_743 (.A(net1109));
 sg13g2_antennanp ANTENNA_744 (.A(net1109));
 sg13g2_antennanp ANTENNA_745 (.A(net1109));
 sg13g2_antennanp ANTENNA_746 (.A(net1109));
 sg13g2_antennanp ANTENNA_747 (.A(net1109));
 sg13g2_antennanp ANTENNA_748 (.A(net1109));
 sg13g2_antennanp ANTENNA_749 (.A(net1109));
 sg13g2_antennanp ANTENNA_750 (.A(net1109));
 sg13g2_antennanp ANTENNA_751 (.A(net1109));
 sg13g2_antennanp ANTENNA_752 (.A(net1109));
 sg13g2_antennanp ANTENNA_753 (.A(net1109));
 sg13g2_antennanp ANTENNA_754 (.A(net1109));
 sg13g2_antennanp ANTENNA_755 (.A(net1109));
 sg13g2_antennanp ANTENNA_756 (.A(net1109));
 sg13g2_antennanp ANTENNA_757 (.A(net1109));
 sg13g2_antennanp ANTENNA_758 (.A(net1109));
 sg13g2_antennanp ANTENNA_759 (.A(net1109));
 sg13g2_antennanp ANTENNA_760 (.A(net1110));
 sg13g2_antennanp ANTENNA_761 (.A(net1110));
 sg13g2_antennanp ANTENNA_762 (.A(net1110));
 sg13g2_antennanp ANTENNA_763 (.A(net1110));
 sg13g2_antennanp ANTENNA_764 (.A(net1110));
 sg13g2_antennanp ANTENNA_765 (.A(net1110));
 sg13g2_antennanp ANTENNA_766 (.A(net1110));
 sg13g2_antennanp ANTENNA_767 (.A(net1110));
 sg13g2_antennanp ANTENNA_768 (.A(net1110));
 sg13g2_antennanp ANTENNA_769 (.A(net1110));
 sg13g2_antennanp ANTENNA_770 (.A(net1110));
 sg13g2_antennanp ANTENNA_771 (.A(net1110));
 sg13g2_antennanp ANTENNA_772 (.A(net1110));
 sg13g2_antennanp ANTENNA_773 (.A(net1113));
 sg13g2_antennanp ANTENNA_774 (.A(net1113));
 sg13g2_antennanp ANTENNA_775 (.A(net1113));
 sg13g2_antennanp ANTENNA_776 (.A(net1113));
 sg13g2_antennanp ANTENNA_777 (.A(net1113));
 sg13g2_antennanp ANTENNA_778 (.A(net1113));
 sg13g2_antennanp ANTENNA_779 (.A(net1113));
 sg13g2_antennanp ANTENNA_780 (.A(net1113));
 sg13g2_antennanp ANTENNA_781 (.A(net1113));
 sg13g2_antennanp ANTENNA_782 (.A(net1150));
 sg13g2_antennanp ANTENNA_783 (.A(net1150));
 sg13g2_antennanp ANTENNA_784 (.A(net1150));
 sg13g2_antennanp ANTENNA_785 (.A(net1150));
 sg13g2_antennanp ANTENNA_786 (.A(net1150));
 sg13g2_antennanp ANTENNA_787 (.A(net1150));
 sg13g2_antennanp ANTENNA_788 (.A(net1150));
 sg13g2_antennanp ANTENNA_789 (.A(net1150));
 sg13g2_antennanp ANTENNA_790 (.A(net1150));
 sg13g2_antennanp ANTENNA_791 (.A(net1150));
 sg13g2_antennanp ANTENNA_792 (.A(net1150));
 sg13g2_antennanp ANTENNA_793 (.A(net1150));
 sg13g2_antennanp ANTENNA_794 (.A(net1150));
 sg13g2_antennanp ANTENNA_795 (.A(_00000_));
 sg13g2_antennanp ANTENNA_796 (.A(_00000_));
 sg13g2_antennanp ANTENNA_797 (.A(_00230_));
 sg13g2_antennanp ANTENNA_798 (.A(_00237_));
 sg13g2_antennanp ANTENNA_799 (.A(_00237_));
 sg13g2_antennanp ANTENNA_800 (.A(_00237_));
 sg13g2_antennanp ANTENNA_801 (.A(_00752_));
 sg13g2_antennanp ANTENNA_802 (.A(_00800_));
 sg13g2_antennanp ANTENNA_803 (.A(_00800_));
 sg13g2_antennanp ANTENNA_804 (.A(_01061_));
 sg13g2_antennanp ANTENNA_805 (.A(_01063_));
 sg13g2_antennanp ANTENNA_806 (.A(_01066_));
 sg13g2_antennanp ANTENNA_807 (.A(_02909_));
 sg13g2_antennanp ANTENNA_808 (.A(_02909_));
 sg13g2_antennanp ANTENNA_809 (.A(_02909_));
 sg13g2_antennanp ANTENNA_810 (.A(_02909_));
 sg13g2_antennanp ANTENNA_811 (.A(_02909_));
 sg13g2_antennanp ANTENNA_812 (.A(_02909_));
 sg13g2_antennanp ANTENNA_813 (.A(_02909_));
 sg13g2_antennanp ANTENNA_814 (.A(_02909_));
 sg13g2_antennanp ANTENNA_815 (.A(_02909_));
 sg13g2_antennanp ANTENNA_816 (.A(_02918_));
 sg13g2_antennanp ANTENNA_817 (.A(_02918_));
 sg13g2_antennanp ANTENNA_818 (.A(_02918_));
 sg13g2_antennanp ANTENNA_819 (.A(_02918_));
 sg13g2_antennanp ANTENNA_820 (.A(_02918_));
 sg13g2_antennanp ANTENNA_821 (.A(_02918_));
 sg13g2_antennanp ANTENNA_822 (.A(_02918_));
 sg13g2_antennanp ANTENNA_823 (.A(_02918_));
 sg13g2_antennanp ANTENNA_824 (.A(_02918_));
 sg13g2_antennanp ANTENNA_825 (.A(_02922_));
 sg13g2_antennanp ANTENNA_826 (.A(_02922_));
 sg13g2_antennanp ANTENNA_827 (.A(_02922_));
 sg13g2_antennanp ANTENNA_828 (.A(_02922_));
 sg13g2_antennanp ANTENNA_829 (.A(_02922_));
 sg13g2_antennanp ANTENNA_830 (.A(_02922_));
 sg13g2_antennanp ANTENNA_831 (.A(_02922_));
 sg13g2_antennanp ANTENNA_832 (.A(_02922_));
 sg13g2_antennanp ANTENNA_833 (.A(_02922_));
 sg13g2_antennanp ANTENNA_834 (.A(_02933_));
 sg13g2_antennanp ANTENNA_835 (.A(_02933_));
 sg13g2_antennanp ANTENNA_836 (.A(_02933_));
 sg13g2_antennanp ANTENNA_837 (.A(_02933_));
 sg13g2_antennanp ANTENNA_838 (.A(_02933_));
 sg13g2_antennanp ANTENNA_839 (.A(_02933_));
 sg13g2_antennanp ANTENNA_840 (.A(_02933_));
 sg13g2_antennanp ANTENNA_841 (.A(_02933_));
 sg13g2_antennanp ANTENNA_842 (.A(_02933_));
 sg13g2_antennanp ANTENNA_843 (.A(_03020_));
 sg13g2_antennanp ANTENNA_844 (.A(_03020_));
 sg13g2_antennanp ANTENNA_845 (.A(_03020_));
 sg13g2_antennanp ANTENNA_846 (.A(_03161_));
 sg13g2_antennanp ANTENNA_847 (.A(_03535_));
 sg13g2_antennanp ANTENNA_848 (.A(_03535_));
 sg13g2_antennanp ANTENNA_849 (.A(_03535_));
 sg13g2_antennanp ANTENNA_850 (.A(_03535_));
 sg13g2_antennanp ANTENNA_851 (.A(_03535_));
 sg13g2_antennanp ANTENNA_852 (.A(_03535_));
 sg13g2_antennanp ANTENNA_853 (.A(_03535_));
 sg13g2_antennanp ANTENNA_854 (.A(_03535_));
 sg13g2_antennanp ANTENNA_855 (.A(_03535_));
 sg13g2_antennanp ANTENNA_856 (.A(_03535_));
 sg13g2_antennanp ANTENNA_857 (.A(_03535_));
 sg13g2_antennanp ANTENNA_858 (.A(_03535_));
 sg13g2_antennanp ANTENNA_859 (.A(_03535_));
 sg13g2_antennanp ANTENNA_860 (.A(_03535_));
 sg13g2_antennanp ANTENNA_861 (.A(_04843_));
 sg13g2_antennanp ANTENNA_862 (.A(_04890_));
 sg13g2_antennanp ANTENNA_863 (.A(_04890_));
 sg13g2_antennanp ANTENNA_864 (.A(_04890_));
 sg13g2_antennanp ANTENNA_865 (.A(_04890_));
 sg13g2_antennanp ANTENNA_866 (.A(_04914_));
 sg13g2_antennanp ANTENNA_867 (.A(_04954_));
 sg13g2_antennanp ANTENNA_868 (.A(_05005_));
 sg13g2_antennanp ANTENNA_869 (.A(_05175_));
 sg13g2_antennanp ANTENNA_870 (.A(_05207_));
 sg13g2_antennanp ANTENNA_871 (.A(_05231_));
 sg13g2_antennanp ANTENNA_872 (.A(_05267_));
 sg13g2_antennanp ANTENNA_873 (.A(_05282_));
 sg13g2_antennanp ANTENNA_874 (.A(_05293_));
 sg13g2_antennanp ANTENNA_875 (.A(_05293_));
 sg13g2_antennanp ANTENNA_876 (.A(_05293_));
 sg13g2_antennanp ANTENNA_877 (.A(_05373_));
 sg13g2_antennanp ANTENNA_878 (.A(_05437_));
 sg13g2_antennanp ANTENNA_879 (.A(_05437_));
 sg13g2_antennanp ANTENNA_880 (.A(_05577_));
 sg13g2_antennanp ANTENNA_881 (.A(_05649_));
 sg13g2_antennanp ANTENNA_882 (.A(_05722_));
 sg13g2_antennanp ANTENNA_883 (.A(_05737_));
 sg13g2_antennanp ANTENNA_884 (.A(_05783_));
 sg13g2_antennanp ANTENNA_885 (.A(_05789_));
 sg13g2_antennanp ANTENNA_886 (.A(_05792_));
 sg13g2_antennanp ANTENNA_887 (.A(_05795_));
 sg13g2_antennanp ANTENNA_888 (.A(_05800_));
 sg13g2_antennanp ANTENNA_889 (.A(_05800_));
 sg13g2_antennanp ANTENNA_890 (.A(_05800_));
 sg13g2_antennanp ANTENNA_891 (.A(_05838_));
 sg13g2_antennanp ANTENNA_892 (.A(_05838_));
 sg13g2_antennanp ANTENNA_893 (.A(_05838_));
 sg13g2_antennanp ANTENNA_894 (.A(_05838_));
 sg13g2_antennanp ANTENNA_895 (.A(_05838_));
 sg13g2_antennanp ANTENNA_896 (.A(_05838_));
 sg13g2_antennanp ANTENNA_897 (.A(_05838_));
 sg13g2_antennanp ANTENNA_898 (.A(_05838_));
 sg13g2_antennanp ANTENNA_899 (.A(_05838_));
 sg13g2_antennanp ANTENNA_900 (.A(_05838_));
 sg13g2_antennanp ANTENNA_901 (.A(_06038_));
 sg13g2_antennanp ANTENNA_902 (.A(_06479_));
 sg13g2_antennanp ANTENNA_903 (.A(_06479_));
 sg13g2_antennanp ANTENNA_904 (.A(_06479_));
 sg13g2_antennanp ANTENNA_905 (.A(_06479_));
 sg13g2_antennanp ANTENNA_906 (.A(_06479_));
 sg13g2_antennanp ANTENNA_907 (.A(_06479_));
 sg13g2_antennanp ANTENNA_908 (.A(_06479_));
 sg13g2_antennanp ANTENNA_909 (.A(_06479_));
 sg13g2_antennanp ANTENNA_910 (.A(_06479_));
 sg13g2_antennanp ANTENNA_911 (.A(_06822_));
 sg13g2_antennanp ANTENNA_912 (.A(_06856_));
 sg13g2_antennanp ANTENNA_913 (.A(_06905_));
 sg13g2_antennanp ANTENNA_914 (.A(_06978_));
 sg13g2_antennanp ANTENNA_915 (.A(_07663_));
 sg13g2_antennanp ANTENNA_916 (.A(_07663_));
 sg13g2_antennanp ANTENNA_917 (.A(_07663_));
 sg13g2_antennanp ANTENNA_918 (.A(_07663_));
 sg13g2_antennanp ANTENNA_919 (.A(_07663_));
 sg13g2_antennanp ANTENNA_920 (.A(_07663_));
 sg13g2_antennanp ANTENNA_921 (.A(_07663_));
 sg13g2_antennanp ANTENNA_922 (.A(_07663_));
 sg13g2_antennanp ANTENNA_923 (.A(_07663_));
 sg13g2_antennanp ANTENNA_924 (.A(_07663_));
 sg13g2_antennanp ANTENNA_925 (.A(_08377_));
 sg13g2_antennanp ANTENNA_926 (.A(_08377_));
 sg13g2_antennanp ANTENNA_927 (.A(_08377_));
 sg13g2_antennanp ANTENNA_928 (.A(_08411_));
 sg13g2_antennanp ANTENNA_929 (.A(_08411_));
 sg13g2_antennanp ANTENNA_930 (.A(_08411_));
 sg13g2_antennanp ANTENNA_931 (.A(_08411_));
 sg13g2_antennanp ANTENNA_932 (.A(_08443_));
 sg13g2_antennanp ANTENNA_933 (.A(_08443_));
 sg13g2_antennanp ANTENNA_934 (.A(_08443_));
 sg13g2_antennanp ANTENNA_935 (.A(_08486_));
 sg13g2_antennanp ANTENNA_936 (.A(_08556_));
 sg13g2_antennanp ANTENNA_937 (.A(_08556_));
 sg13g2_antennanp ANTENNA_938 (.A(_08556_));
 sg13g2_antennanp ANTENNA_939 (.A(_08565_));
 sg13g2_antennanp ANTENNA_940 (.A(_08565_));
 sg13g2_antennanp ANTENNA_941 (.A(_08565_));
 sg13g2_antennanp ANTENNA_942 (.A(_08565_));
 sg13g2_antennanp ANTENNA_943 (.A(_08565_));
 sg13g2_antennanp ANTENNA_944 (.A(_08565_));
 sg13g2_antennanp ANTENNA_945 (.A(_08669_));
 sg13g2_antennanp ANTENNA_946 (.A(_08691_));
 sg13g2_antennanp ANTENNA_947 (.A(_08691_));
 sg13g2_antennanp ANTENNA_948 (.A(_08691_));
 sg13g2_antennanp ANTENNA_949 (.A(_08804_));
 sg13g2_antennanp ANTENNA_950 (.A(_08839_));
 sg13g2_antennanp ANTENNA_951 (.A(_08839_));
 sg13g2_antennanp ANTENNA_952 (.A(_08839_));
 sg13g2_antennanp ANTENNA_953 (.A(_08894_));
 sg13g2_antennanp ANTENNA_954 (.A(_08894_));
 sg13g2_antennanp ANTENNA_955 (.A(_08894_));
 sg13g2_antennanp ANTENNA_956 (.A(_08940_));
 sg13g2_antennanp ANTENNA_957 (.A(_08940_));
 sg13g2_antennanp ANTENNA_958 (.A(_08976_));
 sg13g2_antennanp ANTENNA_959 (.A(_09068_));
 sg13g2_antennanp ANTENNA_960 (.A(_09223_));
 sg13g2_antennanp ANTENNA_961 (.A(_09223_));
 sg13g2_antennanp ANTENNA_962 (.A(_09223_));
 sg13g2_antennanp ANTENNA_963 (.A(_09223_));
 sg13g2_antennanp ANTENNA_964 (.A(_09225_));
 sg13g2_antennanp ANTENNA_965 (.A(_09225_));
 sg13g2_antennanp ANTENNA_966 (.A(_09225_));
 sg13g2_antennanp ANTENNA_967 (.A(_09225_));
 sg13g2_antennanp ANTENNA_968 (.A(_09227_));
 sg13g2_antennanp ANTENNA_969 (.A(_09227_));
 sg13g2_antennanp ANTENNA_970 (.A(_09227_));
 sg13g2_antennanp ANTENNA_971 (.A(_09227_));
 sg13g2_antennanp ANTENNA_972 (.A(_09227_));
 sg13g2_antennanp ANTENNA_973 (.A(_09227_));
 sg13g2_antennanp ANTENNA_974 (.A(_09240_));
 sg13g2_antennanp ANTENNA_975 (.A(_09240_));
 sg13g2_antennanp ANTENNA_976 (.A(_09240_));
 sg13g2_antennanp ANTENNA_977 (.A(_09240_));
 sg13g2_antennanp ANTENNA_978 (.A(_09240_));
 sg13g2_antennanp ANTENNA_979 (.A(_09240_));
 sg13g2_antennanp ANTENNA_980 (.A(_09282_));
 sg13g2_antennanp ANTENNA_981 (.A(_09282_));
 sg13g2_antennanp ANTENNA_982 (.A(_09282_));
 sg13g2_antennanp ANTENNA_983 (.A(_09282_));
 sg13g2_antennanp ANTENNA_984 (.A(_09284_));
 sg13g2_antennanp ANTENNA_985 (.A(_09284_));
 sg13g2_antennanp ANTENNA_986 (.A(_09284_));
 sg13g2_antennanp ANTENNA_987 (.A(_09284_));
 sg13g2_antennanp ANTENNA_988 (.A(_09310_));
 sg13g2_antennanp ANTENNA_989 (.A(_09310_));
 sg13g2_antennanp ANTENNA_990 (.A(_09310_));
 sg13g2_antennanp ANTENNA_991 (.A(_09363_));
 sg13g2_antennanp ANTENNA_992 (.A(_09363_));
 sg13g2_antennanp ANTENNA_993 (.A(_09363_));
 sg13g2_antennanp ANTENNA_994 (.A(_09365_));
 sg13g2_antennanp ANTENNA_995 (.A(_09365_));
 sg13g2_antennanp ANTENNA_996 (.A(_09365_));
 sg13g2_antennanp ANTENNA_997 (.A(_09365_));
 sg13g2_antennanp ANTENNA_998 (.A(_09435_));
 sg13g2_antennanp ANTENNA_999 (.A(_09435_));
 sg13g2_antennanp ANTENNA_1000 (.A(_09435_));
 sg13g2_antennanp ANTENNA_1001 (.A(_09512_));
 sg13g2_antennanp ANTENNA_1002 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1003 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1004 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1005 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1006 (.A(_09588_));
 sg13g2_antennanp ANTENNA_1007 (.A(_09639_));
 sg13g2_antennanp ANTENNA_1008 (.A(_09700_));
 sg13g2_antennanp ANTENNA_1009 (.A(_09854_));
 sg13g2_antennanp ANTENNA_1010 (.A(_09897_));
 sg13g2_antennanp ANTENNA_1011 (.A(_09897_));
 sg13g2_antennanp ANTENNA_1012 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1013 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1014 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1015 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1016 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1017 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1018 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1019 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1020 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1021 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1022 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1023 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1024 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1025 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1026 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1027 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1028 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1029 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1030 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1031 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1032 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1033 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1034 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1035 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1036 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1037 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1038 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1039 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1040 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1041 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1042 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1043 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1044 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1045 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1046 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1047 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1048 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1049 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1050 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1051 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1052 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1053 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1054 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1055 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1056 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1057 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1058 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1059 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1060 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1061 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1062 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1063 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1064 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1065 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1066 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1067 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1068 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1069 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1070 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1071 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1072 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1073 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1074 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1075 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1076 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1077 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1078 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1079 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1080 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1081 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1082 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1083 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1084 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1085 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1086 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1087 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1088 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1089 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1090 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1091 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1092 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1093 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1094 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1095 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1096 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1097 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1098 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1099 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1100 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1101 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1102 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1103 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1104 (.A(_12255_));
 sg13g2_antennanp ANTENNA_1105 (.A(_12255_));
 sg13g2_antennanp ANTENNA_1106 (.A(_12255_));
 sg13g2_antennanp ANTENNA_1107 (.A(clk));
 sg13g2_antennanp ANTENNA_1108 (.A(clk));
 sg13g2_antennanp ANTENNA_1109 (.A(\cpu.d_flush_all ));
 sg13g2_antennanp ANTENNA_1110 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1111 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_1112 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_1113 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1114 (.A(net1));
 sg13g2_antennanp ANTENNA_1115 (.A(net1));
 sg13g2_antennanp ANTENNA_1116 (.A(net1));
 sg13g2_antennanp ANTENNA_1117 (.A(net1));
 sg13g2_antennanp ANTENNA_1118 (.A(net1));
 sg13g2_antennanp ANTENNA_1119 (.A(net1));
 sg13g2_antennanp ANTENNA_1120 (.A(net1));
 sg13g2_antennanp ANTENNA_1121 (.A(net1));
 sg13g2_antennanp ANTENNA_1122 (.A(net3));
 sg13g2_antennanp ANTENNA_1123 (.A(net3));
 sg13g2_antennanp ANTENNA_1124 (.A(net11));
 sg13g2_antennanp ANTENNA_1125 (.A(net11));
 sg13g2_antennanp ANTENNA_1126 (.A(net12));
 sg13g2_antennanp ANTENNA_1127 (.A(net12));
 sg13g2_antennanp ANTENNA_1128 (.A(net14));
 sg13g2_antennanp ANTENNA_1129 (.A(net14));
 sg13g2_antennanp ANTENNA_1130 (.A(net484));
 sg13g2_antennanp ANTENNA_1131 (.A(net484));
 sg13g2_antennanp ANTENNA_1132 (.A(net484));
 sg13g2_antennanp ANTENNA_1133 (.A(net484));
 sg13g2_antennanp ANTENNA_1134 (.A(net484));
 sg13g2_antennanp ANTENNA_1135 (.A(net484));
 sg13g2_antennanp ANTENNA_1136 (.A(net484));
 sg13g2_antennanp ANTENNA_1137 (.A(net484));
 sg13g2_antennanp ANTENNA_1138 (.A(net484));
 sg13g2_antennanp ANTENNA_1139 (.A(net520));
 sg13g2_antennanp ANTENNA_1140 (.A(net520));
 sg13g2_antennanp ANTENNA_1141 (.A(net520));
 sg13g2_antennanp ANTENNA_1142 (.A(net520));
 sg13g2_antennanp ANTENNA_1143 (.A(net520));
 sg13g2_antennanp ANTENNA_1144 (.A(net520));
 sg13g2_antennanp ANTENNA_1145 (.A(net520));
 sg13g2_antennanp ANTENNA_1146 (.A(net520));
 sg13g2_antennanp ANTENNA_1147 (.A(net544));
 sg13g2_antennanp ANTENNA_1148 (.A(net544));
 sg13g2_antennanp ANTENNA_1149 (.A(net544));
 sg13g2_antennanp ANTENNA_1150 (.A(net544));
 sg13g2_antennanp ANTENNA_1151 (.A(net544));
 sg13g2_antennanp ANTENNA_1152 (.A(net544));
 sg13g2_antennanp ANTENNA_1153 (.A(net544));
 sg13g2_antennanp ANTENNA_1154 (.A(net544));
 sg13g2_antennanp ANTENNA_1155 (.A(net544));
 sg13g2_antennanp ANTENNA_1156 (.A(net544));
 sg13g2_antennanp ANTENNA_1157 (.A(net544));
 sg13g2_antennanp ANTENNA_1158 (.A(net544));
 sg13g2_antennanp ANTENNA_1159 (.A(net544));
 sg13g2_antennanp ANTENNA_1160 (.A(net544));
 sg13g2_antennanp ANTENNA_1161 (.A(net653));
 sg13g2_antennanp ANTENNA_1162 (.A(net653));
 sg13g2_antennanp ANTENNA_1163 (.A(net653));
 sg13g2_antennanp ANTENNA_1164 (.A(net653));
 sg13g2_antennanp ANTENNA_1165 (.A(net653));
 sg13g2_antennanp ANTENNA_1166 (.A(net653));
 sg13g2_antennanp ANTENNA_1167 (.A(net653));
 sg13g2_antennanp ANTENNA_1168 (.A(net653));
 sg13g2_antennanp ANTENNA_1169 (.A(net653));
 sg13g2_antennanp ANTENNA_1170 (.A(net653));
 sg13g2_antennanp ANTENNA_1171 (.A(net653));
 sg13g2_antennanp ANTENNA_1172 (.A(net653));
 sg13g2_antennanp ANTENNA_1173 (.A(net653));
 sg13g2_antennanp ANTENNA_1174 (.A(net653));
 sg13g2_antennanp ANTENNA_1175 (.A(net653));
 sg13g2_antennanp ANTENNA_1176 (.A(net653));
 sg13g2_antennanp ANTENNA_1177 (.A(net653));
 sg13g2_antennanp ANTENNA_1178 (.A(net653));
 sg13g2_antennanp ANTENNA_1179 (.A(net728));
 sg13g2_antennanp ANTENNA_1180 (.A(net728));
 sg13g2_antennanp ANTENNA_1181 (.A(net728));
 sg13g2_antennanp ANTENNA_1182 (.A(net728));
 sg13g2_antennanp ANTENNA_1183 (.A(net728));
 sg13g2_antennanp ANTENNA_1184 (.A(net728));
 sg13g2_antennanp ANTENNA_1185 (.A(net728));
 sg13g2_antennanp ANTENNA_1186 (.A(net728));
 sg13g2_antennanp ANTENNA_1187 (.A(net797));
 sg13g2_antennanp ANTENNA_1188 (.A(net797));
 sg13g2_antennanp ANTENNA_1189 (.A(net797));
 sg13g2_antennanp ANTENNA_1190 (.A(net797));
 sg13g2_antennanp ANTENNA_1191 (.A(net797));
 sg13g2_antennanp ANTENNA_1192 (.A(net797));
 sg13g2_antennanp ANTENNA_1193 (.A(net797));
 sg13g2_antennanp ANTENNA_1194 (.A(net797));
 sg13g2_antennanp ANTENNA_1195 (.A(net797));
 sg13g2_antennanp ANTENNA_1196 (.A(net812));
 sg13g2_antennanp ANTENNA_1197 (.A(net812));
 sg13g2_antennanp ANTENNA_1198 (.A(net812));
 sg13g2_antennanp ANTENNA_1199 (.A(net812));
 sg13g2_antennanp ANTENNA_1200 (.A(net812));
 sg13g2_antennanp ANTENNA_1201 (.A(net812));
 sg13g2_antennanp ANTENNA_1202 (.A(net812));
 sg13g2_antennanp ANTENNA_1203 (.A(net812));
 sg13g2_antennanp ANTENNA_1204 (.A(net812));
 sg13g2_antennanp ANTENNA_1205 (.A(net812));
 sg13g2_antennanp ANTENNA_1206 (.A(net812));
 sg13g2_antennanp ANTENNA_1207 (.A(net812));
 sg13g2_antennanp ANTENNA_1208 (.A(net812));
 sg13g2_antennanp ANTENNA_1209 (.A(net812));
 sg13g2_antennanp ANTENNA_1210 (.A(net812));
 sg13g2_antennanp ANTENNA_1211 (.A(net812));
 sg13g2_antennanp ANTENNA_1212 (.A(net812));
 sg13g2_antennanp ANTENNA_1213 (.A(net812));
 sg13g2_antennanp ANTENNA_1214 (.A(net812));
 sg13g2_antennanp ANTENNA_1215 (.A(net812));
 sg13g2_antennanp ANTENNA_1216 (.A(net861));
 sg13g2_antennanp ANTENNA_1217 (.A(net861));
 sg13g2_antennanp ANTENNA_1218 (.A(net861));
 sg13g2_antennanp ANTENNA_1219 (.A(net861));
 sg13g2_antennanp ANTENNA_1220 (.A(net861));
 sg13g2_antennanp ANTENNA_1221 (.A(net861));
 sg13g2_antennanp ANTENNA_1222 (.A(net861));
 sg13g2_antennanp ANTENNA_1223 (.A(net861));
 sg13g2_antennanp ANTENNA_1224 (.A(net861));
 sg13g2_antennanp ANTENNA_1225 (.A(net861));
 sg13g2_antennanp ANTENNA_1226 (.A(net861));
 sg13g2_antennanp ANTENNA_1227 (.A(net861));
 sg13g2_antennanp ANTENNA_1228 (.A(net861));
 sg13g2_antennanp ANTENNA_1229 (.A(net861));
 sg13g2_antennanp ANTENNA_1230 (.A(net861));
 sg13g2_antennanp ANTENNA_1231 (.A(net861));
 sg13g2_antennanp ANTENNA_1232 (.A(net862));
 sg13g2_antennanp ANTENNA_1233 (.A(net862));
 sg13g2_antennanp ANTENNA_1234 (.A(net862));
 sg13g2_antennanp ANTENNA_1235 (.A(net862));
 sg13g2_antennanp ANTENNA_1236 (.A(net862));
 sg13g2_antennanp ANTENNA_1237 (.A(net862));
 sg13g2_antennanp ANTENNA_1238 (.A(net862));
 sg13g2_antennanp ANTENNA_1239 (.A(net862));
 sg13g2_antennanp ANTENNA_1240 (.A(net862));
 sg13g2_antennanp ANTENNA_1241 (.A(net862));
 sg13g2_antennanp ANTENNA_1242 (.A(net862));
 sg13g2_antennanp ANTENNA_1243 (.A(net862));
 sg13g2_antennanp ANTENNA_1244 (.A(net862));
 sg13g2_antennanp ANTENNA_1245 (.A(net862));
 sg13g2_antennanp ANTENNA_1246 (.A(net862));
 sg13g2_antennanp ANTENNA_1247 (.A(net862));
 sg13g2_antennanp ANTENNA_1248 (.A(net862));
 sg13g2_antennanp ANTENNA_1249 (.A(net862));
 sg13g2_antennanp ANTENNA_1250 (.A(net862));
 sg13g2_antennanp ANTENNA_1251 (.A(net862));
 sg13g2_antennanp ANTENNA_1252 (.A(net862));
 sg13g2_antennanp ANTENNA_1253 (.A(net862));
 sg13g2_antennanp ANTENNA_1254 (.A(net862));
 sg13g2_antennanp ANTENNA_1255 (.A(net862));
 sg13g2_antennanp ANTENNA_1256 (.A(net862));
 sg13g2_antennanp ANTENNA_1257 (.A(net862));
 sg13g2_antennanp ANTENNA_1258 (.A(net862));
 sg13g2_antennanp ANTENNA_1259 (.A(net862));
 sg13g2_antennanp ANTENNA_1260 (.A(net862));
 sg13g2_antennanp ANTENNA_1261 (.A(net862));
 sg13g2_antennanp ANTENNA_1262 (.A(net907));
 sg13g2_antennanp ANTENNA_1263 (.A(net907));
 sg13g2_antennanp ANTENNA_1264 (.A(net907));
 sg13g2_antennanp ANTENNA_1265 (.A(net907));
 sg13g2_antennanp ANTENNA_1266 (.A(net907));
 sg13g2_antennanp ANTENNA_1267 (.A(net907));
 sg13g2_antennanp ANTENNA_1268 (.A(net907));
 sg13g2_antennanp ANTENNA_1269 (.A(net907));
 sg13g2_antennanp ANTENNA_1270 (.A(net907));
 sg13g2_antennanp ANTENNA_1271 (.A(net907));
 sg13g2_antennanp ANTENNA_1272 (.A(net907));
 sg13g2_antennanp ANTENNA_1273 (.A(net907));
 sg13g2_antennanp ANTENNA_1274 (.A(net907));
 sg13g2_antennanp ANTENNA_1275 (.A(net907));
 sg13g2_antennanp ANTENNA_1276 (.A(net907));
 sg13g2_antennanp ANTENNA_1277 (.A(net916));
 sg13g2_antennanp ANTENNA_1278 (.A(net916));
 sg13g2_antennanp ANTENNA_1279 (.A(net916));
 sg13g2_antennanp ANTENNA_1280 (.A(net916));
 sg13g2_antennanp ANTENNA_1281 (.A(net916));
 sg13g2_antennanp ANTENNA_1282 (.A(net916));
 sg13g2_antennanp ANTENNA_1283 (.A(net916));
 sg13g2_antennanp ANTENNA_1284 (.A(net916));
 sg13g2_antennanp ANTENNA_1285 (.A(net916));
 sg13g2_antennanp ANTENNA_1286 (.A(net916));
 sg13g2_antennanp ANTENNA_1287 (.A(net916));
 sg13g2_antennanp ANTENNA_1288 (.A(net916));
 sg13g2_antennanp ANTENNA_1289 (.A(net916));
 sg13g2_antennanp ANTENNA_1290 (.A(net916));
 sg13g2_antennanp ANTENNA_1291 (.A(net916));
 sg13g2_antennanp ANTENNA_1292 (.A(net916));
 sg13g2_antennanp ANTENNA_1293 (.A(net993));
 sg13g2_antennanp ANTENNA_1294 (.A(net993));
 sg13g2_antennanp ANTENNA_1295 (.A(net993));
 sg13g2_antennanp ANTENNA_1296 (.A(net993));
 sg13g2_antennanp ANTENNA_1297 (.A(net993));
 sg13g2_antennanp ANTENNA_1298 (.A(net993));
 sg13g2_antennanp ANTENNA_1299 (.A(net993));
 sg13g2_antennanp ANTENNA_1300 (.A(net993));
 sg13g2_antennanp ANTENNA_1301 (.A(net993));
 sg13g2_antennanp ANTENNA_1302 (.A(net993));
 sg13g2_antennanp ANTENNA_1303 (.A(net993));
 sg13g2_antennanp ANTENNA_1304 (.A(net993));
 sg13g2_antennanp ANTENNA_1305 (.A(net993));
 sg13g2_antennanp ANTENNA_1306 (.A(net993));
 sg13g2_antennanp ANTENNA_1307 (.A(net993));
 sg13g2_antennanp ANTENNA_1308 (.A(net993));
 sg13g2_antennanp ANTENNA_1309 (.A(net1020));
 sg13g2_antennanp ANTENNA_1310 (.A(net1020));
 sg13g2_antennanp ANTENNA_1311 (.A(net1020));
 sg13g2_antennanp ANTENNA_1312 (.A(net1020));
 sg13g2_antennanp ANTENNA_1313 (.A(net1020));
 sg13g2_antennanp ANTENNA_1314 (.A(net1020));
 sg13g2_antennanp ANTENNA_1315 (.A(net1020));
 sg13g2_antennanp ANTENNA_1316 (.A(net1020));
 sg13g2_antennanp ANTENNA_1317 (.A(net1020));
 sg13g2_antennanp ANTENNA_1318 (.A(net1021));
 sg13g2_antennanp ANTENNA_1319 (.A(net1021));
 sg13g2_antennanp ANTENNA_1320 (.A(net1021));
 sg13g2_antennanp ANTENNA_1321 (.A(net1021));
 sg13g2_antennanp ANTENNA_1322 (.A(net1021));
 sg13g2_antennanp ANTENNA_1323 (.A(net1021));
 sg13g2_antennanp ANTENNA_1324 (.A(net1021));
 sg13g2_antennanp ANTENNA_1325 (.A(net1021));
 sg13g2_antennanp ANTENNA_1326 (.A(net1021));
 sg13g2_antennanp ANTENNA_1327 (.A(net1021));
 sg13g2_antennanp ANTENNA_1328 (.A(net1021));
 sg13g2_antennanp ANTENNA_1329 (.A(net1021));
 sg13g2_antennanp ANTENNA_1330 (.A(net1021));
 sg13g2_antennanp ANTENNA_1331 (.A(net1021));
 sg13g2_antennanp ANTENNA_1332 (.A(net1070));
 sg13g2_antennanp ANTENNA_1333 (.A(net1070));
 sg13g2_antennanp ANTENNA_1334 (.A(net1070));
 sg13g2_antennanp ANTENNA_1335 (.A(net1070));
 sg13g2_antennanp ANTENNA_1336 (.A(net1070));
 sg13g2_antennanp ANTENNA_1337 (.A(net1070));
 sg13g2_antennanp ANTENNA_1338 (.A(net1070));
 sg13g2_antennanp ANTENNA_1339 (.A(net1070));
 sg13g2_antennanp ANTENNA_1340 (.A(net1071));
 sg13g2_antennanp ANTENNA_1341 (.A(net1071));
 sg13g2_antennanp ANTENNA_1342 (.A(net1071));
 sg13g2_antennanp ANTENNA_1343 (.A(net1071));
 sg13g2_antennanp ANTENNA_1344 (.A(net1071));
 sg13g2_antennanp ANTENNA_1345 (.A(net1071));
 sg13g2_antennanp ANTENNA_1346 (.A(net1071));
 sg13g2_antennanp ANTENNA_1347 (.A(net1071));
 sg13g2_antennanp ANTENNA_1348 (.A(net1071));
 sg13g2_antennanp ANTENNA_1349 (.A(net1109));
 sg13g2_antennanp ANTENNA_1350 (.A(net1109));
 sg13g2_antennanp ANTENNA_1351 (.A(net1109));
 sg13g2_antennanp ANTENNA_1352 (.A(net1109));
 sg13g2_antennanp ANTENNA_1353 (.A(net1109));
 sg13g2_antennanp ANTENNA_1354 (.A(net1109));
 sg13g2_antennanp ANTENNA_1355 (.A(net1109));
 sg13g2_antennanp ANTENNA_1356 (.A(net1109));
 sg13g2_antennanp ANTENNA_1357 (.A(net1109));
 sg13g2_antennanp ANTENNA_1358 (.A(net1109));
 sg13g2_antennanp ANTENNA_1359 (.A(net1109));
 sg13g2_antennanp ANTENNA_1360 (.A(net1109));
 sg13g2_antennanp ANTENNA_1361 (.A(net1109));
 sg13g2_antennanp ANTENNA_1362 (.A(net1109));
 sg13g2_antennanp ANTENNA_1363 (.A(net1109));
 sg13g2_antennanp ANTENNA_1364 (.A(net1109));
 sg13g2_antennanp ANTENNA_1365 (.A(net1109));
 sg13g2_antennanp ANTENNA_1366 (.A(net1109));
 sg13g2_antennanp ANTENNA_1367 (.A(net1109));
 sg13g2_antennanp ANTENNA_1368 (.A(net1109));
 sg13g2_antennanp ANTENNA_1369 (.A(net1109));
 sg13g2_antennanp ANTENNA_1370 (.A(net1109));
 sg13g2_antennanp ANTENNA_1371 (.A(net1109));
 sg13g2_antennanp ANTENNA_1372 (.A(net1109));
 sg13g2_antennanp ANTENNA_1373 (.A(net1109));
 sg13g2_antennanp ANTENNA_1374 (.A(net1109));
 sg13g2_antennanp ANTENNA_1375 (.A(net1109));
 sg13g2_antennanp ANTENNA_1376 (.A(net1109));
 sg13g2_antennanp ANTENNA_1377 (.A(net1109));
 sg13g2_antennanp ANTENNA_1378 (.A(net1109));
 sg13g2_antennanp ANTENNA_1379 (.A(net1111));
 sg13g2_antennanp ANTENNA_1380 (.A(net1111));
 sg13g2_antennanp ANTENNA_1381 (.A(net1111));
 sg13g2_antennanp ANTENNA_1382 (.A(net1111));
 sg13g2_antennanp ANTENNA_1383 (.A(net1111));
 sg13g2_antennanp ANTENNA_1384 (.A(net1111));
 sg13g2_antennanp ANTENNA_1385 (.A(net1111));
 sg13g2_antennanp ANTENNA_1386 (.A(net1111));
 sg13g2_antennanp ANTENNA_1387 (.A(net1111));
 sg13g2_antennanp ANTENNA_1388 (.A(net1111));
 sg13g2_antennanp ANTENNA_1389 (.A(net1111));
 sg13g2_antennanp ANTENNA_1390 (.A(net1111));
 sg13g2_antennanp ANTENNA_1391 (.A(net1111));
 sg13g2_antennanp ANTENNA_1392 (.A(net1111));
 sg13g2_antennanp ANTENNA_1393 (.A(net1113));
 sg13g2_antennanp ANTENNA_1394 (.A(net1113));
 sg13g2_antennanp ANTENNA_1395 (.A(net1113));
 sg13g2_antennanp ANTENNA_1396 (.A(net1113));
 sg13g2_antennanp ANTENNA_1397 (.A(net1113));
 sg13g2_antennanp ANTENNA_1398 (.A(net1113));
 sg13g2_antennanp ANTENNA_1399 (.A(net1113));
 sg13g2_antennanp ANTENNA_1400 (.A(net1113));
 sg13g2_antennanp ANTENNA_1401 (.A(net1113));
 sg13g2_antennanp ANTENNA_1402 (.A(net1114));
 sg13g2_antennanp ANTENNA_1403 (.A(net1114));
 sg13g2_antennanp ANTENNA_1404 (.A(net1114));
 sg13g2_antennanp ANTENNA_1405 (.A(net1114));
 sg13g2_antennanp ANTENNA_1406 (.A(net1114));
 sg13g2_antennanp ANTENNA_1407 (.A(net1114));
 sg13g2_antennanp ANTENNA_1408 (.A(net1114));
 sg13g2_antennanp ANTENNA_1409 (.A(net1114));
 sg13g2_antennanp ANTENNA_1410 (.A(net1114));
 sg13g2_antennanp ANTENNA_1411 (.A(net1150));
 sg13g2_antennanp ANTENNA_1412 (.A(net1150));
 sg13g2_antennanp ANTENNA_1413 (.A(net1150));
 sg13g2_antennanp ANTENNA_1414 (.A(net1150));
 sg13g2_antennanp ANTENNA_1415 (.A(net1150));
 sg13g2_antennanp ANTENNA_1416 (.A(net1150));
 sg13g2_antennanp ANTENNA_1417 (.A(net1150));
 sg13g2_antennanp ANTENNA_1418 (.A(net1150));
 sg13g2_antennanp ANTENNA_1419 (.A(net1150));
 sg13g2_antennanp ANTENNA_1420 (.A(net1150));
 sg13g2_antennanp ANTENNA_1421 (.A(net1150));
 sg13g2_antennanp ANTENNA_1422 (.A(net1150));
 sg13g2_antennanp ANTENNA_1423 (.A(net1150));
 sg13g2_antennanp ANTENNA_1424 (.A(_00000_));
 sg13g2_antennanp ANTENNA_1425 (.A(_00000_));
 sg13g2_antennanp ANTENNA_1426 (.A(_00230_));
 sg13g2_antennanp ANTENNA_1427 (.A(_00752_));
 sg13g2_antennanp ANTENNA_1428 (.A(_00800_));
 sg13g2_antennanp ANTENNA_1429 (.A(_00800_));
 sg13g2_antennanp ANTENNA_1430 (.A(_01063_));
 sg13g2_antennanp ANTENNA_1431 (.A(_01066_));
 sg13g2_antennanp ANTENNA_1432 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1433 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1434 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1435 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1436 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1437 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1438 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1439 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1440 (.A(_02909_));
 sg13g2_antennanp ANTENNA_1441 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1442 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1443 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1444 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1445 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1446 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1447 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1448 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1449 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1450 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1451 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1452 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1453 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1454 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1455 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1456 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1457 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1458 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1459 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1460 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1461 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1462 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1463 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1464 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1465 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1466 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1467 (.A(_02933_));
 sg13g2_antennanp ANTENNA_1468 (.A(_03020_));
 sg13g2_antennanp ANTENNA_1469 (.A(_03020_));
 sg13g2_antennanp ANTENNA_1470 (.A(_03020_));
 sg13g2_antennanp ANTENNA_1471 (.A(_03161_));
 sg13g2_antennanp ANTENNA_1472 (.A(_03161_));
 sg13g2_antennanp ANTENNA_1473 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1474 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1475 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1476 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1477 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1478 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1479 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1480 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1481 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1482 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1483 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1484 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1485 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1486 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1487 (.A(_04843_));
 sg13g2_antennanp ANTENNA_1488 (.A(_04890_));
 sg13g2_antennanp ANTENNA_1489 (.A(_04890_));
 sg13g2_antennanp ANTENNA_1490 (.A(_04890_));
 sg13g2_antennanp ANTENNA_1491 (.A(_04890_));
 sg13g2_antennanp ANTENNA_1492 (.A(_04914_));
 sg13g2_antennanp ANTENNA_1493 (.A(_04954_));
 sg13g2_antennanp ANTENNA_1494 (.A(_05005_));
 sg13g2_antennanp ANTENNA_1495 (.A(_05175_));
 sg13g2_antennanp ANTENNA_1496 (.A(_05231_));
 sg13g2_antennanp ANTENNA_1497 (.A(_05267_));
 sg13g2_antennanp ANTENNA_1498 (.A(_05282_));
 sg13g2_antennanp ANTENNA_1499 (.A(_05293_));
 sg13g2_antennanp ANTENNA_1500 (.A(_05293_));
 sg13g2_antennanp ANTENNA_1501 (.A(_05293_));
 sg13g2_antennanp ANTENNA_1502 (.A(_05373_));
 sg13g2_antennanp ANTENNA_1503 (.A(_05437_));
 sg13g2_antennanp ANTENNA_1504 (.A(_05437_));
 sg13g2_antennanp ANTENNA_1505 (.A(_05577_));
 sg13g2_antennanp ANTENNA_1506 (.A(_05649_));
 sg13g2_antennanp ANTENNA_1507 (.A(_05722_));
 sg13g2_antennanp ANTENNA_1508 (.A(_05737_));
 sg13g2_antennanp ANTENNA_1509 (.A(_05783_));
 sg13g2_antennanp ANTENNA_1510 (.A(_05787_));
 sg13g2_antennanp ANTENNA_1511 (.A(_05787_));
 sg13g2_antennanp ANTENNA_1512 (.A(_05789_));
 sg13g2_antennanp ANTENNA_1513 (.A(_05792_));
 sg13g2_antennanp ANTENNA_1514 (.A(_05795_));
 sg13g2_antennanp ANTENNA_1515 (.A(_05800_));
 sg13g2_antennanp ANTENNA_1516 (.A(_05800_));
 sg13g2_antennanp ANTENNA_1517 (.A(_05800_));
 sg13g2_antennanp ANTENNA_1518 (.A(_05838_));
 sg13g2_antennanp ANTENNA_1519 (.A(_05838_));
 sg13g2_antennanp ANTENNA_1520 (.A(_05838_));
 sg13g2_antennanp ANTENNA_1521 (.A(_06038_));
 sg13g2_antennanp ANTENNA_1522 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1523 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1524 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1525 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1526 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1527 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1528 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1529 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1530 (.A(_06479_));
 sg13g2_antennanp ANTENNA_1531 (.A(_06822_));
 sg13g2_antennanp ANTENNA_1532 (.A(_06856_));
 sg13g2_antennanp ANTENNA_1533 (.A(_06905_));
 sg13g2_antennanp ANTENNA_1534 (.A(_06978_));
 sg13g2_antennanp ANTENNA_1535 (.A(_08377_));
 sg13g2_antennanp ANTENNA_1536 (.A(_08377_));
 sg13g2_antennanp ANTENNA_1537 (.A(_08377_));
 sg13g2_antennanp ANTENNA_1538 (.A(_08411_));
 sg13g2_antennanp ANTENNA_1539 (.A(_08411_));
 sg13g2_antennanp ANTENNA_1540 (.A(_08411_));
 sg13g2_antennanp ANTENNA_1541 (.A(_08411_));
 sg13g2_antennanp ANTENNA_1542 (.A(_08443_));
 sg13g2_antennanp ANTENNA_1543 (.A(_08443_));
 sg13g2_antennanp ANTENNA_1544 (.A(_08443_));
 sg13g2_antennanp ANTENNA_1545 (.A(_08486_));
 sg13g2_antennanp ANTENNA_1546 (.A(_08556_));
 sg13g2_antennanp ANTENNA_1547 (.A(_08556_));
 sg13g2_antennanp ANTENNA_1548 (.A(_08556_));
 sg13g2_antennanp ANTENNA_1549 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1550 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1551 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1552 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1553 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1554 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1555 (.A(_08669_));
 sg13g2_antennanp ANTENNA_1556 (.A(_08804_));
 sg13g2_antennanp ANTENNA_1557 (.A(_08839_));
 sg13g2_antennanp ANTENNA_1558 (.A(_08839_));
 sg13g2_antennanp ANTENNA_1559 (.A(_08839_));
 sg13g2_antennanp ANTENNA_1560 (.A(_08940_));
 sg13g2_antennanp ANTENNA_1561 (.A(_08940_));
 sg13g2_antennanp ANTENNA_1562 (.A(_08976_));
 sg13g2_antennanp ANTENNA_1563 (.A(_09068_));
 sg13g2_antennanp ANTENNA_1564 (.A(_09225_));
 sg13g2_antennanp ANTENNA_1565 (.A(_09225_));
 sg13g2_antennanp ANTENNA_1566 (.A(_09225_));
 sg13g2_antennanp ANTENNA_1567 (.A(_09225_));
 sg13g2_antennanp ANTENNA_1568 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1569 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1570 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1571 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1572 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1573 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1574 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1575 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1576 (.A(_09240_));
 sg13g2_antennanp ANTENNA_1577 (.A(_09282_));
 sg13g2_antennanp ANTENNA_1578 (.A(_09282_));
 sg13g2_antennanp ANTENNA_1579 (.A(_09282_));
 sg13g2_antennanp ANTENNA_1580 (.A(_09282_));
 sg13g2_antennanp ANTENNA_1581 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1582 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1583 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1584 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1585 (.A(_09310_));
 sg13g2_antennanp ANTENNA_1586 (.A(_09310_));
 sg13g2_antennanp ANTENNA_1587 (.A(_09310_));
 sg13g2_antennanp ANTENNA_1588 (.A(_09363_));
 sg13g2_antennanp ANTENNA_1589 (.A(_09363_));
 sg13g2_antennanp ANTENNA_1590 (.A(_09363_));
 sg13g2_antennanp ANTENNA_1591 (.A(_09435_));
 sg13g2_antennanp ANTENNA_1592 (.A(_09435_));
 sg13g2_antennanp ANTENNA_1593 (.A(_09435_));
 sg13g2_antennanp ANTENNA_1594 (.A(_09512_));
 sg13g2_antennanp ANTENNA_1595 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1596 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1597 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1598 (.A(_09558_));
 sg13g2_antennanp ANTENNA_1599 (.A(_09588_));
 sg13g2_antennanp ANTENNA_1600 (.A(_09639_));
 sg13g2_antennanp ANTENNA_1601 (.A(_09639_));
 sg13g2_antennanp ANTENNA_1602 (.A(_09700_));
 sg13g2_antennanp ANTENNA_1603 (.A(_09854_));
 sg13g2_antennanp ANTENNA_1604 (.A(_09897_));
 sg13g2_antennanp ANTENNA_1605 (.A(_09897_));
 sg13g2_antennanp ANTENNA_1606 (.A(_09899_));
 sg13g2_antennanp ANTENNA_1607 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1608 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1609 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1610 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1611 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1612 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1613 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1614 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1615 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1616 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1617 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1618 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1619 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1620 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1621 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1622 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1623 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1624 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1625 (.A(_10137_));
 sg13g2_antennanp ANTENNA_1626 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1627 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1628 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1629 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1630 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1631 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1632 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1633 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1634 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1635 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1636 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1637 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1638 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1639 (.A(_10210_));
 sg13g2_antennanp ANTENNA_1640 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1641 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1642 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1643 (.A(_10383_));
 sg13g2_antennanp ANTENNA_1644 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1645 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1646 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1647 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1648 (.A(_10721_));
 sg13g2_antennanp ANTENNA_1649 (.A(_11086_));
 sg13g2_antennanp ANTENNA_1650 (.A(_11086_));
 sg13g2_antennanp ANTENNA_1651 (.A(_11086_));
 sg13g2_antennanp ANTENNA_1652 (.A(_11086_));
 sg13g2_antennanp ANTENNA_1653 (.A(_11086_));
 sg13g2_antennanp ANTENNA_1654 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1655 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1656 (.A(_12000_));
 sg13g2_antennanp ANTENNA_1657 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1658 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1659 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1660 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1661 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1662 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1663 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1664 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1665 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1666 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1667 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1668 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1669 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1670 (.A(_12010_));
 sg13g2_antennanp ANTENNA_1671 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1672 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1673 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1674 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1675 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1676 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1677 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1678 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1679 (.A(_12052_));
 sg13g2_antennanp ANTENNA_1680 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1681 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1682 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1683 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1684 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1685 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1686 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1687 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1688 (.A(_12087_));
 sg13g2_antennanp ANTENNA_1689 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1690 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1691 (.A(_12201_));
 sg13g2_antennanp ANTENNA_1692 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1693 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1694 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1695 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1696 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1697 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1698 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1699 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1700 (.A(_12209_));
 sg13g2_antennanp ANTENNA_1701 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1702 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1703 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1704 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1705 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1706 (.A(_12216_));
 sg13g2_antennanp ANTENNA_1707 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1708 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1709 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1710 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1711 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1712 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1713 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1714 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1715 (.A(_12220_));
 sg13g2_antennanp ANTENNA_1716 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1717 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1718 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1719 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1720 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1721 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1722 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1723 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1724 (.A(_12227_));
 sg13g2_antennanp ANTENNA_1725 (.A(clk));
 sg13g2_antennanp ANTENNA_1726 (.A(clk));
 sg13g2_antennanp ANTENNA_1727 (.A(\cpu.d_flush_all ));
 sg13g2_antennanp ANTENNA_1728 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1729 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_1730 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_1731 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1732 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1733 (.A(net1));
 sg13g2_antennanp ANTENNA_1734 (.A(net1));
 sg13g2_antennanp ANTENNA_1735 (.A(net1));
 sg13g2_antennanp ANTENNA_1736 (.A(net1));
 sg13g2_antennanp ANTENNA_1737 (.A(net1));
 sg13g2_antennanp ANTENNA_1738 (.A(net1));
 sg13g2_antennanp ANTENNA_1739 (.A(net1));
 sg13g2_antennanp ANTENNA_1740 (.A(net1));
 sg13g2_antennanp ANTENNA_1741 (.A(net3));
 sg13g2_antennanp ANTENNA_1742 (.A(net3));
 sg13g2_antennanp ANTENNA_1743 (.A(net11));
 sg13g2_antennanp ANTENNA_1744 (.A(net11));
 sg13g2_antennanp ANTENNA_1745 (.A(net12));
 sg13g2_antennanp ANTENNA_1746 (.A(net12));
 sg13g2_antennanp ANTENNA_1747 (.A(net14));
 sg13g2_antennanp ANTENNA_1748 (.A(net14));
 sg13g2_antennanp ANTENNA_1749 (.A(net484));
 sg13g2_antennanp ANTENNA_1750 (.A(net484));
 sg13g2_antennanp ANTENNA_1751 (.A(net484));
 sg13g2_antennanp ANTENNA_1752 (.A(net484));
 sg13g2_antennanp ANTENNA_1753 (.A(net484));
 sg13g2_antennanp ANTENNA_1754 (.A(net484));
 sg13g2_antennanp ANTENNA_1755 (.A(net484));
 sg13g2_antennanp ANTENNA_1756 (.A(net484));
 sg13g2_antennanp ANTENNA_1757 (.A(net484));
 sg13g2_antennanp ANTENNA_1758 (.A(net520));
 sg13g2_antennanp ANTENNA_1759 (.A(net520));
 sg13g2_antennanp ANTENNA_1760 (.A(net520));
 sg13g2_antennanp ANTENNA_1761 (.A(net520));
 sg13g2_antennanp ANTENNA_1762 (.A(net520));
 sg13g2_antennanp ANTENNA_1763 (.A(net520));
 sg13g2_antennanp ANTENNA_1764 (.A(net520));
 sg13g2_antennanp ANTENNA_1765 (.A(net520));
 sg13g2_antennanp ANTENNA_1766 (.A(net520));
 sg13g2_antennanp ANTENNA_1767 (.A(net520));
 sg13g2_antennanp ANTENNA_1768 (.A(net520));
 sg13g2_antennanp ANTENNA_1769 (.A(net520));
 sg13g2_antennanp ANTENNA_1770 (.A(net544));
 sg13g2_antennanp ANTENNA_1771 (.A(net544));
 sg13g2_antennanp ANTENNA_1772 (.A(net544));
 sg13g2_antennanp ANTENNA_1773 (.A(net544));
 sg13g2_antennanp ANTENNA_1774 (.A(net544));
 sg13g2_antennanp ANTENNA_1775 (.A(net544));
 sg13g2_antennanp ANTENNA_1776 (.A(net544));
 sg13g2_antennanp ANTENNA_1777 (.A(net544));
 sg13g2_antennanp ANTENNA_1778 (.A(net653));
 sg13g2_antennanp ANTENNA_1779 (.A(net653));
 sg13g2_antennanp ANTENNA_1780 (.A(net653));
 sg13g2_antennanp ANTENNA_1781 (.A(net653));
 sg13g2_antennanp ANTENNA_1782 (.A(net653));
 sg13g2_antennanp ANTENNA_1783 (.A(net653));
 sg13g2_antennanp ANTENNA_1784 (.A(net653));
 sg13g2_antennanp ANTENNA_1785 (.A(net653));
 sg13g2_antennanp ANTENNA_1786 (.A(net653));
 sg13g2_antennanp ANTENNA_1787 (.A(net797));
 sg13g2_antennanp ANTENNA_1788 (.A(net797));
 sg13g2_antennanp ANTENNA_1789 (.A(net797));
 sg13g2_antennanp ANTENNA_1790 (.A(net797));
 sg13g2_antennanp ANTENNA_1791 (.A(net797));
 sg13g2_antennanp ANTENNA_1792 (.A(net797));
 sg13g2_antennanp ANTENNA_1793 (.A(net797));
 sg13g2_antennanp ANTENNA_1794 (.A(net797));
 sg13g2_antennanp ANTENNA_1795 (.A(net797));
 sg13g2_antennanp ANTENNA_1796 (.A(net797));
 sg13g2_antennanp ANTENNA_1797 (.A(net797));
 sg13g2_antennanp ANTENNA_1798 (.A(net797));
 sg13g2_antennanp ANTENNA_1799 (.A(net797));
 sg13g2_antennanp ANTENNA_1800 (.A(net797));
 sg13g2_antennanp ANTENNA_1801 (.A(net797));
 sg13g2_antennanp ANTENNA_1802 (.A(net797));
 sg13g2_antennanp ANTENNA_1803 (.A(net797));
 sg13g2_antennanp ANTENNA_1804 (.A(net797));
 sg13g2_antennanp ANTENNA_1805 (.A(net861));
 sg13g2_antennanp ANTENNA_1806 (.A(net861));
 sg13g2_antennanp ANTENNA_1807 (.A(net861));
 sg13g2_antennanp ANTENNA_1808 (.A(net861));
 sg13g2_antennanp ANTENNA_1809 (.A(net861));
 sg13g2_antennanp ANTENNA_1810 (.A(net861));
 sg13g2_antennanp ANTENNA_1811 (.A(net861));
 sg13g2_antennanp ANTENNA_1812 (.A(net861));
 sg13g2_antennanp ANTENNA_1813 (.A(net861));
 sg13g2_antennanp ANTENNA_1814 (.A(net861));
 sg13g2_antennanp ANTENNA_1815 (.A(net861));
 sg13g2_antennanp ANTENNA_1816 (.A(net861));
 sg13g2_antennanp ANTENNA_1817 (.A(net861));
 sg13g2_antennanp ANTENNA_1818 (.A(net861));
 sg13g2_antennanp ANTENNA_1819 (.A(net861));
 sg13g2_antennanp ANTENNA_1820 (.A(net861));
 sg13g2_antennanp ANTENNA_1821 (.A(net862));
 sg13g2_antennanp ANTENNA_1822 (.A(net862));
 sg13g2_antennanp ANTENNA_1823 (.A(net862));
 sg13g2_antennanp ANTENNA_1824 (.A(net862));
 sg13g2_antennanp ANTENNA_1825 (.A(net862));
 sg13g2_antennanp ANTENNA_1826 (.A(net862));
 sg13g2_antennanp ANTENNA_1827 (.A(net862));
 sg13g2_antennanp ANTENNA_1828 (.A(net862));
 sg13g2_antennanp ANTENNA_1829 (.A(net862));
 sg13g2_antennanp ANTENNA_1830 (.A(net862));
 sg13g2_antennanp ANTENNA_1831 (.A(net862));
 sg13g2_antennanp ANTENNA_1832 (.A(net862));
 sg13g2_antennanp ANTENNA_1833 (.A(net862));
 sg13g2_antennanp ANTENNA_1834 (.A(net862));
 sg13g2_antennanp ANTENNA_1835 (.A(net862));
 sg13g2_antennanp ANTENNA_1836 (.A(net862));
 sg13g2_antennanp ANTENNA_1837 (.A(net862));
 sg13g2_antennanp ANTENNA_1838 (.A(net862));
 sg13g2_antennanp ANTENNA_1839 (.A(net862));
 sg13g2_antennanp ANTENNA_1840 (.A(net862));
 sg13g2_antennanp ANTENNA_1841 (.A(net862));
 sg13g2_antennanp ANTENNA_1842 (.A(net862));
 sg13g2_antennanp ANTENNA_1843 (.A(net862));
 sg13g2_antennanp ANTENNA_1844 (.A(net862));
 sg13g2_antennanp ANTENNA_1845 (.A(net862));
 sg13g2_antennanp ANTENNA_1846 (.A(net862));
 sg13g2_antennanp ANTENNA_1847 (.A(net862));
 sg13g2_antennanp ANTENNA_1848 (.A(net862));
 sg13g2_antennanp ANTENNA_1849 (.A(net862));
 sg13g2_antennanp ANTENNA_1850 (.A(net907));
 sg13g2_antennanp ANTENNA_1851 (.A(net907));
 sg13g2_antennanp ANTENNA_1852 (.A(net907));
 sg13g2_antennanp ANTENNA_1853 (.A(net907));
 sg13g2_antennanp ANTENNA_1854 (.A(net907));
 sg13g2_antennanp ANTENNA_1855 (.A(net907));
 sg13g2_antennanp ANTENNA_1856 (.A(net907));
 sg13g2_antennanp ANTENNA_1857 (.A(net907));
 sg13g2_antennanp ANTENNA_1858 (.A(net916));
 sg13g2_antennanp ANTENNA_1859 (.A(net916));
 sg13g2_antennanp ANTENNA_1860 (.A(net916));
 sg13g2_antennanp ANTENNA_1861 (.A(net916));
 sg13g2_antennanp ANTENNA_1862 (.A(net916));
 sg13g2_antennanp ANTENNA_1863 (.A(net916));
 sg13g2_antennanp ANTENNA_1864 (.A(net916));
 sg13g2_antennanp ANTENNA_1865 (.A(net916));
 sg13g2_antennanp ANTENNA_1866 (.A(net916));
 sg13g2_antennanp ANTENNA_1867 (.A(net916));
 sg13g2_antennanp ANTENNA_1868 (.A(net916));
 sg13g2_antennanp ANTENNA_1869 (.A(net916));
 sg13g2_antennanp ANTENNA_1870 (.A(net916));
 sg13g2_antennanp ANTENNA_1871 (.A(net916));
 sg13g2_antennanp ANTENNA_1872 (.A(net916));
 sg13g2_antennanp ANTENNA_1873 (.A(net916));
 sg13g2_antennanp ANTENNA_1874 (.A(net916));
 sg13g2_antennanp ANTENNA_1875 (.A(net916));
 sg13g2_antennanp ANTENNA_1876 (.A(net916));
 sg13g2_antennanp ANTENNA_1877 (.A(net916));
 sg13g2_antennanp ANTENNA_1878 (.A(net916));
 sg13g2_antennanp ANTENNA_1879 (.A(net916));
 sg13g2_antennanp ANTENNA_1880 (.A(net916));
 sg13g2_antennanp ANTENNA_1881 (.A(net933));
 sg13g2_antennanp ANTENNA_1882 (.A(net933));
 sg13g2_antennanp ANTENNA_1883 (.A(net933));
 sg13g2_antennanp ANTENNA_1884 (.A(net933));
 sg13g2_antennanp ANTENNA_1885 (.A(net933));
 sg13g2_antennanp ANTENNA_1886 (.A(net933));
 sg13g2_antennanp ANTENNA_1887 (.A(net933));
 sg13g2_antennanp ANTENNA_1888 (.A(net933));
 sg13g2_antennanp ANTENNA_1889 (.A(net933));
 sg13g2_antennanp ANTENNA_1890 (.A(net993));
 sg13g2_antennanp ANTENNA_1891 (.A(net993));
 sg13g2_antennanp ANTENNA_1892 (.A(net993));
 sg13g2_antennanp ANTENNA_1893 (.A(net993));
 sg13g2_antennanp ANTENNA_1894 (.A(net993));
 sg13g2_antennanp ANTENNA_1895 (.A(net993));
 sg13g2_antennanp ANTENNA_1896 (.A(net993));
 sg13g2_antennanp ANTENNA_1897 (.A(net993));
 sg13g2_antennanp ANTENNA_1898 (.A(net993));
 sg13g2_antennanp ANTENNA_1899 (.A(net993));
 sg13g2_antennanp ANTENNA_1900 (.A(net993));
 sg13g2_antennanp ANTENNA_1901 (.A(net993));
 sg13g2_antennanp ANTENNA_1902 (.A(net993));
 sg13g2_antennanp ANTENNA_1903 (.A(net993));
 sg13g2_antennanp ANTENNA_1904 (.A(net993));
 sg13g2_antennanp ANTENNA_1905 (.A(net993));
 sg13g2_antennanp ANTENNA_1906 (.A(net993));
 sg13g2_antennanp ANTENNA_1907 (.A(net993));
 sg13g2_antennanp ANTENNA_1908 (.A(net993));
 sg13g2_antennanp ANTENNA_1909 (.A(net993));
 sg13g2_antennanp ANTENNA_1910 (.A(net993));
 sg13g2_antennanp ANTENNA_1911 (.A(net993));
 sg13g2_antennanp ANTENNA_1912 (.A(net993));
 sg13g2_antennanp ANTENNA_1913 (.A(net993));
 sg13g2_antennanp ANTENNA_1914 (.A(net993));
 sg13g2_antennanp ANTENNA_1915 (.A(net1020));
 sg13g2_antennanp ANTENNA_1916 (.A(net1020));
 sg13g2_antennanp ANTENNA_1917 (.A(net1020));
 sg13g2_antennanp ANTENNA_1918 (.A(net1020));
 sg13g2_antennanp ANTENNA_1919 (.A(net1020));
 sg13g2_antennanp ANTENNA_1920 (.A(net1020));
 sg13g2_antennanp ANTENNA_1921 (.A(net1020));
 sg13g2_antennanp ANTENNA_1922 (.A(net1020));
 sg13g2_antennanp ANTENNA_1923 (.A(net1020));
 sg13g2_antennanp ANTENNA_1924 (.A(net1020));
 sg13g2_antennanp ANTENNA_1925 (.A(net1020));
 sg13g2_antennanp ANTENNA_1926 (.A(net1020));
 sg13g2_antennanp ANTENNA_1927 (.A(net1020));
 sg13g2_antennanp ANTENNA_1928 (.A(net1020));
 sg13g2_antennanp ANTENNA_1929 (.A(net1020));
 sg13g2_antennanp ANTENNA_1930 (.A(net1020));
 sg13g2_antennanp ANTENNA_1931 (.A(net1020));
 sg13g2_antennanp ANTENNA_1932 (.A(net1020));
 sg13g2_antennanp ANTENNA_1933 (.A(net1020));
 sg13g2_antennanp ANTENNA_1934 (.A(net1020));
 sg13g2_antennanp ANTENNA_1935 (.A(net1021));
 sg13g2_antennanp ANTENNA_1936 (.A(net1021));
 sg13g2_antennanp ANTENNA_1937 (.A(net1021));
 sg13g2_antennanp ANTENNA_1938 (.A(net1021));
 sg13g2_antennanp ANTENNA_1939 (.A(net1021));
 sg13g2_antennanp ANTENNA_1940 (.A(net1021));
 sg13g2_antennanp ANTENNA_1941 (.A(net1021));
 sg13g2_antennanp ANTENNA_1942 (.A(net1021));
 sg13g2_antennanp ANTENNA_1943 (.A(net1021));
 sg13g2_antennanp ANTENNA_1944 (.A(net1066));
 sg13g2_antennanp ANTENNA_1945 (.A(net1066));
 sg13g2_antennanp ANTENNA_1946 (.A(net1066));
 sg13g2_antennanp ANTENNA_1947 (.A(net1066));
 sg13g2_antennanp ANTENNA_1948 (.A(net1066));
 sg13g2_antennanp ANTENNA_1949 (.A(net1066));
 sg13g2_antennanp ANTENNA_1950 (.A(net1066));
 sg13g2_antennanp ANTENNA_1951 (.A(net1066));
 sg13g2_antennanp ANTENNA_1952 (.A(net1066));
 sg13g2_antennanp ANTENNA_1953 (.A(net1066));
 sg13g2_antennanp ANTENNA_1954 (.A(net1066));
 sg13g2_antennanp ANTENNA_1955 (.A(net1066));
 sg13g2_antennanp ANTENNA_1956 (.A(net1066));
 sg13g2_antennanp ANTENNA_1957 (.A(net1066));
 sg13g2_antennanp ANTENNA_1958 (.A(net1066));
 sg13g2_antennanp ANTENNA_1959 (.A(net1069));
 sg13g2_antennanp ANTENNA_1960 (.A(net1069));
 sg13g2_antennanp ANTENNA_1961 (.A(net1069));
 sg13g2_antennanp ANTENNA_1962 (.A(net1069));
 sg13g2_antennanp ANTENNA_1963 (.A(net1069));
 sg13g2_antennanp ANTENNA_1964 (.A(net1069));
 sg13g2_antennanp ANTENNA_1965 (.A(net1069));
 sg13g2_antennanp ANTENNA_1966 (.A(net1069));
 sg13g2_antennanp ANTENNA_1967 (.A(net1070));
 sg13g2_antennanp ANTENNA_1968 (.A(net1070));
 sg13g2_antennanp ANTENNA_1969 (.A(net1070));
 sg13g2_antennanp ANTENNA_1970 (.A(net1070));
 sg13g2_antennanp ANTENNA_1971 (.A(net1070));
 sg13g2_antennanp ANTENNA_1972 (.A(net1070));
 sg13g2_antennanp ANTENNA_1973 (.A(net1070));
 sg13g2_antennanp ANTENNA_1974 (.A(net1070));
 sg13g2_antennanp ANTENNA_1975 (.A(net1071));
 sg13g2_antennanp ANTENNA_1976 (.A(net1071));
 sg13g2_antennanp ANTENNA_1977 (.A(net1071));
 sg13g2_antennanp ANTENNA_1978 (.A(net1071));
 sg13g2_antennanp ANTENNA_1979 (.A(net1071));
 sg13g2_antennanp ANTENNA_1980 (.A(net1071));
 sg13g2_antennanp ANTENNA_1981 (.A(net1071));
 sg13g2_antennanp ANTENNA_1982 (.A(net1071));
 sg13g2_antennanp ANTENNA_1983 (.A(net1071));
 sg13g2_antennanp ANTENNA_1984 (.A(net1109));
 sg13g2_antennanp ANTENNA_1985 (.A(net1109));
 sg13g2_antennanp ANTENNA_1986 (.A(net1109));
 sg13g2_antennanp ANTENNA_1987 (.A(net1109));
 sg13g2_antennanp ANTENNA_1988 (.A(net1109));
 sg13g2_antennanp ANTENNA_1989 (.A(net1109));
 sg13g2_antennanp ANTENNA_1990 (.A(net1109));
 sg13g2_antennanp ANTENNA_1991 (.A(net1109));
 sg13g2_antennanp ANTENNA_1992 (.A(net1109));
 sg13g2_antennanp ANTENNA_1993 (.A(net1109));
 sg13g2_antennanp ANTENNA_1994 (.A(net1109));
 sg13g2_antennanp ANTENNA_1995 (.A(net1109));
 sg13g2_antennanp ANTENNA_1996 (.A(net1109));
 sg13g2_antennanp ANTENNA_1997 (.A(net1109));
 sg13g2_antennanp ANTENNA_1998 (.A(net1109));
 sg13g2_antennanp ANTENNA_1999 (.A(net1109));
 sg13g2_antennanp ANTENNA_2000 (.A(net1109));
 sg13g2_antennanp ANTENNA_2001 (.A(net1109));
 sg13g2_antennanp ANTENNA_2002 (.A(net1109));
 sg13g2_antennanp ANTENNA_2003 (.A(net1109));
 sg13g2_antennanp ANTENNA_2004 (.A(net1109));
 sg13g2_antennanp ANTENNA_2005 (.A(net1109));
 sg13g2_antennanp ANTENNA_2006 (.A(net1109));
 sg13g2_antennanp ANTENNA_2007 (.A(net1109));
 sg13g2_antennanp ANTENNA_2008 (.A(net1109));
 sg13g2_antennanp ANTENNA_2009 (.A(net1109));
 sg13g2_antennanp ANTENNA_2010 (.A(net1109));
 sg13g2_antennanp ANTENNA_2011 (.A(net1109));
 sg13g2_antennanp ANTENNA_2012 (.A(net1109));
 sg13g2_antennanp ANTENNA_2013 (.A(net1109));
 sg13g2_antennanp ANTENNA_2014 (.A(net1150));
 sg13g2_antennanp ANTENNA_2015 (.A(net1150));
 sg13g2_antennanp ANTENNA_2016 (.A(net1150));
 sg13g2_antennanp ANTENNA_2017 (.A(net1150));
 sg13g2_antennanp ANTENNA_2018 (.A(net1150));
 sg13g2_antennanp ANTENNA_2019 (.A(net1150));
 sg13g2_antennanp ANTENNA_2020 (.A(net1150));
 sg13g2_antennanp ANTENNA_2021 (.A(net1150));
 sg13g2_antennanp ANTENNA_2022 (.A(net1150));
 sg13g2_antennanp ANTENNA_2023 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2024 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2025 (.A(_00230_));
 sg13g2_antennanp ANTENNA_2026 (.A(_00752_));
 sg13g2_antennanp ANTENNA_2027 (.A(_00800_));
 sg13g2_antennanp ANTENNA_2028 (.A(_00800_));
 sg13g2_antennanp ANTENNA_2029 (.A(_01063_));
 sg13g2_antennanp ANTENNA_2030 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2031 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2032 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2033 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2034 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2035 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2036 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2037 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2038 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2039 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2040 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2041 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2042 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2043 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2044 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2045 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2046 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2047 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2048 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2049 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2050 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2051 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2052 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2053 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2054 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2055 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2056 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2057 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2058 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2059 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2060 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2061 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2062 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2063 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2064 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2065 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2066 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2067 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2068 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2069 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2070 (.A(_03161_));
 sg13g2_antennanp ANTENNA_2071 (.A(_03161_));
 sg13g2_antennanp ANTENNA_2072 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2073 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2074 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2075 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2076 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2077 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2078 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2079 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2080 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2081 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2082 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2083 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2084 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2085 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2086 (.A(_04843_));
 sg13g2_antennanp ANTENNA_2087 (.A(_04914_));
 sg13g2_antennanp ANTENNA_2088 (.A(_04954_));
 sg13g2_antennanp ANTENNA_2089 (.A(_05005_));
 sg13g2_antennanp ANTENNA_2090 (.A(_05175_));
 sg13g2_antennanp ANTENNA_2091 (.A(_05207_));
 sg13g2_antennanp ANTENNA_2092 (.A(_05231_));
 sg13g2_antennanp ANTENNA_2093 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2094 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2095 (.A(_05282_));
 sg13g2_antennanp ANTENNA_2096 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2097 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2098 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2099 (.A(_05373_));
 sg13g2_antennanp ANTENNA_2100 (.A(_05577_));
 sg13g2_antennanp ANTENNA_2101 (.A(_05649_));
 sg13g2_antennanp ANTENNA_2102 (.A(_05722_));
 sg13g2_antennanp ANTENNA_2103 (.A(_05737_));
 sg13g2_antennanp ANTENNA_2104 (.A(_05783_));
 sg13g2_antennanp ANTENNA_2105 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2106 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2107 (.A(_05789_));
 sg13g2_antennanp ANTENNA_2108 (.A(_05792_));
 sg13g2_antennanp ANTENNA_2109 (.A(_05795_));
 sg13g2_antennanp ANTENNA_2110 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2111 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2112 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2113 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2114 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2115 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2116 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2117 (.A(_06038_));
 sg13g2_antennanp ANTENNA_2118 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2119 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2120 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2121 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2122 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2123 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2124 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2125 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2126 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2127 (.A(_06822_));
 sg13g2_antennanp ANTENNA_2128 (.A(_06856_));
 sg13g2_antennanp ANTENNA_2129 (.A(_06905_));
 sg13g2_antennanp ANTENNA_2130 (.A(_06978_));
 sg13g2_antennanp ANTENNA_2131 (.A(_08220_));
 sg13g2_antennanp ANTENNA_2132 (.A(_08220_));
 sg13g2_antennanp ANTENNA_2133 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2134 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2135 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2136 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2137 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2138 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2139 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2140 (.A(_08443_));
 sg13g2_antennanp ANTENNA_2141 (.A(_08443_));
 sg13g2_antennanp ANTENNA_2142 (.A(_08443_));
 sg13g2_antennanp ANTENNA_2143 (.A(_08486_));
 sg13g2_antennanp ANTENNA_2144 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2145 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2146 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2147 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2148 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2149 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2150 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2151 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2152 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2153 (.A(_08669_));
 sg13g2_antennanp ANTENNA_2154 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2155 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2156 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2157 (.A(_08804_));
 sg13g2_antennanp ANTENNA_2158 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2159 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2160 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2161 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2162 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2163 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2164 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2165 (.A(_08940_));
 sg13g2_antennanp ANTENNA_2166 (.A(_08940_));
 sg13g2_antennanp ANTENNA_2167 (.A(_08976_));
 sg13g2_antennanp ANTENNA_2168 (.A(_09068_));
 sg13g2_antennanp ANTENNA_2169 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2170 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2171 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2172 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2173 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2174 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2175 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2176 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2177 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2178 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2179 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2180 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2181 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2182 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2183 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2184 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2185 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2186 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2187 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2188 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2189 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2190 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2191 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2192 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2193 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2194 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2195 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2196 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2197 (.A(_09512_));
 sg13g2_antennanp ANTENNA_2198 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2199 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2200 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2201 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2202 (.A(_09588_));
 sg13g2_antennanp ANTENNA_2203 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2204 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2205 (.A(_09700_));
 sg13g2_antennanp ANTENNA_2206 (.A(_09854_));
 sg13g2_antennanp ANTENNA_2207 (.A(_09854_));
 sg13g2_antennanp ANTENNA_2208 (.A(_09897_));
 sg13g2_antennanp ANTENNA_2209 (.A(_09897_));
 sg13g2_antennanp ANTENNA_2210 (.A(_09899_));
 sg13g2_antennanp ANTENNA_2211 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2212 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2213 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2214 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2215 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2216 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2217 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2218 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2219 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2220 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2221 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2222 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2223 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2224 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2225 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2226 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2227 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2228 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2229 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2230 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2231 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2232 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2233 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2234 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2235 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2236 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2237 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2238 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2239 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2240 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2241 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2242 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2243 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2244 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2245 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2246 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2247 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2248 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2249 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2250 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2251 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2252 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2253 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2254 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2255 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2256 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2257 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2258 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2259 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2260 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2261 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2262 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2263 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2264 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2265 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2266 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2267 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2268 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2269 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2270 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2271 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2272 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2273 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2274 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2275 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2276 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2277 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2278 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2279 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2280 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2281 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2282 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2283 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2284 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2285 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2286 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2287 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2288 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2289 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2290 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2291 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2292 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2293 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2294 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2295 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2296 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2297 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2298 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2299 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2300 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2301 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2302 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2303 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2304 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2305 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2306 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2307 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2308 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2309 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2310 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2311 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2312 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2313 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2314 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2315 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2316 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2317 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2318 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2319 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2320 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2321 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2322 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2323 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2324 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2325 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2326 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2327 (.A(clk));
 sg13g2_antennanp ANTENNA_2328 (.A(clk));
 sg13g2_antennanp ANTENNA_2329 (.A(\cpu.d_flush_all ));
 sg13g2_antennanp ANTENNA_2330 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2331 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_2332 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_2333 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2334 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2335 (.A(net1));
 sg13g2_antennanp ANTENNA_2336 (.A(net1));
 sg13g2_antennanp ANTENNA_2337 (.A(net1));
 sg13g2_antennanp ANTENNA_2338 (.A(net1));
 sg13g2_antennanp ANTENNA_2339 (.A(net1));
 sg13g2_antennanp ANTENNA_2340 (.A(net1));
 sg13g2_antennanp ANTENNA_2341 (.A(net1));
 sg13g2_antennanp ANTENNA_2342 (.A(net1));
 sg13g2_antennanp ANTENNA_2343 (.A(net11));
 sg13g2_antennanp ANTENNA_2344 (.A(net11));
 sg13g2_antennanp ANTENNA_2345 (.A(net12));
 sg13g2_antennanp ANTENNA_2346 (.A(net12));
 sg13g2_antennanp ANTENNA_2347 (.A(net14));
 sg13g2_antennanp ANTENNA_2348 (.A(net14));
 sg13g2_antennanp ANTENNA_2349 (.A(net484));
 sg13g2_antennanp ANTENNA_2350 (.A(net484));
 sg13g2_antennanp ANTENNA_2351 (.A(net484));
 sg13g2_antennanp ANTENNA_2352 (.A(net484));
 sg13g2_antennanp ANTENNA_2353 (.A(net484));
 sg13g2_antennanp ANTENNA_2354 (.A(net484));
 sg13g2_antennanp ANTENNA_2355 (.A(net484));
 sg13g2_antennanp ANTENNA_2356 (.A(net484));
 sg13g2_antennanp ANTENNA_2357 (.A(net484));
 sg13g2_antennanp ANTENNA_2358 (.A(net544));
 sg13g2_antennanp ANTENNA_2359 (.A(net544));
 sg13g2_antennanp ANTENNA_2360 (.A(net544));
 sg13g2_antennanp ANTENNA_2361 (.A(net544));
 sg13g2_antennanp ANTENNA_2362 (.A(net544));
 sg13g2_antennanp ANTENNA_2363 (.A(net544));
 sg13g2_antennanp ANTENNA_2364 (.A(net544));
 sg13g2_antennanp ANTENNA_2365 (.A(net544));
 sg13g2_antennanp ANTENNA_2366 (.A(net653));
 sg13g2_antennanp ANTENNA_2367 (.A(net653));
 sg13g2_antennanp ANTENNA_2368 (.A(net653));
 sg13g2_antennanp ANTENNA_2369 (.A(net653));
 sg13g2_antennanp ANTENNA_2370 (.A(net653));
 sg13g2_antennanp ANTENNA_2371 (.A(net653));
 sg13g2_antennanp ANTENNA_2372 (.A(net653));
 sg13g2_antennanp ANTENNA_2373 (.A(net653));
 sg13g2_antennanp ANTENNA_2374 (.A(net653));
 sg13g2_antennanp ANTENNA_2375 (.A(net797));
 sg13g2_antennanp ANTENNA_2376 (.A(net797));
 sg13g2_antennanp ANTENNA_2377 (.A(net797));
 sg13g2_antennanp ANTENNA_2378 (.A(net797));
 sg13g2_antennanp ANTENNA_2379 (.A(net797));
 sg13g2_antennanp ANTENNA_2380 (.A(net797));
 sg13g2_antennanp ANTENNA_2381 (.A(net797));
 sg13g2_antennanp ANTENNA_2382 (.A(net797));
 sg13g2_antennanp ANTENNA_2383 (.A(net797));
 sg13g2_antennanp ANTENNA_2384 (.A(net797));
 sg13g2_antennanp ANTENNA_2385 (.A(net797));
 sg13g2_antennanp ANTENNA_2386 (.A(net797));
 sg13g2_antennanp ANTENNA_2387 (.A(net797));
 sg13g2_antennanp ANTENNA_2388 (.A(net797));
 sg13g2_antennanp ANTENNA_2389 (.A(net797));
 sg13g2_antennanp ANTENNA_2390 (.A(net797));
 sg13g2_antennanp ANTENNA_2391 (.A(net797));
 sg13g2_antennanp ANTENNA_2392 (.A(net861));
 sg13g2_antennanp ANTENNA_2393 (.A(net861));
 sg13g2_antennanp ANTENNA_2394 (.A(net861));
 sg13g2_antennanp ANTENNA_2395 (.A(net861));
 sg13g2_antennanp ANTENNA_2396 (.A(net861));
 sg13g2_antennanp ANTENNA_2397 (.A(net861));
 sg13g2_antennanp ANTENNA_2398 (.A(net861));
 sg13g2_antennanp ANTENNA_2399 (.A(net861));
 sg13g2_antennanp ANTENNA_2400 (.A(net861));
 sg13g2_antennanp ANTENNA_2401 (.A(net861));
 sg13g2_antennanp ANTENNA_2402 (.A(net861));
 sg13g2_antennanp ANTENNA_2403 (.A(net861));
 sg13g2_antennanp ANTENNA_2404 (.A(net861));
 sg13g2_antennanp ANTENNA_2405 (.A(net861));
 sg13g2_antennanp ANTENNA_2406 (.A(net861));
 sg13g2_antennanp ANTENNA_2407 (.A(net861));
 sg13g2_antennanp ANTENNA_2408 (.A(net861));
 sg13g2_antennanp ANTENNA_2409 (.A(net861));
 sg13g2_antennanp ANTENNA_2410 (.A(net861));
 sg13g2_antennanp ANTENNA_2411 (.A(net861));
 sg13g2_antennanp ANTENNA_2412 (.A(net861));
 sg13g2_antennanp ANTENNA_2413 (.A(net861));
 sg13g2_antennanp ANTENNA_2414 (.A(net861));
 sg13g2_antennanp ANTENNA_2415 (.A(net861));
 sg13g2_antennanp ANTENNA_2416 (.A(net916));
 sg13g2_antennanp ANTENNA_2417 (.A(net916));
 sg13g2_antennanp ANTENNA_2418 (.A(net916));
 sg13g2_antennanp ANTENNA_2419 (.A(net916));
 sg13g2_antennanp ANTENNA_2420 (.A(net916));
 sg13g2_antennanp ANTENNA_2421 (.A(net916));
 sg13g2_antennanp ANTENNA_2422 (.A(net916));
 sg13g2_antennanp ANTENNA_2423 (.A(net916));
 sg13g2_antennanp ANTENNA_2424 (.A(net916));
 sg13g2_antennanp ANTENNA_2425 (.A(net916));
 sg13g2_antennanp ANTENNA_2426 (.A(net916));
 sg13g2_antennanp ANTENNA_2427 (.A(net916));
 sg13g2_antennanp ANTENNA_2428 (.A(net916));
 sg13g2_antennanp ANTENNA_2429 (.A(net916));
 sg13g2_antennanp ANTENNA_2430 (.A(net916));
 sg13g2_antennanp ANTENNA_2431 (.A(net916));
 sg13g2_antennanp ANTENNA_2432 (.A(net993));
 sg13g2_antennanp ANTENNA_2433 (.A(net993));
 sg13g2_antennanp ANTENNA_2434 (.A(net993));
 sg13g2_antennanp ANTENNA_2435 (.A(net993));
 sg13g2_antennanp ANTENNA_2436 (.A(net993));
 sg13g2_antennanp ANTENNA_2437 (.A(net993));
 sg13g2_antennanp ANTENNA_2438 (.A(net993));
 sg13g2_antennanp ANTENNA_2439 (.A(net993));
 sg13g2_antennanp ANTENNA_2440 (.A(net993));
 sg13g2_antennanp ANTENNA_2441 (.A(net993));
 sg13g2_antennanp ANTENNA_2442 (.A(net993));
 sg13g2_antennanp ANTENNA_2443 (.A(net993));
 sg13g2_antennanp ANTENNA_2444 (.A(net993));
 sg13g2_antennanp ANTENNA_2445 (.A(net993));
 sg13g2_antennanp ANTENNA_2446 (.A(net993));
 sg13g2_antennanp ANTENNA_2447 (.A(net993));
 sg13g2_antennanp ANTENNA_2448 (.A(net993));
 sg13g2_antennanp ANTENNA_2449 (.A(net993));
 sg13g2_antennanp ANTENNA_2450 (.A(net993));
 sg13g2_antennanp ANTENNA_2451 (.A(net993));
 sg13g2_antennanp ANTENNA_2452 (.A(net993));
 sg13g2_antennanp ANTENNA_2453 (.A(net993));
 sg13g2_antennanp ANTENNA_2454 (.A(net993));
 sg13g2_antennanp ANTENNA_2455 (.A(net993));
 sg13g2_antennanp ANTENNA_2456 (.A(net993));
 sg13g2_antennanp ANTENNA_2457 (.A(net1066));
 sg13g2_antennanp ANTENNA_2458 (.A(net1066));
 sg13g2_antennanp ANTENNA_2459 (.A(net1066));
 sg13g2_antennanp ANTENNA_2460 (.A(net1066));
 sg13g2_antennanp ANTENNA_2461 (.A(net1066));
 sg13g2_antennanp ANTENNA_2462 (.A(net1066));
 sg13g2_antennanp ANTENNA_2463 (.A(net1066));
 sg13g2_antennanp ANTENNA_2464 (.A(net1066));
 sg13g2_antennanp ANTENNA_2465 (.A(net1066));
 sg13g2_antennanp ANTENNA_2466 (.A(net1069));
 sg13g2_antennanp ANTENNA_2467 (.A(net1069));
 sg13g2_antennanp ANTENNA_2468 (.A(net1069));
 sg13g2_antennanp ANTENNA_2469 (.A(net1069));
 sg13g2_antennanp ANTENNA_2470 (.A(net1069));
 sg13g2_antennanp ANTENNA_2471 (.A(net1069));
 sg13g2_antennanp ANTENNA_2472 (.A(net1069));
 sg13g2_antennanp ANTENNA_2473 (.A(net1069));
 sg13g2_antennanp ANTENNA_2474 (.A(net1071));
 sg13g2_antennanp ANTENNA_2475 (.A(net1071));
 sg13g2_antennanp ANTENNA_2476 (.A(net1071));
 sg13g2_antennanp ANTENNA_2477 (.A(net1071));
 sg13g2_antennanp ANTENNA_2478 (.A(net1071));
 sg13g2_antennanp ANTENNA_2479 (.A(net1071));
 sg13g2_antennanp ANTENNA_2480 (.A(net1071));
 sg13g2_antennanp ANTENNA_2481 (.A(net1071));
 sg13g2_antennanp ANTENNA_2482 (.A(net1071));
 sg13g2_antennanp ANTENNA_2483 (.A(net1113));
 sg13g2_antennanp ANTENNA_2484 (.A(net1113));
 sg13g2_antennanp ANTENNA_2485 (.A(net1113));
 sg13g2_antennanp ANTENNA_2486 (.A(net1113));
 sg13g2_antennanp ANTENNA_2487 (.A(net1113));
 sg13g2_antennanp ANTENNA_2488 (.A(net1113));
 sg13g2_antennanp ANTENNA_2489 (.A(net1113));
 sg13g2_antennanp ANTENNA_2490 (.A(net1113));
 sg13g2_antennanp ANTENNA_2491 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2492 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2493 (.A(_00230_));
 sg13g2_antennanp ANTENNA_2494 (.A(_00752_));
 sg13g2_antennanp ANTENNA_2495 (.A(_00800_));
 sg13g2_antennanp ANTENNA_2496 (.A(_00800_));
 sg13g2_antennanp ANTENNA_2497 (.A(_01063_));
 sg13g2_antennanp ANTENNA_2498 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2499 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2500 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2501 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2502 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2503 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2504 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2505 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2506 (.A(_02909_));
 sg13g2_antennanp ANTENNA_2507 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2508 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2509 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2510 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2511 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2512 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2513 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2514 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2515 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2516 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2517 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2518 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2519 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2520 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2521 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2522 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2523 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2524 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2525 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2526 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2527 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2528 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2529 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2530 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2531 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2532 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2533 (.A(_02933_));
 sg13g2_antennanp ANTENNA_2534 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2535 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2536 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2537 (.A(_03020_));
 sg13g2_antennanp ANTENNA_2538 (.A(_03161_));
 sg13g2_antennanp ANTENNA_2539 (.A(_03161_));
 sg13g2_antennanp ANTENNA_2540 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2541 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2542 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2543 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2544 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2545 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2546 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2547 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2548 (.A(_03535_));
 sg13g2_antennanp ANTENNA_2549 (.A(_04843_));
 sg13g2_antennanp ANTENNA_2550 (.A(_04914_));
 sg13g2_antennanp ANTENNA_2551 (.A(_04954_));
 sg13g2_antennanp ANTENNA_2552 (.A(_05005_));
 sg13g2_antennanp ANTENNA_2553 (.A(_05175_));
 sg13g2_antennanp ANTENNA_2554 (.A(_05207_));
 sg13g2_antennanp ANTENNA_2555 (.A(_05207_));
 sg13g2_antennanp ANTENNA_2556 (.A(_05231_));
 sg13g2_antennanp ANTENNA_2557 (.A(_05267_));
 sg13g2_antennanp ANTENNA_2558 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2559 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2560 (.A(_05293_));
 sg13g2_antennanp ANTENNA_2561 (.A(_05373_));
 sg13g2_antennanp ANTENNA_2562 (.A(_05577_));
 sg13g2_antennanp ANTENNA_2563 (.A(_05649_));
 sg13g2_antennanp ANTENNA_2564 (.A(_05722_));
 sg13g2_antennanp ANTENNA_2565 (.A(_05737_));
 sg13g2_antennanp ANTENNA_2566 (.A(_05783_));
 sg13g2_antennanp ANTENNA_2567 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2568 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2569 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2570 (.A(_05787_));
 sg13g2_antennanp ANTENNA_2571 (.A(_05789_));
 sg13g2_antennanp ANTENNA_2572 (.A(_05792_));
 sg13g2_antennanp ANTENNA_2573 (.A(_05795_));
 sg13g2_antennanp ANTENNA_2574 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2575 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2576 (.A(_05800_));
 sg13g2_antennanp ANTENNA_2577 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2578 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2579 (.A(_05838_));
 sg13g2_antennanp ANTENNA_2580 (.A(_06038_));
 sg13g2_antennanp ANTENNA_2581 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2582 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2583 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2584 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2585 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2586 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2587 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2588 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2589 (.A(_06479_));
 sg13g2_antennanp ANTENNA_2590 (.A(_06822_));
 sg13g2_antennanp ANTENNA_2591 (.A(_06856_));
 sg13g2_antennanp ANTENNA_2592 (.A(_06905_));
 sg13g2_antennanp ANTENNA_2593 (.A(_06978_));
 sg13g2_antennanp ANTENNA_2594 (.A(_08220_));
 sg13g2_antennanp ANTENNA_2595 (.A(_08220_));
 sg13g2_antennanp ANTENNA_2596 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2597 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2598 (.A(_08377_));
 sg13g2_antennanp ANTENNA_2599 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2600 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2601 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2602 (.A(_08411_));
 sg13g2_antennanp ANTENNA_2603 (.A(_08486_));
 sg13g2_antennanp ANTENNA_2604 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2605 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2606 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2607 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2608 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2609 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2610 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2611 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2612 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2613 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2614 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2615 (.A(_08691_));
 sg13g2_antennanp ANTENNA_2616 (.A(_08804_));
 sg13g2_antennanp ANTENNA_2617 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2618 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2619 (.A(_08839_));
 sg13g2_antennanp ANTENNA_2620 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2621 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2622 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2623 (.A(_08894_));
 sg13g2_antennanp ANTENNA_2624 (.A(_08940_));
 sg13g2_antennanp ANTENNA_2625 (.A(_08940_));
 sg13g2_antennanp ANTENNA_2626 (.A(_08976_));
 sg13g2_antennanp ANTENNA_2627 (.A(_09068_));
 sg13g2_antennanp ANTENNA_2628 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2629 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2630 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2631 (.A(_09225_));
 sg13g2_antennanp ANTENNA_2632 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2633 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2634 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2635 (.A(_09282_));
 sg13g2_antennanp ANTENNA_2636 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2637 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2638 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2639 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2640 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2641 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2642 (.A(_09310_));
 sg13g2_antennanp ANTENNA_2643 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2644 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2645 (.A(_09363_));
 sg13g2_antennanp ANTENNA_2646 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2647 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2648 (.A(_09435_));
 sg13g2_antennanp ANTENNA_2649 (.A(_09512_));
 sg13g2_antennanp ANTENNA_2650 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2651 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2652 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2653 (.A(_09558_));
 sg13g2_antennanp ANTENNA_2654 (.A(_09588_));
 sg13g2_antennanp ANTENNA_2655 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2656 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2657 (.A(_09700_));
 sg13g2_antennanp ANTENNA_2658 (.A(_09854_));
 sg13g2_antennanp ANTENNA_2659 (.A(_09897_));
 sg13g2_antennanp ANTENNA_2660 (.A(_09897_));
 sg13g2_antennanp ANTENNA_2661 (.A(_09899_));
 sg13g2_antennanp ANTENNA_2662 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2663 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2664 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2665 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2666 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2667 (.A(_10027_));
 sg13g2_antennanp ANTENNA_2668 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2669 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2670 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2671 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2672 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2673 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2674 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2675 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2676 (.A(_10137_));
 sg13g2_antennanp ANTENNA_2677 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2678 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2679 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2680 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2681 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2682 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2683 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2684 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2685 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2686 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2687 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2688 (.A(_10210_));
 sg13g2_antennanp ANTENNA_2689 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2690 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2691 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2692 (.A(_10383_));
 sg13g2_antennanp ANTENNA_2693 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2694 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2695 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2696 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2697 (.A(_10721_));
 sg13g2_antennanp ANTENNA_2698 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2699 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2700 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2701 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2702 (.A(_11086_));
 sg13g2_antennanp ANTENNA_2703 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2704 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2705 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2706 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2707 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2708 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2709 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2710 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2711 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2712 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2713 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2714 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2715 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2716 (.A(_12010_));
 sg13g2_antennanp ANTENNA_2717 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2718 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2719 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2720 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2721 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2722 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2723 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2724 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2725 (.A(_12052_));
 sg13g2_antennanp ANTENNA_2726 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2727 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2728 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2729 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2730 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2731 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2732 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2733 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2734 (.A(_12087_));
 sg13g2_antennanp ANTENNA_2735 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2736 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2737 (.A(_12201_));
 sg13g2_antennanp ANTENNA_2738 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2739 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2740 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2741 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2742 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2743 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2744 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2745 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2746 (.A(_12209_));
 sg13g2_antennanp ANTENNA_2747 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2748 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2749 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2750 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2751 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2752 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2753 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2754 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2755 (.A(_12216_));
 sg13g2_antennanp ANTENNA_2756 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2757 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2758 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2759 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2760 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2761 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2762 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2763 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2764 (.A(_12227_));
 sg13g2_antennanp ANTENNA_2765 (.A(\cpu.d_flush_all ));
 sg13g2_antennanp ANTENNA_2766 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2767 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_2768 (.A(\cpu.qspi.c_wstrobe_d ));
 sg13g2_antennanp ANTENNA_2769 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2770 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2771 (.A(net1));
 sg13g2_antennanp ANTENNA_2772 (.A(net1));
 sg13g2_antennanp ANTENNA_2773 (.A(net1));
 sg13g2_antennanp ANTENNA_2774 (.A(net1));
 sg13g2_antennanp ANTENNA_2775 (.A(net1));
 sg13g2_antennanp ANTENNA_2776 (.A(net1));
 sg13g2_antennanp ANTENNA_2777 (.A(net1));
 sg13g2_antennanp ANTENNA_2778 (.A(net1));
 sg13g2_antennanp ANTENNA_2779 (.A(net11));
 sg13g2_antennanp ANTENNA_2780 (.A(net11));
 sg13g2_antennanp ANTENNA_2781 (.A(net12));
 sg13g2_antennanp ANTENNA_2782 (.A(net12));
 sg13g2_antennanp ANTENNA_2783 (.A(net13));
 sg13g2_antennanp ANTENNA_2784 (.A(net13));
 sg13g2_antennanp ANTENNA_2785 (.A(net14));
 sg13g2_antennanp ANTENNA_2786 (.A(net14));
 sg13g2_antennanp ANTENNA_2787 (.A(net484));
 sg13g2_antennanp ANTENNA_2788 (.A(net484));
 sg13g2_antennanp ANTENNA_2789 (.A(net484));
 sg13g2_antennanp ANTENNA_2790 (.A(net484));
 sg13g2_antennanp ANTENNA_2791 (.A(net484));
 sg13g2_antennanp ANTENNA_2792 (.A(net484));
 sg13g2_antennanp ANTENNA_2793 (.A(net484));
 sg13g2_antennanp ANTENNA_2794 (.A(net484));
 sg13g2_antennanp ANTENNA_2795 (.A(net484));
 sg13g2_antennanp ANTENNA_2796 (.A(net544));
 sg13g2_antennanp ANTENNA_2797 (.A(net544));
 sg13g2_antennanp ANTENNA_2798 (.A(net544));
 sg13g2_antennanp ANTENNA_2799 (.A(net544));
 sg13g2_antennanp ANTENNA_2800 (.A(net544));
 sg13g2_antennanp ANTENNA_2801 (.A(net544));
 sg13g2_antennanp ANTENNA_2802 (.A(net544));
 sg13g2_antennanp ANTENNA_2803 (.A(net544));
 sg13g2_antennanp ANTENNA_2804 (.A(net797));
 sg13g2_antennanp ANTENNA_2805 (.A(net797));
 sg13g2_antennanp ANTENNA_2806 (.A(net797));
 sg13g2_antennanp ANTENNA_2807 (.A(net797));
 sg13g2_antennanp ANTENNA_2808 (.A(net797));
 sg13g2_antennanp ANTENNA_2809 (.A(net797));
 sg13g2_antennanp ANTENNA_2810 (.A(net797));
 sg13g2_antennanp ANTENNA_2811 (.A(net797));
 sg13g2_antennanp ANTENNA_2812 (.A(net797));
 sg13g2_antennanp ANTENNA_2813 (.A(net797));
 sg13g2_antennanp ANTENNA_2814 (.A(net797));
 sg13g2_antennanp ANTENNA_2815 (.A(net797));
 sg13g2_antennanp ANTENNA_2816 (.A(net797));
 sg13g2_antennanp ANTENNA_2817 (.A(net797));
 sg13g2_antennanp ANTENNA_2818 (.A(net797));
 sg13g2_antennanp ANTENNA_2819 (.A(net797));
 sg13g2_antennanp ANTENNA_2820 (.A(net797));
 sg13g2_antennanp ANTENNA_2821 (.A(net861));
 sg13g2_antennanp ANTENNA_2822 (.A(net861));
 sg13g2_antennanp ANTENNA_2823 (.A(net861));
 sg13g2_antennanp ANTENNA_2824 (.A(net861));
 sg13g2_antennanp ANTENNA_2825 (.A(net861));
 sg13g2_antennanp ANTENNA_2826 (.A(net861));
 sg13g2_antennanp ANTENNA_2827 (.A(net861));
 sg13g2_antennanp ANTENNA_2828 (.A(net861));
 sg13g2_antennanp ANTENNA_2829 (.A(net861));
 sg13g2_antennanp ANTENNA_2830 (.A(net861));
 sg13g2_antennanp ANTENNA_2831 (.A(net861));
 sg13g2_antennanp ANTENNA_2832 (.A(net861));
 sg13g2_antennanp ANTENNA_2833 (.A(net861));
 sg13g2_antennanp ANTENNA_2834 (.A(net861));
 sg13g2_antennanp ANTENNA_2835 (.A(net861));
 sg13g2_antennanp ANTENNA_2836 (.A(net861));
 sg13g2_antennanp ANTENNA_2837 (.A(net861));
 sg13g2_antennanp ANTENNA_2838 (.A(net861));
 sg13g2_antennanp ANTENNA_2839 (.A(net861));
 sg13g2_antennanp ANTENNA_2840 (.A(net861));
 sg13g2_antennanp ANTENNA_2841 (.A(net861));
 sg13g2_antennanp ANTENNA_2842 (.A(net861));
 sg13g2_antennanp ANTENNA_2843 (.A(net861));
 sg13g2_antennanp ANTENNA_2844 (.A(net861));
 sg13g2_antennanp ANTENNA_2845 (.A(net916));
 sg13g2_antennanp ANTENNA_2846 (.A(net916));
 sg13g2_antennanp ANTENNA_2847 (.A(net916));
 sg13g2_antennanp ANTENNA_2848 (.A(net916));
 sg13g2_antennanp ANTENNA_2849 (.A(net916));
 sg13g2_antennanp ANTENNA_2850 (.A(net916));
 sg13g2_antennanp ANTENNA_2851 (.A(net916));
 sg13g2_antennanp ANTENNA_2852 (.A(net916));
 sg13g2_antennanp ANTENNA_2853 (.A(net916));
 sg13g2_antennanp ANTENNA_2854 (.A(net916));
 sg13g2_antennanp ANTENNA_2855 (.A(net916));
 sg13g2_antennanp ANTENNA_2856 (.A(net916));
 sg13g2_antennanp ANTENNA_2857 (.A(net916));
 sg13g2_antennanp ANTENNA_2858 (.A(net916));
 sg13g2_antennanp ANTENNA_2859 (.A(net916));
 sg13g2_antennanp ANTENNA_2860 (.A(net916));
 sg13g2_antennanp ANTENNA_2861 (.A(net993));
 sg13g2_antennanp ANTENNA_2862 (.A(net993));
 sg13g2_antennanp ANTENNA_2863 (.A(net993));
 sg13g2_antennanp ANTENNA_2864 (.A(net993));
 sg13g2_antennanp ANTENNA_2865 (.A(net993));
 sg13g2_antennanp ANTENNA_2866 (.A(net993));
 sg13g2_antennanp ANTENNA_2867 (.A(net993));
 sg13g2_antennanp ANTENNA_2868 (.A(net993));
 sg13g2_antennanp ANTENNA_2869 (.A(net993));
 sg13g2_antennanp ANTENNA_2870 (.A(net993));
 sg13g2_antennanp ANTENNA_2871 (.A(net993));
 sg13g2_antennanp ANTENNA_2872 (.A(net993));
 sg13g2_antennanp ANTENNA_2873 (.A(net993));
 sg13g2_antennanp ANTENNA_2874 (.A(net993));
 sg13g2_antennanp ANTENNA_2875 (.A(net993));
 sg13g2_antennanp ANTENNA_2876 (.A(net993));
 sg13g2_antennanp ANTENNA_2877 (.A(net993));
 sg13g2_antennanp ANTENNA_2878 (.A(net993));
 sg13g2_antennanp ANTENNA_2879 (.A(net993));
 sg13g2_antennanp ANTENNA_2880 (.A(net993));
 sg13g2_antennanp ANTENNA_2881 (.A(net993));
 sg13g2_antennanp ANTENNA_2882 (.A(net993));
 sg13g2_antennanp ANTENNA_2883 (.A(net993));
 sg13g2_antennanp ANTENNA_2884 (.A(net993));
 sg13g2_antennanp ANTENNA_2885 (.A(net993));
 sg13g2_antennanp ANTENNA_2886 (.A(net1066));
 sg13g2_antennanp ANTENNA_2887 (.A(net1066));
 sg13g2_antennanp ANTENNA_2888 (.A(net1066));
 sg13g2_antennanp ANTENNA_2889 (.A(net1066));
 sg13g2_antennanp ANTENNA_2890 (.A(net1066));
 sg13g2_antennanp ANTENNA_2891 (.A(net1066));
 sg13g2_antennanp ANTENNA_2892 (.A(net1066));
 sg13g2_antennanp ANTENNA_2893 (.A(net1066));
 sg13g2_antennanp ANTENNA_2894 (.A(net1066));
 sg13g2_antennanp ANTENNA_2895 (.A(net1066));
 sg13g2_antennanp ANTENNA_2896 (.A(net1066));
 sg13g2_antennanp ANTENNA_2897 (.A(net1066));
 sg13g2_antennanp ANTENNA_2898 (.A(net1066));
 sg13g2_antennanp ANTENNA_2899 (.A(net1066));
 sg13g2_antennanp ANTENNA_2900 (.A(net1066));
 sg13g2_antennanp ANTENNA_2901 (.A(net1066));
 sg13g2_antennanp ANTENNA_2902 (.A(net1066));
 sg13g2_antennanp ANTENNA_2903 (.A(net1066));
 sg13g2_antennanp ANTENNA_2904 (.A(net1071));
 sg13g2_antennanp ANTENNA_2905 (.A(net1071));
 sg13g2_antennanp ANTENNA_2906 (.A(net1071));
 sg13g2_antennanp ANTENNA_2907 (.A(net1071));
 sg13g2_antennanp ANTENNA_2908 (.A(net1071));
 sg13g2_antennanp ANTENNA_2909 (.A(net1071));
 sg13g2_antennanp ANTENNA_2910 (.A(net1071));
 sg13g2_antennanp ANTENNA_2911 (.A(net1071));
 sg13g2_antennanp ANTENNA_2912 (.A(net1071));
 sg13g2_antennanp ANTENNA_2913 (.A(net1071));
 sg13g2_antennanp ANTENNA_2914 (.A(net1071));
 sg13g2_antennanp ANTENNA_2915 (.A(net1071));
 sg13g2_antennanp ANTENNA_2916 (.A(net1071));
 sg13g2_antennanp ANTENNA_2917 (.A(net1071));
 sg13g2_antennanp ANTENNA_2918 (.A(net1071));
 sg13g2_antennanp ANTENNA_2919 (.A(net1071));
 sg13g2_antennanp ANTENNA_2920 (.A(net1071));
 sg13g2_antennanp ANTENNA_2921 (.A(net1071));
 sg13g2_antennanp ANTENNA_2922 (.A(net1071));
 sg13g2_antennanp ANTENNA_2923 (.A(net1071));
 sg13g2_antennanp ANTENNA_2924 (.A(net1071));
 sg13g2_antennanp ANTENNA_2925 (.A(net1071));
 sg13g2_antennanp ANTENNA_2926 (.A(net1071));
 sg13g2_antennanp ANTENNA_2927 (.A(net1071));
 sg13g2_antennanp ANTENNA_2928 (.A(net1071));
 sg13g2_antennanp ANTENNA_2929 (.A(net1071));
 sg13g2_antennanp ANTENNA_2930 (.A(net1071));
 sg13g2_antennanp ANTENNA_2931 (.A(net1071));
 sg13g2_antennanp ANTENNA_2932 (.A(net1071));
 sg13g2_antennanp ANTENNA_2933 (.A(net1071));
 sg13g2_antennanp ANTENNA_2934 (.A(net1071));
 sg13g2_antennanp ANTENNA_2935 (.A(net1071));
 sg13g2_antennanp ANTENNA_2936 (.A(net1071));
 sg13g2_antennanp ANTENNA_2937 (.A(net1071));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_fill_2 FILLER_0_42 ();
 sg13g2_fill_1 FILLER_0_44 ();
 sg13g2_decap_8 FILLER_0_71 ();
 sg13g2_decap_4 FILLER_0_78 ();
 sg13g2_decap_8 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_100 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_fill_1 FILLER_0_128 ();
 sg13g2_decap_4 FILLER_0_155 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_fill_2 FILLER_0_242 ();
 sg13g2_fill_1 FILLER_0_244 ();
 sg13g2_fill_2 FILLER_0_249 ();
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_fill_2 FILLER_0_257 ();
 sg13g2_fill_1 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_fill_1 FILLER_0_285 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_fill_1 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_fill_1 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_4 FILLER_0_395 ();
 sg13g2_fill_1 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_fill_1 FILLER_0_425 ();
 sg13g2_decap_4 FILLER_0_482 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_fill_2 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_fill_2 FILLER_0_567 ();
 sg13g2_fill_1 FILLER_0_569 ();
 sg13g2_decap_4 FILLER_0_596 ();
 sg13g2_fill_1 FILLER_0_600 ();
 sg13g2_fill_1 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_fill_2 FILLER_0_647 ();
 sg13g2_fill_1 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_fill_1 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_fill_1 FILLER_0_718 ();
 sg13g2_fill_1 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_fill_2 FILLER_0_787 ();
 sg13g2_decap_4 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_4 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_839 ();
 sg13g2_decap_8 FILLER_0_846 ();
 sg13g2_decap_8 FILLER_0_853 ();
 sg13g2_decap_8 FILLER_0_860 ();
 sg13g2_decap_4 FILLER_0_881 ();
 sg13g2_fill_1 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_fill_1 FILLER_0_903 ();
 sg13g2_fill_2 FILLER_0_918 ();
 sg13g2_fill_1 FILLER_0_920 ();
 sg13g2_fill_2 FILLER_0_960 ();
 sg13g2_fill_1 FILLER_0_962 ();
 sg13g2_fill_2 FILLER_0_967 ();
 sg13g2_fill_2 FILLER_0_979 ();
 sg13g2_fill_1 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_fill_1 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1034 ();
 sg13g2_fill_2 FILLER_0_1041 ();
 sg13g2_fill_1 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1074 ();
 sg13g2_decap_8 FILLER_0_1081 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_8 FILLER_0_1095 ();
 sg13g2_decap_8 FILLER_0_1112 ();
 sg13g2_decap_8 FILLER_0_1119 ();
 sg13g2_decap_8 FILLER_0_1126 ();
 sg13g2_fill_2 FILLER_0_1133 ();
 sg13g2_fill_1 FILLER_0_1135 ();
 sg13g2_decap_8 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1153 ();
 sg13g2_decap_8 FILLER_0_1160 ();
 sg13g2_decap_8 FILLER_0_1167 ();
 sg13g2_decap_8 FILLER_0_1174 ();
 sg13g2_decap_8 FILLER_0_1181 ();
 sg13g2_decap_8 FILLER_0_1188 ();
 sg13g2_fill_2 FILLER_0_1195 ();
 sg13g2_fill_1 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1234 ();
 sg13g2_decap_4 FILLER_0_1241 ();
 sg13g2_fill_1 FILLER_0_1245 ();
 sg13g2_decap_4 FILLER_0_1300 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_4 FILLER_0_1344 ();
 sg13g2_fill_1 FILLER_0_1352 ();
 sg13g2_decap_8 FILLER_0_1357 ();
 sg13g2_decap_8 FILLER_0_1364 ();
 sg13g2_decap_8 FILLER_0_1371 ();
 sg13g2_decap_4 FILLER_0_1378 ();
 sg13g2_fill_2 FILLER_0_1382 ();
 sg13g2_decap_4 FILLER_0_1420 ();
 sg13g2_fill_1 FILLER_0_1424 ();
 sg13g2_decap_8 FILLER_0_1451 ();
 sg13g2_decap_8 FILLER_0_1458 ();
 sg13g2_decap_8 FILLER_0_1465 ();
 sg13g2_decap_4 FILLER_0_1472 ();
 sg13g2_fill_2 FILLER_0_1480 ();
 sg13g2_fill_2 FILLER_0_1496 ();
 sg13g2_fill_1 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1513 ();
 sg13g2_decap_8 FILLER_0_1520 ();
 sg13g2_decap_8 FILLER_0_1527 ();
 sg13g2_decap_8 FILLER_0_1534 ();
 sg13g2_decap_8 FILLER_0_1541 ();
 sg13g2_decap_8 FILLER_0_1548 ();
 sg13g2_decap_8 FILLER_0_1555 ();
 sg13g2_decap_4 FILLER_0_1562 ();
 sg13g2_fill_1 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1571 ();
 sg13g2_decap_8 FILLER_0_1578 ();
 sg13g2_fill_1 FILLER_0_1585 ();
 sg13g2_fill_2 FILLER_0_1624 ();
 sg13g2_fill_1 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_4 FILLER_0_1678 ();
 sg13g2_fill_1 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1709 ();
 sg13g2_decap_4 FILLER_0_1716 ();
 sg13g2_fill_1 FILLER_0_1720 ();
 sg13g2_decap_4 FILLER_0_1725 ();
 sg13g2_fill_1 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1738 ();
 sg13g2_decap_8 FILLER_0_1745 ();
 sg13g2_decap_8 FILLER_0_1752 ();
 sg13g2_decap_8 FILLER_0_1759 ();
 sg13g2_decap_8 FILLER_0_1776 ();
 sg13g2_decap_8 FILLER_0_1783 ();
 sg13g2_decap_8 FILLER_0_1790 ();
 sg13g2_decap_8 FILLER_0_1797 ();
 sg13g2_fill_1 FILLER_0_1804 ();
 sg13g2_decap_8 FILLER_0_1819 ();
 sg13g2_decap_8 FILLER_0_1826 ();
 sg13g2_decap_8 FILLER_0_1833 ();
 sg13g2_fill_2 FILLER_0_1840 ();
 sg13g2_decap_8 FILLER_0_1846 ();
 sg13g2_decap_8 FILLER_0_1853 ();
 sg13g2_decap_8 FILLER_0_1860 ();
 sg13g2_fill_1 FILLER_0_1867 ();
 sg13g2_decap_8 FILLER_0_1882 ();
 sg13g2_decap_8 FILLER_0_1889 ();
 sg13g2_decap_8 FILLER_0_1896 ();
 sg13g2_decap_8 FILLER_0_1903 ();
 sg13g2_fill_2 FILLER_0_1910 ();
 sg13g2_fill_1 FILLER_0_1912 ();
 sg13g2_decap_8 FILLER_0_1965 ();
 sg13g2_decap_8 FILLER_0_1972 ();
 sg13g2_decap_8 FILLER_0_1979 ();
 sg13g2_decap_8 FILLER_0_1986 ();
 sg13g2_decap_8 FILLER_0_1993 ();
 sg13g2_decap_4 FILLER_0_2000 ();
 sg13g2_fill_1 FILLER_0_2004 ();
 sg13g2_decap_8 FILLER_0_2043 ();
 sg13g2_decap_8 FILLER_0_2050 ();
 sg13g2_decap_8 FILLER_0_2057 ();
 sg13g2_fill_2 FILLER_0_2064 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2099 ();
 sg13g2_decap_8 FILLER_0_2142 ();
 sg13g2_decap_8 FILLER_0_2149 ();
 sg13g2_decap_4 FILLER_0_2182 ();
 sg13g2_fill_2 FILLER_0_2186 ();
 sg13g2_decap_8 FILLER_0_2196 ();
 sg13g2_decap_8 FILLER_0_2203 ();
 sg13g2_decap_8 FILLER_0_2210 ();
 sg13g2_decap_8 FILLER_0_2217 ();
 sg13g2_decap_8 FILLER_0_2224 ();
 sg13g2_decap_8 FILLER_0_2231 ();
 sg13g2_fill_2 FILLER_0_2238 ();
 sg13g2_decap_8 FILLER_0_2266 ();
 sg13g2_decap_4 FILLER_0_2273 ();
 sg13g2_fill_1 FILLER_0_2277 ();
 sg13g2_decap_8 FILLER_0_2312 ();
 sg13g2_decap_8 FILLER_0_2319 ();
 sg13g2_decap_8 FILLER_0_2326 ();
 sg13g2_decap_8 FILLER_0_2333 ();
 sg13g2_decap_8 FILLER_0_2340 ();
 sg13g2_fill_2 FILLER_0_2347 ();
 sg13g2_fill_1 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2418 ();
 sg13g2_decap_8 FILLER_0_2425 ();
 sg13g2_decap_4 FILLER_0_2432 ();
 sg13g2_fill_1 FILLER_0_2436 ();
 sg13g2_fill_2 FILLER_0_2473 ();
 sg13g2_decap_8 FILLER_0_2516 ();
 sg13g2_decap_8 FILLER_0_2523 ();
 sg13g2_decap_8 FILLER_0_2530 ();
 sg13g2_decap_8 FILLER_0_2537 ();
 sg13g2_decap_8 FILLER_0_2544 ();
 sg13g2_decap_8 FILLER_0_2551 ();
 sg13g2_decap_8 FILLER_0_2558 ();
 sg13g2_decap_8 FILLER_0_2565 ();
 sg13g2_decap_8 FILLER_0_2572 ();
 sg13g2_decap_8 FILLER_0_2579 ();
 sg13g2_decap_8 FILLER_0_2586 ();
 sg13g2_decap_8 FILLER_0_2593 ();
 sg13g2_decap_8 FILLER_0_2600 ();
 sg13g2_decap_8 FILLER_0_2607 ();
 sg13g2_decap_8 FILLER_0_2614 ();
 sg13g2_decap_8 FILLER_0_2621 ();
 sg13g2_decap_8 FILLER_0_2628 ();
 sg13g2_decap_8 FILLER_0_2635 ();
 sg13g2_decap_8 FILLER_0_2642 ();
 sg13g2_decap_8 FILLER_0_2649 ();
 sg13g2_decap_8 FILLER_0_2656 ();
 sg13g2_decap_8 FILLER_0_2663 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_34 ();
 sg13g2_decap_8 FILLER_1_41 ();
 sg13g2_fill_2 FILLER_1_86 ();
 sg13g2_decap_8 FILLER_1_114 ();
 sg13g2_decap_4 FILLER_1_121 ();
 sg13g2_fill_2 FILLER_1_129 ();
 sg13g2_fill_2 FILLER_1_164 ();
 sg13g2_fill_1 FILLER_1_248 ();
 sg13g2_fill_1 FILLER_1_275 ();
 sg13g2_decap_4 FILLER_1_280 ();
 sg13g2_fill_1 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_333 ();
 sg13g2_fill_2 FILLER_1_340 ();
 sg13g2_fill_1 FILLER_1_342 ();
 sg13g2_fill_1 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_4 FILLER_1_359 ();
 sg13g2_fill_2 FILLER_1_436 ();
 sg13g2_fill_2 FILLER_1_464 ();
 sg13g2_fill_1 FILLER_1_466 ();
 sg13g2_decap_4 FILLER_1_471 ();
 sg13g2_fill_2 FILLER_1_475 ();
 sg13g2_decap_8 FILLER_1_503 ();
 sg13g2_fill_2 FILLER_1_510 ();
 sg13g2_fill_2 FILLER_1_535 ();
 sg13g2_fill_1 FILLER_1_537 ();
 sg13g2_decap_8 FILLER_1_568 ();
 sg13g2_decap_8 FILLER_1_575 ();
 sg13g2_fill_2 FILLER_1_623 ();
 sg13g2_fill_1 FILLER_1_629 ();
 sg13g2_fill_2 FILLER_1_656 ();
 sg13g2_decap_4 FILLER_1_694 ();
 sg13g2_fill_2 FILLER_1_698 ();
 sg13g2_fill_2 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_4 FILLER_1_777 ();
 sg13g2_fill_2 FILLER_1_815 ();
 sg13g2_fill_1 FILLER_1_822 ();
 sg13g2_decap_8 FILLER_1_849 ();
 sg13g2_fill_1 FILLER_1_856 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_fill_2 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_fill_2 FILLER_1_907 ();
 sg13g2_fill_1 FILLER_1_940 ();
 sg13g2_fill_2 FILLER_1_1029 ();
 sg13g2_fill_2 FILLER_1_1055 ();
 sg13g2_fill_1 FILLER_1_1083 ();
 sg13g2_decap_4 FILLER_1_1088 ();
 sg13g2_fill_1 FILLER_1_1092 ();
 sg13g2_fill_2 FILLER_1_1110 ();
 sg13g2_decap_8 FILLER_1_1178 ();
 sg13g2_decap_4 FILLER_1_1185 ();
 sg13g2_fill_2 FILLER_1_1203 ();
 sg13g2_fill_1 FILLER_1_1205 ();
 sg13g2_decap_8 FILLER_1_1220 ();
 sg13g2_fill_1 FILLER_1_1227 ();
 sg13g2_decap_4 FILLER_1_1238 ();
 sg13g2_fill_2 FILLER_1_1242 ();
 sg13g2_fill_2 FILLER_1_1304 ();
 sg13g2_fill_1 FILLER_1_1306 ();
 sg13g2_fill_2 FILLER_1_1333 ();
 sg13g2_fill_1 FILLER_1_1345 ();
 sg13g2_decap_4 FILLER_1_1372 ();
 sg13g2_decap_8 FILLER_1_1390 ();
 sg13g2_decap_8 FILLER_1_1427 ();
 sg13g2_decap_4 FILLER_1_1434 ();
 sg13g2_fill_2 FILLER_1_1472 ();
 sg13g2_fill_2 FILLER_1_1500 ();
 sg13g2_fill_1 FILLER_1_1502 ();
 sg13g2_fill_1 FILLER_1_1507 ();
 sg13g2_decap_8 FILLER_1_1534 ();
 sg13g2_decap_8 FILLER_1_1541 ();
 sg13g2_fill_2 FILLER_1_1548 ();
 sg13g2_decap_4 FILLER_1_1631 ();
 sg13g2_fill_2 FILLER_1_1635 ();
 sg13g2_fill_2 FILLER_1_1641 ();
 sg13g2_fill_1 FILLER_1_1643 ();
 sg13g2_decap_4 FILLER_1_1748 ();
 sg13g2_fill_1 FILLER_1_1752 ();
 sg13g2_decap_4 FILLER_1_1789 ();
 sg13g2_fill_1 FILLER_1_1793 ();
 sg13g2_decap_4 FILLER_1_1830 ();
 sg13g2_fill_1 FILLER_1_1834 ();
 sg13g2_decap_4 FILLER_1_1861 ();
 sg13g2_fill_2 FILLER_1_1865 ();
 sg13g2_decap_8 FILLER_1_1893 ();
 sg13g2_fill_2 FILLER_1_1900 ();
 sg13g2_fill_1 FILLER_1_1902 ();
 sg13g2_fill_2 FILLER_1_1907 ();
 sg13g2_decap_4 FILLER_1_1969 ();
 sg13g2_fill_2 FILLER_1_2075 ();
 sg13g2_decap_8 FILLER_1_2100 ();
 sg13g2_fill_1 FILLER_1_2107 ();
 sg13g2_decap_4 FILLER_1_2129 ();
 sg13g2_fill_1 FILLER_1_2133 ();
 sg13g2_fill_2 FILLER_1_2154 ();
 sg13g2_decap_4 FILLER_1_2166 ();
 sg13g2_fill_1 FILLER_1_2170 ();
 sg13g2_decap_4 FILLER_1_2211 ();
 sg13g2_fill_2 FILLER_1_2215 ();
 sg13g2_decap_4 FILLER_1_2243 ();
 sg13g2_fill_2 FILLER_1_2247 ();
 sg13g2_fill_1 FILLER_1_2300 ();
 sg13g2_decap_4 FILLER_1_2337 ();
 sg13g2_fill_1 FILLER_1_2341 ();
 sg13g2_fill_1 FILLER_1_2392 ();
 sg13g2_fill_2 FILLER_1_2419 ();
 sg13g2_fill_1 FILLER_1_2421 ();
 sg13g2_fill_2 FILLER_1_2426 ();
 sg13g2_fill_1 FILLER_1_2428 ();
 sg13g2_fill_2 FILLER_1_2459 ();
 sg13g2_fill_1 FILLER_1_2461 ();
 sg13g2_decap_8 FILLER_1_2537 ();
 sg13g2_decap_8 FILLER_1_2544 ();
 sg13g2_decap_8 FILLER_1_2551 ();
 sg13g2_decap_8 FILLER_1_2558 ();
 sg13g2_decap_8 FILLER_1_2565 ();
 sg13g2_decap_8 FILLER_1_2572 ();
 sg13g2_decap_8 FILLER_1_2579 ();
 sg13g2_decap_8 FILLER_1_2586 ();
 sg13g2_decap_8 FILLER_1_2593 ();
 sg13g2_decap_8 FILLER_1_2600 ();
 sg13g2_decap_8 FILLER_1_2607 ();
 sg13g2_decap_8 FILLER_1_2614 ();
 sg13g2_decap_8 FILLER_1_2621 ();
 sg13g2_decap_8 FILLER_1_2628 ();
 sg13g2_decap_8 FILLER_1_2635 ();
 sg13g2_decap_8 FILLER_1_2642 ();
 sg13g2_decap_8 FILLER_1_2649 ();
 sg13g2_decap_8 FILLER_1_2656 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_fill_1 FILLER_2_110 ();
 sg13g2_fill_2 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_fill_2 FILLER_2_197 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_fill_2 FILLER_2_223 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_353 ();
 sg13g2_fill_1 FILLER_2_364 ();
 sg13g2_decap_4 FILLER_2_386 ();
 sg13g2_fill_1 FILLER_2_390 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_fill_1 FILLER_2_481 ();
 sg13g2_fill_1 FILLER_2_518 ();
 sg13g2_fill_1 FILLER_2_549 ();
 sg13g2_fill_1 FILLER_2_576 ();
 sg13g2_fill_1 FILLER_2_603 ();
 sg13g2_fill_2 FILLER_2_635 ();
 sg13g2_fill_1 FILLER_2_637 ();
 sg13g2_fill_1 FILLER_2_669 ();
 sg13g2_fill_2 FILLER_2_696 ();
 sg13g2_fill_2 FILLER_2_729 ();
 sg13g2_fill_2 FILLER_2_819 ();
 sg13g2_fill_1 FILLER_2_821 ();
 sg13g2_fill_2 FILLER_2_853 ();
 sg13g2_decap_4 FILLER_2_907 ();
 sg13g2_decap_4 FILLER_2_941 ();
 sg13g2_decap_8 FILLER_2_996 ();
 sg13g2_fill_1 FILLER_2_1003 ();
 sg13g2_decap_4 FILLER_2_1133 ();
 sg13g2_fill_1 FILLER_2_1163 ();
 sg13g2_decap_4 FILLER_2_1204 ();
 sg13g2_fill_2 FILLER_2_1242 ();
 sg13g2_decap_4 FILLER_2_1270 ();
 sg13g2_fill_2 FILLER_2_1274 ();
 sg13g2_decap_4 FILLER_2_1299 ();
 sg13g2_fill_2 FILLER_2_1303 ();
 sg13g2_decap_8 FILLER_2_1393 ();
 sg13g2_fill_2 FILLER_2_1400 ();
 sg13g2_fill_2 FILLER_2_1607 ();
 sg13g2_fill_1 FILLER_2_1609 ();
 sg13g2_fill_2 FILLER_2_1645 ();
 sg13g2_fill_2 FILLER_2_1657 ();
 sg13g2_decap_4 FILLER_2_1689 ();
 sg13g2_fill_2 FILLER_2_1697 ();
 sg13g2_fill_1 FILLER_2_1699 ();
 sg13g2_fill_1 FILLER_2_1714 ();
 sg13g2_fill_2 FILLER_2_1720 ();
 sg13g2_fill_1 FILLER_2_1722 ();
 sg13g2_fill_2 FILLER_2_1749 ();
 sg13g2_fill_1 FILLER_2_1751 ();
 sg13g2_decap_4 FILLER_2_1788 ();
 sg13g2_fill_2 FILLER_2_1857 ();
 sg13g2_fill_1 FILLER_2_1859 ();
 sg13g2_fill_1 FILLER_2_1912 ();
 sg13g2_fill_1 FILLER_2_1933 ();
 sg13g2_fill_1 FILLER_2_1938 ();
 sg13g2_fill_1 FILLER_2_1943 ();
 sg13g2_fill_2 FILLER_2_1969 ();
 sg13g2_fill_1 FILLER_2_1971 ();
 sg13g2_fill_2 FILLER_2_2008 ();
 sg13g2_fill_2 FILLER_2_2054 ();
 sg13g2_fill_1 FILLER_2_2056 ();
 sg13g2_decap_8 FILLER_2_2097 ();
 sg13g2_fill_1 FILLER_2_2130 ();
 sg13g2_fill_1 FILLER_2_2157 ();
 sg13g2_fill_2 FILLER_2_2194 ();
 sg13g2_fill_2 FILLER_2_2222 ();
 sg13g2_fill_1 FILLER_2_2228 ();
 sg13g2_fill_2 FILLER_2_2322 ();
 sg13g2_decap_4 FILLER_2_2328 ();
 sg13g2_fill_1 FILLER_2_2332 ();
 sg13g2_fill_2 FILLER_2_2369 ();
 sg13g2_fill_1 FILLER_2_2371 ();
 sg13g2_decap_4 FILLER_2_2421 ();
 sg13g2_decap_4 FILLER_2_2455 ();
 sg13g2_fill_2 FILLER_2_2459 ();
 sg13g2_fill_2 FILLER_2_2531 ();
 sg13g2_fill_1 FILLER_2_2533 ();
 sg13g2_decap_8 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2545 ();
 sg13g2_decap_8 FILLER_2_2552 ();
 sg13g2_decap_8 FILLER_2_2559 ();
 sg13g2_decap_8 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2573 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_decap_8 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2601 ();
 sg13g2_decap_8 FILLER_2_2608 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_decap_8 FILLER_2_2622 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_decap_8 FILLER_2_2636 ();
 sg13g2_decap_8 FILLER_2_2643 ();
 sg13g2_decap_8 FILLER_2_2650 ();
 sg13g2_decap_8 FILLER_2_2657 ();
 sg13g2_decap_4 FILLER_2_2664 ();
 sg13g2_fill_2 FILLER_2_2668 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_4 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_32 ();
 sg13g2_decap_4 FILLER_3_37 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_2 FILLER_3_95 ();
 sg13g2_fill_1 FILLER_3_111 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_141 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_4 FILLER_3_209 ();
 sg13g2_fill_1 FILLER_3_213 ();
 sg13g2_fill_2 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_259 ();
 sg13g2_fill_2 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_fill_2 FILLER_3_330 ();
 sg13g2_decap_4 FILLER_3_368 ();
 sg13g2_fill_2 FILLER_3_382 ();
 sg13g2_fill_2 FILLER_3_441 ();
 sg13g2_fill_2 FILLER_3_453 ();
 sg13g2_fill_1 FILLER_3_455 ();
 sg13g2_fill_1 FILLER_3_466 ();
 sg13g2_fill_1 FILLER_3_477 ();
 sg13g2_decap_4 FILLER_3_497 ();
 sg13g2_fill_2 FILLER_3_501 ();
 sg13g2_fill_1 FILLER_3_529 ();
 sg13g2_fill_2 FILLER_3_580 ();
 sg13g2_fill_2 FILLER_3_629 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_fill_1 FILLER_3_698 ();
 sg13g2_fill_1 FILLER_3_773 ();
 sg13g2_fill_1 FILLER_3_782 ();
 sg13g2_fill_1 FILLER_3_788 ();
 sg13g2_decap_4 FILLER_3_854 ();
 sg13g2_fill_2 FILLER_3_858 ();
 sg13g2_fill_2 FILLER_3_907 ();
 sg13g2_fill_1 FILLER_3_909 ();
 sg13g2_fill_1 FILLER_3_936 ();
 sg13g2_fill_1 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_1000 ();
 sg13g2_fill_1 FILLER_3_1007 ();
 sg13g2_fill_1 FILLER_3_1048 ();
 sg13g2_decap_8 FILLER_3_1079 ();
 sg13g2_fill_1 FILLER_3_1086 ();
 sg13g2_decap_8 FILLER_3_1131 ();
 sg13g2_fill_2 FILLER_3_1138 ();
 sg13g2_fill_1 FILLER_3_1140 ();
 sg13g2_fill_2 FILLER_3_1159 ();
 sg13g2_fill_1 FILLER_3_1200 ();
 sg13g2_decap_4 FILLER_3_1227 ();
 sg13g2_fill_1 FILLER_3_1231 ();
 sg13g2_decap_4 FILLER_3_1258 ();
 sg13g2_fill_1 FILLER_3_1262 ();
 sg13g2_fill_2 FILLER_3_1309 ();
 sg13g2_fill_2 FILLER_3_1323 ();
 sg13g2_fill_2 FILLER_3_1335 ();
 sg13g2_fill_1 FILLER_3_1340 ();
 sg13g2_fill_2 FILLER_3_1377 ();
 sg13g2_fill_2 FILLER_3_1441 ();
 sg13g2_fill_1 FILLER_3_1443 ();
 sg13g2_fill_2 FILLER_3_1470 ();
 sg13g2_fill_1 FILLER_3_1511 ();
 sg13g2_fill_1 FILLER_3_1538 ();
 sg13g2_fill_1 FILLER_3_1543 ();
 sg13g2_fill_2 FILLER_3_1570 ();
 sg13g2_fill_1 FILLER_3_1578 ();
 sg13g2_fill_1 FILLER_3_1600 ();
 sg13g2_fill_1 FILLER_3_1618 ();
 sg13g2_fill_1 FILLER_3_1625 ();
 sg13g2_decap_4 FILLER_3_1673 ();
 sg13g2_fill_1 FILLER_3_1677 ();
 sg13g2_fill_1 FILLER_3_1682 ();
 sg13g2_fill_1 FILLER_3_1718 ();
 sg13g2_decap_8 FILLER_3_1725 ();
 sg13g2_fill_2 FILLER_3_1732 ();
 sg13g2_decap_8 FILLER_3_1738 ();
 sg13g2_decap_8 FILLER_3_1745 ();
 sg13g2_decap_4 FILLER_3_1795 ();
 sg13g2_fill_1 FILLER_3_1803 ();
 sg13g2_fill_1 FILLER_3_1830 ();
 sg13g2_decap_4 FILLER_3_1857 ();
 sg13g2_decap_8 FILLER_3_1874 ();
 sg13g2_fill_1 FILLER_3_1881 ();
 sg13g2_fill_2 FILLER_3_1903 ();
 sg13g2_decap_8 FILLER_3_1909 ();
 sg13g2_decap_8 FILLER_3_1916 ();
 sg13g2_decap_4 FILLER_3_1923 ();
 sg13g2_fill_2 FILLER_3_1964 ();
 sg13g2_fill_1 FILLER_3_1966 ();
 sg13g2_fill_1 FILLER_3_2028 ();
 sg13g2_decap_8 FILLER_3_2058 ();
 sg13g2_decap_8 FILLER_3_2065 ();
 sg13g2_fill_2 FILLER_3_2072 ();
 sg13g2_fill_1 FILLER_3_2074 ();
 sg13g2_fill_2 FILLER_3_2105 ();
 sg13g2_fill_1 FILLER_3_2107 ();
 sg13g2_fill_1 FILLER_3_2138 ();
 sg13g2_fill_2 FILLER_3_2192 ();
 sg13g2_fill_1 FILLER_3_2230 ();
 sg13g2_fill_1 FILLER_3_2241 ();
 sg13g2_fill_1 FILLER_3_2246 ();
 sg13g2_fill_2 FILLER_3_2283 ();
 sg13g2_fill_2 FILLER_3_2305 ();
 sg13g2_decap_4 FILLER_3_2333 ();
 sg13g2_fill_2 FILLER_3_2337 ();
 sg13g2_fill_1 FILLER_3_2349 ();
 sg13g2_fill_2 FILLER_3_2376 ();
 sg13g2_fill_1 FILLER_3_2399 ();
 sg13g2_decap_4 FILLER_3_2451 ();
 sg13g2_fill_1 FILLER_3_2455 ();
 sg13g2_decap_4 FILLER_3_2496 ();
 sg13g2_fill_2 FILLER_3_2500 ();
 sg13g2_decap_8 FILLER_3_2542 ();
 sg13g2_decap_8 FILLER_3_2549 ();
 sg13g2_decap_8 FILLER_3_2556 ();
 sg13g2_decap_8 FILLER_3_2563 ();
 sg13g2_decap_8 FILLER_3_2570 ();
 sg13g2_decap_8 FILLER_3_2577 ();
 sg13g2_decap_8 FILLER_3_2584 ();
 sg13g2_decap_8 FILLER_3_2591 ();
 sg13g2_decap_8 FILLER_3_2598 ();
 sg13g2_decap_8 FILLER_3_2605 ();
 sg13g2_decap_8 FILLER_3_2612 ();
 sg13g2_decap_8 FILLER_3_2619 ();
 sg13g2_decap_8 FILLER_3_2626 ();
 sg13g2_decap_8 FILLER_3_2633 ();
 sg13g2_decap_8 FILLER_3_2640 ();
 sg13g2_decap_8 FILLER_3_2647 ();
 sg13g2_decap_8 FILLER_3_2654 ();
 sg13g2_decap_8 FILLER_3_2661 ();
 sg13g2_fill_2 FILLER_3_2668 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_36 ();
 sg13g2_fill_2 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_111 ();
 sg13g2_fill_1 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_144 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_fill_1 FILLER_4_164 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_fill_1 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_fill_1 FILLER_4_247 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_261 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_fill_2 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_4 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_348 ();
 sg13g2_fill_2 FILLER_4_359 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_fill_2 FILLER_4_383 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_2 FILLER_4_429 ();
 sg13g2_fill_2 FILLER_4_461 ();
 sg13g2_fill_1 FILLER_4_463 ();
 sg13g2_fill_1 FILLER_4_490 ();
 sg13g2_fill_2 FILLER_4_539 ();
 sg13g2_fill_1 FILLER_4_541 ();
 sg13g2_fill_2 FILLER_4_556 ();
 sg13g2_fill_1 FILLER_4_558 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_4 FILLER_4_587 ();
 sg13g2_fill_1 FILLER_4_591 ();
 sg13g2_fill_2 FILLER_4_614 ();
 sg13g2_fill_2 FILLER_4_628 ();
 sg13g2_decap_4 FILLER_4_635 ();
 sg13g2_fill_1 FILLER_4_643 ();
 sg13g2_fill_2 FILLER_4_649 ();
 sg13g2_fill_1 FILLER_4_665 ();
 sg13g2_fill_2 FILLER_4_670 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_4 FILLER_4_700 ();
 sg13g2_fill_2 FILLER_4_734 ();
 sg13g2_fill_1 FILLER_4_736 ();
 sg13g2_fill_1 FILLER_4_773 ();
 sg13g2_fill_2 FILLER_4_788 ();
 sg13g2_fill_1 FILLER_4_790 ();
 sg13g2_fill_1 FILLER_4_795 ();
 sg13g2_fill_1 FILLER_4_821 ();
 sg13g2_fill_2 FILLER_4_835 ();
 sg13g2_decap_8 FILLER_4_845 ();
 sg13g2_fill_1 FILLER_4_852 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_fill_2 FILLER_4_881 ();
 sg13g2_fill_2 FILLER_4_901 ();
 sg13g2_fill_1 FILLER_4_913 ();
 sg13g2_fill_1 FILLER_4_918 ();
 sg13g2_fill_2 FILLER_4_961 ();
 sg13g2_fill_1 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_4 FILLER_4_992 ();
 sg13g2_fill_2 FILLER_4_996 ();
 sg13g2_fill_1 FILLER_4_1006 ();
 sg13g2_fill_2 FILLER_4_1063 ();
 sg13g2_decap_8 FILLER_4_1077 ();
 sg13g2_decap_4 FILLER_4_1084 ();
 sg13g2_fill_2 FILLER_4_1088 ();
 sg13g2_decap_8 FILLER_4_1098 ();
 sg13g2_decap_8 FILLER_4_1105 ();
 sg13g2_decap_4 FILLER_4_1122 ();
 sg13g2_fill_1 FILLER_4_1198 ();
 sg13g2_fill_2 FILLER_4_1209 ();
 sg13g2_fill_1 FILLER_4_1211 ();
 sg13g2_decap_4 FILLER_4_1216 ();
 sg13g2_fill_2 FILLER_4_1246 ();
 sg13g2_fill_2 FILLER_4_1274 ();
 sg13g2_decap_8 FILLER_4_1310 ();
 sg13g2_decap_8 FILLER_4_1317 ();
 sg13g2_decap_4 FILLER_4_1324 ();
 sg13g2_fill_2 FILLER_4_1328 ();
 sg13g2_decap_8 FILLER_4_1334 ();
 sg13g2_decap_4 FILLER_4_1341 ();
 sg13g2_fill_2 FILLER_4_1345 ();
 sg13g2_fill_1 FILLER_4_1357 ();
 sg13g2_fill_1 FILLER_4_1362 ();
 sg13g2_decap_8 FILLER_4_1373 ();
 sg13g2_fill_1 FILLER_4_1380 ();
 sg13g2_fill_1 FILLER_4_1421 ();
 sg13g2_decap_4 FILLER_4_1446 ();
 sg13g2_decap_8 FILLER_4_1454 ();
 sg13g2_decap_8 FILLER_4_1461 ();
 sg13g2_decap_8 FILLER_4_1468 ();
 sg13g2_fill_2 FILLER_4_1475 ();
 sg13g2_fill_2 FILLER_4_1489 ();
 sg13g2_fill_1 FILLER_4_1491 ();
 sg13g2_decap_4 FILLER_4_1495 ();
 sg13g2_fill_1 FILLER_4_1509 ();
 sg13g2_decap_8 FILLER_4_1528 ();
 sg13g2_fill_2 FILLER_4_1535 ();
 sg13g2_decap_4 FILLER_4_1541 ();
 sg13g2_fill_1 FILLER_4_1545 ();
 sg13g2_fill_2 FILLER_4_1550 ();
 sg13g2_fill_2 FILLER_4_1563 ();
 sg13g2_fill_2 FILLER_4_1585 ();
 sg13g2_fill_1 FILLER_4_1593 ();
 sg13g2_fill_1 FILLER_4_1610 ();
 sg13g2_fill_2 FILLER_4_1616 ();
 sg13g2_fill_1 FILLER_4_1623 ();
 sg13g2_decap_4 FILLER_4_1665 ();
 sg13g2_fill_2 FILLER_4_1669 ();
 sg13g2_fill_1 FILLER_4_1687 ();
 sg13g2_fill_2 FILLER_4_1699 ();
 sg13g2_fill_1 FILLER_4_1760 ();
 sg13g2_decap_4 FILLER_4_1773 ();
 sg13g2_fill_1 FILLER_4_1781 ();
 sg13g2_fill_2 FILLER_4_1838 ();
 sg13g2_decap_8 FILLER_4_1844 ();
 sg13g2_fill_2 FILLER_4_1851 ();
 sg13g2_fill_1 FILLER_4_1853 ();
 sg13g2_fill_2 FILLER_4_1955 ();
 sg13g2_fill_1 FILLER_4_1957 ();
 sg13g2_fill_1 FILLER_4_1990 ();
 sg13g2_fill_1 FILLER_4_2017 ();
 sg13g2_fill_1 FILLER_4_2028 ();
 sg13g2_decap_8 FILLER_4_2101 ();
 sg13g2_fill_1 FILLER_4_2122 ();
 sg13g2_decap_8 FILLER_4_2137 ();
 sg13g2_decap_4 FILLER_4_2144 ();
 sg13g2_decap_4 FILLER_4_2152 ();
 sg13g2_fill_1 FILLER_4_2156 ();
 sg13g2_fill_1 FILLER_4_2192 ();
 sg13g2_fill_2 FILLER_4_2229 ();
 sg13g2_fill_1 FILLER_4_2231 ();
 sg13g2_fill_2 FILLER_4_2242 ();
 sg13g2_fill_1 FILLER_4_2244 ();
 sg13g2_decap_4 FILLER_4_2276 ();
 sg13g2_fill_2 FILLER_4_2280 ();
 sg13g2_decap_8 FILLER_4_2286 ();
 sg13g2_decap_8 FILLER_4_2293 ();
 sg13g2_decap_4 FILLER_4_2300 ();
 sg13g2_fill_2 FILLER_4_2314 ();
 sg13g2_decap_8 FILLER_4_2342 ();
 sg13g2_decap_4 FILLER_4_2349 ();
 sg13g2_fill_1 FILLER_4_2353 ();
 sg13g2_decap_4 FILLER_4_2409 ();
 sg13g2_fill_1 FILLER_4_2413 ();
 sg13g2_decap_8 FILLER_4_2457 ();
 sg13g2_fill_2 FILLER_4_2495 ();
 sg13g2_decap_8 FILLER_4_2518 ();
 sg13g2_decap_8 FILLER_4_2525 ();
 sg13g2_decap_8 FILLER_4_2532 ();
 sg13g2_decap_8 FILLER_4_2539 ();
 sg13g2_decap_8 FILLER_4_2546 ();
 sg13g2_decap_8 FILLER_4_2553 ();
 sg13g2_decap_8 FILLER_4_2560 ();
 sg13g2_decap_8 FILLER_4_2567 ();
 sg13g2_decap_8 FILLER_4_2574 ();
 sg13g2_decap_8 FILLER_4_2581 ();
 sg13g2_decap_8 FILLER_4_2588 ();
 sg13g2_decap_8 FILLER_4_2595 ();
 sg13g2_decap_8 FILLER_4_2602 ();
 sg13g2_decap_8 FILLER_4_2609 ();
 sg13g2_decap_8 FILLER_4_2616 ();
 sg13g2_decap_8 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_4 FILLER_4_2665 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_decap_8 FILLER_5_52 ();
 sg13g2_fill_2 FILLER_5_71 ();
 sg13g2_fill_1 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_191 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_235 ();
 sg13g2_decap_4 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_4 FILLER_5_329 ();
 sg13g2_fill_2 FILLER_5_333 ();
 sg13g2_fill_2 FILLER_5_361 ();
 sg13g2_decap_4 FILLER_5_389 ();
 sg13g2_fill_1 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_5_425 ();
 sg13g2_fill_2 FILLER_5_432 ();
 sg13g2_fill_1 FILLER_5_434 ();
 sg13g2_fill_2 FILLER_5_439 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_505 ();
 sg13g2_decap_4 FILLER_5_510 ();
 sg13g2_fill_2 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_533 ();
 sg13g2_decap_8 FILLER_5_540 ();
 sg13g2_decap_4 FILLER_5_547 ();
 sg13g2_decap_4 FILLER_5_561 ();
 sg13g2_fill_2 FILLER_5_565 ();
 sg13g2_fill_2 FILLER_5_572 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_4 FILLER_5_599 ();
 sg13g2_fill_1 FILLER_5_607 ();
 sg13g2_fill_1 FILLER_5_617 ();
 sg13g2_fill_2 FILLER_5_644 ();
 sg13g2_fill_2 FILLER_5_677 ();
 sg13g2_fill_1 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_684 ();
 sg13g2_decap_8 FILLER_5_691 ();
 sg13g2_fill_2 FILLER_5_698 ();
 sg13g2_fill_2 FILLER_5_781 ();
 sg13g2_decap_4 FILLER_5_788 ();
 sg13g2_fill_1 FILLER_5_792 ();
 sg13g2_fill_2 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_fill_2 FILLER_5_819 ();
 sg13g2_fill_1 FILLER_5_826 ();
 sg13g2_fill_2 FILLER_5_876 ();
 sg13g2_fill_2 FILLER_5_902 ();
 sg13g2_fill_1 FILLER_5_904 ();
 sg13g2_fill_2 FILLER_5_909 ();
 sg13g2_fill_1 FILLER_5_968 ();
 sg13g2_fill_1 FILLER_5_973 ();
 sg13g2_fill_2 FILLER_5_979 ();
 sg13g2_fill_1 FILLER_5_981 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_8 FILLER_5_997 ();
 sg13g2_fill_2 FILLER_5_1004 ();
 sg13g2_fill_1 FILLER_5_1020 ();
 sg13g2_fill_2 FILLER_5_1065 ();
 sg13g2_fill_1 FILLER_5_1067 ();
 sg13g2_fill_1 FILLER_5_1155 ();
 sg13g2_fill_2 FILLER_5_1182 ();
 sg13g2_fill_1 FILLER_5_1210 ();
 sg13g2_fill_1 FILLER_5_1215 ();
 sg13g2_fill_1 FILLER_5_1230 ();
 sg13g2_fill_1 FILLER_5_1241 ();
 sg13g2_fill_2 FILLER_5_1258 ();
 sg13g2_decap_8 FILLER_5_1296 ();
 sg13g2_decap_8 FILLER_5_1303 ();
 sg13g2_decap_8 FILLER_5_1310 ();
 sg13g2_decap_4 FILLER_5_1317 ();
 sg13g2_fill_2 FILLER_5_1321 ();
 sg13g2_decap_4 FILLER_5_1349 ();
 sg13g2_fill_1 FILLER_5_1363 ();
 sg13g2_decap_8 FILLER_5_1368 ();
 sg13g2_fill_2 FILLER_5_1375 ();
 sg13g2_fill_1 FILLER_5_1421 ();
 sg13g2_fill_1 FILLER_5_1432 ();
 sg13g2_fill_2 FILLER_5_1459 ();
 sg13g2_decap_8 FILLER_5_1471 ();
 sg13g2_decap_8 FILLER_5_1478 ();
 sg13g2_fill_2 FILLER_5_1485 ();
 sg13g2_decap_8 FILLER_5_1537 ();
 sg13g2_decap_4 FILLER_5_1544 ();
 sg13g2_fill_2 FILLER_5_1548 ();
 sg13g2_decap_4 FILLER_5_1554 ();
 sg13g2_fill_1 FILLER_5_1558 ();
 sg13g2_fill_1 FILLER_5_1597 ();
 sg13g2_fill_1 FILLER_5_1603 ();
 sg13g2_fill_1 FILLER_5_1609 ();
 sg13g2_fill_2 FILLER_5_1622 ();
 sg13g2_fill_1 FILLER_5_1624 ();
 sg13g2_fill_2 FILLER_5_1630 ();
 sg13g2_fill_2 FILLER_5_1638 ();
 sg13g2_fill_1 FILLER_5_1650 ();
 sg13g2_decap_8 FILLER_5_1657 ();
 sg13g2_fill_1 FILLER_5_1664 ();
 sg13g2_fill_1 FILLER_5_1676 ();
 sg13g2_decap_4 FILLER_5_1685 ();
 sg13g2_fill_1 FILLER_5_1693 ();
 sg13g2_fill_1 FILLER_5_1698 ();
 sg13g2_fill_2 FILLER_5_1724 ();
 sg13g2_decap_8 FILLER_5_1750 ();
 sg13g2_decap_8 FILLER_5_1757 ();
 sg13g2_fill_1 FILLER_5_1764 ();
 sg13g2_decap_4 FILLER_5_1773 ();
 sg13g2_fill_2 FILLER_5_1787 ();
 sg13g2_fill_1 FILLER_5_1793 ();
 sg13g2_decap_8 FILLER_5_1804 ();
 sg13g2_fill_2 FILLER_5_1815 ();
 sg13g2_decap_8 FILLER_5_1847 ();
 sg13g2_decap_8 FILLER_5_1854 ();
 sg13g2_fill_2 FILLER_5_1861 ();
 sg13g2_fill_1 FILLER_5_1863 ();
 sg13g2_fill_2 FILLER_5_1868 ();
 sg13g2_fill_1 FILLER_5_1870 ();
 sg13g2_decap_8 FILLER_5_1895 ();
 sg13g2_decap_8 FILLER_5_1902 ();
 sg13g2_decap_8 FILLER_5_1909 ();
 sg13g2_decap_4 FILLER_5_1916 ();
 sg13g2_fill_1 FILLER_5_1920 ();
 sg13g2_fill_2 FILLER_5_1935 ();
 sg13g2_fill_1 FILLER_5_1937 ();
 sg13g2_fill_2 FILLER_5_1972 ();
 sg13g2_fill_1 FILLER_5_1974 ();
 sg13g2_fill_2 FILLER_5_1999 ();
 sg13g2_fill_1 FILLER_5_2001 ();
 sg13g2_fill_2 FILLER_5_2006 ();
 sg13g2_fill_1 FILLER_5_2026 ();
 sg13g2_fill_2 FILLER_5_2086 ();
 sg13g2_fill_2 FILLER_5_2109 ();
 sg13g2_fill_1 FILLER_5_2111 ();
 sg13g2_decap_8 FILLER_5_2122 ();
 sg13g2_decap_8 FILLER_5_2139 ();
 sg13g2_decap_8 FILLER_5_2146 ();
 sg13g2_decap_8 FILLER_5_2153 ();
 sg13g2_decap_8 FILLER_5_2160 ();
 sg13g2_decap_8 FILLER_5_2171 ();
 sg13g2_decap_8 FILLER_5_2178 ();
 sg13g2_fill_1 FILLER_5_2185 ();
 sg13g2_decap_8 FILLER_5_2226 ();
 sg13g2_decap_4 FILLER_5_2233 ();
 sg13g2_fill_1 FILLER_5_2237 ();
 sg13g2_fill_2 FILLER_5_2263 ();
 sg13g2_fill_1 FILLER_5_2301 ();
 sg13g2_fill_1 FILLER_5_2312 ();
 sg13g2_fill_1 FILLER_5_2339 ();
 sg13g2_fill_2 FILLER_5_2350 ();
 sg13g2_fill_1 FILLER_5_2362 ();
 sg13g2_decap_4 FILLER_5_2393 ();
 sg13g2_decap_4 FILLER_5_2423 ();
 sg13g2_fill_2 FILLER_5_2437 ();
 sg13g2_fill_1 FILLER_5_2439 ();
 sg13g2_decap_8 FILLER_5_2461 ();
 sg13g2_decap_4 FILLER_5_2468 ();
 sg13g2_fill_1 FILLER_5_2472 ();
 sg13g2_decap_4 FILLER_5_2481 ();
 sg13g2_fill_2 FILLER_5_2495 ();
 sg13g2_fill_1 FILLER_5_2497 ();
 sg13g2_decap_4 FILLER_5_2528 ();
 sg13g2_decap_8 FILLER_5_2557 ();
 sg13g2_decap_8 FILLER_5_2564 ();
 sg13g2_decap_8 FILLER_5_2571 ();
 sg13g2_decap_8 FILLER_5_2578 ();
 sg13g2_decap_8 FILLER_5_2585 ();
 sg13g2_decap_8 FILLER_5_2592 ();
 sg13g2_decap_8 FILLER_5_2599 ();
 sg13g2_decap_8 FILLER_5_2606 ();
 sg13g2_decap_8 FILLER_5_2613 ();
 sg13g2_decap_8 FILLER_5_2620 ();
 sg13g2_decap_8 FILLER_5_2627 ();
 sg13g2_decap_8 FILLER_5_2634 ();
 sg13g2_decap_8 FILLER_5_2641 ();
 sg13g2_decap_8 FILLER_5_2648 ();
 sg13g2_decap_8 FILLER_5_2655 ();
 sg13g2_decap_8 FILLER_5_2662 ();
 sg13g2_fill_1 FILLER_5_2669 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_1 FILLER_6_29 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_fill_2 FILLER_6_149 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_2 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_decap_4 FILLER_6_216 ();
 sg13g2_fill_2 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_4 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_fill_2 FILLER_6_316 ();
 sg13g2_fill_2 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_fill_2 FILLER_6_403 ();
 sg13g2_fill_1 FILLER_6_405 ();
 sg13g2_fill_1 FILLER_6_442 ();
 sg13g2_fill_2 FILLER_6_482 ();
 sg13g2_decap_8 FILLER_6_492 ();
 sg13g2_decap_8 FILLER_6_499 ();
 sg13g2_decap_8 FILLER_6_506 ();
 sg13g2_fill_2 FILLER_6_513 ();
 sg13g2_fill_1 FILLER_6_541 ();
 sg13g2_fill_1 FILLER_6_546 ();
 sg13g2_decap_4 FILLER_6_551 ();
 sg13g2_fill_1 FILLER_6_555 ();
 sg13g2_fill_2 FILLER_6_603 ();
 sg13g2_fill_1 FILLER_6_605 ();
 sg13g2_decap_4 FILLER_6_637 ();
 sg13g2_fill_2 FILLER_6_646 ();
 sg13g2_fill_2 FILLER_6_652 ();
 sg13g2_fill_2 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_fill_2 FILLER_6_725 ();
 sg13g2_fill_2 FILLER_6_777 ();
 sg13g2_fill_1 FILLER_6_779 ();
 sg13g2_fill_1 FILLER_6_784 ();
 sg13g2_fill_2 FILLER_6_819 ();
 sg13g2_fill_1 FILLER_6_821 ();
 sg13g2_fill_2 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_864 ();
 sg13g2_fill_2 FILLER_6_923 ();
 sg13g2_fill_1 FILLER_6_925 ();
 sg13g2_fill_1 FILLER_6_949 ();
 sg13g2_fill_1 FILLER_6_976 ();
 sg13g2_fill_1 FILLER_6_1081 ();
 sg13g2_decap_4 FILLER_6_1086 ();
 sg13g2_decap_4 FILLER_6_1126 ();
 sg13g2_fill_2 FILLER_6_1130 ();
 sg13g2_fill_2 FILLER_6_1146 ();
 sg13g2_fill_1 FILLER_6_1148 ();
 sg13g2_fill_2 FILLER_6_1173 ();
 sg13g2_fill_1 FILLER_6_1175 ();
 sg13g2_fill_2 FILLER_6_1196 ();
 sg13g2_fill_1 FILLER_6_1198 ();
 sg13g2_decap_8 FILLER_6_1225 ();
 sg13g2_fill_2 FILLER_6_1232 ();
 sg13g2_fill_1 FILLER_6_1247 ();
 sg13g2_decap_8 FILLER_6_1276 ();
 sg13g2_fill_2 FILLER_6_1283 ();
 sg13g2_fill_1 FILLER_6_1285 ();
 sg13g2_fill_1 FILLER_6_1316 ();
 sg13g2_fill_1 FILLER_6_1321 ();
 sg13g2_fill_1 FILLER_6_1392 ();
 sg13g2_decap_8 FILLER_6_1410 ();
 sg13g2_fill_1 FILLER_6_1417 ();
 sg13g2_decap_4 FILLER_6_1428 ();
 sg13g2_fill_2 FILLER_6_1432 ();
 sg13g2_decap_8 FILLER_6_1460 ();
 sg13g2_decap_4 FILLER_6_1503 ();
 sg13g2_decap_4 FILLER_6_1511 ();
 sg13g2_fill_2 FILLER_6_1515 ();
 sg13g2_fill_2 FILLER_6_1578 ();
 sg13g2_fill_1 FILLER_6_1594 ();
 sg13g2_fill_1 FILLER_6_1604 ();
 sg13g2_fill_1 FILLER_6_1609 ();
 sg13g2_fill_1 FILLER_6_1692 ();
 sg13g2_fill_2 FILLER_6_1725 ();
 sg13g2_decap_4 FILLER_6_1753 ();
 sg13g2_fill_2 FILLER_6_1762 ();
 sg13g2_decap_4 FILLER_6_1781 ();
 sg13g2_fill_1 FILLER_6_1785 ();
 sg13g2_decap_8 FILLER_6_1795 ();
 sg13g2_fill_2 FILLER_6_1802 ();
 sg13g2_fill_1 FILLER_6_1804 ();
 sg13g2_fill_2 FILLER_6_1809 ();
 sg13g2_fill_1 FILLER_6_1811 ();
 sg13g2_fill_1 FILLER_6_1816 ();
 sg13g2_decap_4 FILLER_6_1848 ();
 sg13g2_fill_1 FILLER_6_1882 ();
 sg13g2_decap_8 FILLER_6_1904 ();
 sg13g2_fill_1 FILLER_6_1911 ();
 sg13g2_fill_1 FILLER_6_2003 ();
 sg13g2_fill_1 FILLER_6_2030 ();
 sg13g2_decap_4 FILLER_6_2079 ();
 sg13g2_fill_1 FILLER_6_2083 ();
 sg13g2_decap_8 FILLER_6_2092 ();
 sg13g2_decap_8 FILLER_6_2099 ();
 sg13g2_decap_4 FILLER_6_2106 ();
 sg13g2_fill_2 FILLER_6_2110 ();
 sg13g2_fill_1 FILLER_6_2122 ();
 sg13g2_decap_8 FILLER_6_2174 ();
 sg13g2_decap_8 FILLER_6_2181 ();
 sg13g2_decap_4 FILLER_6_2188 ();
 sg13g2_fill_2 FILLER_6_2192 ();
 sg13g2_decap_8 FILLER_6_2215 ();
 sg13g2_fill_2 FILLER_6_2222 ();
 sg13g2_fill_1 FILLER_6_2224 ();
 sg13g2_fill_1 FILLER_6_2235 ();
 sg13g2_decap_4 FILLER_6_2272 ();
 sg13g2_fill_1 FILLER_6_2276 ();
 sg13g2_decap_8 FILLER_6_2290 ();
 sg13g2_fill_2 FILLER_6_2297 ();
 sg13g2_fill_1 FILLER_6_2332 ();
 sg13g2_fill_1 FILLER_6_2337 ();
 sg13g2_fill_2 FILLER_6_2364 ();
 sg13g2_fill_2 FILLER_6_2379 ();
 sg13g2_fill_2 FILLER_6_2394 ();
 sg13g2_decap_8 FILLER_6_2406 ();
 sg13g2_decap_8 FILLER_6_2413 ();
 sg13g2_decap_8 FILLER_6_2420 ();
 sg13g2_decap_8 FILLER_6_2460 ();
 sg13g2_decap_8 FILLER_6_2467 ();
 sg13g2_decap_8 FILLER_6_2474 ();
 sg13g2_decap_8 FILLER_6_2481 ();
 sg13g2_decap_4 FILLER_6_2488 ();
 sg13g2_fill_2 FILLER_6_2528 ();
 sg13g2_decap_8 FILLER_6_2566 ();
 sg13g2_decap_8 FILLER_6_2573 ();
 sg13g2_decap_8 FILLER_6_2580 ();
 sg13g2_decap_8 FILLER_6_2587 ();
 sg13g2_decap_8 FILLER_6_2594 ();
 sg13g2_decap_8 FILLER_6_2601 ();
 sg13g2_decap_8 FILLER_6_2608 ();
 sg13g2_decap_8 FILLER_6_2615 ();
 sg13g2_decap_8 FILLER_6_2622 ();
 sg13g2_decap_8 FILLER_6_2629 ();
 sg13g2_decap_8 FILLER_6_2636 ();
 sg13g2_decap_8 FILLER_6_2643 ();
 sg13g2_decap_8 FILLER_6_2650 ();
 sg13g2_decap_8 FILLER_6_2657 ();
 sg13g2_decap_4 FILLER_6_2664 ();
 sg13g2_fill_2 FILLER_6_2668 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_97 ();
 sg13g2_fill_1 FILLER_7_123 ();
 sg13g2_fill_2 FILLER_7_145 ();
 sg13g2_fill_2 FILLER_7_160 ();
 sg13g2_fill_2 FILLER_7_181 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_fill_1 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_230 ();
 sg13g2_fill_2 FILLER_7_237 ();
 sg13g2_decap_4 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_400 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_417 ();
 sg13g2_decap_4 FILLER_7_428 ();
 sg13g2_fill_2 FILLER_7_432 ();
 sg13g2_decap_4 FILLER_7_460 ();
 sg13g2_fill_2 FILLER_7_495 ();
 sg13g2_decap_4 FILLER_7_506 ();
 sg13g2_fill_2 FILLER_7_566 ();
 sg13g2_fill_1 FILLER_7_620 ();
 sg13g2_fill_2 FILLER_7_647 ();
 sg13g2_fill_1 FILLER_7_714 ();
 sg13g2_fill_1 FILLER_7_723 ();
 sg13g2_fill_1 FILLER_7_741 ();
 sg13g2_fill_1 FILLER_7_768 ();
 sg13g2_fill_1 FILLER_7_795 ();
 sg13g2_fill_1 FILLER_7_848 ();
 sg13g2_fill_1 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_923 ();
 sg13g2_fill_2 FILLER_7_960 ();
 sg13g2_fill_1 FILLER_7_962 ();
 sg13g2_fill_1 FILLER_7_999 ();
 sg13g2_fill_1 FILLER_7_1021 ();
 sg13g2_fill_1 FILLER_7_1032 ();
 sg13g2_fill_2 FILLER_7_1038 ();
 sg13g2_fill_2 FILLER_7_1070 ();
 sg13g2_fill_1 FILLER_7_1072 ();
 sg13g2_fill_2 FILLER_7_1093 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_fill_1 FILLER_7_1113 ();
 sg13g2_decap_4 FILLER_7_1118 ();
 sg13g2_fill_2 FILLER_7_1122 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_fill_2 FILLER_7_1135 ();
 sg13g2_decap_8 FILLER_7_1147 ();
 sg13g2_decap_4 FILLER_7_1154 ();
 sg13g2_fill_1 FILLER_7_1184 ();
 sg13g2_decap_4 FILLER_7_1247 ();
 sg13g2_fill_1 FILLER_7_1251 ();
 sg13g2_decap_8 FILLER_7_1269 ();
 sg13g2_decap_8 FILLER_7_1276 ();
 sg13g2_decap_8 FILLER_7_1283 ();
 sg13g2_decap_4 FILLER_7_1290 ();
 sg13g2_fill_2 FILLER_7_1294 ();
 sg13g2_fill_1 FILLER_7_1306 ();
 sg13g2_fill_2 FILLER_7_1333 ();
 sg13g2_fill_2 FILLER_7_1339 ();
 sg13g2_decap_4 FILLER_7_1351 ();
 sg13g2_decap_8 FILLER_7_1372 ();
 sg13g2_decap_8 FILLER_7_1379 ();
 sg13g2_fill_2 FILLER_7_1386 ();
 sg13g2_fill_2 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1423 ();
 sg13g2_fill_1 FILLER_7_1430 ();
 sg13g2_fill_2 FILLER_7_1471 ();
 sg13g2_decap_4 FILLER_7_1529 ();
 sg13g2_fill_1 FILLER_7_1537 ();
 sg13g2_fill_2 FILLER_7_1598 ();
 sg13g2_fill_1 FILLER_7_1616 ();
 sg13g2_fill_2 FILLER_7_1657 ();
 sg13g2_fill_1 FILLER_7_1664 ();
 sg13g2_fill_1 FILLER_7_1670 ();
 sg13g2_fill_1 FILLER_7_1676 ();
 sg13g2_fill_2 FILLER_7_1703 ();
 sg13g2_fill_2 FILLER_7_1710 ();
 sg13g2_fill_2 FILLER_7_1736 ();
 sg13g2_fill_1 FILLER_7_1738 ();
 sg13g2_fill_2 FILLER_7_1780 ();
 sg13g2_fill_1 FILLER_7_1782 ();
 sg13g2_fill_2 FILLER_7_1809 ();
 sg13g2_fill_1 FILLER_7_1841 ();
 sg13g2_fill_2 FILLER_7_1868 ();
 sg13g2_fill_1 FILLER_7_1896 ();
 sg13g2_decap_8 FILLER_7_1923 ();
 sg13g2_fill_2 FILLER_7_1930 ();
 sg13g2_fill_2 FILLER_7_1965 ();
 sg13g2_fill_1 FILLER_7_1967 ();
 sg13g2_fill_1 FILLER_7_1994 ();
 sg13g2_decap_4 FILLER_7_1999 ();
 sg13g2_fill_2 FILLER_7_2015 ();
 sg13g2_fill_1 FILLER_7_2027 ();
 sg13g2_fill_2 FILLER_7_2065 ();
 sg13g2_fill_1 FILLER_7_2067 ();
 sg13g2_decap_8 FILLER_7_2082 ();
 sg13g2_decap_8 FILLER_7_2089 ();
 sg13g2_decap_8 FILLER_7_2165 ();
 sg13g2_fill_2 FILLER_7_2172 ();
 sg13g2_decap_8 FILLER_7_2204 ();
 sg13g2_decap_8 FILLER_7_2211 ();
 sg13g2_fill_1 FILLER_7_2218 ();
 sg13g2_decap_8 FILLER_7_2300 ();
 sg13g2_decap_4 FILLER_7_2317 ();
 sg13g2_fill_2 FILLER_7_2321 ();
 sg13g2_decap_8 FILLER_7_2385 ();
 sg13g2_fill_1 FILLER_7_2392 ();
 sg13g2_decap_8 FILLER_7_2414 ();
 sg13g2_fill_1 FILLER_7_2421 ();
 sg13g2_decap_8 FILLER_7_2588 ();
 sg13g2_decap_8 FILLER_7_2595 ();
 sg13g2_decap_8 FILLER_7_2602 ();
 sg13g2_decap_8 FILLER_7_2609 ();
 sg13g2_decap_8 FILLER_7_2616 ();
 sg13g2_decap_8 FILLER_7_2623 ();
 sg13g2_decap_8 FILLER_7_2630 ();
 sg13g2_decap_8 FILLER_7_2637 ();
 sg13g2_decap_8 FILLER_7_2644 ();
 sg13g2_decap_8 FILLER_7_2651 ();
 sg13g2_decap_8 FILLER_7_2658 ();
 sg13g2_decap_4 FILLER_7_2665 ();
 sg13g2_fill_1 FILLER_7_2669 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_8 ();
 sg13g2_fill_2 FILLER_8_13 ();
 sg13g2_fill_2 FILLER_8_41 ();
 sg13g2_fill_2 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_58 ();
 sg13g2_fill_2 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_92 ();
 sg13g2_decap_4 FILLER_8_99 ();
 sg13g2_fill_2 FILLER_8_103 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_177 ();
 sg13g2_fill_2 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_fill_2 FILLER_8_361 ();
 sg13g2_decap_4 FILLER_8_377 ();
 sg13g2_fill_2 FILLER_8_411 ();
 sg13g2_fill_1 FILLER_8_413 ();
 sg13g2_fill_2 FILLER_8_471 ();
 sg13g2_fill_1 FILLER_8_473 ();
 sg13g2_fill_2 FILLER_8_556 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_fill_1 FILLER_8_569 ();
 sg13g2_fill_1 FILLER_8_630 ();
 sg13g2_fill_1 FILLER_8_656 ();
 sg13g2_fill_1 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_667 ();
 sg13g2_fill_1 FILLER_8_678 ();
 sg13g2_fill_2 FILLER_8_705 ();
 sg13g2_fill_1 FILLER_8_707 ();
 sg13g2_decap_4 FILLER_8_767 ();
 sg13g2_fill_2 FILLER_8_771 ();
 sg13g2_fill_1 FILLER_8_803 ();
 sg13g2_fill_1 FILLER_8_809 ();
 sg13g2_decap_4 FILLER_8_814 ();
 sg13g2_fill_1 FILLER_8_818 ();
 sg13g2_fill_1 FILLER_8_845 ();
 sg13g2_fill_2 FILLER_8_859 ();
 sg13g2_fill_2 FILLER_8_871 ();
 sg13g2_decap_4 FILLER_8_877 ();
 sg13g2_fill_1 FILLER_8_916 ();
 sg13g2_fill_2 FILLER_8_927 ();
 sg13g2_fill_1 FILLER_8_959 ();
 sg13g2_fill_2 FILLER_8_1043 ();
 sg13g2_fill_2 FILLER_8_1049 ();
 sg13g2_fill_2 FILLER_8_1064 ();
 sg13g2_fill_1 FILLER_8_1066 ();
 sg13g2_decap_8 FILLER_8_1097 ();
 sg13g2_decap_8 FILLER_8_1104 ();
 sg13g2_fill_2 FILLER_8_1111 ();
 sg13g2_fill_2 FILLER_8_1162 ();
 sg13g2_fill_2 FILLER_8_1198 ();
 sg13g2_fill_1 FILLER_8_1200 ();
 sg13g2_decap_8 FILLER_8_1205 ();
 sg13g2_decap_4 FILLER_8_1212 ();
 sg13g2_fill_1 FILLER_8_1216 ();
 sg13g2_decap_8 FILLER_8_1221 ();
 sg13g2_decap_4 FILLER_8_1228 ();
 sg13g2_decap_4 FILLER_8_1235 ();
 sg13g2_fill_2 FILLER_8_1264 ();
 sg13g2_fill_1 FILLER_8_1266 ();
 sg13g2_fill_1 FILLER_8_1274 ();
 sg13g2_decap_8 FILLER_8_1282 ();
 sg13g2_decap_4 FILLER_8_1289 ();
 sg13g2_fill_2 FILLER_8_1293 ();
 sg13g2_fill_1 FILLER_8_1309 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_8_1341 ();
 sg13g2_fill_1 FILLER_8_1348 ();
 sg13g2_decap_8 FILLER_8_1359 ();
 sg13g2_fill_1 FILLER_8_1366 ();
 sg13g2_decap_4 FILLER_8_1372 ();
 sg13g2_fill_2 FILLER_8_1376 ();
 sg13g2_fill_2 FILLER_8_1430 ();
 sg13g2_fill_1 FILLER_8_1432 ();
 sg13g2_decap_4 FILLER_8_1445 ();
 sg13g2_fill_2 FILLER_8_1449 ();
 sg13g2_fill_1 FILLER_8_1461 ();
 sg13g2_fill_1 FILLER_8_1472 ();
 sg13g2_fill_1 FILLER_8_1484 ();
 sg13g2_decap_4 FILLER_8_1495 ();
 sg13g2_fill_2 FILLER_8_1499 ();
 sg13g2_decap_8 FILLER_8_1528 ();
 sg13g2_fill_1 FILLER_8_1535 ();
 sg13g2_fill_2 FILLER_8_1584 ();
 sg13g2_fill_2 FILLER_8_1660 ();
 sg13g2_fill_1 FILLER_8_1662 ();
 sg13g2_fill_1 FILLER_8_1694 ();
 sg13g2_fill_2 FILLER_8_1705 ();
 sg13g2_fill_2 FILLER_8_1733 ();
 sg13g2_fill_1 FILLER_8_1735 ();
 sg13g2_decap_4 FILLER_8_1740 ();
 sg13g2_fill_2 FILLER_8_1744 ();
 sg13g2_decap_4 FILLER_8_1750 ();
 sg13g2_fill_2 FILLER_8_1754 ();
 sg13g2_fill_1 FILLER_8_1761 ();
 sg13g2_fill_1 FILLER_8_1779 ();
 sg13g2_decap_4 FILLER_8_1834 ();
 sg13g2_fill_1 FILLER_8_1838 ();
 sg13g2_fill_2 FILLER_8_1852 ();
 sg13g2_fill_1 FILLER_8_1858 ();
 sg13g2_fill_2 FILLER_8_1869 ();
 sg13g2_decap_4 FILLER_8_1901 ();
 sg13g2_fill_1 FILLER_8_1905 ();
 sg13g2_decap_8 FILLER_8_1910 ();
 sg13g2_fill_2 FILLER_8_1917 ();
 sg13g2_fill_1 FILLER_8_2056 ();
 sg13g2_decap_4 FILLER_8_2109 ();
 sg13g2_fill_1 FILLER_8_2113 ();
 sg13g2_decap_4 FILLER_8_2206 ();
 sg13g2_fill_1 FILLER_8_2210 ();
 sg13g2_fill_2 FILLER_8_2224 ();
 sg13g2_fill_1 FILLER_8_2243 ();
 sg13g2_decap_4 FILLER_8_2318 ();
 sg13g2_fill_2 FILLER_8_2363 ();
 sg13g2_fill_1 FILLER_8_2365 ();
 sg13g2_fill_1 FILLER_8_2370 ();
 sg13g2_fill_1 FILLER_8_2407 ();
 sg13g2_fill_1 FILLER_8_2467 ();
 sg13g2_fill_1 FILLER_8_2472 ();
 sg13g2_fill_1 FILLER_8_2520 ();
 sg13g2_decap_8 FILLER_8_2570 ();
 sg13g2_decap_8 FILLER_8_2577 ();
 sg13g2_decap_8 FILLER_8_2584 ();
 sg13g2_decap_8 FILLER_8_2591 ();
 sg13g2_decap_8 FILLER_8_2598 ();
 sg13g2_decap_8 FILLER_8_2605 ();
 sg13g2_decap_8 FILLER_8_2612 ();
 sg13g2_decap_8 FILLER_8_2619 ();
 sg13g2_decap_8 FILLER_8_2626 ();
 sg13g2_decap_8 FILLER_8_2633 ();
 sg13g2_decap_8 FILLER_8_2640 ();
 sg13g2_decap_8 FILLER_8_2647 ();
 sg13g2_decap_8 FILLER_8_2654 ();
 sg13g2_decap_8 FILLER_8_2661 ();
 sg13g2_fill_2 FILLER_8_2668 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_31 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_4 FILLER_9_46 ();
 sg13g2_decap_4 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_decap_8 FILLER_9_79 ();
 sg13g2_decap_8 FILLER_9_86 ();
 sg13g2_decap_8 FILLER_9_93 ();
 sg13g2_decap_4 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_180 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_285 ();
 sg13g2_decap_4 FILLER_9_292 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_327 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_4 FILLER_9_359 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_decap_4 FILLER_9_416 ();
 sg13g2_fill_2 FILLER_9_456 ();
 sg13g2_fill_1 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_4 FILLER_9_476 ();
 sg13g2_fill_1 FILLER_9_480 ();
 sg13g2_fill_2 FILLER_9_544 ();
 sg13g2_fill_2 FILLER_9_581 ();
 sg13g2_fill_2 FILLER_9_587 ();
 sg13g2_decap_4 FILLER_9_593 ();
 sg13g2_fill_1 FILLER_9_597 ();
 sg13g2_decap_4 FILLER_9_602 ();
 sg13g2_fill_2 FILLER_9_606 ();
 sg13g2_fill_1 FILLER_9_612 ();
 sg13g2_fill_2 FILLER_9_618 ();
 sg13g2_fill_1 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_fill_2 FILLER_9_654 ();
 sg13g2_decap_4 FILLER_9_665 ();
 sg13g2_fill_1 FILLER_9_669 ();
 sg13g2_decap_4 FILLER_9_701 ();
 sg13g2_fill_2 FILLER_9_705 ();
 sg13g2_fill_1 FILLER_9_747 ();
 sg13g2_fill_1 FILLER_9_752 ();
 sg13g2_decap_4 FILLER_9_779 ();
 sg13g2_fill_2 FILLER_9_796 ();
 sg13g2_decap_4 FILLER_9_819 ();
 sg13g2_fill_1 FILLER_9_831 ();
 sg13g2_decap_4 FILLER_9_842 ();
 sg13g2_fill_2 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_915 ();
 sg13g2_fill_1 FILLER_9_922 ();
 sg13g2_fill_2 FILLER_9_983 ();
 sg13g2_fill_1 FILLER_9_985 ();
 sg13g2_fill_2 FILLER_9_1048 ();
 sg13g2_fill_2 FILLER_9_1058 ();
 sg13g2_fill_2 FILLER_9_1064 ();
 sg13g2_fill_2 FILLER_9_1071 ();
 sg13g2_fill_2 FILLER_9_1103 ();
 sg13g2_fill_1 FILLER_9_1105 ();
 sg13g2_fill_1 FILLER_9_1111 ();
 sg13g2_fill_1 FILLER_9_1177 ();
 sg13g2_fill_2 FILLER_9_1192 ();
 sg13g2_fill_2 FILLER_9_1271 ();
 sg13g2_decap_8 FILLER_9_1284 ();
 sg13g2_decap_8 FILLER_9_1291 ();
 sg13g2_fill_1 FILLER_9_1306 ();
 sg13g2_fill_1 FILLER_9_1317 ();
 sg13g2_fill_1 FILLER_9_1333 ();
 sg13g2_decap_8 FILLER_9_1338 ();
 sg13g2_fill_2 FILLER_9_1359 ();
 sg13g2_fill_1 FILLER_9_1361 ();
 sg13g2_fill_1 FILLER_9_1372 ();
 sg13g2_fill_2 FILLER_9_1377 ();
 sg13g2_fill_2 FILLER_9_1389 ();
 sg13g2_fill_1 FILLER_9_1397 ();
 sg13g2_fill_1 FILLER_9_1408 ();
 sg13g2_fill_2 FILLER_9_1414 ();
 sg13g2_fill_1 FILLER_9_1416 ();
 sg13g2_fill_2 FILLER_9_1456 ();
 sg13g2_fill_1 FILLER_9_1458 ();
 sg13g2_decap_8 FILLER_9_1464 ();
 sg13g2_decap_8 FILLER_9_1471 ();
 sg13g2_decap_8 FILLER_9_1478 ();
 sg13g2_decap_8 FILLER_9_1485 ();
 sg13g2_decap_4 FILLER_9_1492 ();
 sg13g2_fill_1 FILLER_9_1515 ();
 sg13g2_fill_2 FILLER_9_1527 ();
 sg13g2_fill_1 FILLER_9_1529 ();
 sg13g2_fill_2 FILLER_9_1567 ();
 sg13g2_fill_2 FILLER_9_1577 ();
 sg13g2_fill_1 FILLER_9_1604 ();
 sg13g2_fill_1 FILLER_9_1610 ();
 sg13g2_fill_2 FILLER_9_1654 ();
 sg13g2_fill_1 FILLER_9_1720 ();
 sg13g2_fill_2 FILLER_9_1747 ();
 sg13g2_fill_1 FILLER_9_1749 ();
 sg13g2_fill_2 FILLER_9_1796 ();
 sg13g2_fill_2 FILLER_9_1808 ();
 sg13g2_fill_1 FILLER_9_1814 ();
 sg13g2_decap_8 FILLER_9_1859 ();
 sg13g2_decap_8 FILLER_9_1866 ();
 sg13g2_fill_2 FILLER_9_1873 ();
 sg13g2_fill_1 FILLER_9_1875 ();
 sg13g2_fill_1 FILLER_9_1880 ();
 sg13g2_fill_1 FILLER_9_1891 ();
 sg13g2_fill_2 FILLER_9_1902 ();
 sg13g2_fill_1 FILLER_9_1913 ();
 sg13g2_fill_2 FILLER_9_1924 ();
 sg13g2_fill_1 FILLER_9_1926 ();
 sg13g2_decap_8 FILLER_9_1936 ();
 sg13g2_fill_2 FILLER_9_1943 ();
 sg13g2_fill_1 FILLER_9_2047 ();
 sg13g2_decap_8 FILLER_9_2118 ();
 sg13g2_fill_1 FILLER_9_2125 ();
 sg13g2_decap_8 FILLER_9_2143 ();
 sg13g2_decap_4 FILLER_9_2150 ();
 sg13g2_fill_1 FILLER_9_2154 ();
 sg13g2_fill_1 FILLER_9_2165 ();
 sg13g2_fill_2 FILLER_9_2219 ();
 sg13g2_fill_1 FILLER_9_2221 ();
 sg13g2_decap_4 FILLER_9_2226 ();
 sg13g2_fill_2 FILLER_9_2243 ();
 sg13g2_fill_2 FILLER_9_2298 ();
 sg13g2_fill_2 FILLER_9_2321 ();
 sg13g2_fill_1 FILLER_9_2343 ();
 sg13g2_decap_4 FILLER_9_2365 ();
 sg13g2_fill_2 FILLER_9_2395 ();
 sg13g2_fill_1 FILLER_9_2441 ();
 sg13g2_fill_1 FILLER_9_2468 ();
 sg13g2_fill_2 FILLER_9_2479 ();
 sg13g2_fill_2 FILLER_9_2485 ();
 sg13g2_fill_1 FILLER_9_2487 ();
 sg13g2_fill_2 FILLER_9_2498 ();
 sg13g2_fill_1 FILLER_9_2500 ();
 sg13g2_fill_2 FILLER_9_2511 ();
 sg13g2_decap_8 FILLER_9_2517 ();
 sg13g2_decap_8 FILLER_9_2524 ();
 sg13g2_decap_8 FILLER_9_2531 ();
 sg13g2_decap_8 FILLER_9_2574 ();
 sg13g2_decap_8 FILLER_9_2581 ();
 sg13g2_decap_8 FILLER_9_2588 ();
 sg13g2_decap_8 FILLER_9_2595 ();
 sg13g2_decap_8 FILLER_9_2602 ();
 sg13g2_decap_8 FILLER_9_2609 ();
 sg13g2_decap_8 FILLER_9_2616 ();
 sg13g2_decap_8 FILLER_9_2623 ();
 sg13g2_decap_8 FILLER_9_2630 ();
 sg13g2_decap_8 FILLER_9_2637 ();
 sg13g2_decap_8 FILLER_9_2644 ();
 sg13g2_decap_8 FILLER_9_2651 ();
 sg13g2_decap_8 FILLER_9_2658 ();
 sg13g2_decap_4 FILLER_9_2665 ();
 sg13g2_fill_1 FILLER_9_2669 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_41 ();
 sg13g2_decap_8 FILLER_10_48 ();
 sg13g2_decap_8 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_decap_4 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_74 ();
 sg13g2_fill_2 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_82 ();
 sg13g2_decap_8 FILLER_10_87 ();
 sg13g2_fill_2 FILLER_10_94 ();
 sg13g2_decap_4 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_110 ();
 sg13g2_fill_1 FILLER_10_121 ();
 sg13g2_decap_4 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_153 ();
 sg13g2_fill_2 FILLER_10_159 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_fill_1 FILLER_10_218 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_4 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_4 FILLER_10_363 ();
 sg13g2_fill_2 FILLER_10_429 ();
 sg13g2_fill_2 FILLER_10_444 ();
 sg13g2_fill_1 FILLER_10_446 ();
 sg13g2_fill_2 FILLER_10_513 ();
 sg13g2_fill_1 FILLER_10_515 ();
 sg13g2_fill_1 FILLER_10_528 ();
 sg13g2_fill_2 FILLER_10_549 ();
 sg13g2_fill_1 FILLER_10_555 ();
 sg13g2_fill_2 FILLER_10_560 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_fill_2 FILLER_10_616 ();
 sg13g2_fill_1 FILLER_10_631 ();
 sg13g2_fill_1 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_fill_1 FILLER_10_653 ();
 sg13g2_decap_4 FILLER_10_692 ();
 sg13g2_fill_2 FILLER_10_696 ();
 sg13g2_fill_2 FILLER_10_702 ();
 sg13g2_fill_2 FILLER_10_713 ();
 sg13g2_fill_2 FILLER_10_723 ();
 sg13g2_fill_1 FILLER_10_730 ();
 sg13g2_decap_4 FILLER_10_735 ();
 sg13g2_fill_2 FILLER_10_739 ();
 sg13g2_fill_1 FILLER_10_745 ();
 sg13g2_decap_4 FILLER_10_763 ();
 sg13g2_fill_2 FILLER_10_767 ();
 sg13g2_fill_2 FILLER_10_777 ();
 sg13g2_fill_1 FILLER_10_792 ();
 sg13g2_decap_8 FILLER_10_824 ();
 sg13g2_decap_4 FILLER_10_831 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_fill_1 FILLER_10_868 ();
 sg13g2_fill_1 FILLER_10_889 ();
 sg13g2_decap_4 FILLER_10_915 ();
 sg13g2_fill_2 FILLER_10_919 ();
 sg13g2_fill_2 FILLER_10_929 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_fill_1 FILLER_10_942 ();
 sg13g2_fill_2 FILLER_10_1017 ();
 sg13g2_fill_1 FILLER_10_1019 ();
 sg13g2_fill_1 FILLER_10_1034 ();
 sg13g2_fill_2 FILLER_10_1040 ();
 sg13g2_fill_2 FILLER_10_1052 ();
 sg13g2_fill_2 FILLER_10_1090 ();
 sg13g2_fill_2 FILLER_10_1102 ();
 sg13g2_fill_2 FILLER_10_1130 ();
 sg13g2_fill_1 FILLER_10_1158 ();
 sg13g2_fill_2 FILLER_10_1169 ();
 sg13g2_decap_8 FILLER_10_1175 ();
 sg13g2_decap_4 FILLER_10_1182 ();
 sg13g2_fill_2 FILLER_10_1186 ();
 sg13g2_fill_2 FILLER_10_1198 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_fill_1 FILLER_10_1211 ();
 sg13g2_fill_2 FILLER_10_1225 ();
 sg13g2_fill_1 FILLER_10_1232 ();
 sg13g2_decap_4 FILLER_10_1281 ();
 sg13g2_fill_2 FILLER_10_1285 ();
 sg13g2_fill_2 FILLER_10_1297 ();
 sg13g2_fill_1 FILLER_10_1299 ();
 sg13g2_fill_1 FILLER_10_1317 ();
 sg13g2_fill_1 FILLER_10_1328 ();
 sg13g2_fill_1 FILLER_10_1334 ();
 sg13g2_fill_2 FILLER_10_1361 ();
 sg13g2_fill_1 FILLER_10_1363 ();
 sg13g2_fill_1 FILLER_10_1384 ();
 sg13g2_fill_1 FILLER_10_1406 ();
 sg13g2_fill_2 FILLER_10_1425 ();
 sg13g2_fill_2 FILLER_10_1442 ();
 sg13g2_fill_2 FILLER_10_1454 ();
 sg13g2_decap_4 FILLER_10_1460 ();
 sg13g2_decap_8 FILLER_10_1472 ();
 sg13g2_fill_1 FILLER_10_1489 ();
 sg13g2_fill_2 FILLER_10_1547 ();
 sg13g2_fill_1 FILLER_10_1608 ();
 sg13g2_fill_2 FILLER_10_1614 ();
 sg13g2_fill_2 FILLER_10_1629 ();
 sg13g2_decap_4 FILLER_10_1660 ();
 sg13g2_fill_1 FILLER_10_1664 ();
 sg13g2_fill_1 FILLER_10_1674 ();
 sg13g2_fill_1 FILLER_10_1683 ();
 sg13g2_fill_2 FILLER_10_1688 ();
 sg13g2_decap_8 FILLER_10_1741 ();
 sg13g2_decap_4 FILLER_10_1748 ();
 sg13g2_fill_2 FILLER_10_1752 ();
 sg13g2_fill_1 FILLER_10_1769 ();
 sg13g2_fill_1 FILLER_10_1774 ();
 sg13g2_decap_4 FILLER_10_1788 ();
 sg13g2_fill_2 FILLER_10_1796 ();
 sg13g2_fill_1 FILLER_10_1798 ();
 sg13g2_decap_8 FILLER_10_1808 ();
 sg13g2_fill_2 FILLER_10_1819 ();
 sg13g2_fill_2 FILLER_10_1825 ();
 sg13g2_decap_4 FILLER_10_1857 ();
 sg13g2_decap_8 FILLER_10_1865 ();
 sg13g2_fill_2 FILLER_10_1872 ();
 sg13g2_fill_1 FILLER_10_1874 ();
 sg13g2_decap_8 FILLER_10_1931 ();
 sg13g2_decap_8 FILLER_10_1948 ();
 sg13g2_decap_8 FILLER_10_1955 ();
 sg13g2_decap_4 FILLER_10_1962 ();
 sg13g2_fill_2 FILLER_10_1987 ();
 sg13g2_fill_1 FILLER_10_2041 ();
 sg13g2_fill_2 FILLER_10_2111 ();
 sg13g2_fill_2 FILLER_10_2155 ();
 sg13g2_decap_8 FILLER_10_2203 ();
 sg13g2_fill_2 FILLER_10_2210 ();
 sg13g2_fill_1 FILLER_10_2259 ();
 sg13g2_fill_2 FILLER_10_2268 ();
 sg13g2_fill_1 FILLER_10_2288 ();
 sg13g2_fill_2 FILLER_10_2349 ();
 sg13g2_fill_2 FILLER_10_2369 ();
 sg13g2_fill_2 FILLER_10_2417 ();
 sg13g2_decap_8 FILLER_10_2422 ();
 sg13g2_fill_2 FILLER_10_2429 ();
 sg13g2_decap_8 FILLER_10_2434 ();
 sg13g2_decap_8 FILLER_10_2441 ();
 sg13g2_fill_2 FILLER_10_2448 ();
 sg13g2_fill_1 FILLER_10_2450 ();
 sg13g2_fill_2 FILLER_10_2485 ();
 sg13g2_fill_1 FILLER_10_2487 ();
 sg13g2_decap_8 FILLER_10_2492 ();
 sg13g2_decap_4 FILLER_10_2499 ();
 sg13g2_decap_8 FILLER_10_2524 ();
 sg13g2_decap_8 FILLER_10_2531 ();
 sg13g2_fill_2 FILLER_10_2538 ();
 sg13g2_fill_1 FILLER_10_2540 ();
 sg13g2_decap_8 FILLER_10_2562 ();
 sg13g2_decap_8 FILLER_10_2569 ();
 sg13g2_decap_8 FILLER_10_2576 ();
 sg13g2_decap_8 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2590 ();
 sg13g2_decap_8 FILLER_10_2597 ();
 sg13g2_decap_8 FILLER_10_2604 ();
 sg13g2_decap_8 FILLER_10_2611 ();
 sg13g2_decap_8 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2625 ();
 sg13g2_decap_8 FILLER_10_2632 ();
 sg13g2_decap_8 FILLER_10_2639 ();
 sg13g2_decap_8 FILLER_10_2646 ();
 sg13g2_decap_8 FILLER_10_2653 ();
 sg13g2_decap_8 FILLER_10_2660 ();
 sg13g2_fill_2 FILLER_10_2667 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_decap_4 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_fill_1 FILLER_11_262 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_decap_4 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_decap_4 FILLER_11_428 ();
 sg13g2_decap_4 FILLER_11_440 ();
 sg13g2_fill_2 FILLER_11_444 ();
 sg13g2_decap_4 FILLER_11_460 ();
 sg13g2_fill_1 FILLER_11_464 ();
 sg13g2_fill_2 FILLER_11_475 ();
 sg13g2_fill_2 FILLER_11_487 ();
 sg13g2_fill_1 FILLER_11_489 ();
 sg13g2_fill_2 FILLER_11_516 ();
 sg13g2_fill_1 FILLER_11_518 ();
 sg13g2_fill_2 FILLER_11_524 ();
 sg13g2_fill_1 FILLER_11_526 ();
 sg13g2_fill_2 FILLER_11_553 ();
 sg13g2_fill_1 FILLER_11_560 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_decap_4 FILLER_11_575 ();
 sg13g2_fill_2 FILLER_11_579 ();
 sg13g2_fill_1 FILLER_11_636 ();
 sg13g2_fill_2 FILLER_11_672 ();
 sg13g2_fill_1 FILLER_11_674 ();
 sg13g2_fill_1 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_fill_1 FILLER_11_789 ();
 sg13g2_fill_1 FILLER_11_794 ();
 sg13g2_decap_4 FILLER_11_825 ();
 sg13g2_fill_2 FILLER_11_829 ();
 sg13g2_decap_4 FILLER_11_835 ();
 sg13g2_fill_2 FILLER_11_839 ();
 sg13g2_decap_4 FILLER_11_845 ();
 sg13g2_fill_1 FILLER_11_849 ();
 sg13g2_fill_2 FILLER_11_906 ();
 sg13g2_fill_1 FILLER_11_908 ();
 sg13g2_decap_8 FILLER_11_913 ();
 sg13g2_decap_4 FILLER_11_920 ();
 sg13g2_fill_2 FILLER_11_947 ();
 sg13g2_fill_1 FILLER_11_949 ();
 sg13g2_decap_4 FILLER_11_976 ();
 sg13g2_fill_1 FILLER_11_1014 ();
 sg13g2_fill_2 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1030 ();
 sg13g2_fill_1 FILLER_11_1061 ();
 sg13g2_decap_4 FILLER_11_1067 ();
 sg13g2_fill_2 FILLER_11_1071 ();
 sg13g2_fill_2 FILLER_11_1119 ();
 sg13g2_fill_1 FILLER_11_1121 ();
 sg13g2_fill_2 FILLER_11_1126 ();
 sg13g2_decap_4 FILLER_11_1146 ();
 sg13g2_decap_4 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1190 ();
 sg13g2_decap_8 FILLER_11_1197 ();
 sg13g2_fill_2 FILLER_11_1204 ();
 sg13g2_fill_1 FILLER_11_1206 ();
 sg13g2_fill_2 FILLER_11_1240 ();
 sg13g2_fill_2 FILLER_11_1272 ();
 sg13g2_fill_2 FILLER_11_1350 ();
 sg13g2_fill_1 FILLER_11_1352 ();
 sg13g2_decap_4 FILLER_11_1371 ();
 sg13g2_fill_1 FILLER_11_1375 ();
 sg13g2_fill_1 FILLER_11_1394 ();
 sg13g2_fill_2 FILLER_11_1401 ();
 sg13g2_fill_2 FILLER_11_1413 ();
 sg13g2_fill_2 FILLER_11_1446 ();
 sg13g2_fill_1 FILLER_11_1524 ();
 sg13g2_fill_1 FILLER_11_1535 ();
 sg13g2_fill_1 FILLER_11_1541 ();
 sg13g2_fill_1 FILLER_11_1548 ();
 sg13g2_fill_2 FILLER_11_1553 ();
 sg13g2_fill_2 FILLER_11_1579 ();
 sg13g2_fill_1 FILLER_11_1590 ();
 sg13g2_fill_1 FILLER_11_1595 ();
 sg13g2_fill_1 FILLER_11_1625 ();
 sg13g2_fill_2 FILLER_11_1631 ();
 sg13g2_fill_2 FILLER_11_1642 ();
 sg13g2_fill_2 FILLER_11_1649 ();
 sg13g2_fill_1 FILLER_11_1651 ();
 sg13g2_decap_4 FILLER_11_1665 ();
 sg13g2_fill_2 FILLER_11_1673 ();
 sg13g2_fill_2 FILLER_11_1701 ();
 sg13g2_fill_1 FILLER_11_1703 ();
 sg13g2_fill_2 FILLER_11_1730 ();
 sg13g2_fill_2 FILLER_11_1736 ();
 sg13g2_fill_1 FILLER_11_1738 ();
 sg13g2_decap_4 FILLER_11_1749 ();
 sg13g2_decap_8 FILLER_11_1794 ();
 sg13g2_decap_8 FILLER_11_1801 ();
 sg13g2_decap_8 FILLER_11_1808 ();
 sg13g2_decap_8 FILLER_11_1845 ();
 sg13g2_fill_2 FILLER_11_1852 ();
 sg13g2_decap_4 FILLER_11_1880 ();
 sg13g2_fill_2 FILLER_11_1965 ();
 sg13g2_decap_4 FILLER_11_1971 ();
 sg13g2_decap_8 FILLER_11_1983 ();
 sg13g2_fill_2 FILLER_11_1994 ();
 sg13g2_fill_2 FILLER_11_2014 ();
 sg13g2_fill_2 FILLER_11_2026 ();
 sg13g2_fill_1 FILLER_11_2028 ();
 sg13g2_decap_4 FILLER_11_2055 ();
 sg13g2_fill_2 FILLER_11_2068 ();
 sg13g2_fill_2 FILLER_11_2080 ();
 sg13g2_fill_2 FILLER_11_2086 ();
 sg13g2_fill_1 FILLER_11_2088 ();
 sg13g2_fill_1 FILLER_11_2099 ();
 sg13g2_fill_1 FILLER_11_2104 ();
 sg13g2_fill_1 FILLER_11_2141 ();
 sg13g2_decap_8 FILLER_11_2146 ();
 sg13g2_fill_2 FILLER_11_2153 ();
 sg13g2_fill_1 FILLER_11_2155 ();
 sg13g2_decap_4 FILLER_11_2161 ();
 sg13g2_fill_1 FILLER_11_2187 ();
 sg13g2_decap_4 FILLER_11_2206 ();
 sg13g2_fill_2 FILLER_11_2254 ();
 sg13g2_decap_4 FILLER_11_2305 ();
 sg13g2_decap_8 FILLER_11_2330 ();
 sg13g2_fill_1 FILLER_11_2337 ();
 sg13g2_fill_1 FILLER_11_2385 ();
 sg13g2_fill_1 FILLER_11_2435 ();
 sg13g2_decap_8 FILLER_11_2462 ();
 sg13g2_fill_2 FILLER_11_2469 ();
 sg13g2_decap_4 FILLER_11_2528 ();
 sg13g2_fill_1 FILLER_11_2532 ();
 sg13g2_fill_1 FILLER_11_2543 ();
 sg13g2_decap_8 FILLER_11_2574 ();
 sg13g2_decap_8 FILLER_11_2581 ();
 sg13g2_decap_8 FILLER_11_2588 ();
 sg13g2_decap_8 FILLER_11_2595 ();
 sg13g2_decap_8 FILLER_11_2602 ();
 sg13g2_decap_8 FILLER_11_2609 ();
 sg13g2_decap_8 FILLER_11_2616 ();
 sg13g2_decap_8 FILLER_11_2623 ();
 sg13g2_decap_8 FILLER_11_2630 ();
 sg13g2_decap_8 FILLER_11_2637 ();
 sg13g2_decap_8 FILLER_11_2644 ();
 sg13g2_decap_8 FILLER_11_2651 ();
 sg13g2_decap_8 FILLER_11_2658 ();
 sg13g2_decap_4 FILLER_11_2665 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_decap_8 FILLER_12_22 ();
 sg13g2_fill_1 FILLER_12_29 ();
 sg13g2_decap_4 FILLER_12_34 ();
 sg13g2_fill_1 FILLER_12_38 ();
 sg13g2_decap_4 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_118 ();
 sg13g2_fill_2 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_fill_1 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_decap_4 FILLER_12_432 ();
 sg13g2_fill_2 FILLER_12_509 ();
 sg13g2_fill_1 FILLER_12_541 ();
 sg13g2_decap_8 FILLER_12_568 ();
 sg13g2_decap_8 FILLER_12_575 ();
 sg13g2_fill_2 FILLER_12_591 ();
 sg13g2_fill_1 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_675 ();
 sg13g2_fill_1 FILLER_12_682 ();
 sg13g2_fill_2 FILLER_12_709 ();
 sg13g2_fill_1 FILLER_12_711 ();
 sg13g2_fill_1 FILLER_12_725 ();
 sg13g2_fill_2 FILLER_12_752 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_fill_1 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_fill_1 FILLER_12_813 ();
 sg13g2_decap_4 FILLER_12_840 ();
 sg13g2_fill_1 FILLER_12_844 ();
 sg13g2_fill_1 FILLER_12_875 ();
 sg13g2_fill_1 FILLER_12_884 ();
 sg13g2_fill_1 FILLER_12_911 ();
 sg13g2_fill_1 FILLER_12_916 ();
 sg13g2_fill_1 FILLER_12_940 ();
 sg13g2_fill_2 FILLER_12_972 ();
 sg13g2_decap_4 FILLER_12_984 ();
 sg13g2_fill_2 FILLER_12_988 ();
 sg13g2_fill_2 FILLER_12_1024 ();
 sg13g2_fill_1 FILLER_12_1026 ();
 sg13g2_fill_2 FILLER_12_1053 ();
 sg13g2_fill_2 FILLER_12_1107 ();
 sg13g2_fill_1 FILLER_12_1109 ();
 sg13g2_decap_4 FILLER_12_1130 ();
 sg13g2_fill_2 FILLER_12_1134 ();
 sg13g2_decap_4 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1170 ();
 sg13g2_decap_4 FILLER_12_1177 ();
 sg13g2_decap_8 FILLER_12_1185 ();
 sg13g2_fill_1 FILLER_12_1192 ();
 sg13g2_fill_2 FILLER_12_1207 ();
 sg13g2_fill_1 FILLER_12_1209 ();
 sg13g2_decap_8 FILLER_12_1219 ();
 sg13g2_decap_8 FILLER_12_1226 ();
 sg13g2_decap_8 FILLER_12_1233 ();
 sg13g2_decap_4 FILLER_12_1240 ();
 sg13g2_fill_1 FILLER_12_1244 ();
 sg13g2_fill_2 FILLER_12_1250 ();
 sg13g2_fill_1 FILLER_12_1252 ();
 sg13g2_fill_2 FILLER_12_1268 ();
 sg13g2_fill_1 FILLER_12_1270 ();
 sg13g2_fill_1 FILLER_12_1276 ();
 sg13g2_decap_4 FILLER_12_1327 ();
 sg13g2_fill_1 FILLER_12_1331 ();
 sg13g2_fill_1 FILLER_12_1372 ();
 sg13g2_fill_1 FILLER_12_1408 ();
 sg13g2_fill_1 FILLER_12_1414 ();
 sg13g2_fill_2 FILLER_12_1422 ();
 sg13g2_fill_1 FILLER_12_1430 ();
 sg13g2_fill_2 FILLER_12_1436 ();
 sg13g2_fill_2 FILLER_12_1486 ();
 sg13g2_fill_1 FILLER_12_1549 ();
 sg13g2_fill_1 FILLER_12_1581 ();
 sg13g2_decap_4 FILLER_12_1673 ();
 sg13g2_fill_2 FILLER_12_1677 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_4 FILLER_12_1701 ();
 sg13g2_fill_2 FILLER_12_1709 ();
 sg13g2_decap_4 FILLER_12_1715 ();
 sg13g2_fill_1 FILLER_12_1719 ();
 sg13g2_fill_1 FILLER_12_1724 ();
 sg13g2_decap_8 FILLER_12_1751 ();
 sg13g2_fill_2 FILLER_12_1758 ();
 sg13g2_fill_1 FILLER_12_1760 ();
 sg13g2_fill_2 FILLER_12_1791 ();
 sg13g2_fill_1 FILLER_12_1922 ();
 sg13g2_fill_2 FILLER_12_1949 ();
 sg13g2_fill_1 FILLER_12_1951 ();
 sg13g2_fill_1 FILLER_12_1978 ();
 sg13g2_fill_1 FILLER_12_2021 ();
 sg13g2_fill_1 FILLER_12_2037 ();
 sg13g2_decap_4 FILLER_12_2042 ();
 sg13g2_fill_2 FILLER_12_2046 ();
 sg13g2_fill_1 FILLER_12_2083 ();
 sg13g2_fill_1 FILLER_12_2120 ();
 sg13g2_decap_4 FILLER_12_2129 ();
 sg13g2_decap_4 FILLER_12_2159 ();
 sg13g2_decap_4 FILLER_12_2167 ();
 sg13g2_fill_1 FILLER_12_2171 ();
 sg13g2_decap_4 FILLER_12_2248 ();
 sg13g2_fill_1 FILLER_12_2252 ();
 sg13g2_decap_8 FILLER_12_2274 ();
 sg13g2_fill_1 FILLER_12_2281 ();
 sg13g2_decap_8 FILLER_12_2302 ();
 sg13g2_decap_8 FILLER_12_2309 ();
 sg13g2_decap_8 FILLER_12_2316 ();
 sg13g2_decap_8 FILLER_12_2323 ();
 sg13g2_decap_4 FILLER_12_2330 ();
 sg13g2_fill_2 FILLER_12_2334 ();
 sg13g2_fill_1 FILLER_12_2362 ();
 sg13g2_decap_4 FILLER_12_2376 ();
 sg13g2_fill_2 FILLER_12_2380 ();
 sg13g2_fill_1 FILLER_12_2396 ();
 sg13g2_fill_2 FILLER_12_2402 ();
 sg13g2_fill_1 FILLER_12_2404 ();
 sg13g2_fill_1 FILLER_12_2434 ();
 sg13g2_decap_8 FILLER_12_2565 ();
 sg13g2_decap_8 FILLER_12_2572 ();
 sg13g2_decap_8 FILLER_12_2579 ();
 sg13g2_decap_8 FILLER_12_2586 ();
 sg13g2_decap_8 FILLER_12_2593 ();
 sg13g2_decap_8 FILLER_12_2600 ();
 sg13g2_decap_8 FILLER_12_2607 ();
 sg13g2_decap_8 FILLER_12_2614 ();
 sg13g2_decap_8 FILLER_12_2621 ();
 sg13g2_decap_8 FILLER_12_2628 ();
 sg13g2_decap_8 FILLER_12_2635 ();
 sg13g2_decap_8 FILLER_12_2642 ();
 sg13g2_decap_8 FILLER_12_2649 ();
 sg13g2_decap_8 FILLER_12_2656 ();
 sg13g2_decap_8 FILLER_12_2663 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_1 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_95 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_fill_2 FILLER_13_382 ();
 sg13g2_fill_2 FILLER_13_410 ();
 sg13g2_fill_2 FILLER_13_438 ();
 sg13g2_fill_1 FILLER_13_440 ();
 sg13g2_fill_2 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_483 ();
 sg13g2_fill_1 FILLER_13_494 ();
 sg13g2_fill_1 FILLER_13_499 ();
 sg13g2_fill_1 FILLER_13_572 ();
 sg13g2_fill_1 FILLER_13_577 ();
 sg13g2_fill_2 FILLER_13_586 ();
 sg13g2_fill_1 FILLER_13_588 ();
 sg13g2_fill_2 FILLER_13_662 ();
 sg13g2_decap_4 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_693 ();
 sg13g2_decap_4 FILLER_13_699 ();
 sg13g2_fill_2 FILLER_13_755 ();
 sg13g2_fill_1 FILLER_13_757 ();
 sg13g2_decap_4 FILLER_13_788 ();
 sg13g2_decap_4 FILLER_13_818 ();
 sg13g2_fill_1 FILLER_13_822 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_fill_1 FILLER_13_834 ();
 sg13g2_fill_2 FILLER_13_840 ();
 sg13g2_fill_1 FILLER_13_842 ();
 sg13g2_fill_1 FILLER_13_871 ();
 sg13g2_fill_1 FILLER_13_897 ();
 sg13g2_decap_8 FILLER_13_902 ();
 sg13g2_decap_8 FILLER_13_909 ();
 sg13g2_decap_4 FILLER_13_916 ();
 sg13g2_fill_1 FILLER_13_920 ();
 sg13g2_decap_4 FILLER_13_925 ();
 sg13g2_fill_1 FILLER_13_929 ();
 sg13g2_decap_8 FILLER_13_985 ();
 sg13g2_fill_2 FILLER_13_992 ();
 sg13g2_fill_1 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_fill_1 FILLER_13_1012 ();
 sg13g2_fill_2 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1033 ();
 sg13g2_fill_2 FILLER_13_1047 ();
 sg13g2_fill_2 FILLER_13_1055 ();
 sg13g2_fill_1 FILLER_13_1057 ();
 sg13g2_fill_2 FILLER_13_1062 ();
 sg13g2_fill_1 FILLER_13_1064 ();
 sg13g2_fill_2 FILLER_13_1069 ();
 sg13g2_fill_1 FILLER_13_1075 ();
 sg13g2_fill_2 FILLER_13_1131 ();
 sg13g2_fill_1 FILLER_13_1163 ();
 sg13g2_fill_1 FILLER_13_1200 ();
 sg13g2_decap_8 FILLER_13_1212 ();
 sg13g2_decap_8 FILLER_13_1219 ();
 sg13g2_fill_2 FILLER_13_1226 ();
 sg13g2_fill_2 FILLER_13_1240 ();
 sg13g2_decap_4 FILLER_13_1255 ();
 sg13g2_fill_1 FILLER_13_1259 ();
 sg13g2_fill_2 FILLER_13_1291 ();
 sg13g2_decap_4 FILLER_13_1308 ();
 sg13g2_fill_1 FILLER_13_1312 ();
 sg13g2_fill_1 FILLER_13_1333 ();
 sg13g2_decap_4 FILLER_13_1340 ();
 sg13g2_fill_1 FILLER_13_1355 ();
 sg13g2_fill_2 FILLER_13_1361 ();
 sg13g2_fill_1 FILLER_13_1408 ();
 sg13g2_decap_4 FILLER_13_1430 ();
 sg13g2_decap_4 FILLER_13_1449 ();
 sg13g2_fill_1 FILLER_13_1453 ();
 sg13g2_fill_2 FILLER_13_1464 ();
 sg13g2_fill_1 FILLER_13_1466 ();
 sg13g2_fill_1 FILLER_13_1512 ();
 sg13g2_fill_1 FILLER_13_1518 ();
 sg13g2_fill_2 FILLER_13_1523 ();
 sg13g2_fill_1 FILLER_13_1525 ();
 sg13g2_fill_2 FILLER_13_1537 ();
 sg13g2_fill_2 FILLER_13_1545 ();
 sg13g2_fill_2 FILLER_13_1620 ();
 sg13g2_fill_2 FILLER_13_1634 ();
 sg13g2_fill_1 FILLER_13_1636 ();
 sg13g2_fill_2 FILLER_13_1663 ();
 sg13g2_fill_2 FILLER_13_1670 ();
 sg13g2_fill_2 FILLER_13_1698 ();
 sg13g2_decap_8 FILLER_13_1752 ();
 sg13g2_decap_8 FILLER_13_1759 ();
 sg13g2_fill_1 FILLER_13_1766 ();
 sg13g2_decap_4 FILLER_13_1806 ();
 sg13g2_fill_1 FILLER_13_1810 ();
 sg13g2_fill_1 FILLER_13_1815 ();
 sg13g2_fill_1 FILLER_13_1826 ();
 sg13g2_decap_8 FILLER_13_1831 ();
 sg13g2_decap_8 FILLER_13_1838 ();
 sg13g2_decap_4 FILLER_13_1845 ();
 sg13g2_decap_4 FILLER_13_1967 ();
 sg13g2_fill_1 FILLER_13_1971 ();
 sg13g2_fill_2 FILLER_13_2006 ();
 sg13g2_fill_2 FILLER_13_2016 ();
 sg13g2_fill_1 FILLER_13_2018 ();
 sg13g2_fill_1 FILLER_13_2029 ();
 sg13g2_fill_1 FILLER_13_2035 ();
 sg13g2_fill_1 FILLER_13_2046 ();
 sg13g2_fill_1 FILLER_13_2073 ();
 sg13g2_fill_1 FILLER_13_2100 ();
 sg13g2_decap_8 FILLER_13_2202 ();
 sg13g2_fill_2 FILLER_13_2209 ();
 sg13g2_fill_1 FILLER_13_2211 ();
 sg13g2_fill_1 FILLER_13_2216 ();
 sg13g2_decap_8 FILLER_13_2222 ();
 sg13g2_decap_4 FILLER_13_2229 ();
 sg13g2_decap_4 FILLER_13_2241 ();
 sg13g2_fill_1 FILLER_13_2245 ();
 sg13g2_decap_8 FILLER_13_2267 ();
 sg13g2_decap_4 FILLER_13_2274 ();
 sg13g2_fill_2 FILLER_13_2278 ();
 sg13g2_decap_4 FILLER_13_2290 ();
 sg13g2_decap_8 FILLER_13_2315 ();
 sg13g2_decap_4 FILLER_13_2322 ();
 sg13g2_fill_2 FILLER_13_2326 ();
 sg13g2_fill_2 FILLER_13_2379 ();
 sg13g2_fill_2 FILLER_13_2422 ();
 sg13g2_fill_2 FILLER_13_2509 ();
 sg13g2_fill_2 FILLER_13_2577 ();
 sg13g2_decap_8 FILLER_13_2583 ();
 sg13g2_decap_8 FILLER_13_2590 ();
 sg13g2_decap_8 FILLER_13_2597 ();
 sg13g2_decap_8 FILLER_13_2604 ();
 sg13g2_decap_8 FILLER_13_2611 ();
 sg13g2_decap_8 FILLER_13_2618 ();
 sg13g2_decap_8 FILLER_13_2625 ();
 sg13g2_decap_8 FILLER_13_2632 ();
 sg13g2_decap_8 FILLER_13_2639 ();
 sg13g2_decap_8 FILLER_13_2646 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_fill_2 FILLER_13_2667 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_36 ();
 sg13g2_fill_2 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_4 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_4 FILLER_14_377 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_fill_2 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_443 ();
 sg13g2_fill_2 FILLER_14_484 ();
 sg13g2_fill_1 FILLER_14_531 ();
 sg13g2_fill_2 FILLER_14_549 ();
 sg13g2_fill_2 FILLER_14_555 ();
 sg13g2_fill_2 FILLER_14_562 ();
 sg13g2_fill_1 FILLER_14_564 ();
 sg13g2_fill_1 FILLER_14_636 ();
 sg13g2_fill_2 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_4 FILLER_14_679 ();
 sg13g2_fill_2 FILLER_14_683 ();
 sg13g2_fill_2 FILLER_14_721 ();
 sg13g2_decap_4 FILLER_14_752 ();
 sg13g2_fill_1 FILLER_14_756 ();
 sg13g2_decap_4 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_769 ();
 sg13g2_fill_2 FILLER_14_776 ();
 sg13g2_decap_8 FILLER_14_787 ();
 sg13g2_decap_4 FILLER_14_794 ();
 sg13g2_decap_4 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_4 FILLER_14_824 ();
 sg13g2_fill_2 FILLER_14_828 ();
 sg13g2_decap_4 FILLER_14_874 ();
 sg13g2_fill_2 FILLER_14_888 ();
 sg13g2_decap_8 FILLER_14_899 ();
 sg13g2_decap_4 FILLER_14_910 ();
 sg13g2_fill_1 FILLER_14_918 ();
 sg13g2_fill_1 FILLER_14_923 ();
 sg13g2_fill_2 FILLER_14_928 ();
 sg13g2_fill_2 FILLER_14_957 ();
 sg13g2_fill_1 FILLER_14_968 ();
 sg13g2_fill_1 FILLER_14_973 ();
 sg13g2_fill_2 FILLER_14_1020 ();
 sg13g2_fill_1 FILLER_14_1037 ();
 sg13g2_decap_8 FILLER_14_1047 ();
 sg13g2_fill_2 FILLER_14_1054 ();
 sg13g2_fill_1 FILLER_14_1056 ();
 sg13g2_fill_1 FILLER_14_1061 ();
 sg13g2_fill_2 FILLER_14_1067 ();
 sg13g2_fill_2 FILLER_14_1082 ();
 sg13g2_fill_1 FILLER_14_1139 ();
 sg13g2_fill_1 FILLER_14_1145 ();
 sg13g2_fill_1 FILLER_14_1150 ();
 sg13g2_fill_1 FILLER_14_1177 ();
 sg13g2_decap_8 FILLER_14_1188 ();
 sg13g2_fill_1 FILLER_14_1195 ();
 sg13g2_fill_1 FILLER_14_1201 ();
 sg13g2_fill_1 FILLER_14_1230 ();
 sg13g2_fill_2 FILLER_14_1257 ();
 sg13g2_fill_1 FILLER_14_1264 ();
 sg13g2_fill_1 FILLER_14_1269 ();
 sg13g2_fill_2 FILLER_14_1276 ();
 sg13g2_fill_1 FILLER_14_1278 ();
 sg13g2_decap_8 FILLER_14_1290 ();
 sg13g2_fill_1 FILLER_14_1303 ();
 sg13g2_fill_1 FILLER_14_1312 ();
 sg13g2_fill_2 FILLER_14_1317 ();
 sg13g2_fill_1 FILLER_14_1319 ();
 sg13g2_decap_8 FILLER_14_1325 ();
 sg13g2_fill_2 FILLER_14_1332 ();
 sg13g2_fill_1 FILLER_14_1334 ();
 sg13g2_fill_2 FILLER_14_1377 ();
 sg13g2_fill_2 FILLER_14_1394 ();
 sg13g2_fill_1 FILLER_14_1396 ();
 sg13g2_decap_8 FILLER_14_1440 ();
 sg13g2_decap_8 FILLER_14_1447 ();
 sg13g2_fill_1 FILLER_14_1454 ();
 sg13g2_decap_8 FILLER_14_1474 ();
 sg13g2_fill_2 FILLER_14_1481 ();
 sg13g2_fill_1 FILLER_14_1483 ();
 sg13g2_decap_8 FILLER_14_1488 ();
 sg13g2_decap_4 FILLER_14_1499 ();
 sg13g2_fill_2 FILLER_14_1503 ();
 sg13g2_fill_2 FILLER_14_1510 ();
 sg13g2_fill_2 FILLER_14_1516 ();
 sg13g2_fill_1 FILLER_14_1518 ();
 sg13g2_fill_2 FILLER_14_1533 ();
 sg13g2_fill_1 FILLER_14_1556 ();
 sg13g2_fill_1 FILLER_14_1601 ();
 sg13g2_fill_1 FILLER_14_1623 ();
 sg13g2_fill_2 FILLER_14_1653 ();
 sg13g2_fill_1 FILLER_14_1655 ();
 sg13g2_fill_2 FILLER_14_1671 ();
 sg13g2_decap_4 FILLER_14_1699 ();
 sg13g2_fill_2 FILLER_14_1708 ();
 sg13g2_fill_1 FILLER_14_1710 ();
 sg13g2_fill_2 FILLER_14_1721 ();
 sg13g2_fill_2 FILLER_14_1736 ();
 sg13g2_fill_1 FILLER_14_1738 ();
 sg13g2_decap_8 FILLER_14_1753 ();
 sg13g2_decap_8 FILLER_14_1760 ();
 sg13g2_fill_2 FILLER_14_1767 ();
 sg13g2_fill_1 FILLER_14_1769 ();
 sg13g2_decap_8 FILLER_14_1809 ();
 sg13g2_decap_8 FILLER_14_1816 ();
 sg13g2_fill_2 FILLER_14_1823 ();
 sg13g2_fill_1 FILLER_14_1825 ();
 sg13g2_decap_8 FILLER_14_1836 ();
 sg13g2_decap_8 FILLER_14_1843 ();
 sg13g2_decap_8 FILLER_14_1850 ();
 sg13g2_fill_2 FILLER_14_1880 ();
 sg13g2_fill_1 FILLER_14_1882 ();
 sg13g2_fill_1 FILLER_14_1926 ();
 sg13g2_decap_4 FILLER_14_1941 ();
 sg13g2_fill_1 FILLER_14_1945 ();
 sg13g2_decap_8 FILLER_14_1956 ();
 sg13g2_decap_8 FILLER_14_1963 ();
 sg13g2_decap_8 FILLER_14_1970 ();
 sg13g2_fill_2 FILLER_14_1977 ();
 sg13g2_fill_2 FILLER_14_1989 ();
 sg13g2_fill_1 FILLER_14_2104 ();
 sg13g2_decap_4 FILLER_14_2122 ();
 sg13g2_fill_1 FILLER_14_2182 ();
 sg13g2_fill_2 FILLER_14_2209 ();
 sg13g2_fill_2 FILLER_14_2221 ();
 sg13g2_fill_2 FILLER_14_2327 ();
 sg13g2_fill_2 FILLER_14_2420 ();
 sg13g2_fill_2 FILLER_14_2429 ();
 sg13g2_fill_2 FILLER_14_2450 ();
 sg13g2_fill_1 FILLER_14_2452 ();
 sg13g2_fill_1 FILLER_14_2463 ();
 sg13g2_decap_8 FILLER_14_2485 ();
 sg13g2_decap_8 FILLER_14_2492 ();
 sg13g2_fill_1 FILLER_14_2499 ();
 sg13g2_fill_2 FILLER_14_2514 ();
 sg13g2_decap_8 FILLER_14_2524 ();
 sg13g2_fill_2 FILLER_14_2531 ();
 sg13g2_fill_1 FILLER_14_2533 ();
 sg13g2_fill_2 FILLER_14_2557 ();
 sg13g2_decap_8 FILLER_14_2585 ();
 sg13g2_decap_8 FILLER_14_2592 ();
 sg13g2_decap_8 FILLER_14_2599 ();
 sg13g2_decap_8 FILLER_14_2606 ();
 sg13g2_decap_8 FILLER_14_2613 ();
 sg13g2_decap_8 FILLER_14_2620 ();
 sg13g2_decap_8 FILLER_14_2627 ();
 sg13g2_decap_8 FILLER_14_2634 ();
 sg13g2_decap_8 FILLER_14_2641 ();
 sg13g2_decap_8 FILLER_14_2648 ();
 sg13g2_decap_8 FILLER_14_2655 ();
 sg13g2_decap_8 FILLER_14_2662 ();
 sg13g2_fill_1 FILLER_14_2669 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_54 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_decap_4 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_419 ();
 sg13g2_decap_8 FILLER_15_433 ();
 sg13g2_decap_8 FILLER_15_440 ();
 sg13g2_fill_2 FILLER_15_447 ();
 sg13g2_decap_4 FILLER_15_461 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_decap_4 FILLER_15_506 ();
 sg13g2_fill_1 FILLER_15_510 ();
 sg13g2_fill_1 FILLER_15_520 ();
 sg13g2_fill_1 FILLER_15_591 ();
 sg13g2_fill_1 FILLER_15_604 ();
 sg13g2_decap_4 FILLER_15_667 ();
 sg13g2_fill_1 FILLER_15_675 ();
 sg13g2_fill_2 FILLER_15_746 ();
 sg13g2_fill_1 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_4 FILLER_15_826 ();
 sg13g2_fill_1 FILLER_15_830 ();
 sg13g2_fill_2 FILLER_15_843 ();
 sg13g2_fill_1 FILLER_15_845 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_fill_2 FILLER_15_883 ();
 sg13g2_fill_1 FILLER_15_885 ();
 sg13g2_fill_1 FILLER_15_890 ();
 sg13g2_fill_2 FILLER_15_895 ();
 sg13g2_fill_1 FILLER_15_897 ();
 sg13g2_fill_1 FILLER_15_938 ();
 sg13g2_fill_2 FILLER_15_965 ();
 sg13g2_fill_2 FILLER_15_1035 ();
 sg13g2_fill_1 FILLER_15_1055 ();
 sg13g2_fill_2 FILLER_15_1082 ();
 sg13g2_fill_2 FILLER_15_1104 ();
 sg13g2_fill_2 FILLER_15_1114 ();
 sg13g2_decap_4 FILLER_15_1120 ();
 sg13g2_decap_4 FILLER_15_1128 ();
 sg13g2_fill_2 FILLER_15_1158 ();
 sg13g2_fill_1 FILLER_15_1160 ();
 sg13g2_fill_1 FILLER_15_1187 ();
 sg13g2_fill_2 FILLER_15_1198 ();
 sg13g2_fill_1 FILLER_15_1203 ();
 sg13g2_fill_1 FILLER_15_1220 ();
 sg13g2_fill_1 FILLER_15_1231 ();
 sg13g2_fill_2 FILLER_15_1250 ();
 sg13g2_fill_1 FILLER_15_1268 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_fill_2 FILLER_15_1305 ();
 sg13g2_fill_1 FILLER_15_1307 ();
 sg13g2_decap_8 FILLER_15_1318 ();
 sg13g2_fill_1 FILLER_15_1325 ();
 sg13g2_fill_2 FILLER_15_1337 ();
 sg13g2_fill_1 FILLER_15_1351 ();
 sg13g2_decap_4 FILLER_15_1377 ();
 sg13g2_decap_8 FILLER_15_1386 ();
 sg13g2_decap_4 FILLER_15_1393 ();
 sg13g2_fill_2 FILLER_15_1410 ();
 sg13g2_fill_1 FILLER_15_1423 ();
 sg13g2_decap_4 FILLER_15_1445 ();
 sg13g2_fill_1 FILLER_15_1463 ();
 sg13g2_decap_8 FILLER_15_1494 ();
 sg13g2_decap_4 FILLER_15_1501 ();
 sg13g2_fill_2 FILLER_15_1539 ();
 sg13g2_fill_1 FILLER_15_1547 ();
 sg13g2_fill_1 FILLER_15_1562 ();
 sg13g2_fill_1 FILLER_15_1589 ();
 sg13g2_fill_1 FILLER_15_1600 ();
 sg13g2_fill_1 FILLER_15_1622 ();
 sg13g2_fill_1 FILLER_15_1675 ();
 sg13g2_fill_1 FILLER_15_1692 ();
 sg13g2_decap_4 FILLER_15_1745 ();
 sg13g2_fill_1 FILLER_15_1749 ();
 sg13g2_fill_1 FILLER_15_1784 ();
 sg13g2_fill_1 FILLER_15_1800 ();
 sg13g2_fill_2 FILLER_15_1805 ();
 sg13g2_fill_1 FILLER_15_1811 ();
 sg13g2_fill_1 FILLER_15_1838 ();
 sg13g2_fill_1 FILLER_15_1860 ();
 sg13g2_fill_2 FILLER_15_1865 ();
 sg13g2_fill_1 FILLER_15_1897 ();
 sg13g2_fill_1 FILLER_15_1908 ();
 sg13g2_fill_2 FILLER_15_1921 ();
 sg13g2_fill_2 FILLER_15_1990 ();
 sg13g2_fill_1 FILLER_15_2023 ();
 sg13g2_fill_1 FILLER_15_2041 ();
 sg13g2_fill_1 FILLER_15_2092 ();
 sg13g2_fill_1 FILLER_15_2112 ();
 sg13g2_fill_1 FILLER_15_2165 ();
 sg13g2_fill_1 FILLER_15_2233 ();
 sg13g2_fill_1 FILLER_15_2283 ();
 sg13g2_decap_4 FILLER_15_2322 ();
 sg13g2_fill_2 FILLER_15_2326 ();
 sg13g2_fill_2 FILLER_15_2338 ();
 sg13g2_decap_8 FILLER_15_2358 ();
 sg13g2_fill_2 FILLER_15_2365 ();
 sg13g2_fill_2 FILLER_15_2377 ();
 sg13g2_fill_1 FILLER_15_2379 ();
 sg13g2_fill_1 FILLER_15_2393 ();
 sg13g2_fill_2 FILLER_15_2424 ();
 sg13g2_fill_1 FILLER_15_2473 ();
 sg13g2_decap_8 FILLER_15_2500 ();
 sg13g2_decap_8 FILLER_15_2507 ();
 sg13g2_fill_1 FILLER_15_2514 ();
 sg13g2_decap_8 FILLER_15_2565 ();
 sg13g2_decap_8 FILLER_15_2572 ();
 sg13g2_decap_8 FILLER_15_2579 ();
 sg13g2_decap_8 FILLER_15_2586 ();
 sg13g2_decap_8 FILLER_15_2593 ();
 sg13g2_decap_8 FILLER_15_2600 ();
 sg13g2_decap_8 FILLER_15_2607 ();
 sg13g2_decap_8 FILLER_15_2614 ();
 sg13g2_decap_8 FILLER_15_2621 ();
 sg13g2_decap_8 FILLER_15_2628 ();
 sg13g2_decap_8 FILLER_15_2635 ();
 sg13g2_decap_8 FILLER_15_2642 ();
 sg13g2_decap_8 FILLER_15_2649 ();
 sg13g2_decap_8 FILLER_15_2656 ();
 sg13g2_decap_8 FILLER_15_2663 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_15 ();
 sg13g2_fill_1 FILLER_16_31 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_2 FILLER_16_72 ();
 sg13g2_decap_4 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_186 ();
 sg13g2_fill_2 FILLER_16_190 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_4 FILLER_16_378 ();
 sg13g2_fill_1 FILLER_16_415 ();
 sg13g2_fill_2 FILLER_16_447 ();
 sg13g2_decap_8 FILLER_16_463 ();
 sg13g2_fill_1 FILLER_16_470 ();
 sg13g2_fill_2 FILLER_16_481 ();
 sg13g2_fill_1 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_505 ();
 sg13g2_fill_2 FILLER_16_512 ();
 sg13g2_fill_2 FILLER_16_549 ();
 sg13g2_fill_1 FILLER_16_551 ();
 sg13g2_fill_1 FILLER_16_615 ();
 sg13g2_fill_1 FILLER_16_626 ();
 sg13g2_fill_1 FILLER_16_645 ();
 sg13g2_fill_2 FILLER_16_701 ();
 sg13g2_decap_4 FILLER_16_718 ();
 sg13g2_fill_1 FILLER_16_748 ();
 sg13g2_decap_4 FILLER_16_796 ();
 sg13g2_decap_4 FILLER_16_834 ();
 sg13g2_fill_1 FILLER_16_890 ();
 sg13g2_fill_1 FILLER_16_895 ();
 sg13g2_fill_1 FILLER_16_906 ();
 sg13g2_fill_2 FILLER_16_937 ();
 sg13g2_fill_1 FILLER_16_939 ();
 sg13g2_fill_1 FILLER_16_999 ();
 sg13g2_decap_4 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1030 ();
 sg13g2_fill_2 FILLER_16_1047 ();
 sg13g2_fill_1 FILLER_16_1049 ();
 sg13g2_fill_1 FILLER_16_1084 ();
 sg13g2_decap_8 FILLER_16_1118 ();
 sg13g2_decap_4 FILLER_16_1129 ();
 sg13g2_decap_8 FILLER_16_1142 ();
 sg13g2_decap_8 FILLER_16_1149 ();
 sg13g2_decap_8 FILLER_16_1156 ();
 sg13g2_fill_2 FILLER_16_1163 ();
 sg13g2_fill_1 FILLER_16_1202 ();
 sg13g2_fill_2 FILLER_16_1218 ();
 sg13g2_fill_2 FILLER_16_1230 ();
 sg13g2_fill_1 FILLER_16_1232 ();
 sg13g2_decap_4 FILLER_16_1268 ();
 sg13g2_fill_2 FILLER_16_1272 ();
 sg13g2_decap_8 FILLER_16_1302 ();
 sg13g2_decap_4 FILLER_16_1309 ();
 sg13g2_fill_1 FILLER_16_1313 ();
 sg13g2_decap_4 FILLER_16_1319 ();
 sg13g2_fill_1 FILLER_16_1323 ();
 sg13g2_decap_4 FILLER_16_1337 ();
 sg13g2_fill_2 FILLER_16_1341 ();
 sg13g2_decap_8 FILLER_16_1354 ();
 sg13g2_decap_4 FILLER_16_1361 ();
 sg13g2_fill_2 FILLER_16_1365 ();
 sg13g2_decap_8 FILLER_16_1386 ();
 sg13g2_fill_2 FILLER_16_1393 ();
 sg13g2_fill_1 FILLER_16_1395 ();
 sg13g2_decap_8 FILLER_16_1435 ();
 sg13g2_fill_1 FILLER_16_1442 ();
 sg13g2_fill_2 FILLER_16_1479 ();
 sg13g2_fill_1 FILLER_16_1481 ();
 sg13g2_fill_2 FILLER_16_1525 ();
 sg13g2_fill_1 FILLER_16_1541 ();
 sg13g2_fill_2 FILLER_16_1553 ();
 sg13g2_fill_2 FILLER_16_1563 ();
 sg13g2_fill_1 FILLER_16_1578 ();
 sg13g2_fill_2 FILLER_16_1583 ();
 sg13g2_fill_2 FILLER_16_1614 ();
 sg13g2_fill_2 FILLER_16_1658 ();
 sg13g2_fill_1 FILLER_16_1660 ();
 sg13g2_fill_1 FILLER_16_1665 ();
 sg13g2_fill_1 FILLER_16_1681 ();
 sg13g2_fill_2 FILLER_16_1690 ();
 sg13g2_fill_1 FILLER_16_1748 ();
 sg13g2_fill_2 FILLER_16_1753 ();
 sg13g2_fill_1 FILLER_16_1763 ();
 sg13g2_fill_1 FILLER_16_1768 ();
 sg13g2_fill_1 FILLER_16_1779 ();
 sg13g2_fill_2 FILLER_16_1837 ();
 sg13g2_fill_2 FILLER_16_1849 ();
 sg13g2_fill_1 FILLER_16_1851 ();
 sg13g2_fill_1 FILLER_16_1878 ();
 sg13g2_fill_2 FILLER_16_1949 ();
 sg13g2_fill_1 FILLER_16_1951 ();
 sg13g2_fill_1 FILLER_16_1956 ();
 sg13g2_fill_2 FILLER_16_1999 ();
 sg13g2_fill_2 FILLER_16_2068 ();
 sg13g2_fill_2 FILLER_16_2098 ();
 sg13g2_fill_1 FILLER_16_2134 ();
 sg13g2_decap_4 FILLER_16_2149 ();
 sg13g2_fill_1 FILLER_16_2153 ();
 sg13g2_fill_1 FILLER_16_2158 ();
 sg13g2_decap_4 FILLER_16_2174 ();
 sg13g2_fill_2 FILLER_16_2178 ();
 sg13g2_decap_8 FILLER_16_2184 ();
 sg13g2_decap_8 FILLER_16_2191 ();
 sg13g2_decap_4 FILLER_16_2198 ();
 sg13g2_fill_1 FILLER_16_2202 ();
 sg13g2_fill_2 FILLER_16_2207 ();
 sg13g2_fill_2 FILLER_16_2318 ();
 sg13g2_fill_1 FILLER_16_2320 ();
 sg13g2_decap_8 FILLER_16_2325 ();
 sg13g2_decap_4 FILLER_16_2332 ();
 sg13g2_fill_1 FILLER_16_2336 ();
 sg13g2_decap_8 FILLER_16_2341 ();
 sg13g2_fill_1 FILLER_16_2348 ();
 sg13g2_fill_2 FILLER_16_2353 ();
 sg13g2_decap_8 FILLER_16_2365 ();
 sg13g2_fill_1 FILLER_16_2372 ();
 sg13g2_fill_1 FILLER_16_2399 ();
 sg13g2_fill_1 FILLER_16_2463 ();
 sg13g2_decap_8 FILLER_16_2510 ();
 sg13g2_fill_1 FILLER_16_2517 ();
 sg13g2_decap_8 FILLER_16_2543 ();
 sg13g2_fill_1 FILLER_16_2550 ();
 sg13g2_decap_8 FILLER_16_2581 ();
 sg13g2_decap_8 FILLER_16_2588 ();
 sg13g2_decap_8 FILLER_16_2595 ();
 sg13g2_decap_8 FILLER_16_2602 ();
 sg13g2_decap_8 FILLER_16_2609 ();
 sg13g2_decap_8 FILLER_16_2616 ();
 sg13g2_decap_8 FILLER_16_2623 ();
 sg13g2_decap_8 FILLER_16_2630 ();
 sg13g2_decap_8 FILLER_16_2637 ();
 sg13g2_decap_8 FILLER_16_2644 ();
 sg13g2_decap_8 FILLER_16_2651 ();
 sg13g2_decap_8 FILLER_16_2658 ();
 sg13g2_decap_4 FILLER_16_2665 ();
 sg13g2_fill_1 FILLER_16_2669 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_57 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_2 FILLER_17_250 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_decap_4 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_fill_1 FILLER_17_409 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_fill_1 FILLER_17_441 ();
 sg13g2_fill_2 FILLER_17_524 ();
 sg13g2_fill_1 FILLER_17_526 ();
 sg13g2_decap_8 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_600 ();
 sg13g2_fill_1 FILLER_17_634 ();
 sg13g2_fill_2 FILLER_17_685 ();
 sg13g2_fill_1 FILLER_17_687 ();
 sg13g2_fill_2 FILLER_17_714 ();
 sg13g2_fill_1 FILLER_17_716 ();
 sg13g2_fill_1 FILLER_17_726 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_fill_1 FILLER_17_789 ();
 sg13g2_fill_1 FILLER_17_803 ();
 sg13g2_fill_2 FILLER_17_863 ();
 sg13g2_fill_2 FILLER_17_936 ();
 sg13g2_fill_1 FILLER_17_938 ();
 sg13g2_fill_1 FILLER_17_965 ();
 sg13g2_fill_1 FILLER_17_969 ();
 sg13g2_fill_1 FILLER_17_982 ();
 sg13g2_decap_4 FILLER_17_987 ();
 sg13g2_fill_2 FILLER_17_991 ();
 sg13g2_fill_2 FILLER_17_1007 ();
 sg13g2_decap_4 FILLER_17_1013 ();
 sg13g2_fill_2 FILLER_17_1017 ();
 sg13g2_fill_2 FILLER_17_1028 ();
 sg13g2_fill_2 FILLER_17_1042 ();
 sg13g2_fill_1 FILLER_17_1044 ();
 sg13g2_fill_2 FILLER_17_1055 ();
 sg13g2_fill_1 FILLER_17_1057 ();
 sg13g2_fill_2 FILLER_17_1063 ();
 sg13g2_fill_2 FILLER_17_1085 ();
 sg13g2_decap_4 FILLER_17_1121 ();
 sg13g2_fill_1 FILLER_17_1125 ();
 sg13g2_decap_8 FILLER_17_1140 ();
 sg13g2_decap_8 FILLER_17_1147 ();
 sg13g2_decap_8 FILLER_17_1154 ();
 sg13g2_fill_2 FILLER_17_1161 ();
 sg13g2_fill_1 FILLER_17_1193 ();
 sg13g2_fill_1 FILLER_17_1204 ();
 sg13g2_fill_1 FILLER_17_1211 ();
 sg13g2_fill_2 FILLER_17_1218 ();
 sg13g2_fill_1 FILLER_17_1220 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_fill_1 FILLER_17_1266 ();
 sg13g2_decap_4 FILLER_17_1273 ();
 sg13g2_fill_2 FILLER_17_1294 ();
 sg13g2_decap_4 FILLER_17_1305 ();
 sg13g2_fill_1 FILLER_17_1309 ();
 sg13g2_fill_2 FILLER_17_1315 ();
 sg13g2_fill_1 FILLER_17_1321 ();
 sg13g2_decap_4 FILLER_17_1332 ();
 sg13g2_decap_8 FILLER_17_1350 ();
 sg13g2_decap_8 FILLER_17_1357 ();
 sg13g2_fill_2 FILLER_17_1364 ();
 sg13g2_fill_1 FILLER_17_1366 ();
 sg13g2_decap_4 FILLER_17_1371 ();
 sg13g2_fill_2 FILLER_17_1375 ();
 sg13g2_fill_1 FILLER_17_1382 ();
 sg13g2_decap_8 FILLER_17_1387 ();
 sg13g2_fill_2 FILLER_17_1394 ();
 sg13g2_fill_2 FILLER_17_1428 ();
 sg13g2_fill_1 FILLER_17_1471 ();
 sg13g2_fill_1 FILLER_17_1517 ();
 sg13g2_fill_1 FILLER_17_1529 ();
 sg13g2_fill_1 FILLER_17_1540 ();
 sg13g2_fill_1 FILLER_17_1553 ();
 sg13g2_fill_1 FILLER_17_1561 ();
 sg13g2_fill_1 FILLER_17_1572 ();
 sg13g2_fill_2 FILLER_17_1609 ();
 sg13g2_decap_8 FILLER_17_1650 ();
 sg13g2_decap_8 FILLER_17_1657 ();
 sg13g2_fill_1 FILLER_17_1699 ();
 sg13g2_fill_1 FILLER_17_1706 ();
 sg13g2_fill_2 FILLER_17_1711 ();
 sg13g2_fill_2 FILLER_17_1734 ();
 sg13g2_fill_1 FILLER_17_1736 ();
 sg13g2_fill_2 FILLER_17_1743 ();
 sg13g2_fill_1 FILLER_17_1745 ();
 sg13g2_fill_2 FILLER_17_1751 ();
 sg13g2_fill_2 FILLER_17_1758 ();
 sg13g2_fill_2 FILLER_17_1786 ();
 sg13g2_fill_1 FILLER_17_1788 ();
 sg13g2_fill_2 FILLER_17_1807 ();
 sg13g2_fill_1 FILLER_17_1809 ();
 sg13g2_fill_2 FILLER_17_1824 ();
 sg13g2_fill_1 FILLER_17_1826 ();
 sg13g2_fill_1 FILLER_17_1863 ();
 sg13g2_decap_8 FILLER_17_1868 ();
 sg13g2_decap_4 FILLER_17_1875 ();
 sg13g2_fill_1 FILLER_17_1904 ();
 sg13g2_fill_1 FILLER_17_1909 ();
 sg13g2_fill_1 FILLER_17_1922 ();
 sg13g2_fill_2 FILLER_17_1930 ();
 sg13g2_fill_2 FILLER_17_1940 ();
 sg13g2_fill_1 FILLER_17_1942 ();
 sg13g2_fill_1 FILLER_17_1947 ();
 sg13g2_fill_1 FILLER_17_1995 ();
 sg13g2_fill_2 FILLER_17_2105 ();
 sg13g2_decap_4 FILLER_17_2143 ();
 sg13g2_decap_8 FILLER_17_2209 ();
 sg13g2_decap_4 FILLER_17_2216 ();
 sg13g2_fill_1 FILLER_17_2246 ();
 sg13g2_fill_2 FILLER_17_2277 ();
 sg13g2_decap_8 FILLER_17_2294 ();
 sg13g2_decap_8 FILLER_17_2301 ();
 sg13g2_fill_2 FILLER_17_2308 ();
 sg13g2_fill_1 FILLER_17_2310 ();
 sg13g2_fill_2 FILLER_17_2314 ();
 sg13g2_fill_2 FILLER_17_2344 ();
 sg13g2_fill_1 FILLER_17_2396 ();
 sg13g2_decap_4 FILLER_17_2425 ();
 sg13g2_fill_1 FILLER_17_2429 ();
 sg13g2_fill_2 FILLER_17_2436 ();
 sg13g2_fill_1 FILLER_17_2438 ();
 sg13g2_decap_8 FILLER_17_2442 ();
 sg13g2_fill_2 FILLER_17_2449 ();
 sg13g2_fill_2 FILLER_17_2481 ();
 sg13g2_decap_4 FILLER_17_2487 ();
 sg13g2_decap_8 FILLER_17_2517 ();
 sg13g2_fill_1 FILLER_17_2524 ();
 sg13g2_fill_1 FILLER_17_2535 ();
 sg13g2_decap_8 FILLER_17_2576 ();
 sg13g2_decap_8 FILLER_17_2583 ();
 sg13g2_decap_8 FILLER_17_2590 ();
 sg13g2_decap_8 FILLER_17_2597 ();
 sg13g2_decap_8 FILLER_17_2604 ();
 sg13g2_decap_8 FILLER_17_2611 ();
 sg13g2_decap_8 FILLER_17_2618 ();
 sg13g2_decap_8 FILLER_17_2625 ();
 sg13g2_decap_8 FILLER_17_2632 ();
 sg13g2_decap_8 FILLER_17_2639 ();
 sg13g2_decap_8 FILLER_17_2646 ();
 sg13g2_decap_8 FILLER_17_2653 ();
 sg13g2_decap_8 FILLER_17_2660 ();
 sg13g2_fill_2 FILLER_17_2667 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_18 ();
 sg13g2_decap_4 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_33 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_59 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_fill_2 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_258 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_fill_2 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_538 ();
 sg13g2_fill_2 FILLER_18_545 ();
 sg13g2_fill_2 FILLER_18_608 ();
 sg13g2_fill_2 FILLER_18_628 ();
 sg13g2_fill_1 FILLER_18_630 ();
 sg13g2_decap_4 FILLER_18_664 ();
 sg13g2_fill_1 FILLER_18_668 ();
 sg13g2_decap_4 FILLER_18_705 ();
 sg13g2_fill_1 FILLER_18_709 ();
 sg13g2_fill_2 FILLER_18_736 ();
 sg13g2_fill_1 FILLER_18_738 ();
 sg13g2_fill_2 FILLER_18_760 ();
 sg13g2_fill_1 FILLER_18_762 ();
 sg13g2_fill_2 FILLER_18_786 ();
 sg13g2_decap_4 FILLER_18_844 ();
 sg13g2_fill_2 FILLER_18_848 ();
 sg13g2_fill_2 FILLER_18_871 ();
 sg13g2_fill_1 FILLER_18_873 ();
 sg13g2_fill_1 FILLER_18_878 ();
 sg13g2_fill_2 FILLER_18_889 ();
 sg13g2_fill_2 FILLER_18_900 ();
 sg13g2_fill_1 FILLER_18_928 ();
 sg13g2_fill_2 FILLER_18_944 ();
 sg13g2_fill_1 FILLER_18_960 ();
 sg13g2_fill_1 FILLER_18_965 ();
 sg13g2_decap_8 FILLER_18_969 ();
 sg13g2_decap_8 FILLER_18_976 ();
 sg13g2_decap_8 FILLER_18_983 ();
 sg13g2_fill_1 FILLER_18_990 ();
 sg13g2_fill_2 FILLER_18_1006 ();
 sg13g2_fill_1 FILLER_18_1018 ();
 sg13g2_fill_2 FILLER_18_1023 ();
 sg13g2_fill_2 FILLER_18_1051 ();
 sg13g2_fill_1 FILLER_18_1053 ();
 sg13g2_fill_1 FILLER_18_1058 ();
 sg13g2_fill_1 FILLER_18_1075 ();
 sg13g2_fill_1 FILLER_18_1098 ();
 sg13g2_fill_1 FILLER_18_1107 ();
 sg13g2_fill_2 FILLER_18_1113 ();
 sg13g2_fill_1 FILLER_18_1115 ();
 sg13g2_fill_2 FILLER_18_1120 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_decap_8 FILLER_18_1127 ();
 sg13g2_fill_2 FILLER_18_1134 ();
 sg13g2_fill_1 FILLER_18_1136 ();
 sg13g2_decap_4 FILLER_18_1172 ();
 sg13g2_decap_4 FILLER_18_1180 ();
 sg13g2_fill_2 FILLER_18_1184 ();
 sg13g2_fill_1 FILLER_18_1198 ();
 sg13g2_decap_4 FILLER_18_1221 ();
 sg13g2_decap_4 FILLER_18_1235 ();
 sg13g2_fill_1 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1248 ();
 sg13g2_fill_1 FILLER_18_1255 ();
 sg13g2_fill_2 FILLER_18_1265 ();
 sg13g2_fill_2 FILLER_18_1306 ();
 sg13g2_fill_1 FILLER_18_1326 ();
 sg13g2_fill_1 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1350 ();
 sg13g2_decap_4 FILLER_18_1357 ();
 sg13g2_fill_2 FILLER_18_1361 ();
 sg13g2_decap_8 FILLER_18_1370 ();
 sg13g2_decap_8 FILLER_18_1377 ();
 sg13g2_decap_4 FILLER_18_1384 ();
 sg13g2_fill_1 FILLER_18_1416 ();
 sg13g2_fill_2 FILLER_18_1421 ();
 sg13g2_fill_1 FILLER_18_1423 ();
 sg13g2_fill_1 FILLER_18_1429 ();
 sg13g2_fill_2 FILLER_18_1436 ();
 sg13g2_fill_2 FILLER_18_1476 ();
 sg13g2_fill_1 FILLER_18_1478 ();
 sg13g2_fill_2 FILLER_18_1527 ();
 sg13g2_decap_4 FILLER_18_1537 ();
 sg13g2_fill_2 FILLER_18_1584 ();
 sg13g2_fill_2 FILLER_18_1598 ();
 sg13g2_fill_1 FILLER_18_1605 ();
 sg13g2_fill_2 FILLER_18_1627 ();
 sg13g2_fill_2 FILLER_18_1637 ();
 sg13g2_fill_1 FILLER_18_1652 ();
 sg13g2_fill_2 FILLER_18_1662 ();
 sg13g2_fill_1 FILLER_18_1664 ();
 sg13g2_fill_1 FILLER_18_1725 ();
 sg13g2_decap_8 FILLER_18_1730 ();
 sg13g2_fill_2 FILLER_18_1737 ();
 sg13g2_decap_4 FILLER_18_1743 ();
 sg13g2_fill_1 FILLER_18_1751 ();
 sg13g2_fill_2 FILLER_18_1761 ();
 sg13g2_fill_1 FILLER_18_1768 ();
 sg13g2_fill_2 FILLER_18_1824 ();
 sg13g2_fill_1 FILLER_18_1826 ();
 sg13g2_decap_4 FILLER_18_1848 ();
 sg13g2_decap_8 FILLER_18_1856 ();
 sg13g2_decap_8 FILLER_18_1863 ();
 sg13g2_fill_1 FILLER_18_1870 ();
 sg13g2_decap_8 FILLER_18_1902 ();
 sg13g2_decap_8 FILLER_18_1909 ();
 sg13g2_decap_4 FILLER_18_1916 ();
 sg13g2_fill_1 FILLER_18_1920 ();
 sg13g2_fill_2 FILLER_18_1965 ();
 sg13g2_fill_1 FILLER_18_2035 ();
 sg13g2_fill_1 FILLER_18_2066 ();
 sg13g2_fill_1 FILLER_18_2088 ();
 sg13g2_fill_2 FILLER_18_2093 ();
 sg13g2_fill_1 FILLER_18_2128 ();
 sg13g2_fill_2 FILLER_18_2196 ();
 sg13g2_fill_1 FILLER_18_2198 ();
 sg13g2_decap_8 FILLER_18_2203 ();
 sg13g2_decap_8 FILLER_18_2210 ();
 sg13g2_decap_8 FILLER_18_2217 ();
 sg13g2_fill_2 FILLER_18_2224 ();
 sg13g2_fill_1 FILLER_18_2226 ();
 sg13g2_decap_8 FILLER_18_2262 ();
 sg13g2_decap_4 FILLER_18_2269 ();
 sg13g2_fill_1 FILLER_18_2273 ();
 sg13g2_fill_2 FILLER_18_2279 ();
 sg13g2_decap_8 FILLER_18_2294 ();
 sg13g2_fill_2 FILLER_18_2338 ();
 sg13g2_fill_1 FILLER_18_2340 ();
 sg13g2_decap_4 FILLER_18_2367 ();
 sg13g2_fill_2 FILLER_18_2457 ();
 sg13g2_fill_1 FILLER_18_2459 ();
 sg13g2_fill_2 FILLER_18_2507 ();
 sg13g2_fill_2 FILLER_18_2526 ();
 sg13g2_fill_1 FILLER_18_2528 ();
 sg13g2_decap_8 FILLER_18_2569 ();
 sg13g2_decap_8 FILLER_18_2576 ();
 sg13g2_decap_8 FILLER_18_2583 ();
 sg13g2_decap_8 FILLER_18_2590 ();
 sg13g2_decap_8 FILLER_18_2597 ();
 sg13g2_decap_8 FILLER_18_2604 ();
 sg13g2_decap_8 FILLER_18_2611 ();
 sg13g2_decap_8 FILLER_18_2618 ();
 sg13g2_decap_8 FILLER_18_2625 ();
 sg13g2_decap_8 FILLER_18_2632 ();
 sg13g2_decap_8 FILLER_18_2639 ();
 sg13g2_decap_8 FILLER_18_2646 ();
 sg13g2_decap_8 FILLER_18_2653 ();
 sg13g2_decap_8 FILLER_18_2660 ();
 sg13g2_fill_2 FILLER_18_2667 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_13 ();
 sg13g2_fill_1 FILLER_19_20 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_106 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_222 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_360 ();
 sg13g2_fill_2 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_fill_2 FILLER_19_473 ();
 sg13g2_decap_8 FILLER_19_479 ();
 sg13g2_decap_4 FILLER_19_486 ();
 sg13g2_decap_4 FILLER_19_494 ();
 sg13g2_decap_4 FILLER_19_511 ();
 sg13g2_fill_2 FILLER_19_550 ();
 sg13g2_fill_1 FILLER_19_552 ();
 sg13g2_decap_8 FILLER_19_614 ();
 sg13g2_fill_1 FILLER_19_621 ();
 sg13g2_fill_1 FILLER_19_650 ();
 sg13g2_fill_2 FILLER_19_662 ();
 sg13g2_fill_2 FILLER_19_671 ();
 sg13g2_fill_1 FILLER_19_673 ();
 sg13g2_decap_8 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_fill_2 FILLER_19_713 ();
 sg13g2_fill_2 FILLER_19_770 ();
 sg13g2_fill_1 FILLER_19_772 ();
 sg13g2_fill_2 FILLER_19_812 ();
 sg13g2_decap_4 FILLER_19_840 ();
 sg13g2_fill_1 FILLER_19_849 ();
 sg13g2_fill_1 FILLER_19_860 ();
 sg13g2_fill_1 FILLER_19_890 ();
 sg13g2_decap_8 FILLER_19_900 ();
 sg13g2_fill_2 FILLER_19_907 ();
 sg13g2_fill_1 FILLER_19_909 ();
 sg13g2_fill_1 FILLER_19_914 ();
 sg13g2_decap_8 FILLER_19_919 ();
 sg13g2_fill_1 FILLER_19_926 ();
 sg13g2_fill_2 FILLER_19_939 ();
 sg13g2_decap_8 FILLER_19_981 ();
 sg13g2_decap_4 FILLER_19_988 ();
 sg13g2_fill_1 FILLER_19_992 ();
 sg13g2_decap_8 FILLER_19_997 ();
 sg13g2_fill_2 FILLER_19_1004 ();
 sg13g2_fill_1 FILLER_19_1014 ();
 sg13g2_fill_1 FILLER_19_1020 ();
 sg13g2_decap_4 FILLER_19_1046 ();
 sg13g2_fill_2 FILLER_19_1050 ();
 sg13g2_fill_1 FILLER_19_1056 ();
 sg13g2_fill_1 FILLER_19_1061 ();
 sg13g2_fill_2 FILLER_19_1067 ();
 sg13g2_decap_4 FILLER_19_1187 ();
 sg13g2_fill_1 FILLER_19_1191 ();
 sg13g2_fill_2 FILLER_19_1213 ();
 sg13g2_fill_1 FILLER_19_1215 ();
 sg13g2_decap_4 FILLER_19_1239 ();
 sg13g2_decap_8 FILLER_19_1248 ();
 sg13g2_decap_4 FILLER_19_1259 ();
 sg13g2_fill_2 FILLER_19_1271 ();
 sg13g2_fill_1 FILLER_19_1273 ();
 sg13g2_fill_1 FILLER_19_1285 ();
 sg13g2_fill_2 FILLER_19_1296 ();
 sg13g2_fill_1 FILLER_19_1309 ();
 sg13g2_fill_2 FILLER_19_1337 ();
 sg13g2_fill_1 FILLER_19_1343 ();
 sg13g2_fill_2 FILLER_19_1355 ();
 sg13g2_fill_2 FILLER_19_1370 ();
 sg13g2_fill_1 FILLER_19_1377 ();
 sg13g2_fill_2 FILLER_19_1383 ();
 sg13g2_fill_2 FILLER_19_1394 ();
 sg13g2_fill_1 FILLER_19_1396 ();
 sg13g2_decap_4 FILLER_19_1459 ();
 sg13g2_fill_1 FILLER_19_1463 ();
 sg13g2_fill_2 FILLER_19_1468 ();
 sg13g2_fill_1 FILLER_19_1470 ();
 sg13g2_fill_1 FILLER_19_1475 ();
 sg13g2_fill_2 FILLER_19_1491 ();
 sg13g2_fill_2 FILLER_19_1497 ();
 sg13g2_fill_1 FILLER_19_1499 ();
 sg13g2_fill_1 FILLER_19_1545 ();
 sg13g2_fill_1 FILLER_19_1564 ();
 sg13g2_fill_2 FILLER_19_1581 ();
 sg13g2_fill_1 FILLER_19_1615 ();
 sg13g2_fill_1 FILLER_19_1620 ();
 sg13g2_fill_1 FILLER_19_1625 ();
 sg13g2_fill_1 FILLER_19_1638 ();
 sg13g2_fill_2 FILLER_19_1645 ();
 sg13g2_decap_4 FILLER_19_1658 ();
 sg13g2_decap_4 FILLER_19_1696 ();
 sg13g2_fill_2 FILLER_19_1700 ();
 sg13g2_decap_8 FILLER_19_1706 ();
 sg13g2_decap_8 FILLER_19_1713 ();
 sg13g2_decap_8 FILLER_19_1720 ();
 sg13g2_decap_4 FILLER_19_1727 ();
 sg13g2_fill_2 FILLER_19_1731 ();
 sg13g2_fill_1 FILLER_19_1765 ();
 sg13g2_fill_1 FILLER_19_1796 ();
 sg13g2_fill_1 FILLER_19_1844 ();
 sg13g2_decap_8 FILLER_19_1849 ();
 sg13g2_decap_8 FILLER_19_1856 ();
 sg13g2_fill_2 FILLER_19_1863 ();
 sg13g2_fill_1 FILLER_19_1865 ();
 sg13g2_decap_8 FILLER_19_1906 ();
 sg13g2_decap_8 FILLER_19_1913 ();
 sg13g2_decap_8 FILLER_19_1920 ();
 sg13g2_decap_4 FILLER_19_1927 ();
 sg13g2_fill_2 FILLER_19_1971 ();
 sg13g2_fill_2 FILLER_19_1983 ();
 sg13g2_fill_1 FILLER_19_2002 ();
 sg13g2_fill_2 FILLER_19_2080 ();
 sg13g2_fill_2 FILLER_19_2092 ();
 sg13g2_fill_1 FILLER_19_2114 ();
 sg13g2_decap_4 FILLER_19_2146 ();
 sg13g2_fill_1 FILLER_19_2215 ();
 sg13g2_decap_4 FILLER_19_2242 ();
 sg13g2_fill_2 FILLER_19_2246 ();
 sg13g2_fill_1 FILLER_19_2357 ();
 sg13g2_decap_4 FILLER_19_2362 ();
 sg13g2_fill_2 FILLER_19_2366 ();
 sg13g2_fill_1 FILLER_19_2421 ();
 sg13g2_decap_4 FILLER_19_2432 ();
 sg13g2_fill_1 FILLER_19_2463 ();
 sg13g2_fill_2 FILLER_19_2469 ();
 sg13g2_decap_8 FILLER_19_2475 ();
 sg13g2_decap_4 FILLER_19_2482 ();
 sg13g2_fill_1 FILLER_19_2486 ();
 sg13g2_fill_2 FILLER_19_2497 ();
 sg13g2_decap_8 FILLER_19_2530 ();
 sg13g2_decap_8 FILLER_19_2537 ();
 sg13g2_fill_1 FILLER_19_2544 ();
 sg13g2_decap_8 FILLER_19_2581 ();
 sg13g2_decap_8 FILLER_19_2588 ();
 sg13g2_decap_8 FILLER_19_2595 ();
 sg13g2_decap_8 FILLER_19_2602 ();
 sg13g2_decap_8 FILLER_19_2609 ();
 sg13g2_decap_8 FILLER_19_2616 ();
 sg13g2_decap_8 FILLER_19_2623 ();
 sg13g2_decap_8 FILLER_19_2630 ();
 sg13g2_decap_8 FILLER_19_2637 ();
 sg13g2_decap_8 FILLER_19_2644 ();
 sg13g2_decap_8 FILLER_19_2651 ();
 sg13g2_decap_8 FILLER_19_2658 ();
 sg13g2_decap_4 FILLER_19_2665 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_88 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_fill_1 FILLER_20_444 ();
 sg13g2_fill_2 FILLER_20_457 ();
 sg13g2_fill_1 FILLER_20_471 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_516 ();
 sg13g2_fill_1 FILLER_20_523 ();
 sg13g2_fill_1 FILLER_20_547 ();
 sg13g2_fill_2 FILLER_20_592 ();
 sg13g2_fill_2 FILLER_20_678 ();
 sg13g2_decap_4 FILLER_20_701 ();
 sg13g2_fill_1 FILLER_20_705 ();
 sg13g2_fill_2 FILLER_20_715 ();
 sg13g2_fill_1 FILLER_20_717 ();
 sg13g2_fill_2 FILLER_20_739 ();
 sg13g2_decap_4 FILLER_20_801 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_decap_4 FILLER_20_836 ();
 sg13g2_decap_4 FILLER_20_850 ();
 sg13g2_fill_1 FILLER_20_894 ();
 sg13g2_fill_1 FILLER_20_908 ();
 sg13g2_decap_8 FILLER_20_913 ();
 sg13g2_fill_2 FILLER_20_920 ();
 sg13g2_fill_2 FILLER_20_1023 ();
 sg13g2_fill_1 FILLER_20_1055 ();
 sg13g2_fill_1 FILLER_20_1061 ();
 sg13g2_fill_1 FILLER_20_1093 ();
 sg13g2_fill_1 FILLER_20_1155 ();
 sg13g2_fill_2 FILLER_20_1160 ();
 sg13g2_fill_1 FILLER_20_1162 ();
 sg13g2_fill_1 FILLER_20_1199 ();
 sg13g2_fill_1 FILLER_20_1205 ();
 sg13g2_fill_1 FILLER_20_1222 ();
 sg13g2_decap_4 FILLER_20_1230 ();
 sg13g2_fill_1 FILLER_20_1234 ();
 sg13g2_decap_8 FILLER_20_1262 ();
 sg13g2_decap_8 FILLER_20_1269 ();
 sg13g2_fill_2 FILLER_20_1276 ();
 sg13g2_fill_2 FILLER_20_1283 ();
 sg13g2_fill_1 FILLER_20_1285 ();
 sg13g2_decap_4 FILLER_20_1297 ();
 sg13g2_fill_1 FILLER_20_1301 ();
 sg13g2_fill_1 FILLER_20_1312 ();
 sg13g2_fill_1 FILLER_20_1319 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_fill_1 FILLER_20_1332 ();
 sg13g2_fill_1 FILLER_20_1338 ();
 sg13g2_fill_1 FILLER_20_1351 ();
 sg13g2_decap_4 FILLER_20_1357 ();
 sg13g2_fill_1 FILLER_20_1361 ();
 sg13g2_fill_2 FILLER_20_1369 ();
 sg13g2_fill_1 FILLER_20_1384 ();
 sg13g2_fill_1 FILLER_20_1389 ();
 sg13g2_fill_1 FILLER_20_1425 ();
 sg13g2_decap_8 FILLER_20_1439 ();
 sg13g2_fill_2 FILLER_20_1446 ();
 sg13g2_fill_1 FILLER_20_1448 ();
 sg13g2_decap_8 FILLER_20_1453 ();
 sg13g2_decap_8 FILLER_20_1460 ();
 sg13g2_fill_2 FILLER_20_1467 ();
 sg13g2_fill_2 FILLER_20_1479 ();
 sg13g2_decap_8 FILLER_20_1485 ();
 sg13g2_decap_8 FILLER_20_1492 ();
 sg13g2_decap_4 FILLER_20_1499 ();
 sg13g2_fill_2 FILLER_20_1503 ();
 sg13g2_fill_2 FILLER_20_1516 ();
 sg13g2_fill_2 FILLER_20_1563 ();
 sg13g2_fill_2 FILLER_20_1568 ();
 sg13g2_fill_1 FILLER_20_1585 ();
 sg13g2_fill_1 FILLER_20_1620 ();
 sg13g2_decap_8 FILLER_20_1655 ();
 sg13g2_fill_2 FILLER_20_1662 ();
 sg13g2_fill_1 FILLER_20_1664 ();
 sg13g2_fill_2 FILLER_20_1687 ();
 sg13g2_decap_4 FILLER_20_1715 ();
 sg13g2_fill_1 FILLER_20_1723 ();
 sg13g2_decap_8 FILLER_20_1734 ();
 sg13g2_fill_1 FILLER_20_1741 ();
 sg13g2_decap_4 FILLER_20_1751 ();
 sg13g2_decap_4 FILLER_20_1759 ();
 sg13g2_fill_1 FILLER_20_1763 ();
 sg13g2_decap_4 FILLER_20_1780 ();
 sg13g2_decap_8 FILLER_20_1792 ();
 sg13g2_fill_1 FILLER_20_1799 ();
 sg13g2_decap_8 FILLER_20_1844 ();
 sg13g2_decap_8 FILLER_20_1851 ();
 sg13g2_fill_2 FILLER_20_1858 ();
 sg13g2_fill_1 FILLER_20_1860 ();
 sg13g2_decap_8 FILLER_20_1949 ();
 sg13g2_fill_1 FILLER_20_1989 ();
 sg13g2_fill_1 FILLER_20_2002 ();
 sg13g2_fill_1 FILLER_20_2013 ();
 sg13g2_decap_8 FILLER_20_2142 ();
 sg13g2_decap_8 FILLER_20_2149 ();
 sg13g2_decap_4 FILLER_20_2156 ();
 sg13g2_fill_2 FILLER_20_2160 ();
 sg13g2_fill_2 FILLER_20_2183 ();
 sg13g2_decap_4 FILLER_20_2206 ();
 sg13g2_decap_8 FILLER_20_2260 ();
 sg13g2_decap_8 FILLER_20_2267 ();
 sg13g2_decap_4 FILLER_20_2274 ();
 sg13g2_fill_1 FILLER_20_2278 ();
 sg13g2_decap_4 FILLER_20_2283 ();
 sg13g2_fill_1 FILLER_20_2287 ();
 sg13g2_decap_4 FILLER_20_2347 ();
 sg13g2_fill_1 FILLER_20_2351 ();
 sg13g2_fill_1 FILLER_20_2367 ();
 sg13g2_fill_2 FILLER_20_2398 ();
 sg13g2_fill_2 FILLER_20_2430 ();
 sg13g2_fill_2 FILLER_20_2440 ();
 sg13g2_decap_8 FILLER_20_2446 ();
 sg13g2_decap_4 FILLER_20_2453 ();
 sg13g2_fill_1 FILLER_20_2457 ();
 sg13g2_decap_4 FILLER_20_2509 ();
 sg13g2_decap_8 FILLER_20_2517 ();
 sg13g2_decap_8 FILLER_20_2524 ();
 sg13g2_decap_4 FILLER_20_2531 ();
 sg13g2_fill_1 FILLER_20_2535 ();
 sg13g2_fill_2 FILLER_20_2546 ();
 sg13g2_fill_1 FILLER_20_2548 ();
 sg13g2_decap_4 FILLER_20_2559 ();
 sg13g2_fill_1 FILLER_20_2563 ();
 sg13g2_decap_8 FILLER_20_2568 ();
 sg13g2_decap_8 FILLER_20_2575 ();
 sg13g2_decap_8 FILLER_20_2582 ();
 sg13g2_decap_8 FILLER_20_2589 ();
 sg13g2_decap_8 FILLER_20_2596 ();
 sg13g2_decap_8 FILLER_20_2603 ();
 sg13g2_decap_8 FILLER_20_2610 ();
 sg13g2_decap_8 FILLER_20_2617 ();
 sg13g2_decap_8 FILLER_20_2624 ();
 sg13g2_decap_8 FILLER_20_2631 ();
 sg13g2_decap_8 FILLER_20_2638 ();
 sg13g2_decap_8 FILLER_20_2645 ();
 sg13g2_decap_8 FILLER_20_2652 ();
 sg13g2_decap_8 FILLER_20_2659 ();
 sg13g2_decap_4 FILLER_20_2666 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_52 ();
 sg13g2_decap_8 FILLER_21_57 ();
 sg13g2_fill_2 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_395 ();
 sg13g2_fill_1 FILLER_21_420 ();
 sg13g2_fill_1 FILLER_21_440 ();
 sg13g2_fill_1 FILLER_21_449 ();
 sg13g2_fill_2 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_464 ();
 sg13g2_decap_8 FILLER_21_492 ();
 sg13g2_decap_8 FILLER_21_506 ();
 sg13g2_fill_2 FILLER_21_513 ();
 sg13g2_fill_1 FILLER_21_515 ();
 sg13g2_fill_1 FILLER_21_559 ();
 sg13g2_fill_2 FILLER_21_582 ();
 sg13g2_fill_2 FILLER_21_594 ();
 sg13g2_fill_2 FILLER_21_631 ();
 sg13g2_fill_1 FILLER_21_633 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_decap_4 FILLER_21_682 ();
 sg13g2_fill_1 FILLER_21_764 ();
 sg13g2_fill_2 FILLER_21_775 ();
 sg13g2_fill_1 FILLER_21_777 ();
 sg13g2_fill_1 FILLER_21_804 ();
 sg13g2_fill_1 FILLER_21_810 ();
 sg13g2_fill_1 FILLER_21_841 ();
 sg13g2_fill_1 FILLER_21_894 ();
 sg13g2_fill_2 FILLER_21_931 ();
 sg13g2_fill_1 FILLER_21_943 ();
 sg13g2_fill_2 FILLER_21_970 ();
 sg13g2_fill_2 FILLER_21_1019 ();
 sg13g2_fill_1 FILLER_21_1021 ();
 sg13g2_fill_2 FILLER_21_1032 ();
 sg13g2_fill_1 FILLER_21_1034 ();
 sg13g2_fill_2 FILLER_21_1061 ();
 sg13g2_decap_8 FILLER_21_1115 ();
 sg13g2_fill_2 FILLER_21_1122 ();
 sg13g2_decap_4 FILLER_21_1132 ();
 sg13g2_fill_1 FILLER_21_1136 ();
 sg13g2_decap_4 FILLER_21_1142 ();
 sg13g2_decap_8 FILLER_21_1150 ();
 sg13g2_decap_8 FILLER_21_1157 ();
 sg13g2_decap_8 FILLER_21_1164 ();
 sg13g2_fill_1 FILLER_21_1171 ();
 sg13g2_decap_4 FILLER_21_1186 ();
 sg13g2_fill_2 FILLER_21_1190 ();
 sg13g2_fill_2 FILLER_21_1242 ();
 sg13g2_fill_1 FILLER_21_1244 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_decap_4 FILLER_21_1274 ();
 sg13g2_fill_2 FILLER_21_1288 ();
 sg13g2_fill_2 FILLER_21_1314 ();
 sg13g2_fill_1 FILLER_21_1316 ();
 sg13g2_fill_2 FILLER_21_1404 ();
 sg13g2_decap_4 FILLER_21_1411 ();
 sg13g2_decap_4 FILLER_21_1419 ();
 sg13g2_fill_1 FILLER_21_1423 ();
 sg13g2_decap_8 FILLER_21_1430 ();
 sg13g2_decap_4 FILLER_21_1437 ();
 sg13g2_decap_4 FILLER_21_1445 ();
 sg13g2_decap_4 FILLER_21_1505 ();
 sg13g2_fill_1 FILLER_21_1509 ();
 sg13g2_fill_2 FILLER_21_1560 ();
 sg13g2_fill_1 FILLER_21_1610 ();
 sg13g2_fill_2 FILLER_21_1616 ();
 sg13g2_decap_8 FILLER_21_1656 ();
 sg13g2_fill_2 FILLER_21_1663 ();
 sg13g2_fill_1 FILLER_21_1665 ();
 sg13g2_fill_2 FILLER_21_1704 ();
 sg13g2_fill_1 FILLER_21_1706 ();
 sg13g2_fill_1 FILLER_21_1718 ();
 sg13g2_decap_4 FILLER_21_1728 ();
 sg13g2_fill_2 FILLER_21_1732 ();
 sg13g2_fill_1 FILLER_21_1750 ();
 sg13g2_fill_1 FILLER_21_1759 ();
 sg13g2_fill_2 FILLER_21_1767 ();
 sg13g2_fill_1 FILLER_21_1769 ();
 sg13g2_fill_1 FILLER_21_1778 ();
 sg13g2_decap_8 FILLER_21_1794 ();
 sg13g2_decap_4 FILLER_21_1801 ();
 sg13g2_decap_4 FILLER_21_1809 ();
 sg13g2_fill_1 FILLER_21_1813 ();
 sg13g2_fill_1 FILLER_21_1850 ();
 sg13g2_fill_2 FILLER_21_1885 ();
 sg13g2_fill_2 FILLER_21_1908 ();
 sg13g2_fill_2 FILLER_21_1914 ();
 sg13g2_fill_1 FILLER_21_1926 ();
 sg13g2_fill_1 FILLER_21_1944 ();
 sg13g2_fill_1 FILLER_21_1954 ();
 sg13g2_fill_1 FILLER_21_1976 ();
 sg13g2_fill_2 FILLER_21_1998 ();
 sg13g2_fill_2 FILLER_21_2077 ();
 sg13g2_fill_1 FILLER_21_2128 ();
 sg13g2_decap_8 FILLER_21_2163 ();
 sg13g2_fill_2 FILLER_21_2196 ();
 sg13g2_fill_1 FILLER_21_2198 ();
 sg13g2_decap_4 FILLER_21_2214 ();
 sg13g2_fill_1 FILLER_21_2218 ();
 sg13g2_fill_1 FILLER_21_2223 ();
 sg13g2_decap_4 FILLER_21_2228 ();
 sg13g2_fill_1 FILLER_21_2292 ();
 sg13g2_decap_4 FILLER_21_2334 ();
 sg13g2_fill_1 FILLER_21_2338 ();
 sg13g2_fill_2 FILLER_21_2342 ();
 sg13g2_fill_1 FILLER_21_2344 ();
 sg13g2_fill_2 FILLER_21_2375 ();
 sg13g2_decap_4 FILLER_21_2421 ();
 sg13g2_fill_1 FILLER_21_2425 ();
 sg13g2_decap_8 FILLER_21_2550 ();
 sg13g2_decap_8 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2590 ();
 sg13g2_decap_8 FILLER_21_2597 ();
 sg13g2_decap_8 FILLER_21_2604 ();
 sg13g2_decap_8 FILLER_21_2611 ();
 sg13g2_decap_8 FILLER_21_2618 ();
 sg13g2_decap_8 FILLER_21_2625 ();
 sg13g2_decap_8 FILLER_21_2632 ();
 sg13g2_decap_8 FILLER_21_2639 ();
 sg13g2_decap_8 FILLER_21_2646 ();
 sg13g2_decap_8 FILLER_21_2653 ();
 sg13g2_decap_8 FILLER_21_2660 ();
 sg13g2_fill_2 FILLER_21_2667 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_4 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_467 ();
 sg13g2_fill_2 FILLER_22_471 ();
 sg13g2_decap_4 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_485 ();
 sg13g2_fill_1 FILLER_22_527 ();
 sg13g2_fill_1 FILLER_22_568 ();
 sg13g2_fill_2 FILLER_22_657 ();
 sg13g2_fill_2 FILLER_22_663 ();
 sg13g2_fill_1 FILLER_22_669 ();
 sg13g2_fill_2 FILLER_22_696 ();
 sg13g2_fill_1 FILLER_22_698 ();
 sg13g2_decap_4 FILLER_22_735 ();
 sg13g2_fill_2 FILLER_22_743 ();
 sg13g2_fill_1 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_806 ();
 sg13g2_decap_4 FILLER_22_818 ();
 sg13g2_decap_4 FILLER_22_890 ();
 sg13g2_fill_2 FILLER_22_933 ();
 sg13g2_fill_1 FILLER_22_935 ();
 sg13g2_fill_1 FILLER_22_966 ();
 sg13g2_decap_8 FILLER_22_1046 ();
 sg13g2_decap_8 FILLER_22_1053 ();
 sg13g2_fill_1 FILLER_22_1060 ();
 sg13g2_fill_2 FILLER_22_1070 ();
 sg13g2_decap_8 FILLER_22_1112 ();
 sg13g2_fill_2 FILLER_22_1119 ();
 sg13g2_decap_4 FILLER_22_1125 ();
 sg13g2_fill_2 FILLER_22_1129 ();
 sg13g2_decap_4 FILLER_22_1141 ();
 sg13g2_decap_4 FILLER_22_1149 ();
 sg13g2_fill_2 FILLER_22_1168 ();
 sg13g2_fill_2 FILLER_22_1187 ();
 sg13g2_fill_2 FILLER_22_1208 ();
 sg13g2_fill_1 FILLER_22_1210 ();
 sg13g2_fill_1 FILLER_22_1218 ();
 sg13g2_fill_1 FILLER_22_1224 ();
 sg13g2_fill_2 FILLER_22_1249 ();
 sg13g2_fill_1 FILLER_22_1256 ();
 sg13g2_fill_1 FILLER_22_1261 ();
 sg13g2_fill_2 FILLER_22_1271 ();
 sg13g2_decap_8 FILLER_22_1308 ();
 sg13g2_decap_8 FILLER_22_1315 ();
 sg13g2_decap_8 FILLER_22_1322 ();
 sg13g2_decap_4 FILLER_22_1329 ();
 sg13g2_fill_1 FILLER_22_1350 ();
 sg13g2_fill_1 FILLER_22_1385 ();
 sg13g2_decap_8 FILLER_22_1405 ();
 sg13g2_decap_4 FILLER_22_1412 ();
 sg13g2_fill_1 FILLER_22_1416 ();
 sg13g2_decap_4 FILLER_22_1421 ();
 sg13g2_fill_2 FILLER_22_1425 ();
 sg13g2_decap_8 FILLER_22_1451 ();
 sg13g2_decap_4 FILLER_22_1458 ();
 sg13g2_fill_1 FILLER_22_1462 ();
 sg13g2_decap_4 FILLER_22_1467 ();
 sg13g2_fill_2 FILLER_22_1471 ();
 sg13g2_fill_2 FILLER_22_1513 ();
 sg13g2_fill_1 FILLER_22_1521 ();
 sg13g2_fill_2 FILLER_22_1528 ();
 sg13g2_fill_2 FILLER_22_1534 ();
 sg13g2_fill_1 FILLER_22_1563 ();
 sg13g2_fill_1 FILLER_22_1568 ();
 sg13g2_fill_1 FILLER_22_1576 ();
 sg13g2_decap_4 FILLER_22_1595 ();
 sg13g2_fill_1 FILLER_22_1625 ();
 sg13g2_fill_1 FILLER_22_1635 ();
 sg13g2_fill_2 FILLER_22_1657 ();
 sg13g2_fill_1 FILLER_22_1659 ();
 sg13g2_decap_4 FILLER_22_1665 ();
 sg13g2_fill_1 FILLER_22_1669 ();
 sg13g2_fill_1 FILLER_22_1686 ();
 sg13g2_fill_1 FILLER_22_1692 ();
 sg13g2_fill_1 FILLER_22_1750 ();
 sg13g2_fill_2 FILLER_22_1774 ();
 sg13g2_fill_1 FILLER_22_1776 ();
 sg13g2_fill_2 FILLER_22_1808 ();
 sg13g2_fill_1 FILLER_22_1810 ();
 sg13g2_fill_2 FILLER_22_1825 ();
 sg13g2_fill_1 FILLER_22_1827 ();
 sg13g2_fill_1 FILLER_22_1832 ();
 sg13g2_decap_4 FILLER_22_1837 ();
 sg13g2_fill_1 FILLER_22_1866 ();
 sg13g2_fill_2 FILLER_22_1877 ();
 sg13g2_fill_1 FILLER_22_1929 ();
 sg13g2_fill_1 FILLER_22_1979 ();
 sg13g2_fill_1 FILLER_22_1984 ();
 sg13g2_fill_2 FILLER_22_2023 ();
 sg13g2_fill_2 FILLER_22_2068 ();
 sg13g2_fill_1 FILLER_22_2088 ();
 sg13g2_fill_1 FILLER_22_2102 ();
 sg13g2_decap_8 FILLER_22_2202 ();
 sg13g2_fill_1 FILLER_22_2209 ();
 sg13g2_fill_2 FILLER_22_2240 ();
 sg13g2_fill_1 FILLER_22_2242 ();
 sg13g2_fill_2 FILLER_22_2278 ();
 sg13g2_fill_1 FILLER_22_2280 ();
 sg13g2_decap_4 FILLER_22_2326 ();
 sg13g2_fill_2 FILLER_22_2330 ();
 sg13g2_fill_2 FILLER_22_2429 ();
 sg13g2_fill_1 FILLER_22_2431 ();
 sg13g2_fill_1 FILLER_22_2446 ();
 sg13g2_decap_4 FILLER_22_2507 ();
 sg13g2_fill_2 FILLER_22_2511 ();
 sg13g2_fill_1 FILLER_22_2517 ();
 sg13g2_fill_2 FILLER_22_2558 ();
 sg13g2_fill_1 FILLER_22_2560 ();
 sg13g2_decap_8 FILLER_22_2587 ();
 sg13g2_decap_8 FILLER_22_2594 ();
 sg13g2_decap_8 FILLER_22_2601 ();
 sg13g2_decap_8 FILLER_22_2608 ();
 sg13g2_decap_8 FILLER_22_2615 ();
 sg13g2_decap_8 FILLER_22_2622 ();
 sg13g2_decap_8 FILLER_22_2629 ();
 sg13g2_decap_8 FILLER_22_2636 ();
 sg13g2_decap_8 FILLER_22_2643 ();
 sg13g2_decap_8 FILLER_22_2650 ();
 sg13g2_decap_8 FILLER_22_2657 ();
 sg13g2_decap_4 FILLER_22_2664 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_12 ();
 sg13g2_decap_4 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_22 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_443 ();
 sg13g2_fill_1 FILLER_23_454 ();
 sg13g2_fill_1 FILLER_23_490 ();
 sg13g2_fill_2 FILLER_23_502 ();
 sg13g2_fill_2 FILLER_23_542 ();
 sg13g2_fill_2 FILLER_23_563 ();
 sg13g2_fill_1 FILLER_23_598 ();
 sg13g2_decap_4 FILLER_23_663 ();
 sg13g2_fill_2 FILLER_23_693 ();
 sg13g2_fill_2 FILLER_23_730 ();
 sg13g2_fill_1 FILLER_23_732 ();
 sg13g2_fill_2 FILLER_23_737 ();
 sg13g2_fill_2 FILLER_23_744 ();
 sg13g2_fill_2 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_797 ();
 sg13g2_decap_8 FILLER_23_804 ();
 sg13g2_decap_4 FILLER_23_811 ();
 sg13g2_fill_2 FILLER_23_815 ();
 sg13g2_fill_2 FILLER_23_873 ();
 sg13g2_decap_4 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_888 ();
 sg13g2_fill_1 FILLER_23_895 ();
 sg13g2_decap_8 FILLER_23_955 ();
 sg13g2_fill_2 FILLER_23_962 ();
 sg13g2_fill_1 FILLER_23_964 ();
 sg13g2_fill_1 FILLER_23_985 ();
 sg13g2_fill_2 FILLER_23_1038 ();
 sg13g2_fill_1 FILLER_23_1040 ();
 sg13g2_decap_4 FILLER_23_1045 ();
 sg13g2_fill_2 FILLER_23_1049 ();
 sg13g2_fill_2 FILLER_23_1054 ();
 sg13g2_fill_1 FILLER_23_1056 ();
 sg13g2_fill_1 FILLER_23_1061 ();
 sg13g2_fill_1 FILLER_23_1075 ();
 sg13g2_fill_2 FILLER_23_1080 ();
 sg13g2_fill_2 FILLER_23_1086 ();
 sg13g2_fill_2 FILLER_23_1094 ();
 sg13g2_decap_8 FILLER_23_1138 ();
 sg13g2_fill_2 FILLER_23_1149 ();
 sg13g2_fill_1 FILLER_23_1151 ();
 sg13g2_fill_1 FILLER_23_1178 ();
 sg13g2_decap_4 FILLER_23_1213 ();
 sg13g2_decap_4 FILLER_23_1239 ();
 sg13g2_fill_2 FILLER_23_1248 ();
 sg13g2_fill_2 FILLER_23_1257 ();
 sg13g2_fill_1 FILLER_23_1259 ();
 sg13g2_fill_1 FILLER_23_1275 ();
 sg13g2_decap_8 FILLER_23_1285 ();
 sg13g2_fill_2 FILLER_23_1297 ();
 sg13g2_decap_4 FILLER_23_1308 ();
 sg13g2_fill_1 FILLER_23_1312 ();
 sg13g2_fill_1 FILLER_23_1337 ();
 sg13g2_decap_4 FILLER_23_1342 ();
 sg13g2_fill_1 FILLER_23_1346 ();
 sg13g2_decap_4 FILLER_23_1355 ();
 sg13g2_fill_1 FILLER_23_1373 ();
 sg13g2_fill_2 FILLER_23_1383 ();
 sg13g2_fill_1 FILLER_23_1390 ();
 sg13g2_fill_1 FILLER_23_1396 ();
 sg13g2_fill_1 FILLER_23_1403 ();
 sg13g2_decap_4 FILLER_23_1409 ();
 sg13g2_fill_2 FILLER_23_1422 ();
 sg13g2_fill_1 FILLER_23_1424 ();
 sg13g2_decap_8 FILLER_23_1465 ();
 sg13g2_decap_8 FILLER_23_1472 ();
 sg13g2_decap_4 FILLER_23_1479 ();
 sg13g2_fill_1 FILLER_23_1483 ();
 sg13g2_fill_2 FILLER_23_1520 ();
 sg13g2_fill_2 FILLER_23_1534 ();
 sg13g2_fill_1 FILLER_23_1557 ();
 sg13g2_fill_2 FILLER_23_1586 ();
 sg13g2_fill_2 FILLER_23_1608 ();
 sg13g2_fill_1 FILLER_23_1619 ();
 sg13g2_fill_2 FILLER_23_1663 ();
 sg13g2_fill_1 FILLER_23_1669 ();
 sg13g2_fill_1 FILLER_23_1675 ();
 sg13g2_fill_1 FILLER_23_1680 ();
 sg13g2_fill_1 FILLER_23_1686 ();
 sg13g2_fill_1 FILLER_23_1692 ();
 sg13g2_decap_4 FILLER_23_1698 ();
 sg13g2_fill_2 FILLER_23_1702 ();
 sg13g2_fill_2 FILLER_23_1708 ();
 sg13g2_fill_2 FILLER_23_1714 ();
 sg13g2_fill_1 FILLER_23_1716 ();
 sg13g2_fill_2 FILLER_23_1735 ();
 sg13g2_fill_1 FILLER_23_1747 ();
 sg13g2_fill_2 FILLER_23_1753 ();
 sg13g2_fill_1 FILLER_23_1755 ();
 sg13g2_fill_2 FILLER_23_1760 ();
 sg13g2_fill_1 FILLER_23_1808 ();
 sg13g2_fill_2 FILLER_23_1858 ();
 sg13g2_fill_1 FILLER_23_1860 ();
 sg13g2_fill_2 FILLER_23_1887 ();
 sg13g2_decap_8 FILLER_23_1938 ();
 sg13g2_fill_2 FILLER_23_1945 ();
 sg13g2_fill_1 FILLER_23_1999 ();
 sg13g2_fill_2 FILLER_23_2052 ();
 sg13g2_fill_1 FILLER_23_2064 ();
 sg13g2_fill_1 FILLER_23_2091 ();
 sg13g2_fill_2 FILLER_23_2106 ();
 sg13g2_fill_1 FILLER_23_2132 ();
 sg13g2_fill_1 FILLER_23_2159 ();
 sg13g2_fill_2 FILLER_23_2164 ();
 sg13g2_fill_1 FILLER_23_2176 ();
 sg13g2_fill_2 FILLER_23_2203 ();
 sg13g2_fill_1 FILLER_23_2209 ();
 sg13g2_decap_4 FILLER_23_2223 ();
 sg13g2_fill_2 FILLER_23_2227 ();
 sg13g2_fill_2 FILLER_23_2281 ();
 sg13g2_fill_1 FILLER_23_2345 ();
 sg13g2_fill_1 FILLER_23_2349 ();
 sg13g2_fill_1 FILLER_23_2360 ();
 sg13g2_fill_1 FILLER_23_2387 ();
 sg13g2_fill_1 FILLER_23_2398 ();
 sg13g2_decap_8 FILLER_23_2515 ();
 sg13g2_decap_8 FILLER_23_2522 ();
 sg13g2_decap_8 FILLER_23_2529 ();
 sg13g2_decap_8 FILLER_23_2536 ();
 sg13g2_decap_8 FILLER_23_2543 ();
 sg13g2_decap_4 FILLER_23_2550 ();
 sg13g2_fill_1 FILLER_23_2554 ();
 sg13g2_fill_1 FILLER_23_2569 ();
 sg13g2_decap_8 FILLER_23_2574 ();
 sg13g2_decap_8 FILLER_23_2581 ();
 sg13g2_decap_8 FILLER_23_2588 ();
 sg13g2_decap_8 FILLER_23_2595 ();
 sg13g2_decap_8 FILLER_23_2602 ();
 sg13g2_decap_8 FILLER_23_2609 ();
 sg13g2_decap_8 FILLER_23_2616 ();
 sg13g2_decap_8 FILLER_23_2623 ();
 sg13g2_decap_8 FILLER_23_2630 ();
 sg13g2_decap_8 FILLER_23_2637 ();
 sg13g2_decap_8 FILLER_23_2644 ();
 sg13g2_decap_8 FILLER_23_2651 ();
 sg13g2_decap_8 FILLER_23_2658 ();
 sg13g2_decap_4 FILLER_23_2665 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_30 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_319 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_4 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_369 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_24_422 ();
 sg13g2_fill_2 FILLER_24_433 ();
 sg13g2_fill_1 FILLER_24_465 ();
 sg13g2_fill_1 FILLER_24_528 ();
 sg13g2_fill_2 FILLER_24_568 ();
 sg13g2_fill_1 FILLER_24_611 ();
 sg13g2_fill_2 FILLER_24_638 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_fill_2 FILLER_24_668 ();
 sg13g2_fill_2 FILLER_24_681 ();
 sg13g2_fill_1 FILLER_24_683 ();
 sg13g2_fill_2 FILLER_24_721 ();
 sg13g2_fill_1 FILLER_24_723 ();
 sg13g2_decap_4 FILLER_24_728 ();
 sg13g2_fill_2 FILLER_24_732 ();
 sg13g2_fill_2 FILLER_24_758 ();
 sg13g2_fill_2 FILLER_24_786 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_decap_4 FILLER_24_819 ();
 sg13g2_decap_4 FILLER_24_858 ();
 sg13g2_fill_2 FILLER_24_862 ();
 sg13g2_fill_1 FILLER_24_894 ();
 sg13g2_fill_1 FILLER_24_904 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_4 FILLER_24_961 ();
 sg13g2_fill_1 FILLER_24_965 ();
 sg13g2_fill_1 FILLER_24_975 ();
 sg13g2_fill_2 FILLER_24_985 ();
 sg13g2_fill_1 FILLER_24_987 ();
 sg13g2_fill_1 FILLER_24_1015 ();
 sg13g2_fill_2 FILLER_24_1024 ();
 sg13g2_fill_2 FILLER_24_1040 ();
 sg13g2_fill_1 FILLER_24_1054 ();
 sg13g2_decap_4 FILLER_24_1147 ();
 sg13g2_fill_2 FILLER_24_1151 ();
 sg13g2_fill_1 FILLER_24_1163 ();
 sg13g2_fill_1 FILLER_24_1169 ();
 sg13g2_fill_1 FILLER_24_1175 ();
 sg13g2_fill_2 FILLER_24_1186 ();
 sg13g2_fill_1 FILLER_24_1191 ();
 sg13g2_decap_8 FILLER_24_1199 ();
 sg13g2_decap_4 FILLER_24_1206 ();
 sg13g2_fill_2 FILLER_24_1210 ();
 sg13g2_fill_1 FILLER_24_1217 ();
 sg13g2_decap_4 FILLER_24_1272 ();
 sg13g2_fill_1 FILLER_24_1276 ();
 sg13g2_fill_1 FILLER_24_1282 ();
 sg13g2_decap_8 FILLER_24_1294 ();
 sg13g2_decap_8 FILLER_24_1301 ();
 sg13g2_decap_4 FILLER_24_1308 ();
 sg13g2_fill_2 FILLER_24_1312 ();
 sg13g2_decap_4 FILLER_24_1319 ();
 sg13g2_decap_4 FILLER_24_1327 ();
 sg13g2_fill_1 FILLER_24_1331 ();
 sg13g2_fill_2 FILLER_24_1336 ();
 sg13g2_fill_1 FILLER_24_1338 ();
 sg13g2_fill_2 FILLER_24_1344 ();
 sg13g2_fill_2 FILLER_24_1354 ();
 sg13g2_fill_2 FILLER_24_1360 ();
 sg13g2_fill_1 FILLER_24_1381 ();
 sg13g2_fill_1 FILLER_24_1406 ();
 sg13g2_decap_4 FILLER_24_1446 ();
 sg13g2_fill_2 FILLER_24_1450 ();
 sg13g2_fill_1 FILLER_24_1478 ();
 sg13g2_fill_1 FILLER_24_1503 ();
 sg13g2_fill_1 FILLER_24_1514 ();
 sg13g2_fill_1 FILLER_24_1523 ();
 sg13g2_decap_4 FILLER_24_1534 ();
 sg13g2_fill_2 FILLER_24_1545 ();
 sg13g2_fill_1 FILLER_24_1560 ();
 sg13g2_fill_1 FILLER_24_1571 ();
 sg13g2_fill_1 FILLER_24_1604 ();
 sg13g2_fill_2 FILLER_24_1619 ();
 sg13g2_fill_2 FILLER_24_1733 ();
 sg13g2_fill_2 FILLER_24_1751 ();
 sg13g2_fill_1 FILLER_24_1822 ();
 sg13g2_decap_8 FILLER_24_1853 ();
 sg13g2_fill_2 FILLER_24_1860 ();
 sg13g2_fill_1 FILLER_24_1892 ();
 sg13g2_fill_2 FILLER_24_1925 ();
 sg13g2_fill_2 FILLER_24_1996 ();
 sg13g2_fill_2 FILLER_24_2027 ();
 sg13g2_fill_1 FILLER_24_2045 ();
 sg13g2_fill_2 FILLER_24_2103 ();
 sg13g2_fill_1 FILLER_24_2143 ();
 sg13g2_decap_8 FILLER_24_2161 ();
 sg13g2_decap_8 FILLER_24_2199 ();
 sg13g2_fill_2 FILLER_24_2232 ();
 sg13g2_fill_1 FILLER_24_2234 ();
 sg13g2_fill_1 FILLER_24_2239 ();
 sg13g2_fill_2 FILLER_24_2248 ();
 sg13g2_fill_2 FILLER_24_2275 ();
 sg13g2_decap_4 FILLER_24_2303 ();
 sg13g2_decap_8 FILLER_24_2464 ();
 sg13g2_decap_4 FILLER_24_2471 ();
 sg13g2_decap_8 FILLER_24_2522 ();
 sg13g2_fill_1 FILLER_24_2529 ();
 sg13g2_fill_2 FILLER_24_2540 ();
 sg13g2_fill_2 FILLER_24_2556 ();
 sg13g2_fill_1 FILLER_24_2558 ();
 sg13g2_decap_8 FILLER_24_2595 ();
 sg13g2_decap_8 FILLER_24_2602 ();
 sg13g2_decap_8 FILLER_24_2609 ();
 sg13g2_decap_8 FILLER_24_2616 ();
 sg13g2_decap_8 FILLER_24_2623 ();
 sg13g2_decap_8 FILLER_24_2630 ();
 sg13g2_decap_8 FILLER_24_2637 ();
 sg13g2_decap_8 FILLER_24_2644 ();
 sg13g2_decap_8 FILLER_24_2651 ();
 sg13g2_decap_8 FILLER_24_2658 ();
 sg13g2_decap_4 FILLER_24_2665 ();
 sg13g2_fill_1 FILLER_24_2669 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_decap_4 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_decap_4 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_2 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_333 ();
 sg13g2_fill_2 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_fill_1 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_468 ();
 sg13g2_fill_1 FILLER_25_544 ();
 sg13g2_fill_2 FILLER_25_575 ();
 sg13g2_fill_1 FILLER_25_634 ();
 sg13g2_fill_1 FILLER_25_661 ();
 sg13g2_fill_1 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_decap_4 FILLER_25_698 ();
 sg13g2_fill_2 FILLER_25_702 ();
 sg13g2_fill_2 FILLER_25_739 ();
 sg13g2_fill_1 FILLER_25_741 ();
 sg13g2_fill_2 FILLER_25_746 ();
 sg13g2_fill_2 FILLER_25_760 ();
 sg13g2_fill_2 FILLER_25_766 ();
 sg13g2_fill_2 FILLER_25_780 ();
 sg13g2_decap_4 FILLER_25_826 ();
 sg13g2_fill_1 FILLER_25_834 ();
 sg13g2_fill_2 FILLER_25_849 ();
 sg13g2_fill_1 FILLER_25_886 ();
 sg13g2_fill_2 FILLER_25_923 ();
 sg13g2_fill_1 FILLER_25_925 ();
 sg13g2_fill_2 FILLER_25_944 ();
 sg13g2_decap_4 FILLER_25_950 ();
 sg13g2_fill_1 FILLER_25_954 ();
 sg13g2_fill_2 FILLER_25_990 ();
 sg13g2_fill_1 FILLER_25_1002 ();
 sg13g2_fill_2 FILLER_25_1014 ();
 sg13g2_fill_1 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1025 ();
 sg13g2_decap_4 FILLER_25_1035 ();
 sg13g2_fill_1 FILLER_25_1039 ();
 sg13g2_fill_2 FILLER_25_1123 ();
 sg13g2_decap_4 FILLER_25_1154 ();
 sg13g2_fill_2 FILLER_25_1184 ();
 sg13g2_fill_2 FILLER_25_1193 ();
 sg13g2_fill_2 FILLER_25_1200 ();
 sg13g2_fill_1 FILLER_25_1202 ();
 sg13g2_fill_2 FILLER_25_1240 ();
 sg13g2_fill_1 FILLER_25_1242 ();
 sg13g2_decap_4 FILLER_25_1254 ();
 sg13g2_fill_1 FILLER_25_1258 ();
 sg13g2_decap_8 FILLER_25_1264 ();
 sg13g2_decap_4 FILLER_25_1281 ();
 sg13g2_fill_2 FILLER_25_1285 ();
 sg13g2_fill_1 FILLER_25_1300 ();
 sg13g2_fill_1 FILLER_25_1352 ();
 sg13g2_fill_1 FILLER_25_1358 ();
 sg13g2_fill_1 FILLER_25_1366 ();
 sg13g2_fill_2 FILLER_25_1392 ();
 sg13g2_fill_2 FILLER_25_1402 ();
 sg13g2_fill_2 FILLER_25_1509 ();
 sg13g2_fill_2 FILLER_25_1542 ();
 sg13g2_fill_1 FILLER_25_1552 ();
 sg13g2_fill_1 FILLER_25_1562 ();
 sg13g2_fill_1 FILLER_25_1582 ();
 sg13g2_fill_1 FILLER_25_1614 ();
 sg13g2_fill_1 FILLER_25_1622 ();
 sg13g2_fill_2 FILLER_25_1642 ();
 sg13g2_fill_2 FILLER_25_1649 ();
 sg13g2_fill_1 FILLER_25_1651 ();
 sg13g2_fill_1 FILLER_25_1656 ();
 sg13g2_fill_2 FILLER_25_1687 ();
 sg13g2_fill_1 FILLER_25_1689 ();
 sg13g2_fill_2 FILLER_25_1699 ();
 sg13g2_decap_8 FILLER_25_1727 ();
 sg13g2_decap_8 FILLER_25_1734 ();
 sg13g2_decap_8 FILLER_25_1741 ();
 sg13g2_decap_4 FILLER_25_1765 ();
 sg13g2_fill_2 FILLER_25_1769 ();
 sg13g2_fill_2 FILLER_25_1821 ();
 sg13g2_fill_1 FILLER_25_1823 ();
 sg13g2_decap_4 FILLER_25_1874 ();
 sg13g2_decap_8 FILLER_25_1914 ();
 sg13g2_decap_8 FILLER_25_1921 ();
 sg13g2_decap_4 FILLER_25_1928 ();
 sg13g2_fill_2 FILLER_25_1951 ();
 sg13g2_fill_1 FILLER_25_1953 ();
 sg13g2_fill_1 FILLER_25_1979 ();
 sg13g2_fill_2 FILLER_25_2019 ();
 sg13g2_fill_2 FILLER_25_2034 ();
 sg13g2_decap_4 FILLER_25_2152 ();
 sg13g2_fill_2 FILLER_25_2211 ();
 sg13g2_fill_1 FILLER_25_2213 ();
 sg13g2_fill_2 FILLER_25_2269 ();
 sg13g2_fill_1 FILLER_25_2271 ();
 sg13g2_decap_4 FILLER_25_2280 ();
 sg13g2_fill_2 FILLER_25_2284 ();
 sg13g2_decap_8 FILLER_25_2289 ();
 sg13g2_decap_8 FILLER_25_2296 ();
 sg13g2_fill_1 FILLER_25_2303 ();
 sg13g2_fill_1 FILLER_25_2325 ();
 sg13g2_decap_4 FILLER_25_2334 ();
 sg13g2_fill_2 FILLER_25_2338 ();
 sg13g2_fill_1 FILLER_25_2416 ();
 sg13g2_fill_1 FILLER_25_2446 ();
 sg13g2_fill_1 FILLER_25_2454 ();
 sg13g2_fill_2 FILLER_25_2479 ();
 sg13g2_fill_1 FILLER_25_2493 ();
 sg13g2_fill_2 FILLER_25_2519 ();
 sg13g2_decap_8 FILLER_25_2599 ();
 sg13g2_decap_8 FILLER_25_2606 ();
 sg13g2_decap_8 FILLER_25_2613 ();
 sg13g2_decap_8 FILLER_25_2620 ();
 sg13g2_decap_8 FILLER_25_2627 ();
 sg13g2_decap_8 FILLER_25_2634 ();
 sg13g2_decap_8 FILLER_25_2641 ();
 sg13g2_decap_8 FILLER_25_2648 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_fill_1 FILLER_25_2669 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_fill_2 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_367 ();
 sg13g2_decap_4 FILLER_26_374 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_26_385 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_fill_1 FILLER_26_398 ();
 sg13g2_fill_2 FILLER_26_468 ();
 sg13g2_fill_1 FILLER_26_528 ();
 sg13g2_fill_1 FILLER_26_533 ();
 sg13g2_fill_1 FILLER_26_544 ();
 sg13g2_fill_1 FILLER_26_571 ();
 sg13g2_fill_2 FILLER_26_593 ();
 sg13g2_fill_2 FILLER_26_704 ();
 sg13g2_fill_2 FILLER_26_742 ();
 sg13g2_fill_1 FILLER_26_744 ();
 sg13g2_fill_2 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_fill_2 FILLER_26_858 ();
 sg13g2_fill_1 FILLER_26_860 ();
 sg13g2_decap_4 FILLER_26_886 ();
 sg13g2_fill_1 FILLER_26_890 ();
 sg13g2_fill_2 FILLER_26_923 ();
 sg13g2_decap_8 FILLER_26_960 ();
 sg13g2_fill_1 FILLER_26_993 ();
 sg13g2_fill_1 FILLER_26_1015 ();
 sg13g2_fill_1 FILLER_26_1050 ();
 sg13g2_fill_2 FILLER_26_1099 ();
 sg13g2_fill_2 FILLER_26_1130 ();
 sg13g2_decap_4 FILLER_26_1155 ();
 sg13g2_decap_8 FILLER_26_1167 ();
 sg13g2_fill_1 FILLER_26_1181 ();
 sg13g2_decap_4 FILLER_26_1189 ();
 sg13g2_fill_1 FILLER_26_1193 ();
 sg13g2_decap_8 FILLER_26_1224 ();
 sg13g2_decap_4 FILLER_26_1236 ();
 sg13g2_fill_1 FILLER_26_1240 ();
 sg13g2_decap_4 FILLER_26_1251 ();
 sg13g2_fill_1 FILLER_26_1255 ();
 sg13g2_fill_1 FILLER_26_1269 ();
 sg13g2_fill_2 FILLER_26_1282 ();
 sg13g2_decap_4 FILLER_26_1291 ();
 sg13g2_fill_2 FILLER_26_1305 ();
 sg13g2_fill_2 FILLER_26_1312 ();
 sg13g2_fill_1 FILLER_26_1324 ();
 sg13g2_fill_1 FILLER_26_1331 ();
 sg13g2_fill_2 FILLER_26_1345 ();
 sg13g2_fill_1 FILLER_26_1367 ();
 sg13g2_fill_1 FILLER_26_1382 ();
 sg13g2_fill_1 FILLER_26_1391 ();
 sg13g2_fill_2 FILLER_26_1438 ();
 sg13g2_fill_2 FILLER_26_1473 ();
 sg13g2_decap_4 FILLER_26_1563 ();
 sg13g2_fill_1 FILLER_26_1567 ();
 sg13g2_fill_2 FILLER_26_1611 ();
 sg13g2_fill_2 FILLER_26_1640 ();
 sg13g2_fill_1 FILLER_26_1651 ();
 sg13g2_fill_1 FILLER_26_1657 ();
 sg13g2_fill_2 FILLER_26_1663 ();
 sg13g2_decap_8 FILLER_26_1677 ();
 sg13g2_decap_8 FILLER_26_1684 ();
 sg13g2_fill_2 FILLER_26_1691 ();
 sg13g2_decap_8 FILLER_26_1723 ();
 sg13g2_fill_2 FILLER_26_1730 ();
 sg13g2_fill_1 FILLER_26_1732 ();
 sg13g2_decap_8 FILLER_26_1755 ();
 sg13g2_fill_2 FILLER_26_1762 ();
 sg13g2_decap_8 FILLER_26_1794 ();
 sg13g2_decap_8 FILLER_26_1805 ();
 sg13g2_decap_8 FILLER_26_1812 ();
 sg13g2_decap_8 FILLER_26_1819 ();
 sg13g2_decap_4 FILLER_26_1826 ();
 sg13g2_decap_8 FILLER_26_1834 ();
 sg13g2_fill_1 FILLER_26_1841 ();
 sg13g2_decap_8 FILLER_26_1846 ();
 sg13g2_decap_4 FILLER_26_1853 ();
 sg13g2_decap_8 FILLER_26_1861 ();
 sg13g2_decap_8 FILLER_26_1868 ();
 sg13g2_decap_8 FILLER_26_1875 ();
 sg13g2_decap_8 FILLER_26_1882 ();
 sg13g2_decap_4 FILLER_26_1923 ();
 sg13g2_fill_2 FILLER_26_1927 ();
 sg13g2_fill_1 FILLER_26_1969 ();
 sg13g2_fill_1 FILLER_26_1992 ();
 sg13g2_fill_2 FILLER_26_2027 ();
 sg13g2_fill_2 FILLER_26_2108 ();
 sg13g2_fill_1 FILLER_26_2166 ();
 sg13g2_decap_8 FILLER_26_2193 ();
 sg13g2_fill_2 FILLER_26_2200 ();
 sg13g2_decap_8 FILLER_26_2238 ();
 sg13g2_decap_4 FILLER_26_2245 ();
 sg13g2_fill_2 FILLER_26_2249 ();
 sg13g2_fill_1 FILLER_26_2263 ();
 sg13g2_decap_8 FILLER_26_2276 ();
 sg13g2_fill_2 FILLER_26_2283 ();
 sg13g2_fill_1 FILLER_26_2285 ();
 sg13g2_fill_1 FILLER_26_2290 ();
 sg13g2_fill_2 FILLER_26_2305 ();
 sg13g2_fill_2 FILLER_26_2332 ();
 sg13g2_fill_1 FILLER_26_2334 ();
 sg13g2_fill_2 FILLER_26_2343 ();
 sg13g2_fill_1 FILLER_26_2345 ();
 sg13g2_fill_1 FILLER_26_2354 ();
 sg13g2_fill_1 FILLER_26_2379 ();
 sg13g2_fill_2 FILLER_26_2422 ();
 sg13g2_fill_2 FILLER_26_2445 ();
 sg13g2_fill_1 FILLER_26_2457 ();
 sg13g2_fill_2 FILLER_26_2479 ();
 sg13g2_fill_2 FILLER_26_2502 ();
 sg13g2_fill_2 FILLER_26_2508 ();
 sg13g2_decap_4 FILLER_26_2536 ();
 sg13g2_fill_2 FILLER_26_2546 ();
 sg13g2_fill_2 FILLER_26_2569 ();
 sg13g2_fill_1 FILLER_26_2571 ();
 sg13g2_decap_8 FILLER_26_2598 ();
 sg13g2_decap_8 FILLER_26_2605 ();
 sg13g2_decap_8 FILLER_26_2612 ();
 sg13g2_decap_8 FILLER_26_2619 ();
 sg13g2_decap_8 FILLER_26_2626 ();
 sg13g2_decap_8 FILLER_26_2633 ();
 sg13g2_decap_8 FILLER_26_2640 ();
 sg13g2_decap_8 FILLER_26_2647 ();
 sg13g2_decap_8 FILLER_26_2654 ();
 sg13g2_decap_8 FILLER_26_2661 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_27_411 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_8 FILLER_27_426 ();
 sg13g2_fill_2 FILLER_27_433 ();
 sg13g2_fill_2 FILLER_27_447 ();
 sg13g2_fill_2 FILLER_27_463 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_fill_2 FILLER_27_479 ();
 sg13g2_fill_1 FILLER_27_532 ();
 sg13g2_fill_1 FILLER_27_552 ();
 sg13g2_fill_1 FILLER_27_557 ();
 sg13g2_fill_2 FILLER_27_584 ();
 sg13g2_fill_2 FILLER_27_702 ();
 sg13g2_fill_1 FILLER_27_704 ();
 sg13g2_fill_1 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_fill_1 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_fill_2 FILLER_27_830 ();
 sg13g2_fill_1 FILLER_27_832 ();
 sg13g2_fill_2 FILLER_27_843 ();
 sg13g2_fill_2 FILLER_27_849 ();
 sg13g2_fill_1 FILLER_27_851 ();
 sg13g2_decap_4 FILLER_27_886 ();
 sg13g2_fill_2 FILLER_27_921 ();
 sg13g2_fill_1 FILLER_27_984 ();
 sg13g2_decap_4 FILLER_27_1013 ();
 sg13g2_decap_4 FILLER_27_1022 ();
 sg13g2_fill_1 FILLER_27_1026 ();
 sg13g2_fill_2 FILLER_27_1056 ();
 sg13g2_fill_1 FILLER_27_1058 ();
 sg13g2_decap_8 FILLER_27_1063 ();
 sg13g2_decap_4 FILLER_27_1070 ();
 sg13g2_fill_2 FILLER_27_1074 ();
 sg13g2_fill_1 FILLER_27_1102 ();
 sg13g2_fill_2 FILLER_27_1119 ();
 sg13g2_fill_1 FILLER_27_1180 ();
 sg13g2_fill_1 FILLER_27_1191 ();
 sg13g2_fill_2 FILLER_27_1208 ();
 sg13g2_fill_1 FILLER_27_1210 ();
 sg13g2_fill_2 FILLER_27_1225 ();
 sg13g2_fill_1 FILLER_27_1227 ();
 sg13g2_fill_1 FILLER_27_1241 ();
 sg13g2_fill_1 FILLER_27_1252 ();
 sg13g2_decap_4 FILLER_27_1257 ();
 sg13g2_fill_1 FILLER_27_1261 ();
 sg13g2_decap_8 FILLER_27_1276 ();
 sg13g2_fill_2 FILLER_27_1294 ();
 sg13g2_fill_1 FILLER_27_1296 ();
 sg13g2_fill_1 FILLER_27_1302 ();
 sg13g2_fill_2 FILLER_27_1309 ();
 sg13g2_fill_1 FILLER_27_1311 ();
 sg13g2_fill_2 FILLER_27_1339 ();
 sg13g2_fill_1 FILLER_27_1392 ();
 sg13g2_fill_1 FILLER_27_1398 ();
 sg13g2_decap_4 FILLER_27_1415 ();
 sg13g2_fill_2 FILLER_27_1424 ();
 sg13g2_fill_2 FILLER_27_1436 ();
 sg13g2_fill_1 FILLER_27_1442 ();
 sg13g2_fill_2 FILLER_27_1539 ();
 sg13g2_fill_1 FILLER_27_1541 ();
 sg13g2_fill_2 FILLER_27_1568 ();
 sg13g2_fill_2 FILLER_27_1574 ();
 sg13g2_fill_2 FILLER_27_1602 ();
 sg13g2_fill_1 FILLER_27_1604 ();
 sg13g2_fill_1 FILLER_27_1614 ();
 sg13g2_fill_2 FILLER_27_1624 ();
 sg13g2_fill_1 FILLER_27_1631 ();
 sg13g2_decap_4 FILLER_27_1636 ();
 sg13g2_decap_8 FILLER_27_1656 ();
 sg13g2_fill_1 FILLER_27_1663 ();
 sg13g2_decap_8 FILLER_27_1668 ();
 sg13g2_decap_4 FILLER_27_1675 ();
 sg13g2_decap_4 FILLER_27_1689 ();
 sg13g2_fill_2 FILLER_27_1693 ();
 sg13g2_decap_8 FILLER_27_1699 ();
 sg13g2_fill_2 FILLER_27_1706 ();
 sg13g2_fill_1 FILLER_27_1712 ();
 sg13g2_decap_4 FILLER_27_1731 ();
 sg13g2_decap_8 FILLER_27_1748 ();
 sg13g2_decap_8 FILLER_27_1755 ();
 sg13g2_decap_8 FILLER_27_1762 ();
 sg13g2_fill_1 FILLER_27_1769 ();
 sg13g2_decap_8 FILLER_27_1774 ();
 sg13g2_decap_8 FILLER_27_1781 ();
 sg13g2_decap_8 FILLER_27_1788 ();
 sg13g2_decap_8 FILLER_27_1795 ();
 sg13g2_decap_8 FILLER_27_1802 ();
 sg13g2_decap_8 FILLER_27_1809 ();
 sg13g2_decap_8 FILLER_27_1816 ();
 sg13g2_decap_8 FILLER_27_1823 ();
 sg13g2_decap_4 FILLER_27_1830 ();
 sg13g2_fill_1 FILLER_27_1834 ();
 sg13g2_fill_1 FILLER_27_1839 ();
 sg13g2_fill_1 FILLER_27_1844 ();
 sg13g2_decap_8 FILLER_27_1861 ();
 sg13g2_decap_8 FILLER_27_1868 ();
 sg13g2_decap_8 FILLER_27_1875 ();
 sg13g2_decap_8 FILLER_27_1882 ();
 sg13g2_decap_8 FILLER_27_1889 ();
 sg13g2_decap_4 FILLER_27_1896 ();
 sg13g2_fill_2 FILLER_27_1900 ();
 sg13g2_decap_4 FILLER_27_1933 ();
 sg13g2_fill_1 FILLER_27_1937 ();
 sg13g2_fill_1 FILLER_27_1959 ();
 sg13g2_fill_2 FILLER_27_1988 ();
 sg13g2_fill_2 FILLER_27_1993 ();
 sg13g2_fill_1 FILLER_27_2005 ();
 sg13g2_fill_2 FILLER_27_2011 ();
 sg13g2_fill_2 FILLER_27_2073 ();
 sg13g2_fill_1 FILLER_27_2093 ();
 sg13g2_fill_1 FILLER_27_2177 ();
 sg13g2_fill_1 FILLER_27_2182 ();
 sg13g2_fill_1 FILLER_27_2209 ();
 sg13g2_fill_1 FILLER_27_2224 ();
 sg13g2_fill_1 FILLER_27_2235 ();
 sg13g2_fill_1 FILLER_27_2274 ();
 sg13g2_fill_1 FILLER_27_2301 ();
 sg13g2_decap_8 FILLER_27_2323 ();
 sg13g2_fill_1 FILLER_27_2330 ();
 sg13g2_fill_2 FILLER_27_2357 ();
 sg13g2_fill_1 FILLER_27_2369 ();
 sg13g2_fill_1 FILLER_27_2421 ();
 sg13g2_fill_1 FILLER_27_2448 ();
 sg13g2_fill_1 FILLER_27_2453 ();
 sg13g2_fill_2 FILLER_27_2480 ();
 sg13g2_fill_2 FILLER_27_2511 ();
 sg13g2_fill_2 FILLER_27_2569 ();
 sg13g2_decap_8 FILLER_27_2596 ();
 sg13g2_decap_8 FILLER_27_2603 ();
 sg13g2_decap_8 FILLER_27_2610 ();
 sg13g2_decap_8 FILLER_27_2617 ();
 sg13g2_decap_8 FILLER_27_2624 ();
 sg13g2_decap_8 FILLER_27_2631 ();
 sg13g2_decap_8 FILLER_27_2638 ();
 sg13g2_decap_8 FILLER_27_2645 ();
 sg13g2_decap_8 FILLER_27_2652 ();
 sg13g2_decap_8 FILLER_27_2659 ();
 sg13g2_decap_4 FILLER_27_2666 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_34 ();
 sg13g2_fill_2 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_decap_4 FILLER_28_419 ();
 sg13g2_fill_2 FILLER_28_423 ();
 sg13g2_fill_1 FILLER_28_455 ();
 sg13g2_fill_1 FILLER_28_460 ();
 sg13g2_fill_2 FILLER_28_558 ();
 sg13g2_fill_1 FILLER_28_640 ();
 sg13g2_fill_2 FILLER_28_644 ();
 sg13g2_fill_2 FILLER_28_672 ();
 sg13g2_fill_2 FILLER_28_681 ();
 sg13g2_fill_1 FILLER_28_722 ();
 sg13g2_decap_4 FILLER_28_748 ();
 sg13g2_fill_1 FILLER_28_761 ();
 sg13g2_decap_4 FILLER_28_791 ();
 sg13g2_fill_1 FILLER_28_795 ();
 sg13g2_fill_1 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_fill_1 FILLER_28_835 ();
 sg13g2_fill_1 FILLER_28_862 ();
 sg13g2_fill_1 FILLER_28_889 ();
 sg13g2_fill_1 FILLER_28_1005 ();
 sg13g2_fill_2 FILLER_28_1058 ();
 sg13g2_fill_2 FILLER_28_1084 ();
 sg13g2_fill_1 FILLER_28_1086 ();
 sg13g2_fill_2 FILLER_28_1091 ();
 sg13g2_fill_2 FILLER_28_1106 ();
 sg13g2_fill_1 FILLER_28_1124 ();
 sg13g2_fill_2 FILLER_28_1133 ();
 sg13g2_fill_1 FILLER_28_1141 ();
 sg13g2_fill_1 FILLER_28_1227 ();
 sg13g2_fill_1 FILLER_28_1232 ();
 sg13g2_fill_1 FILLER_28_1252 ();
 sg13g2_decap_8 FILLER_28_1270 ();
 sg13g2_fill_1 FILLER_28_1277 ();
 sg13g2_decap_8 FILLER_28_1288 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_fill_2 FILLER_28_1311 ();
 sg13g2_decap_4 FILLER_28_1317 ();
 sg13g2_fill_2 FILLER_28_1321 ();
 sg13g2_decap_4 FILLER_28_1328 ();
 sg13g2_fill_1 FILLER_28_1332 ();
 sg13g2_fill_2 FILLER_28_1349 ();
 sg13g2_decap_4 FILLER_28_1358 ();
 sg13g2_fill_2 FILLER_28_1381 ();
 sg13g2_decap_4 FILLER_28_1408 ();
 sg13g2_fill_1 FILLER_28_1412 ();
 sg13g2_fill_1 FILLER_28_1434 ();
 sg13g2_fill_2 FILLER_28_1502 ();
 sg13g2_fill_1 FILLER_28_1530 ();
 sg13g2_fill_2 FILLER_28_1562 ();
 sg13g2_decap_8 FILLER_28_1574 ();
 sg13g2_fill_1 FILLER_28_1581 ();
 sg13g2_fill_2 FILLER_28_1586 ();
 sg13g2_decap_8 FILLER_28_1592 ();
 sg13g2_decap_4 FILLER_28_1599 ();
 sg13g2_fill_1 FILLER_28_1603 ();
 sg13g2_fill_1 FILLER_28_1611 ();
 sg13g2_fill_1 FILLER_28_1617 ();
 sg13g2_decap_8 FILLER_28_1628 ();
 sg13g2_fill_2 FILLER_28_1635 ();
 sg13g2_decap_8 FILLER_28_1672 ();
 sg13g2_fill_2 FILLER_28_1689 ();
 sg13g2_decap_8 FILLER_28_1717 ();
 sg13g2_decap_8 FILLER_28_1724 ();
 sg13g2_decap_8 FILLER_28_1731 ();
 sg13g2_decap_8 FILLER_28_1738 ();
 sg13g2_decap_8 FILLER_28_1745 ();
 sg13g2_decap_4 FILLER_28_1752 ();
 sg13g2_decap_8 FILLER_28_1760 ();
 sg13g2_decap_8 FILLER_28_1767 ();
 sg13g2_decap_8 FILLER_28_1774 ();
 sg13g2_decap_8 FILLER_28_1781 ();
 sg13g2_decap_8 FILLER_28_1788 ();
 sg13g2_decap_4 FILLER_28_1795 ();
 sg13g2_fill_1 FILLER_28_1799 ();
 sg13g2_fill_2 FILLER_28_1805 ();
 sg13g2_fill_1 FILLER_28_1807 ();
 sg13g2_decap_4 FILLER_28_1829 ();
 sg13g2_fill_1 FILLER_28_1833 ();
 sg13g2_fill_2 FILLER_28_1844 ();
 sg13g2_fill_1 FILLER_28_1876 ();
 sg13g2_decap_8 FILLER_28_1880 ();
 sg13g2_decap_8 FILLER_28_1891 ();
 sg13g2_decap_8 FILLER_28_1898 ();
 sg13g2_decap_8 FILLER_28_1905 ();
 sg13g2_decap_8 FILLER_28_1912 ();
 sg13g2_fill_2 FILLER_28_1919 ();
 sg13g2_fill_1 FILLER_28_1921 ();
 sg13g2_fill_1 FILLER_28_1997 ();
 sg13g2_fill_2 FILLER_28_2011 ();
 sg13g2_fill_1 FILLER_28_2062 ();
 sg13g2_fill_2 FILLER_28_2102 ();
 sg13g2_fill_2 FILLER_28_2122 ();
 sg13g2_fill_1 FILLER_28_2124 ();
 sg13g2_decap_8 FILLER_28_2160 ();
 sg13g2_decap_8 FILLER_28_2167 ();
 sg13g2_fill_1 FILLER_28_2174 ();
 sg13g2_decap_8 FILLER_28_2193 ();
 sg13g2_decap_8 FILLER_28_2200 ();
 sg13g2_decap_8 FILLER_28_2207 ();
 sg13g2_decap_8 FILLER_28_2214 ();
 sg13g2_fill_1 FILLER_28_2221 ();
 sg13g2_fill_2 FILLER_28_2226 ();
 sg13g2_fill_1 FILLER_28_2228 ();
 sg13g2_decap_4 FILLER_28_2246 ();
 sg13g2_fill_1 FILLER_28_2250 ();
 sg13g2_fill_1 FILLER_28_2270 ();
 sg13g2_fill_1 FILLER_28_2278 ();
 sg13g2_decap_4 FILLER_28_2297 ();
 sg13g2_fill_1 FILLER_28_2301 ();
 sg13g2_fill_1 FILLER_28_2338 ();
 sg13g2_fill_1 FILLER_28_2376 ();
 sg13g2_fill_2 FILLER_28_2420 ();
 sg13g2_fill_2 FILLER_28_2448 ();
 sg13g2_fill_1 FILLER_28_2476 ();
 sg13g2_fill_1 FILLER_28_2487 ();
 sg13g2_fill_1 FILLER_28_2492 ();
 sg13g2_fill_2 FILLER_28_2519 ();
 sg13g2_decap_8 FILLER_28_2594 ();
 sg13g2_decap_8 FILLER_28_2601 ();
 sg13g2_decap_8 FILLER_28_2608 ();
 sg13g2_decap_8 FILLER_28_2615 ();
 sg13g2_decap_8 FILLER_28_2622 ();
 sg13g2_decap_8 FILLER_28_2629 ();
 sg13g2_decap_8 FILLER_28_2636 ();
 sg13g2_decap_8 FILLER_28_2643 ();
 sg13g2_decap_8 FILLER_28_2650 ();
 sg13g2_decap_8 FILLER_28_2657 ();
 sg13g2_decap_4 FILLER_28_2664 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_fill_2 FILLER_29_455 ();
 sg13g2_fill_2 FILLER_29_502 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_fill_2 FILLER_29_560 ();
 sg13g2_fill_2 FILLER_29_572 ();
 sg13g2_fill_1 FILLER_29_624 ();
 sg13g2_fill_1 FILLER_29_665 ();
 sg13g2_fill_1 FILLER_29_677 ();
 sg13g2_fill_2 FILLER_29_686 ();
 sg13g2_fill_1 FILLER_29_691 ();
 sg13g2_fill_2 FILLER_29_711 ();
 sg13g2_fill_2 FILLER_29_718 ();
 sg13g2_fill_1 FILLER_29_720 ();
 sg13g2_fill_1 FILLER_29_725 ();
 sg13g2_fill_1 FILLER_29_730 ();
 sg13g2_fill_1 FILLER_29_757 ();
 sg13g2_fill_2 FILLER_29_792 ();
 sg13g2_decap_8 FILLER_29_820 ();
 sg13g2_fill_1 FILLER_29_827 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_4 FILLER_29_847 ();
 sg13g2_fill_2 FILLER_29_851 ();
 sg13g2_fill_2 FILLER_29_884 ();
 sg13g2_fill_1 FILLER_29_886 ();
 sg13g2_fill_2 FILLER_29_943 ();
 sg13g2_fill_1 FILLER_29_980 ();
 sg13g2_fill_2 FILLER_29_1012 ();
 sg13g2_decap_4 FILLER_29_1044 ();
 sg13g2_fill_1 FILLER_29_1048 ();
 sg13g2_fill_2 FILLER_29_1084 ();
 sg13g2_fill_1 FILLER_29_1086 ();
 sg13g2_fill_2 FILLER_29_1118 ();
 sg13g2_fill_1 FILLER_29_1152 ();
 sg13g2_fill_1 FILLER_29_1157 ();
 sg13g2_fill_1 FILLER_29_1162 ();
 sg13g2_fill_1 FILLER_29_1167 ();
 sg13g2_fill_1 FILLER_29_1171 ();
 sg13g2_fill_1 FILLER_29_1177 ();
 sg13g2_fill_1 FILLER_29_1182 ();
 sg13g2_fill_2 FILLER_29_1201 ();
 sg13g2_fill_1 FILLER_29_1213 ();
 sg13g2_fill_1 FILLER_29_1219 ();
 sg13g2_fill_1 FILLER_29_1236 ();
 sg13g2_fill_2 FILLER_29_1285 ();
 sg13g2_fill_1 FILLER_29_1297 ();
 sg13g2_fill_1 FILLER_29_1303 ();
 sg13g2_fill_1 FILLER_29_1309 ();
 sg13g2_fill_1 FILLER_29_1315 ();
 sg13g2_fill_1 FILLER_29_1326 ();
 sg13g2_decap_4 FILLER_29_1361 ();
 sg13g2_fill_2 FILLER_29_1370 ();
 sg13g2_fill_2 FILLER_29_1410 ();
 sg13g2_fill_1 FILLER_29_1412 ();
 sg13g2_fill_1 FILLER_29_1439 ();
 sg13g2_fill_1 FILLER_29_1500 ();
 sg13g2_fill_2 FILLER_29_1527 ();
 sg13g2_fill_1 FILLER_29_1529 ();
 sg13g2_fill_2 FILLER_29_1543 ();
 sg13g2_fill_1 FILLER_29_1545 ();
 sg13g2_decap_8 FILLER_29_1550 ();
 sg13g2_decap_8 FILLER_29_1557 ();
 sg13g2_decap_8 FILLER_29_1564 ();
 sg13g2_decap_8 FILLER_29_1571 ();
 sg13g2_decap_8 FILLER_29_1578 ();
 sg13g2_decap_8 FILLER_29_1585 ();
 sg13g2_decap_8 FILLER_29_1592 ();
 sg13g2_decap_8 FILLER_29_1599 ();
 sg13g2_fill_1 FILLER_29_1606 ();
 sg13g2_fill_2 FILLER_29_1612 ();
 sg13g2_decap_4 FILLER_29_1625 ();
 sg13g2_decap_4 FILLER_29_1662 ();
 sg13g2_fill_2 FILLER_29_1670 ();
 sg13g2_fill_1 FILLER_29_1672 ();
 sg13g2_fill_1 FILLER_29_1687 ();
 sg13g2_fill_2 FILLER_29_1714 ();
 sg13g2_fill_1 FILLER_29_1716 ();
 sg13g2_decap_8 FILLER_29_1756 ();
 sg13g2_decap_8 FILLER_29_1763 ();
 sg13g2_decap_4 FILLER_29_1770 ();
 sg13g2_fill_1 FILLER_29_1783 ();
 sg13g2_fill_1 FILLER_29_1795 ();
 sg13g2_fill_2 FILLER_29_1815 ();
 sg13g2_fill_2 FILLER_29_1852 ();
 sg13g2_fill_1 FILLER_29_1905 ();
 sg13g2_decap_8 FILLER_29_1910 ();
 sg13g2_decap_4 FILLER_29_1917 ();
 sg13g2_fill_2 FILLER_29_1921 ();
 sg13g2_fill_2 FILLER_29_2019 ();
 sg13g2_fill_2 FILLER_29_2067 ();
 sg13g2_fill_1 FILLER_29_2069 ();
 sg13g2_fill_2 FILLER_29_2073 ();
 sg13g2_fill_1 FILLER_29_2075 ();
 sg13g2_decap_8 FILLER_29_2105 ();
 sg13g2_decap_8 FILLER_29_2112 ();
 sg13g2_decap_8 FILLER_29_2119 ();
 sg13g2_decap_8 FILLER_29_2126 ();
 sg13g2_fill_2 FILLER_29_2151 ();
 sg13g2_fill_1 FILLER_29_2153 ();
 sg13g2_fill_1 FILLER_29_2164 ();
 sg13g2_decap_8 FILLER_29_2190 ();
 sg13g2_decap_8 FILLER_29_2197 ();
 sg13g2_decap_4 FILLER_29_2204 ();
 sg13g2_fill_2 FILLER_29_2208 ();
 sg13g2_decap_8 FILLER_29_2214 ();
 sg13g2_fill_1 FILLER_29_2273 ();
 sg13g2_fill_1 FILLER_29_2300 ();
 sg13g2_fill_1 FILLER_29_2311 ();
 sg13g2_fill_1 FILLER_29_2442 ();
 sg13g2_fill_2 FILLER_29_2453 ();
 sg13g2_fill_2 FILLER_29_2507 ();
 sg13g2_decap_8 FILLER_29_2591 ();
 sg13g2_decap_8 FILLER_29_2598 ();
 sg13g2_decap_8 FILLER_29_2605 ();
 sg13g2_decap_8 FILLER_29_2612 ();
 sg13g2_decap_8 FILLER_29_2619 ();
 sg13g2_decap_8 FILLER_29_2626 ();
 sg13g2_decap_8 FILLER_29_2633 ();
 sg13g2_decap_8 FILLER_29_2640 ();
 sg13g2_decap_8 FILLER_29_2647 ();
 sg13g2_decap_8 FILLER_29_2654 ();
 sg13g2_decap_8 FILLER_29_2661 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_8 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_2 FILLER_30_421 ();
 sg13g2_fill_1 FILLER_30_468 ();
 sg13g2_fill_1 FILLER_30_503 ();
 sg13g2_fill_2 FILLER_30_522 ();
 sg13g2_fill_1 FILLER_30_545 ();
 sg13g2_fill_2 FILLER_30_610 ();
 sg13g2_fill_1 FILLER_30_654 ();
 sg13g2_fill_2 FILLER_30_683 ();
 sg13g2_fill_1 FILLER_30_736 ();
 sg13g2_fill_1 FILLER_30_799 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_fill_1 FILLER_30_866 ();
 sg13g2_decap_4 FILLER_30_876 ();
 sg13g2_fill_2 FILLER_30_880 ();
 sg13g2_fill_1 FILLER_30_892 ();
 sg13g2_decap_4 FILLER_30_903 ();
 sg13g2_fill_2 FILLER_30_921 ();
 sg13g2_fill_2 FILLER_30_928 ();
 sg13g2_fill_2 FILLER_30_947 ();
 sg13g2_fill_2 FILLER_30_980 ();
 sg13g2_fill_1 FILLER_30_982 ();
 sg13g2_fill_2 FILLER_30_993 ();
 sg13g2_fill_1 FILLER_30_995 ();
 sg13g2_fill_1 FILLER_30_1001 ();
 sg13g2_fill_1 FILLER_30_1040 ();
 sg13g2_decap_8 FILLER_30_1163 ();
 sg13g2_decap_4 FILLER_30_1170 ();
 sg13g2_fill_2 FILLER_30_1174 ();
 sg13g2_fill_2 FILLER_30_1181 ();
 sg13g2_fill_1 FILLER_30_1183 ();
 sg13g2_fill_2 FILLER_30_1201 ();
 sg13g2_fill_1 FILLER_30_1203 ();
 sg13g2_fill_2 FILLER_30_1209 ();
 sg13g2_fill_1 FILLER_30_1273 ();
 sg13g2_fill_2 FILLER_30_1286 ();
 sg13g2_fill_1 FILLER_30_1288 ();
 sg13g2_fill_2 FILLER_30_1294 ();
 sg13g2_fill_1 FILLER_30_1296 ();
 sg13g2_fill_1 FILLER_30_1313 ();
 sg13g2_fill_1 FILLER_30_1321 ();
 sg13g2_decap_4 FILLER_30_1347 ();
 sg13g2_fill_1 FILLER_30_1361 ();
 sg13g2_fill_2 FILLER_30_1373 ();
 sg13g2_fill_1 FILLER_30_1375 ();
 sg13g2_fill_1 FILLER_30_1384 ();
 sg13g2_fill_2 FILLER_30_1402 ();
 sg13g2_fill_1 FILLER_30_1425 ();
 sg13g2_decap_4 FILLER_30_1434 ();
 sg13g2_fill_2 FILLER_30_1446 ();
 sg13g2_decap_4 FILLER_30_1452 ();
 sg13g2_fill_2 FILLER_30_1459 ();
 sg13g2_fill_1 FILLER_30_1523 ();
 sg13g2_fill_1 FILLER_30_1528 ();
 sg13g2_decap_8 FILLER_30_1565 ();
 sg13g2_decap_4 FILLER_30_1577 ();
 sg13g2_fill_1 FILLER_30_1581 ();
 sg13g2_fill_1 FILLER_30_1619 ();
 sg13g2_decap_8 FILLER_30_1625 ();
 sg13g2_fill_2 FILLER_30_1632 ();
 sg13g2_fill_1 FILLER_30_1634 ();
 sg13g2_decap_4 FILLER_30_1639 ();
 sg13g2_decap_4 FILLER_30_1703 ();
 sg13g2_fill_2 FILLER_30_1707 ();
 sg13g2_decap_8 FILLER_30_1753 ();
 sg13g2_decap_4 FILLER_30_1760 ();
 sg13g2_fill_1 FILLER_30_1777 ();
 sg13g2_fill_2 FILLER_30_1820 ();
 sg13g2_fill_2 FILLER_30_1861 ();
 sg13g2_fill_1 FILLER_30_1897 ();
 sg13g2_fill_1 FILLER_30_1902 ();
 sg13g2_fill_1 FILLER_30_1907 ();
 sg13g2_fill_2 FILLER_30_1925 ();
 sg13g2_fill_2 FILLER_30_2010 ();
 sg13g2_decap_8 FILLER_30_2081 ();
 sg13g2_decap_8 FILLER_30_2088 ();
 sg13g2_decap_8 FILLER_30_2095 ();
 sg13g2_decap_8 FILLER_30_2102 ();
 sg13g2_decap_4 FILLER_30_2109 ();
 sg13g2_fill_1 FILLER_30_2123 ();
 sg13g2_fill_1 FILLER_30_2150 ();
 sg13g2_fill_1 FILLER_30_2177 ();
 sg13g2_fill_2 FILLER_30_2188 ();
 sg13g2_fill_2 FILLER_30_2194 ();
 sg13g2_fill_1 FILLER_30_2232 ();
 sg13g2_fill_1 FILLER_30_2259 ();
 sg13g2_fill_1 FILLER_30_2286 ();
 sg13g2_fill_1 FILLER_30_2308 ();
 sg13g2_fill_1 FILLER_30_2313 ();
 sg13g2_fill_1 FILLER_30_2340 ();
 sg13g2_decap_8 FILLER_30_2433 ();
 sg13g2_fill_1 FILLER_30_2440 ();
 sg13g2_fill_2 FILLER_30_2466 ();
 sg13g2_decap_4 FILLER_30_2525 ();
 sg13g2_fill_2 FILLER_30_2529 ();
 sg13g2_fill_1 FILLER_30_2541 ();
 sg13g2_decap_8 FILLER_30_2556 ();
 sg13g2_decap_4 FILLER_30_2563 ();
 sg13g2_fill_2 FILLER_30_2567 ();
 sg13g2_decap_8 FILLER_30_2599 ();
 sg13g2_decap_8 FILLER_30_2606 ();
 sg13g2_decap_8 FILLER_30_2613 ();
 sg13g2_decap_8 FILLER_30_2620 ();
 sg13g2_decap_8 FILLER_30_2627 ();
 sg13g2_decap_8 FILLER_30_2634 ();
 sg13g2_decap_8 FILLER_30_2641 ();
 sg13g2_decap_8 FILLER_30_2648 ();
 sg13g2_decap_8 FILLER_30_2655 ();
 sg13g2_decap_8 FILLER_30_2662 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_123 ();
 sg13g2_decap_4 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_4 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_302 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_389 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_decap_4 FILLER_31_424 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_fill_1 FILLER_31_440 ();
 sg13g2_fill_1 FILLER_31_527 ();
 sg13g2_fill_2 FILLER_31_532 ();
 sg13g2_fill_1 FILLER_31_563 ();
 sg13g2_fill_1 FILLER_31_606 ();
 sg13g2_fill_2 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_4 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_8 FILLER_31_857 ();
 sg13g2_decap_8 FILLER_31_864 ();
 sg13g2_fill_2 FILLER_31_875 ();
 sg13g2_fill_1 FILLER_31_877 ();
 sg13g2_decap_8 FILLER_31_908 ();
 sg13g2_decap_4 FILLER_31_915 ();
 sg13g2_fill_1 FILLER_31_924 ();
 sg13g2_fill_1 FILLER_31_933 ();
 sg13g2_fill_1 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_fill_2 FILLER_31_1002 ();
 sg13g2_fill_1 FILLER_31_1004 ();
 sg13g2_fill_1 FILLER_31_1062 ();
 sg13g2_fill_2 FILLER_31_1069 ();
 sg13g2_fill_2 FILLER_31_1078 ();
 sg13g2_fill_1 FILLER_31_1111 ();
 sg13g2_decap_8 FILLER_31_1164 ();
 sg13g2_decap_4 FILLER_31_1171 ();
 sg13g2_fill_1 FILLER_31_1175 ();
 sg13g2_fill_2 FILLER_31_1185 ();
 sg13g2_fill_2 FILLER_31_1245 ();
 sg13g2_fill_2 FILLER_31_1254 ();
 sg13g2_fill_1 FILLER_31_1287 ();
 sg13g2_decap_4 FILLER_31_1300 ();
 sg13g2_fill_2 FILLER_31_1304 ();
 sg13g2_fill_1 FILLER_31_1321 ();
 sg13g2_fill_1 FILLER_31_1327 ();
 sg13g2_fill_1 FILLER_31_1344 ();
 sg13g2_fill_2 FILLER_31_1364 ();
 sg13g2_fill_1 FILLER_31_1366 ();
 sg13g2_fill_2 FILLER_31_1409 ();
 sg13g2_fill_1 FILLER_31_1411 ();
 sg13g2_decap_4 FILLER_31_1442 ();
 sg13g2_fill_1 FILLER_31_1446 ();
 sg13g2_fill_2 FILLER_31_1467 ();
 sg13g2_fill_1 FILLER_31_1479 ();
 sg13g2_fill_1 FILLER_31_1484 ();
 sg13g2_fill_1 FILLER_31_1489 ();
 sg13g2_fill_1 FILLER_31_1493 ();
 sg13g2_fill_1 FILLER_31_1504 ();
 sg13g2_fill_2 FILLER_31_1509 ();
 sg13g2_fill_1 FILLER_31_1515 ();
 sg13g2_decap_4 FILLER_31_1641 ();
 sg13g2_fill_1 FILLER_31_1645 ();
 sg13g2_decap_8 FILLER_31_1666 ();
 sg13g2_decap_4 FILLER_31_1673 ();
 sg13g2_fill_1 FILLER_31_1677 ();
 sg13g2_fill_1 FILLER_31_1682 ();
 sg13g2_decap_8 FILLER_31_1696 ();
 sg13g2_fill_2 FILLER_31_1703 ();
 sg13g2_fill_1 FILLER_31_1705 ();
 sg13g2_fill_1 FILLER_31_1737 ();
 sg13g2_decap_4 FILLER_31_1742 ();
 sg13g2_fill_2 FILLER_31_1746 ();
 sg13g2_fill_2 FILLER_31_1771 ();
 sg13g2_fill_2 FILLER_31_1832 ();
 sg13g2_fill_2 FILLER_31_1838 ();
 sg13g2_fill_2 FILLER_31_1875 ();
 sg13g2_fill_2 FILLER_31_1914 ();
 sg13g2_fill_1 FILLER_31_1921 ();
 sg13g2_fill_1 FILLER_31_1930 ();
 sg13g2_fill_1 FILLER_31_1935 ();
 sg13g2_fill_1 FILLER_31_2028 ();
 sg13g2_fill_2 FILLER_31_2033 ();
 sg13g2_fill_2 FILLER_31_2071 ();
 sg13g2_fill_2 FILLER_31_2099 ();
 sg13g2_fill_1 FILLER_31_2101 ();
 sg13g2_fill_2 FILLER_31_2112 ();
 sg13g2_fill_1 FILLER_31_2114 ();
 sg13g2_fill_2 FILLER_31_2151 ();
 sg13g2_fill_1 FILLER_31_2153 ();
 sg13g2_fill_2 FILLER_31_2180 ();
 sg13g2_fill_1 FILLER_31_2208 ();
 sg13g2_fill_1 FILLER_31_2256 ();
 sg13g2_fill_2 FILLER_31_2326 ();
 sg13g2_fill_2 FILLER_31_2338 ();
 sg13g2_fill_2 FILLER_31_2345 ();
 sg13g2_fill_1 FILLER_31_2347 ();
 sg13g2_fill_1 FILLER_31_2356 ();
 sg13g2_decap_4 FILLER_31_2361 ();
 sg13g2_fill_2 FILLER_31_2451 ();
 sg13g2_decap_8 FILLER_31_2512 ();
 sg13g2_decap_8 FILLER_31_2519 ();
 sg13g2_decap_8 FILLER_31_2526 ();
 sg13g2_decap_8 FILLER_31_2533 ();
 sg13g2_decap_8 FILLER_31_2540 ();
 sg13g2_decap_8 FILLER_31_2547 ();
 sg13g2_decap_8 FILLER_31_2554 ();
 sg13g2_decap_4 FILLER_31_2561 ();
 sg13g2_fill_1 FILLER_31_2565 ();
 sg13g2_fill_1 FILLER_31_2570 ();
 sg13g2_decap_8 FILLER_31_2581 ();
 sg13g2_decap_8 FILLER_31_2588 ();
 sg13g2_decap_8 FILLER_31_2595 ();
 sg13g2_decap_8 FILLER_31_2602 ();
 sg13g2_decap_8 FILLER_31_2609 ();
 sg13g2_decap_8 FILLER_31_2616 ();
 sg13g2_decap_8 FILLER_31_2623 ();
 sg13g2_decap_8 FILLER_31_2630 ();
 sg13g2_decap_8 FILLER_31_2637 ();
 sg13g2_decap_8 FILLER_31_2644 ();
 sg13g2_decap_8 FILLER_31_2651 ();
 sg13g2_decap_8 FILLER_31_2658 ();
 sg13g2_decap_4 FILLER_31_2665 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_354 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_fill_2 FILLER_32_430 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_453 ();
 sg13g2_fill_1 FILLER_32_465 ();
 sg13g2_fill_1 FILLER_32_540 ();
 sg13g2_fill_1 FILLER_32_620 ();
 sg13g2_fill_2 FILLER_32_657 ();
 sg13g2_decap_4 FILLER_32_750 ();
 sg13g2_fill_2 FILLER_32_754 ();
 sg13g2_fill_2 FILLER_32_774 ();
 sg13g2_fill_2 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_4 FILLER_32_796 ();
 sg13g2_fill_2 FILLER_32_800 ();
 sg13g2_fill_2 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_4 FILLER_32_857 ();
 sg13g2_fill_2 FILLER_32_861 ();
 sg13g2_fill_2 FILLER_32_889 ();
 sg13g2_fill_1 FILLER_32_891 ();
 sg13g2_fill_2 FILLER_32_909 ();
 sg13g2_fill_2 FILLER_32_967 ();
 sg13g2_fill_1 FILLER_32_978 ();
 sg13g2_fill_2 FILLER_32_1000 ();
 sg13g2_fill_2 FILLER_32_1012 ();
 sg13g2_fill_1 FILLER_32_1014 ();
 sg13g2_fill_2 FILLER_32_1040 ();
 sg13g2_fill_2 FILLER_32_1095 ();
 sg13g2_fill_1 FILLER_32_1143 ();
 sg13g2_decap_8 FILLER_32_1151 ();
 sg13g2_decap_8 FILLER_32_1158 ();
 sg13g2_decap_8 FILLER_32_1165 ();
 sg13g2_decap_8 FILLER_32_1172 ();
 sg13g2_fill_2 FILLER_32_1209 ();
 sg13g2_fill_2 FILLER_32_1216 ();
 sg13g2_fill_1 FILLER_32_1218 ();
 sg13g2_fill_1 FILLER_32_1224 ();
 sg13g2_fill_2 FILLER_32_1230 ();
 sg13g2_fill_1 FILLER_32_1237 ();
 sg13g2_decap_8 FILLER_32_1268 ();
 sg13g2_decap_8 FILLER_32_1285 ();
 sg13g2_decap_8 FILLER_32_1292 ();
 sg13g2_decap_8 FILLER_32_1299 ();
 sg13g2_decap_8 FILLER_32_1306 ();
 sg13g2_decap_8 FILLER_32_1313 ();
 sg13g2_decap_8 FILLER_32_1320 ();
 sg13g2_decap_8 FILLER_32_1327 ();
 sg13g2_fill_1 FILLER_32_1349 ();
 sg13g2_decap_8 FILLER_32_1355 ();
 sg13g2_fill_2 FILLER_32_1362 ();
 sg13g2_fill_1 FILLER_32_1364 ();
 sg13g2_decap_8 FILLER_32_1377 ();
 sg13g2_decap_8 FILLER_32_1390 ();
 sg13g2_fill_2 FILLER_32_1397 ();
 sg13g2_decap_8 FILLER_32_1466 ();
 sg13g2_decap_8 FILLER_32_1473 ();
 sg13g2_fill_2 FILLER_32_1480 ();
 sg13g2_decap_8 FILLER_32_1487 ();
 sg13g2_decap_4 FILLER_32_1494 ();
 sg13g2_fill_1 FILLER_32_1508 ();
 sg13g2_fill_1 FILLER_32_1513 ();
 sg13g2_decap_8 FILLER_32_1519 ();
 sg13g2_decap_4 FILLER_32_1526 ();
 sg13g2_decap_4 FILLER_32_1534 ();
 sg13g2_fill_1 FILLER_32_1538 ();
 sg13g2_fill_2 FILLER_32_1552 ();
 sg13g2_fill_1 FILLER_32_1554 ();
 sg13g2_fill_2 FILLER_32_1597 ();
 sg13g2_fill_1 FILLER_32_1616 ();
 sg13g2_fill_1 FILLER_32_1624 ();
 sg13g2_fill_1 FILLER_32_1630 ();
 sg13g2_fill_2 FILLER_32_1667 ();
 sg13g2_fill_2 FILLER_32_1695 ();
 sg13g2_decap_8 FILLER_32_1702 ();
 sg13g2_decap_4 FILLER_32_1709 ();
 sg13g2_decap_8 FILLER_32_1721 ();
 sg13g2_fill_1 FILLER_32_1728 ();
 sg13g2_fill_2 FILLER_32_1757 ();
 sg13g2_fill_1 FILLER_32_1766 ();
 sg13g2_fill_1 FILLER_32_1829 ();
 sg13g2_fill_1 FILLER_32_1835 ();
 sg13g2_fill_2 FILLER_32_1840 ();
 sg13g2_fill_2 FILLER_32_1861 ();
 sg13g2_fill_1 FILLER_32_1885 ();
 sg13g2_fill_1 FILLER_32_1896 ();
 sg13g2_fill_2 FILLER_32_1906 ();
 sg13g2_fill_1 FILLER_32_1912 ();
 sg13g2_fill_2 FILLER_32_1918 ();
 sg13g2_fill_2 FILLER_32_1928 ();
 sg13g2_decap_8 FILLER_32_1956 ();
 sg13g2_fill_2 FILLER_32_1963 ();
 sg13g2_fill_1 FILLER_32_2012 ();
 sg13g2_fill_2 FILLER_32_2075 ();
 sg13g2_fill_2 FILLER_32_2164 ();
 sg13g2_fill_2 FILLER_32_2170 ();
 sg13g2_fill_1 FILLER_32_2172 ();
 sg13g2_fill_1 FILLER_32_2177 ();
 sg13g2_fill_1 FILLER_32_2204 ();
 sg13g2_fill_2 FILLER_32_2215 ();
 sg13g2_fill_1 FILLER_32_2221 ();
 sg13g2_decap_8 FILLER_32_2226 ();
 sg13g2_fill_2 FILLER_32_2233 ();
 sg13g2_decap_4 FILLER_32_2252 ();
 sg13g2_fill_1 FILLER_32_2256 ();
 sg13g2_fill_2 FILLER_32_2274 ();
 sg13g2_fill_1 FILLER_32_2276 ();
 sg13g2_fill_2 FILLER_32_2295 ();
 sg13g2_fill_1 FILLER_32_2297 ();
 sg13g2_decap_8 FILLER_32_2302 ();
 sg13g2_decap_8 FILLER_32_2309 ();
 sg13g2_decap_8 FILLER_32_2316 ();
 sg13g2_fill_1 FILLER_32_2323 ();
 sg13g2_decap_4 FILLER_32_2334 ();
 sg13g2_fill_1 FILLER_32_2338 ();
 sg13g2_decap_8 FILLER_32_2343 ();
 sg13g2_decap_8 FILLER_32_2350 ();
 sg13g2_decap_8 FILLER_32_2357 ();
 sg13g2_decap_8 FILLER_32_2364 ();
 sg13g2_decap_8 FILLER_32_2371 ();
 sg13g2_decap_4 FILLER_32_2378 ();
 sg13g2_fill_2 FILLER_32_2415 ();
 sg13g2_decap_4 FILLER_32_2443 ();
 sg13g2_decap_4 FILLER_32_2493 ();
 sg13g2_decap_8 FILLER_32_2501 ();
 sg13g2_decap_8 FILLER_32_2508 ();
 sg13g2_decap_8 FILLER_32_2515 ();
 sg13g2_decap_8 FILLER_32_2522 ();
 sg13g2_decap_4 FILLER_32_2529 ();
 sg13g2_fill_1 FILLER_32_2611 ();
 sg13g2_decap_8 FILLER_32_2630 ();
 sg13g2_decap_8 FILLER_32_2637 ();
 sg13g2_decap_8 FILLER_32_2644 ();
 sg13g2_decap_8 FILLER_32_2651 ();
 sg13g2_decap_8 FILLER_32_2658 ();
 sg13g2_decap_4 FILLER_32_2665 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_115 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_405 ();
 sg13g2_fill_1 FILLER_33_415 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_fill_1 FILLER_33_485 ();
 sg13g2_fill_1 FILLER_33_502 ();
 sg13g2_fill_1 FILLER_33_519 ();
 sg13g2_fill_2 FILLER_33_526 ();
 sg13g2_decap_8 FILLER_33_576 ();
 sg13g2_decap_4 FILLER_33_583 ();
 sg13g2_fill_1 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_640 ();
 sg13g2_fill_1 FILLER_33_698 ();
 sg13g2_decap_4 FILLER_33_729 ();
 sg13g2_fill_1 FILLER_33_733 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_fill_1 FILLER_33_764 ();
 sg13g2_fill_2 FILLER_33_773 ();
 sg13g2_fill_1 FILLER_33_775 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_4 FILLER_33_793 ();
 sg13g2_fill_2 FILLER_33_797 ();
 sg13g2_fill_1 FILLER_33_829 ();
 sg13g2_fill_1 FILLER_33_856 ();
 sg13g2_fill_1 FILLER_33_867 ();
 sg13g2_fill_2 FILLER_33_917 ();
 sg13g2_fill_1 FILLER_33_919 ();
 sg13g2_fill_1 FILLER_33_1006 ();
 sg13g2_fill_2 FILLER_33_1035 ();
 sg13g2_fill_2 FILLER_33_1075 ();
 sg13g2_fill_1 FILLER_33_1095 ();
 sg13g2_fill_2 FILLER_33_1145 ();
 sg13g2_fill_1 FILLER_33_1147 ();
 sg13g2_decap_8 FILLER_33_1177 ();
 sg13g2_decap_8 FILLER_33_1184 ();
 sg13g2_decap_4 FILLER_33_1201 ();
 sg13g2_decap_8 FILLER_33_1210 ();
 sg13g2_fill_1 FILLER_33_1248 ();
 sg13g2_decap_8 FILLER_33_1285 ();
 sg13g2_decap_8 FILLER_33_1292 ();
 sg13g2_decap_4 FILLER_33_1325 ();
 sg13g2_fill_2 FILLER_33_1329 ();
 sg13g2_decap_8 FILLER_33_1403 ();
 sg13g2_fill_1 FILLER_33_1410 ();
 sg13g2_fill_2 FILLER_33_1437 ();
 sg13g2_fill_1 FILLER_33_1439 ();
 sg13g2_fill_2 FILLER_33_1450 ();
 sg13g2_fill_1 FILLER_33_1452 ();
 sg13g2_fill_2 FILLER_33_1463 ();
 sg13g2_fill_1 FILLER_33_1465 ();
 sg13g2_decap_8 FILLER_33_1470 ();
 sg13g2_decap_8 FILLER_33_1477 ();
 sg13g2_fill_2 FILLER_33_1484 ();
 sg13g2_decap_8 FILLER_33_1517 ();
 sg13g2_fill_1 FILLER_33_1524 ();
 sg13g2_decap_8 FILLER_33_1529 ();
 sg13g2_fill_1 FILLER_33_1536 ();
 sg13g2_decap_8 FILLER_33_1568 ();
 sg13g2_fill_1 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1580 ();
 sg13g2_decap_8 FILLER_33_1587 ();
 sg13g2_decap_4 FILLER_33_1594 ();
 sg13g2_fill_1 FILLER_33_1598 ();
 sg13g2_fill_2 FILLER_33_1606 ();
 sg13g2_fill_1 FILLER_33_1608 ();
 sg13g2_fill_1 FILLER_33_1636 ();
 sg13g2_decap_8 FILLER_33_1663 ();
 sg13g2_decap_8 FILLER_33_1670 ();
 sg13g2_fill_2 FILLER_33_1677 ();
 sg13g2_fill_1 FILLER_33_1679 ();
 sg13g2_fill_2 FILLER_33_1688 ();
 sg13g2_fill_1 FILLER_33_1710 ();
 sg13g2_decap_8 FILLER_33_1742 ();
 sg13g2_fill_2 FILLER_33_1749 ();
 sg13g2_fill_1 FILLER_33_1756 ();
 sg13g2_fill_1 FILLER_33_1775 ();
 sg13g2_fill_2 FILLER_33_1785 ();
 sg13g2_fill_2 FILLER_33_1802 ();
 sg13g2_fill_1 FILLER_33_1819 ();
 sg13g2_fill_2 FILLER_33_1824 ();
 sg13g2_fill_2 FILLER_33_1832 ();
 sg13g2_fill_2 FILLER_33_1839 ();
 sg13g2_decap_4 FILLER_33_1846 ();
 sg13g2_fill_2 FILLER_33_1850 ();
 sg13g2_fill_2 FILLER_33_1856 ();
 sg13g2_fill_2 FILLER_33_1882 ();
 sg13g2_fill_1 FILLER_33_1889 ();
 sg13g2_fill_1 FILLER_33_1895 ();
 sg13g2_decap_4 FILLER_33_1903 ();
 sg13g2_fill_1 FILLER_33_1907 ();
 sg13g2_fill_1 FILLER_33_1926 ();
 sg13g2_fill_1 FILLER_33_1932 ();
 sg13g2_decap_8 FILLER_33_1952 ();
 sg13g2_fill_1 FILLER_33_1959 ();
 sg13g2_fill_1 FILLER_33_2000 ();
 sg13g2_fill_1 FILLER_33_2037 ();
 sg13g2_decap_4 FILLER_33_2104 ();
 sg13g2_decap_8 FILLER_33_2144 ();
 sg13g2_decap_4 FILLER_33_2151 ();
 sg13g2_decap_8 FILLER_33_2168 ();
 sg13g2_fill_2 FILLER_33_2175 ();
 sg13g2_fill_1 FILLER_33_2177 ();
 sg13g2_fill_2 FILLER_33_2188 ();
 sg13g2_fill_1 FILLER_33_2190 ();
 sg13g2_decap_8 FILLER_33_2195 ();
 sg13g2_decap_8 FILLER_33_2202 ();
 sg13g2_decap_4 FILLER_33_2209 ();
 sg13g2_decap_4 FILLER_33_2243 ();
 sg13g2_fill_1 FILLER_33_2247 ();
 sg13g2_decap_4 FILLER_33_2252 ();
 sg13g2_fill_1 FILLER_33_2256 ();
 sg13g2_decap_8 FILLER_33_2261 ();
 sg13g2_decap_8 FILLER_33_2268 ();
 sg13g2_fill_2 FILLER_33_2275 ();
 sg13g2_fill_1 FILLER_33_2277 ();
 sg13g2_decap_8 FILLER_33_2282 ();
 sg13g2_decap_8 FILLER_33_2289 ();
 sg13g2_fill_1 FILLER_33_2296 ();
 sg13g2_decap_8 FILLER_33_2323 ();
 sg13g2_fill_2 FILLER_33_2330 ();
 sg13g2_decap_8 FILLER_33_2358 ();
 sg13g2_decap_4 FILLER_33_2365 ();
 sg13g2_fill_2 FILLER_33_2369 ();
 sg13g2_decap_4 FILLER_33_2381 ();
 sg13g2_fill_2 FILLER_33_2385 ();
 sg13g2_fill_2 FILLER_33_2406 ();
 sg13g2_fill_1 FILLER_33_2408 ();
 sg13g2_fill_2 FILLER_33_2421 ();
 sg13g2_decap_4 FILLER_33_2427 ();
 sg13g2_decap_8 FILLER_33_2435 ();
 sg13g2_decap_8 FILLER_33_2442 ();
 sg13g2_fill_1 FILLER_33_2449 ();
 sg13g2_fill_1 FILLER_33_2464 ();
 sg13g2_decap_8 FILLER_33_2483 ();
 sg13g2_decap_8 FILLER_33_2490 ();
 sg13g2_decap_8 FILLER_33_2497 ();
 sg13g2_fill_1 FILLER_33_2504 ();
 sg13g2_decap_8 FILLER_33_2549 ();
 sg13g2_fill_2 FILLER_33_2556 ();
 sg13g2_decap_8 FILLER_33_2636 ();
 sg13g2_decap_8 FILLER_33_2643 ();
 sg13g2_decap_8 FILLER_33_2650 ();
 sg13g2_decap_8 FILLER_33_2657 ();
 sg13g2_decap_4 FILLER_33_2664 ();
 sg13g2_fill_2 FILLER_33_2668 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_23 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_decap_4 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_139 ();
 sg13g2_fill_2 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_34_417 ();
 sg13g2_fill_1 FILLER_34_448 ();
 sg13g2_fill_1 FILLER_34_454 ();
 sg13g2_fill_1 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_495 ();
 sg13g2_fill_1 FILLER_34_511 ();
 sg13g2_fill_1 FILLER_34_521 ();
 sg13g2_fill_2 FILLER_34_532 ();
 sg13g2_fill_1 FILLER_34_537 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_decap_8 FILLER_34_709 ();
 sg13g2_decap_8 FILLER_34_716 ();
 sg13g2_decap_4 FILLER_34_723 ();
 sg13g2_fill_2 FILLER_34_727 ();
 sg13g2_decap_4 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_780 ();
 sg13g2_decap_4 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_fill_2 FILLER_34_808 ();
 sg13g2_fill_1 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_fill_2 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_fill_2 FILLER_34_848 ();
 sg13g2_fill_1 FILLER_34_850 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_fill_1 FILLER_34_945 ();
 sg13g2_fill_2 FILLER_34_986 ();
 sg13g2_fill_1 FILLER_34_992 ();
 sg13g2_fill_2 FILLER_34_1033 ();
 sg13g2_fill_1 FILLER_34_1035 ();
 sg13g2_fill_2 FILLER_34_1077 ();
 sg13g2_fill_1 FILLER_34_1092 ();
 sg13g2_decap_8 FILLER_34_1097 ();
 sg13g2_fill_1 FILLER_34_1104 ();
 sg13g2_fill_1 FILLER_34_1123 ();
 sg13g2_decap_8 FILLER_34_1145 ();
 sg13g2_fill_1 FILLER_34_1152 ();
 sg13g2_fill_1 FILLER_34_1160 ();
 sg13g2_fill_2 FILLER_34_1175 ();
 sg13g2_fill_1 FILLER_34_1181 ();
 sg13g2_fill_1 FILLER_34_1212 ();
 sg13g2_fill_2 FILLER_34_1225 ();
 sg13g2_fill_1 FILLER_34_1227 ();
 sg13g2_fill_2 FILLER_34_1251 ();
 sg13g2_decap_8 FILLER_34_1260 ();
 sg13g2_decap_8 FILLER_34_1273 ();
 sg13g2_decap_4 FILLER_34_1280 ();
 sg13g2_fill_2 FILLER_34_1320 ();
 sg13g2_fill_1 FILLER_34_1332 ();
 sg13g2_fill_1 FILLER_34_1343 ();
 sg13g2_fill_1 FILLER_34_1370 ();
 sg13g2_fill_2 FILLER_34_1397 ();
 sg13g2_fill_2 FILLER_34_1429 ();
 sg13g2_fill_1 FILLER_34_1457 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_decap_8 FILLER_34_1516 ();
 sg13g2_fill_2 FILLER_34_1523 ();
 sg13g2_fill_1 FILLER_34_1525 ();
 sg13g2_fill_1 FILLER_34_1557 ();
 sg13g2_fill_1 FILLER_34_1562 ();
 sg13g2_fill_1 FILLER_34_1589 ();
 sg13g2_fill_2 FILLER_34_1629 ();
 sg13g2_fill_2 FILLER_34_1639 ();
 sg13g2_decap_8 FILLER_34_1652 ();
 sg13g2_decap_8 FILLER_34_1659 ();
 sg13g2_fill_2 FILLER_34_1666 ();
 sg13g2_fill_1 FILLER_34_1668 ();
 sg13g2_fill_1 FILLER_34_1699 ();
 sg13g2_fill_1 FILLER_34_1703 ();
 sg13g2_decap_8 FILLER_34_1727 ();
 sg13g2_decap_8 FILLER_34_1734 ();
 sg13g2_fill_1 FILLER_34_1741 ();
 sg13g2_decap_8 FILLER_34_1747 ();
 sg13g2_fill_2 FILLER_34_1754 ();
 sg13g2_fill_1 FILLER_34_1756 ();
 sg13g2_fill_1 FILLER_34_1763 ();
 sg13g2_fill_1 FILLER_34_1769 ();
 sg13g2_fill_1 FILLER_34_1778 ();
 sg13g2_decap_8 FILLER_34_1784 ();
 sg13g2_fill_2 FILLER_34_1791 ();
 sg13g2_fill_2 FILLER_34_1803 ();
 sg13g2_fill_1 FILLER_34_1805 ();
 sg13g2_fill_1 FILLER_34_1811 ();
 sg13g2_fill_1 FILLER_34_1826 ();
 sg13g2_fill_1 FILLER_34_1832 ();
 sg13g2_fill_1 FILLER_34_1837 ();
 sg13g2_fill_1 FILLER_34_1847 ();
 sg13g2_fill_1 FILLER_34_1858 ();
 sg13g2_fill_1 FILLER_34_1864 ();
 sg13g2_fill_1 FILLER_34_1873 ();
 sg13g2_fill_1 FILLER_34_1879 ();
 sg13g2_fill_1 FILLER_34_1884 ();
 sg13g2_fill_2 FILLER_34_1895 ();
 sg13g2_fill_1 FILLER_34_1901 ();
 sg13g2_fill_2 FILLER_34_1923 ();
 sg13g2_decap_8 FILLER_34_1944 ();
 sg13g2_fill_1 FILLER_34_1951 ();
 sg13g2_decap_8 FILLER_34_1956 ();
 sg13g2_decap_8 FILLER_34_1989 ();
 sg13g2_decap_8 FILLER_34_1996 ();
 sg13g2_decap_8 FILLER_34_2003 ();
 sg13g2_decap_8 FILLER_34_2010 ();
 sg13g2_fill_1 FILLER_34_2017 ();
 sg13g2_decap_4 FILLER_34_2022 ();
 sg13g2_fill_1 FILLER_34_2064 ();
 sg13g2_fill_1 FILLER_34_2075 ();
 sg13g2_fill_2 FILLER_34_2109 ();
 sg13g2_decap_8 FILLER_34_2115 ();
 sg13g2_decap_8 FILLER_34_2130 ();
 sg13g2_decap_8 FILLER_34_2137 ();
 sg13g2_fill_2 FILLER_34_2144 ();
 sg13g2_fill_1 FILLER_34_2146 ();
 sg13g2_decap_8 FILLER_34_2173 ();
 sg13g2_fill_2 FILLER_34_2241 ();
 sg13g2_fill_1 FILLER_34_2243 ();
 sg13g2_fill_2 FILLER_34_2249 ();
 sg13g2_decap_8 FILLER_34_2277 ();
 sg13g2_decap_8 FILLER_34_2284 ();
 sg13g2_fill_2 FILLER_34_2291 ();
 sg13g2_fill_1 FILLER_34_2297 ();
 sg13g2_fill_1 FILLER_34_2324 ();
 sg13g2_fill_1 FILLER_34_2361 ();
 sg13g2_decap_8 FILLER_34_2388 ();
 sg13g2_fill_1 FILLER_34_2395 ();
 sg13g2_fill_1 FILLER_34_2399 ();
 sg13g2_fill_1 FILLER_34_2436 ();
 sg13g2_decap_8 FILLER_34_2477 ();
 sg13g2_decap_4 FILLER_34_2484 ();
 sg13g2_fill_1 FILLER_34_2488 ();
 sg13g2_decap_4 FILLER_34_2529 ();
 sg13g2_fill_2 FILLER_34_2533 ();
 sg13g2_fill_1 FILLER_34_2545 ();
 sg13g2_fill_2 FILLER_34_2566 ();
 sg13g2_fill_2 FILLER_34_2582 ();
 sg13g2_fill_2 FILLER_34_2657 ();
 sg13g2_fill_1 FILLER_34_2659 ();
 sg13g2_decap_4 FILLER_34_2664 ();
 sg13g2_fill_2 FILLER_34_2668 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_40 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_fill_2 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_decap_4 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_417 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_430 ();
 sg13g2_fill_2 FILLER_35_435 ();
 sg13g2_fill_1 FILLER_35_437 ();
 sg13g2_fill_1 FILLER_35_503 ();
 sg13g2_fill_2 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_555 ();
 sg13g2_fill_1 FILLER_35_557 ();
 sg13g2_decap_4 FILLER_35_703 ();
 sg13g2_fill_2 FILLER_35_707 ();
 sg13g2_fill_1 FILLER_35_719 ();
 sg13g2_decap_4 FILLER_35_772 ();
 sg13g2_decap_4 FILLER_35_822 ();
 sg13g2_fill_1 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_862 ();
 sg13g2_fill_2 FILLER_35_869 ();
 sg13g2_decap_4 FILLER_35_889 ();
 sg13g2_fill_1 FILLER_35_893 ();
 sg13g2_fill_1 FILLER_35_924 ();
 sg13g2_decap_4 FILLER_35_929 ();
 sg13g2_fill_2 FILLER_35_933 ();
 sg13g2_decap_4 FILLER_35_961 ();
 sg13g2_fill_1 FILLER_35_995 ();
 sg13g2_fill_2 FILLER_35_1005 ();
 sg13g2_fill_1 FILLER_35_1007 ();
 sg13g2_decap_4 FILLER_35_1012 ();
 sg13g2_decap_4 FILLER_35_1178 ();
 sg13g2_fill_2 FILLER_35_1191 ();
 sg13g2_decap_4 FILLER_35_1208 ();
 sg13g2_fill_1 FILLER_35_1244 ();
 sg13g2_fill_1 FILLER_35_1253 ();
 sg13g2_fill_2 FILLER_35_1299 ();
 sg13g2_fill_2 FILLER_35_1305 ();
 sg13g2_decap_8 FILLER_35_1311 ();
 sg13g2_fill_1 FILLER_35_1318 ();
 sg13g2_fill_2 FILLER_35_1325 ();
 sg13g2_decap_8 FILLER_35_1474 ();
 sg13g2_decap_8 FILLER_35_1481 ();
 sg13g2_decap_4 FILLER_35_1488 ();
 sg13g2_fill_1 FILLER_35_1492 ();
 sg13g2_decap_4 FILLER_35_1514 ();
 sg13g2_decap_4 FILLER_35_1522 ();
 sg13g2_decap_8 FILLER_35_1530 ();
 sg13g2_fill_1 FILLER_35_1537 ();
 sg13g2_decap_4 FILLER_35_1542 ();
 sg13g2_fill_2 FILLER_35_1576 ();
 sg13g2_decap_8 FILLER_35_1582 ();
 sg13g2_decap_8 FILLER_35_1589 ();
 sg13g2_fill_1 FILLER_35_1596 ();
 sg13g2_fill_1 FILLER_35_1631 ();
 sg13g2_decap_8 FILLER_35_1663 ();
 sg13g2_fill_2 FILLER_35_1670 ();
 sg13g2_fill_1 FILLER_35_1676 ();
 sg13g2_decap_8 FILLER_35_1735 ();
 sg13g2_decap_8 FILLER_35_1745 ();
 sg13g2_fill_2 FILLER_35_1752 ();
 sg13g2_fill_2 FILLER_35_1772 ();
 sg13g2_fill_1 FILLER_35_1843 ();
 sg13g2_fill_1 FILLER_35_1859 ();
 sg13g2_fill_1 FILLER_35_1932 ();
 sg13g2_decap_8 FILLER_35_1942 ();
 sg13g2_decap_4 FILLER_35_1949 ();
 sg13g2_fill_2 FILLER_35_1979 ();
 sg13g2_decap_4 FILLER_35_2007 ();
 sg13g2_fill_2 FILLER_35_2037 ();
 sg13g2_fill_1 FILLER_35_2049 ();
 sg13g2_fill_1 FILLER_35_2064 ();
 sg13g2_fill_1 FILLER_35_2086 ();
 sg13g2_fill_2 FILLER_35_2094 ();
 sg13g2_decap_8 FILLER_35_2101 ();
 sg13g2_decap_4 FILLER_35_2108 ();
 sg13g2_decap_4 FILLER_35_2138 ();
 sg13g2_fill_1 FILLER_35_2151 ();
 sg13g2_decap_8 FILLER_35_2178 ();
 sg13g2_fill_1 FILLER_35_2185 ();
 sg13g2_fill_2 FILLER_35_2299 ();
 sg13g2_fill_1 FILLER_35_2315 ();
 sg13g2_decap_4 FILLER_35_2326 ();
 sg13g2_fill_1 FILLER_35_2330 ();
 sg13g2_fill_2 FILLER_35_2370 ();
 sg13g2_fill_2 FILLER_35_2398 ();
 sg13g2_decap_8 FILLER_35_2426 ();
 sg13g2_fill_1 FILLER_35_2433 ();
 sg13g2_decap_4 FILLER_35_2468 ();
 sg13g2_fill_2 FILLER_35_2472 ();
 sg13g2_decap_8 FILLER_35_2562 ();
 sg13g2_fill_1 FILLER_35_2569 ();
 sg13g2_decap_8 FILLER_35_2652 ();
 sg13g2_decap_8 FILLER_35_2659 ();
 sg13g2_decap_4 FILLER_35_2666 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_17 ();
 sg13g2_fill_1 FILLER_36_19 ();
 sg13g2_fill_1 FILLER_36_27 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_decap_4 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_4 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_438 ();
 sg13g2_fill_2 FILLER_36_445 ();
 sg13g2_fill_2 FILLER_36_466 ();
 sg13g2_fill_1 FILLER_36_477 ();
 sg13g2_fill_2 FILLER_36_507 ();
 sg13g2_fill_2 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_1 FILLER_36_596 ();
 sg13g2_decap_4 FILLER_36_623 ();
 sg13g2_fill_2 FILLER_36_627 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_fill_2 FILLER_36_676 ();
 sg13g2_fill_1 FILLER_36_682 ();
 sg13g2_fill_1 FILLER_36_709 ();
 sg13g2_fill_2 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_fill_1 FILLER_36_777 ();
 sg13g2_decap_4 FILLER_36_858 ();
 sg13g2_fill_1 FILLER_36_862 ();
 sg13g2_decap_4 FILLER_36_910 ();
 sg13g2_fill_1 FILLER_36_914 ();
 sg13g2_decap_4 FILLER_36_925 ();
 sg13g2_fill_2 FILLER_36_939 ();
 sg13g2_fill_1 FILLER_36_941 ();
 sg13g2_decap_8 FILLER_36_963 ();
 sg13g2_decap_4 FILLER_36_970 ();
 sg13g2_fill_2 FILLER_36_974 ();
 sg13g2_fill_2 FILLER_36_981 ();
 sg13g2_fill_2 FILLER_36_987 ();
 sg13g2_fill_1 FILLER_36_989 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_fill_2 FILLER_36_1022 ();
 sg13g2_fill_1 FILLER_36_1038 ();
 sg13g2_fill_2 FILLER_36_1083 ();
 sg13g2_fill_1 FILLER_36_1100 ();
 sg13g2_decap_8 FILLER_36_1131 ();
 sg13g2_fill_1 FILLER_36_1138 ();
 sg13g2_fill_1 FILLER_36_1144 ();
 sg13g2_decap_8 FILLER_36_1149 ();
 sg13g2_decap_8 FILLER_36_1156 ();
 sg13g2_fill_2 FILLER_36_1163 ();
 sg13g2_decap_8 FILLER_36_1171 ();
 sg13g2_fill_2 FILLER_36_1178 ();
 sg13g2_fill_1 FILLER_36_1180 ();
 sg13g2_fill_2 FILLER_36_1193 ();
 sg13g2_decap_4 FILLER_36_1201 ();
 sg13g2_fill_1 FILLER_36_1205 ();
 sg13g2_fill_2 FILLER_36_1211 ();
 sg13g2_fill_1 FILLER_36_1213 ();
 sg13g2_fill_1 FILLER_36_1246 ();
 sg13g2_fill_1 FILLER_36_1268 ();
 sg13g2_fill_1 FILLER_36_1322 ();
 sg13g2_fill_2 FILLER_36_1328 ();
 sg13g2_fill_1 FILLER_36_1356 ();
 sg13g2_fill_2 FILLER_36_1361 ();
 sg13g2_fill_2 FILLER_36_1386 ();
 sg13g2_fill_1 FILLER_36_1398 ();
 sg13g2_fill_2 FILLER_36_1438 ();
 sg13g2_decap_4 FILLER_36_1458 ();
 sg13g2_fill_2 FILLER_36_1462 ();
 sg13g2_decap_8 FILLER_36_1490 ();
 sg13g2_decap_8 FILLER_36_1497 ();
 sg13g2_decap_8 FILLER_36_1504 ();
 sg13g2_decap_8 FILLER_36_1511 ();
 sg13g2_fill_1 FILLER_36_1518 ();
 sg13g2_decap_8 FILLER_36_1558 ();
 sg13g2_fill_2 FILLER_36_1565 ();
 sg13g2_fill_1 FILLER_36_1597 ();
 sg13g2_fill_2 FILLER_36_1608 ();
 sg13g2_fill_1 FILLER_36_1610 ();
 sg13g2_fill_1 FILLER_36_1615 ();
 sg13g2_fill_2 FILLER_36_1621 ();
 sg13g2_fill_2 FILLER_36_1672 ();
 sg13g2_fill_1 FILLER_36_1674 ();
 sg13g2_fill_2 FILLER_36_1709 ();
 sg13g2_fill_1 FILLER_36_1737 ();
 sg13g2_fill_1 FILLER_36_1749 ();
 sg13g2_fill_2 FILLER_36_1755 ();
 sg13g2_fill_1 FILLER_36_1762 ();
 sg13g2_fill_1 FILLER_36_1774 ();
 sg13g2_fill_1 FILLER_36_1795 ();
 sg13g2_fill_1 FILLER_36_1801 ();
 sg13g2_fill_1 FILLER_36_1807 ();
 sg13g2_fill_2 FILLER_36_1828 ();
 sg13g2_fill_1 FILLER_36_1871 ();
 sg13g2_fill_2 FILLER_36_1893 ();
 sg13g2_fill_1 FILLER_36_1917 ();
 sg13g2_fill_2 FILLER_36_1946 ();
 sg13g2_fill_1 FILLER_36_1948 ();
 sg13g2_fill_2 FILLER_36_1958 ();
 sg13g2_fill_1 FILLER_36_1978 ();
 sg13g2_fill_2 FILLER_36_2019 ();
 sg13g2_fill_2 FILLER_36_2093 ();
 sg13g2_fill_2 FILLER_36_2126 ();
 sg13g2_fill_1 FILLER_36_2128 ();
 sg13g2_decap_4 FILLER_36_2133 ();
 sg13g2_fill_2 FILLER_36_2142 ();
 sg13g2_fill_1 FILLER_36_2148 ();
 sg13g2_fill_1 FILLER_36_2154 ();
 sg13g2_fill_1 FILLER_36_2159 ();
 sg13g2_fill_1 FILLER_36_2165 ();
 sg13g2_fill_1 FILLER_36_2232 ();
 sg13g2_decap_4 FILLER_36_2278 ();
 sg13g2_fill_2 FILLER_36_2348 ();
 sg13g2_decap_4 FILLER_36_2360 ();
 sg13g2_fill_1 FILLER_36_2364 ();
 sg13g2_decap_8 FILLER_36_2387 ();
 sg13g2_decap_4 FILLER_36_2394 ();
 sg13g2_fill_1 FILLER_36_2398 ();
 sg13g2_fill_2 FILLER_36_2412 ();
 sg13g2_fill_1 FILLER_36_2414 ();
 sg13g2_decap_4 FILLER_36_2425 ();
 sg13g2_fill_1 FILLER_36_2429 ();
 sg13g2_decap_8 FILLER_36_2466 ();
 sg13g2_fill_2 FILLER_36_2473 ();
 sg13g2_fill_1 FILLER_36_2475 ();
 sg13g2_fill_2 FILLER_36_2526 ();
 sg13g2_fill_1 FILLER_36_2528 ();
 sg13g2_decap_4 FILLER_36_2539 ();
 sg13g2_fill_1 FILLER_36_2557 ();
 sg13g2_fill_1 FILLER_36_2576 ();
 sg13g2_decap_4 FILLER_36_2587 ();
 sg13g2_fill_1 FILLER_36_2591 ();
 sg13g2_fill_2 FILLER_36_2597 ();
 sg13g2_fill_2 FILLER_36_2656 ();
 sg13g2_fill_1 FILLER_36_2658 ();
 sg13g2_decap_8 FILLER_36_2663 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_fill_1 FILLER_37_47 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_fill_2 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_430 ();
 sg13g2_fill_1 FILLER_37_432 ();
 sg13g2_decap_8 FILLER_37_438 ();
 sg13g2_decap_4 FILLER_37_445 ();
 sg13g2_fill_1 FILLER_37_449 ();
 sg13g2_fill_2 FILLER_37_469 ();
 sg13g2_fill_1 FILLER_37_494 ();
 sg13g2_fill_1 FILLER_37_513 ();
 sg13g2_fill_1 FILLER_37_519 ();
 sg13g2_fill_2 FILLER_37_530 ();
 sg13g2_decap_4 FILLER_37_562 ();
 sg13g2_decap_4 FILLER_37_574 ();
 sg13g2_fill_2 FILLER_37_578 ();
 sg13g2_fill_1 FILLER_37_600 ();
 sg13g2_fill_2 FILLER_37_605 ();
 sg13g2_fill_2 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_4 FILLER_37_657 ();
 sg13g2_fill_2 FILLER_37_691 ();
 sg13g2_fill_1 FILLER_37_703 ();
 sg13g2_fill_2 FILLER_37_751 ();
 sg13g2_fill_1 FILLER_37_773 ();
 sg13g2_fill_1 FILLER_37_785 ();
 sg13g2_fill_1 FILLER_37_820 ();
 sg13g2_fill_2 FILLER_37_852 ();
 sg13g2_fill_1 FILLER_37_854 ();
 sg13g2_decap_4 FILLER_37_895 ();
 sg13g2_fill_1 FILLER_37_899 ();
 sg13g2_fill_1 FILLER_37_921 ();
 sg13g2_decap_8 FILLER_37_956 ();
 sg13g2_decap_4 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_1002 ();
 sg13g2_fill_2 FILLER_37_1074 ();
 sg13g2_decap_4 FILLER_37_1081 ();
 sg13g2_fill_1 FILLER_37_1095 ();
 sg13g2_decap_4 FILLER_37_1100 ();
 sg13g2_fill_1 FILLER_37_1104 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_fill_2 FILLER_37_1120 ();
 sg13g2_fill_1 FILLER_37_1122 ();
 sg13g2_decap_4 FILLER_37_1133 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_decap_8 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1165 ();
 sg13g2_fill_1 FILLER_37_1177 ();
 sg13g2_fill_1 FILLER_37_1183 ();
 sg13g2_fill_1 FILLER_37_1196 ();
 sg13g2_decap_4 FILLER_37_1222 ();
 sg13g2_decap_4 FILLER_37_1231 ();
 sg13g2_fill_2 FILLER_37_1239 ();
 sg13g2_fill_1 FILLER_37_1241 ();
 sg13g2_fill_2 FILLER_37_1278 ();
 sg13g2_fill_2 FILLER_37_1285 ();
 sg13g2_fill_1 FILLER_37_1333 ();
 sg13g2_fill_2 FILLER_37_1344 ();
 sg13g2_fill_1 FILLER_37_1346 ();
 sg13g2_fill_2 FILLER_37_1381 ();
 sg13g2_fill_1 FILLER_37_1442 ();
 sg13g2_decap_4 FILLER_37_1450 ();
 sg13g2_fill_2 FILLER_37_1454 ();
 sg13g2_decap_8 FILLER_37_1459 ();
 sg13g2_decap_4 FILLER_37_1466 ();
 sg13g2_fill_2 FILLER_37_1470 ();
 sg13g2_decap_4 FILLER_37_1503 ();
 sg13g2_fill_2 FILLER_37_1529 ();
 sg13g2_fill_1 FILLER_37_1531 ();
 sg13g2_fill_1 FILLER_37_1558 ();
 sg13g2_decap_8 FILLER_37_1563 ();
 sg13g2_decap_8 FILLER_37_1570 ();
 sg13g2_decap_8 FILLER_37_1577 ();
 sg13g2_fill_2 FILLER_37_1610 ();
 sg13g2_fill_1 FILLER_37_1679 ();
 sg13g2_fill_1 FILLER_37_1709 ();
 sg13g2_fill_2 FILLER_37_1744 ();
 sg13g2_decap_4 FILLER_37_1801 ();
 sg13g2_fill_1 FILLER_37_1818 ();
 sg13g2_fill_1 FILLER_37_1827 ();
 sg13g2_fill_1 FILLER_37_1853 ();
 sg13g2_fill_2 FILLER_37_1877 ();
 sg13g2_fill_1 FILLER_37_1889 ();
 sg13g2_fill_1 FILLER_37_1930 ();
 sg13g2_decap_8 FILLER_37_1959 ();
 sg13g2_decap_4 FILLER_37_1966 ();
 sg13g2_fill_1 FILLER_37_1970 ();
 sg13g2_fill_1 FILLER_37_1984 ();
 sg13g2_fill_1 FILLER_37_1989 ();
 sg13g2_decap_8 FILLER_37_1994 ();
 sg13g2_decap_4 FILLER_37_2001 ();
 sg13g2_fill_1 FILLER_37_2005 ();
 sg13g2_decap_8 FILLER_37_2019 ();
 sg13g2_decap_8 FILLER_37_2026 ();
 sg13g2_decap_4 FILLER_37_2033 ();
 sg13g2_fill_2 FILLER_37_2037 ();
 sg13g2_decap_8 FILLER_37_2043 ();
 sg13g2_fill_1 FILLER_37_2055 ();
 sg13g2_decap_4 FILLER_37_2086 ();
 sg13g2_fill_1 FILLER_37_2100 ();
 sg13g2_fill_2 FILLER_37_2166 ();
 sg13g2_fill_2 FILLER_37_2177 ();
 sg13g2_fill_1 FILLER_37_2203 ();
 sg13g2_fill_2 FILLER_37_2213 ();
 sg13g2_fill_2 FILLER_37_2226 ();
 sg13g2_fill_2 FILLER_37_2242 ();
 sg13g2_fill_1 FILLER_37_2244 ();
 sg13g2_fill_2 FILLER_37_2267 ();
 sg13g2_fill_2 FILLER_37_2275 ();
 sg13g2_decap_8 FILLER_37_2283 ();
 sg13g2_decap_4 FILLER_37_2290 ();
 sg13g2_fill_1 FILLER_37_2298 ();
 sg13g2_fill_2 FILLER_37_2309 ();
 sg13g2_fill_2 FILLER_37_2316 ();
 sg13g2_fill_1 FILLER_37_2337 ();
 sg13g2_fill_1 FILLER_37_2342 ();
 sg13g2_decap_8 FILLER_37_2385 ();
 sg13g2_fill_2 FILLER_37_2392 ();
 sg13g2_fill_1 FILLER_37_2406 ();
 sg13g2_fill_2 FILLER_37_2411 ();
 sg13g2_fill_1 FILLER_37_2425 ();
 sg13g2_fill_2 FILLER_37_2446 ();
 sg13g2_fill_2 FILLER_37_2452 ();
 sg13g2_fill_1 FILLER_37_2454 ();
 sg13g2_decap_4 FILLER_37_2477 ();
 sg13g2_fill_2 FILLER_37_2481 ();
 sg13g2_fill_2 FILLER_37_2487 ();
 sg13g2_fill_1 FILLER_37_2489 ();
 sg13g2_fill_2 FILLER_37_2520 ();
 sg13g2_decap_8 FILLER_37_2531 ();
 sg13g2_decap_4 FILLER_37_2538 ();
 sg13g2_fill_1 FILLER_37_2542 ();
 sg13g2_fill_1 FILLER_37_2561 ();
 sg13g2_fill_1 FILLER_37_2573 ();
 sg13g2_decap_8 FILLER_37_2584 ();
 sg13g2_fill_1 FILLER_37_2591 ();
 sg13g2_fill_1 FILLER_37_2618 ();
 sg13g2_fill_1 FILLER_37_2629 ();
 sg13g2_decap_8 FILLER_37_2660 ();
 sg13g2_fill_2 FILLER_37_2667 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_decap_4 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_decap_8 FILLER_38_95 ();
 sg13g2_decap_4 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_178 ();
 sg13g2_decap_4 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_4 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_341 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_415 ();
 sg13g2_fill_1 FILLER_38_465 ();
 sg13g2_fill_1 FILLER_38_469 ();
 sg13g2_fill_1 FILLER_38_475 ();
 sg13g2_fill_1 FILLER_38_482 ();
 sg13g2_fill_1 FILLER_38_488 ();
 sg13g2_fill_2 FILLER_38_513 ();
 sg13g2_fill_1 FILLER_38_520 ();
 sg13g2_fill_1 FILLER_38_526 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_fill_2 FILLER_38_545 ();
 sg13g2_decap_4 FILLER_38_552 ();
 sg13g2_fill_2 FILLER_38_556 ();
 sg13g2_fill_1 FILLER_38_605 ();
 sg13g2_decap_4 FILLER_38_706 ();
 sg13g2_fill_1 FILLER_38_710 ();
 sg13g2_decap_4 FILLER_38_746 ();
 sg13g2_fill_2 FILLER_38_774 ();
 sg13g2_fill_1 FILLER_38_805 ();
 sg13g2_decap_4 FILLER_38_827 ();
 sg13g2_fill_2 FILLER_38_867 ();
 sg13g2_fill_1 FILLER_38_869 ();
 sg13g2_fill_2 FILLER_38_917 ();
 sg13g2_fill_2 FILLER_38_967 ();
 sg13g2_fill_1 FILLER_38_973 ();
 sg13g2_fill_1 FILLER_38_1026 ();
 sg13g2_fill_2 FILLER_38_1050 ();
 sg13g2_fill_1 FILLER_38_1084 ();
 sg13g2_fill_1 FILLER_38_1111 ();
 sg13g2_fill_2 FILLER_38_1122 ();
 sg13g2_fill_2 FILLER_38_1128 ();
 sg13g2_decap_4 FILLER_38_1156 ();
 sg13g2_fill_1 FILLER_38_1189 ();
 sg13g2_fill_2 FILLER_38_1209 ();
 sg13g2_fill_1 FILLER_38_1247 ();
 sg13g2_fill_1 FILLER_38_1252 ();
 sg13g2_fill_1 FILLER_38_1265 ();
 sg13g2_fill_2 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_fill_2 FILLER_38_1297 ();
 sg13g2_fill_2 FILLER_38_1339 ();
 sg13g2_fill_1 FILLER_38_1354 ();
 sg13g2_fill_1 FILLER_38_1365 ();
 sg13g2_fill_1 FILLER_38_1409 ();
 sg13g2_fill_1 FILLER_38_1441 ();
 sg13g2_decap_4 FILLER_38_1455 ();
 sg13g2_decap_8 FILLER_38_1464 ();
 sg13g2_decap_4 FILLER_38_1471 ();
 sg13g2_fill_1 FILLER_38_1475 ();
 sg13g2_decap_4 FILLER_38_1481 ();
 sg13g2_fill_1 FILLER_38_1509 ();
 sg13g2_fill_1 FILLER_38_1524 ();
 sg13g2_fill_1 FILLER_38_1533 ();
 sg13g2_fill_2 FILLER_38_1544 ();
 sg13g2_fill_2 FILLER_38_1590 ();
 sg13g2_fill_1 FILLER_38_1592 ();
 sg13g2_decap_4 FILLER_38_1601 ();
 sg13g2_fill_2 FILLER_38_1666 ();
 sg13g2_fill_2 FILLER_38_1694 ();
 sg13g2_decap_4 FILLER_38_1700 ();
 sg13g2_decap_4 FILLER_38_1710 ();
 sg13g2_fill_2 FILLER_38_1718 ();
 sg13g2_fill_1 FILLER_38_1720 ();
 sg13g2_decap_8 FILLER_38_1725 ();
 sg13g2_fill_2 FILLER_38_1732 ();
 sg13g2_fill_1 FILLER_38_1734 ();
 sg13g2_fill_1 FILLER_38_1741 ();
 sg13g2_fill_1 FILLER_38_1752 ();
 sg13g2_fill_2 FILLER_38_1763 ();
 sg13g2_fill_1 FILLER_38_1770 ();
 sg13g2_fill_2 FILLER_38_1776 ();
 sg13g2_fill_2 FILLER_38_1792 ();
 sg13g2_fill_1 FILLER_38_1803 ();
 sg13g2_fill_1 FILLER_38_1885 ();
 sg13g2_fill_1 FILLER_38_1914 ();
 sg13g2_fill_2 FILLER_38_1929 ();
 sg13g2_fill_1 FILLER_38_1931 ();
 sg13g2_fill_1 FILLER_38_1982 ();
 sg13g2_fill_2 FILLER_38_1999 ();
 sg13g2_decap_8 FILLER_38_2008 ();
 sg13g2_decap_8 FILLER_38_2015 ();
 sg13g2_decap_8 FILLER_38_2022 ();
 sg13g2_decap_8 FILLER_38_2029 ();
 sg13g2_decap_8 FILLER_38_2036 ();
 sg13g2_decap_4 FILLER_38_2043 ();
 sg13g2_fill_1 FILLER_38_2047 ();
 sg13g2_decap_4 FILLER_38_2053 ();
 sg13g2_fill_2 FILLER_38_2057 ();
 sg13g2_fill_1 FILLER_38_2068 ();
 sg13g2_fill_2 FILLER_38_2147 ();
 sg13g2_fill_1 FILLER_38_2163 ();
 sg13g2_fill_1 FILLER_38_2170 ();
 sg13g2_fill_1 FILLER_38_2179 ();
 sg13g2_fill_1 FILLER_38_2207 ();
 sg13g2_fill_2 FILLER_38_2218 ();
 sg13g2_decap_4 FILLER_38_2248 ();
 sg13g2_fill_2 FILLER_38_2252 ();
 sg13g2_decap_4 FILLER_38_2263 ();
 sg13g2_fill_1 FILLER_38_2267 ();
 sg13g2_decap_4 FILLER_38_2278 ();
 sg13g2_fill_2 FILLER_38_2282 ();
 sg13g2_fill_1 FILLER_38_2310 ();
 sg13g2_fill_2 FILLER_38_2317 ();
 sg13g2_fill_1 FILLER_38_2329 ();
 sg13g2_fill_1 FILLER_38_2391 ();
 sg13g2_fill_2 FILLER_38_2460 ();
 sg13g2_fill_1 FILLER_38_2462 ();
 sg13g2_decap_8 FILLER_38_2473 ();
 sg13g2_decap_8 FILLER_38_2480 ();
 sg13g2_fill_1 FILLER_38_2487 ();
 sg13g2_fill_1 FILLER_38_2498 ();
 sg13g2_fill_2 FILLER_38_2561 ();
 sg13g2_fill_2 FILLER_38_2583 ();
 sg13g2_fill_1 FILLER_38_2585 ();
 sg13g2_decap_4 FILLER_38_2596 ();
 sg13g2_fill_1 FILLER_38_2600 ();
 sg13g2_decap_8 FILLER_38_2605 ();
 sg13g2_fill_2 FILLER_38_2612 ();
 sg13g2_fill_2 FILLER_38_2624 ();
 sg13g2_decap_8 FILLER_38_2656 ();
 sg13g2_decap_8 FILLER_38_2663 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_fill_2 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_39 ();
 sg13g2_fill_1 FILLER_39_62 ();
 sg13g2_fill_2 FILLER_39_90 ();
 sg13g2_decap_4 FILLER_39_128 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_152 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_decap_4 FILLER_39_172 ();
 sg13g2_fill_2 FILLER_39_176 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_210 ();
 sg13g2_decap_4 FILLER_39_229 ();
 sg13g2_decap_4 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_271 ();
 sg13g2_decap_4 FILLER_39_277 ();
 sg13g2_fill_2 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_4 FILLER_39_301 ();
 sg13g2_fill_2 FILLER_39_430 ();
 sg13g2_fill_1 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_443 ();
 sg13g2_fill_1 FILLER_39_445 ();
 sg13g2_fill_2 FILLER_39_450 ();
 sg13g2_fill_1 FILLER_39_452 ();
 sg13g2_fill_2 FILLER_39_458 ();
 sg13g2_fill_1 FILLER_39_460 ();
 sg13g2_fill_2 FILLER_39_476 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_fill_2 FILLER_39_495 ();
 sg13g2_fill_1 FILLER_39_579 ();
 sg13g2_fill_2 FILLER_39_583 ();
 sg13g2_decap_4 FILLER_39_592 ();
 sg13g2_fill_2 FILLER_39_654 ();
 sg13g2_fill_1 FILLER_39_656 ();
 sg13g2_decap_4 FILLER_39_661 ();
 sg13g2_fill_1 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_748 ();
 sg13g2_fill_1 FILLER_39_753 ();
 sg13g2_fill_2 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_877 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_fill_2 FILLER_39_896 ();
 sg13g2_fill_1 FILLER_39_898 ();
 sg13g2_fill_2 FILLER_39_935 ();
 sg13g2_fill_1 FILLER_39_951 ();
 sg13g2_decap_4 FILLER_39_978 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_fill_1 FILLER_39_1023 ();
 sg13g2_fill_1 FILLER_39_1054 ();
 sg13g2_fill_1 FILLER_39_1065 ();
 sg13g2_fill_1 FILLER_39_1092 ();
 sg13g2_fill_1 FILLER_39_1103 ();
 sg13g2_fill_1 FILLER_39_1114 ();
 sg13g2_fill_2 FILLER_39_1160 ();
 sg13g2_fill_2 FILLER_39_1221 ();
 sg13g2_fill_2 FILLER_39_1283 ();
 sg13g2_fill_1 FILLER_39_1290 ();
 sg13g2_fill_1 FILLER_39_1296 ();
 sg13g2_fill_1 FILLER_39_1314 ();
 sg13g2_fill_2 FILLER_39_1322 ();
 sg13g2_fill_2 FILLER_39_1358 ();
 sg13g2_fill_2 FILLER_39_1365 ();
 sg13g2_fill_1 FILLER_39_1371 ();
 sg13g2_fill_2 FILLER_39_1414 ();
 sg13g2_fill_2 FILLER_39_1424 ();
 sg13g2_fill_2 FILLER_39_1446 ();
 sg13g2_fill_1 FILLER_39_1448 ();
 sg13g2_fill_2 FILLER_39_1512 ();
 sg13g2_fill_2 FILLER_39_1524 ();
 sg13g2_fill_1 FILLER_39_1526 ();
 sg13g2_decap_4 FILLER_39_1574 ();
 sg13g2_fill_2 FILLER_39_1608 ();
 sg13g2_decap_4 FILLER_39_1614 ();
 sg13g2_fill_2 FILLER_39_1618 ();
 sg13g2_fill_1 FILLER_39_1660 ();
 sg13g2_decap_8 FILLER_39_1666 ();
 sg13g2_decap_4 FILLER_39_1691 ();
 sg13g2_fill_2 FILLER_39_1695 ();
 sg13g2_fill_2 FILLER_39_1706 ();
 sg13g2_decap_8 FILLER_39_1734 ();
 sg13g2_decap_8 FILLER_39_1741 ();
 sg13g2_decap_8 FILLER_39_1748 ();
 sg13g2_decap_4 FILLER_39_1755 ();
 sg13g2_fill_1 FILLER_39_1759 ();
 sg13g2_fill_2 FILLER_39_1766 ();
 sg13g2_fill_2 FILLER_39_1772 ();
 sg13g2_fill_1 FILLER_39_1774 ();
 sg13g2_decap_4 FILLER_39_1780 ();
 sg13g2_decap_4 FILLER_39_1788 ();
 sg13g2_decap_4 FILLER_39_1797 ();
 sg13g2_fill_1 FILLER_39_1801 ();
 sg13g2_fill_1 FILLER_39_1810 ();
 sg13g2_fill_1 FILLER_39_1820 ();
 sg13g2_fill_1 FILLER_39_1825 ();
 sg13g2_fill_1 FILLER_39_1831 ();
 sg13g2_fill_1 FILLER_39_1837 ();
 sg13g2_decap_4 FILLER_39_1847 ();
 sg13g2_fill_1 FILLER_39_1914 ();
 sg13g2_fill_2 FILLER_39_1929 ();
 sg13g2_fill_2 FILLER_39_1936 ();
 sg13g2_fill_1 FILLER_39_1947 ();
 sg13g2_decap_8 FILLER_39_1965 ();
 sg13g2_fill_2 FILLER_39_1975 ();
 sg13g2_fill_2 FILLER_39_1986 ();
 sg13g2_decap_8 FILLER_39_1996 ();
 sg13g2_decap_8 FILLER_39_2003 ();
 sg13g2_fill_2 FILLER_39_2010 ();
 sg13g2_fill_1 FILLER_39_2012 ();
 sg13g2_decap_8 FILLER_39_2022 ();
 sg13g2_decap_4 FILLER_39_2029 ();
 sg13g2_decap_4 FILLER_39_2037 ();
 sg13g2_fill_1 FILLER_39_2041 ();
 sg13g2_decap_4 FILLER_39_2086 ();
 sg13g2_fill_2 FILLER_39_2094 ();
 sg13g2_fill_1 FILLER_39_2096 ();
 sg13g2_fill_2 FILLER_39_2153 ();
 sg13g2_fill_2 FILLER_39_2159 ();
 sg13g2_decap_4 FILLER_39_2256 ();
 sg13g2_fill_2 FILLER_39_2309 ();
 sg13g2_fill_2 FILLER_39_2331 ();
 sg13g2_fill_1 FILLER_39_2333 ();
 sg13g2_fill_2 FILLER_39_2346 ();
 sg13g2_fill_1 FILLER_39_2355 ();
 sg13g2_fill_1 FILLER_39_2361 ();
 sg13g2_fill_1 FILLER_39_2377 ();
 sg13g2_fill_1 FILLER_39_2415 ();
 sg13g2_fill_1 FILLER_39_2461 ();
 sg13g2_decap_4 FILLER_39_2469 ();
 sg13g2_fill_2 FILLER_39_2485 ();
 sg13g2_fill_1 FILLER_39_2487 ();
 sg13g2_fill_2 FILLER_39_2536 ();
 sg13g2_fill_1 FILLER_39_2538 ();
 sg13g2_fill_2 FILLER_39_2576 ();
 sg13g2_fill_2 FILLER_39_2609 ();
 sg13g2_fill_2 FILLER_39_2621 ();
 sg13g2_decap_8 FILLER_39_2649 ();
 sg13g2_decap_8 FILLER_39_2656 ();
 sg13g2_decap_8 FILLER_39_2663 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_11 ();
 sg13g2_fill_2 FILLER_40_22 ();
 sg13g2_fill_1 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_51 ();
 sg13g2_fill_2 FILLER_40_60 ();
 sg13g2_fill_1 FILLER_40_115 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_decap_4 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_168 ();
 sg13g2_decap_4 FILLER_40_182 ();
 sg13g2_fill_1 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_212 ();
 sg13g2_decap_4 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_335 ();
 sg13g2_decap_4 FILLER_40_342 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_4 FILLER_40_364 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_decap_4 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_decap_4 FILLER_40_449 ();
 sg13g2_fill_1 FILLER_40_453 ();
 sg13g2_fill_2 FILLER_40_515 ();
 sg13g2_fill_1 FILLER_40_544 ();
 sg13g2_fill_2 FILLER_40_555 ();
 sg13g2_fill_2 FILLER_40_587 ();
 sg13g2_fill_1 FILLER_40_647 ();
 sg13g2_fill_1 FILLER_40_652 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_fill_1 FILLER_40_672 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_fill_1 FILLER_40_689 ();
 sg13g2_fill_1 FILLER_40_786 ();
 sg13g2_fill_1 FILLER_40_790 ();
 sg13g2_fill_2 FILLER_40_827 ();
 sg13g2_decap_8 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_846 ();
 sg13g2_decap_4 FILLER_40_860 ();
 sg13g2_fill_2 FILLER_40_864 ();
 sg13g2_decap_4 FILLER_40_870 ();
 sg13g2_fill_1 FILLER_40_874 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_4 FILLER_40_894 ();
 sg13g2_fill_1 FILLER_40_898 ();
 sg13g2_fill_1 FILLER_40_913 ();
 sg13g2_decap_8 FILLER_40_940 ();
 sg13g2_fill_2 FILLER_40_947 ();
 sg13g2_decap_8 FILLER_40_988 ();
 sg13g2_fill_1 FILLER_40_995 ();
 sg13g2_decap_8 FILLER_40_1004 ();
 sg13g2_fill_2 FILLER_40_1011 ();
 sg13g2_fill_1 FILLER_40_1013 ();
 sg13g2_fill_2 FILLER_40_1024 ();
 sg13g2_fill_1 FILLER_40_1040 ();
 sg13g2_decap_4 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1117 ();
 sg13g2_fill_1 FILLER_40_1137 ();
 sg13g2_fill_2 FILLER_40_1142 ();
 sg13g2_fill_2 FILLER_40_1174 ();
 sg13g2_fill_2 FILLER_40_1183 ();
 sg13g2_fill_1 FILLER_40_1198 ();
 sg13g2_fill_1 FILLER_40_1209 ();
 sg13g2_fill_2 FILLER_40_1234 ();
 sg13g2_fill_1 FILLER_40_1261 ();
 sg13g2_fill_2 FILLER_40_1300 ();
 sg13g2_fill_1 FILLER_40_1363 ();
 sg13g2_fill_2 FILLER_40_1396 ();
 sg13g2_fill_2 FILLER_40_1403 ();
 sg13g2_fill_2 FILLER_40_1435 ();
 sg13g2_fill_2 FILLER_40_1481 ();
 sg13g2_fill_2 FILLER_40_1496 ();
 sg13g2_decap_8 FILLER_40_1507 ();
 sg13g2_fill_1 FILLER_40_1514 ();
 sg13g2_fill_2 FILLER_40_1559 ();
 sg13g2_fill_2 FILLER_40_1569 ();
 sg13g2_decap_4 FILLER_40_1589 ();
 sg13g2_fill_2 FILLER_40_1593 ();
 sg13g2_fill_2 FILLER_40_1600 ();
 sg13g2_fill_1 FILLER_40_1602 ();
 sg13g2_fill_1 FILLER_40_1636 ();
 sg13g2_fill_2 FILLER_40_1641 ();
 sg13g2_fill_1 FILLER_40_1643 ();
 sg13g2_fill_2 FILLER_40_1649 ();
 sg13g2_fill_1 FILLER_40_1651 ();
 sg13g2_decap_8 FILLER_40_1656 ();
 sg13g2_decap_8 FILLER_40_1663 ();
 sg13g2_decap_8 FILLER_40_1670 ();
 sg13g2_fill_2 FILLER_40_1677 ();
 sg13g2_fill_2 FILLER_40_1683 ();
 sg13g2_fill_1 FILLER_40_1685 ();
 sg13g2_fill_1 FILLER_40_1691 ();
 sg13g2_fill_1 FILLER_40_1704 ();
 sg13g2_fill_1 FILLER_40_1710 ();
 sg13g2_decap_8 FILLER_40_1716 ();
 sg13g2_fill_2 FILLER_40_1723 ();
 sg13g2_fill_1 FILLER_40_1725 ();
 sg13g2_decap_8 FILLER_40_1756 ();
 sg13g2_decap_8 FILLER_40_1763 ();
 sg13g2_decap_8 FILLER_40_1770 ();
 sg13g2_fill_2 FILLER_40_1777 ();
 sg13g2_fill_2 FILLER_40_1784 ();
 sg13g2_fill_1 FILLER_40_1786 ();
 sg13g2_decap_4 FILLER_40_1798 ();
 sg13g2_fill_1 FILLER_40_1806 ();
 sg13g2_fill_1 FILLER_40_1811 ();
 sg13g2_fill_1 FILLER_40_1817 ();
 sg13g2_fill_2 FILLER_40_1825 ();
 sg13g2_fill_2 FILLER_40_1854 ();
 sg13g2_fill_1 FILLER_40_1856 ();
 sg13g2_fill_1 FILLER_40_1867 ();
 sg13g2_fill_1 FILLER_40_1874 ();
 sg13g2_fill_2 FILLER_40_1911 ();
 sg13g2_decap_4 FILLER_40_1917 ();
 sg13g2_fill_1 FILLER_40_1921 ();
 sg13g2_decap_8 FILLER_40_1930 ();
 sg13g2_decap_8 FILLER_40_1937 ();
 sg13g2_decap_4 FILLER_40_1944 ();
 sg13g2_decap_8 FILLER_40_1954 ();
 sg13g2_decap_8 FILLER_40_1965 ();
 sg13g2_fill_2 FILLER_40_1972 ();
 sg13g2_decap_8 FILLER_40_1993 ();
 sg13g2_decap_8 FILLER_40_2000 ();
 sg13g2_decap_8 FILLER_40_2007 ();
 sg13g2_decap_8 FILLER_40_2014 ();
 sg13g2_decap_8 FILLER_40_2021 ();
 sg13g2_decap_8 FILLER_40_2028 ();
 sg13g2_decap_8 FILLER_40_2035 ();
 sg13g2_fill_2 FILLER_40_2042 ();
 sg13g2_fill_1 FILLER_40_2044 ();
 sg13g2_decap_4 FILLER_40_2080 ();
 sg13g2_fill_1 FILLER_40_2084 ();
 sg13g2_decap_8 FILLER_40_2095 ();
 sg13g2_decap_8 FILLER_40_2102 ();
 sg13g2_fill_2 FILLER_40_2109 ();
 sg13g2_fill_1 FILLER_40_2111 ();
 sg13g2_fill_1 FILLER_40_2116 ();
 sg13g2_fill_1 FILLER_40_2121 ();
 sg13g2_fill_2 FILLER_40_2134 ();
 sg13g2_fill_1 FILLER_40_2136 ();
 sg13g2_fill_2 FILLER_40_2142 ();
 sg13g2_fill_1 FILLER_40_2175 ();
 sg13g2_fill_1 FILLER_40_2180 ();
 sg13g2_fill_1 FILLER_40_2191 ();
 sg13g2_fill_1 FILLER_40_2201 ();
 sg13g2_fill_1 FILLER_40_2211 ();
 sg13g2_fill_1 FILLER_40_2217 ();
 sg13g2_decap_8 FILLER_40_2275 ();
 sg13g2_decap_8 FILLER_40_2282 ();
 sg13g2_fill_2 FILLER_40_2289 ();
 sg13g2_fill_1 FILLER_40_2291 ();
 sg13g2_fill_1 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2301 ();
 sg13g2_fill_2 FILLER_40_2317 ();
 sg13g2_fill_2 FILLER_40_2325 ();
 sg13g2_fill_1 FILLER_40_2327 ();
 sg13g2_fill_2 FILLER_40_2334 ();
 sg13g2_fill_1 FILLER_40_2336 ();
 sg13g2_fill_2 FILLER_40_2342 ();
 sg13g2_decap_8 FILLER_40_2349 ();
 sg13g2_fill_2 FILLER_40_2356 ();
 sg13g2_fill_2 FILLER_40_2387 ();
 sg13g2_decap_4 FILLER_40_2419 ();
 sg13g2_fill_2 FILLER_40_2423 ();
 sg13g2_fill_2 FILLER_40_2456 ();
 sg13g2_fill_2 FILLER_40_2464 ();
 sg13g2_fill_2 FILLER_40_2492 ();
 sg13g2_fill_1 FILLER_40_2494 ();
 sg13g2_fill_2 FILLER_40_2521 ();
 sg13g2_decap_8 FILLER_40_2532 ();
 sg13g2_decap_4 FILLER_40_2539 ();
 sg13g2_fill_1 FILLER_40_2552 ();
 sg13g2_fill_1 FILLER_40_2579 ();
 sg13g2_decap_4 FILLER_40_2590 ();
 sg13g2_fill_2 FILLER_40_2609 ();
 sg13g2_fill_1 FILLER_40_2611 ();
 sg13g2_fill_1 FILLER_40_2622 ();
 sg13g2_decap_8 FILLER_40_2649 ();
 sg13g2_decap_8 FILLER_40_2656 ();
 sg13g2_decap_8 FILLER_40_2663 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_38 ();
 sg13g2_fill_1 FILLER_41_47 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_125 ();
 sg13g2_decap_8 FILLER_41_132 ();
 sg13g2_decap_8 FILLER_41_139 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_decap_8 FILLER_41_158 ();
 sg13g2_decap_4 FILLER_41_165 ();
 sg13g2_fill_1 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_decap_4 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_202 ();
 sg13g2_decap_4 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_229 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_8 FILLER_41_255 ();
 sg13g2_decap_4 FILLER_41_262 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_288 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_fill_1 FILLER_41_316 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_388 ();
 sg13g2_decap_4 FILLER_41_395 ();
 sg13g2_fill_1 FILLER_41_399 ();
 sg13g2_decap_4 FILLER_41_406 ();
 sg13g2_decap_4 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_461 ();
 sg13g2_decap_4 FILLER_41_468 ();
 sg13g2_fill_2 FILLER_41_506 ();
 sg13g2_fill_1 FILLER_41_516 ();
 sg13g2_fill_1 FILLER_41_522 ();
 sg13g2_fill_1 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_573 ();
 sg13g2_fill_1 FILLER_41_614 ();
 sg13g2_fill_2 FILLER_41_692 ();
 sg13g2_fill_1 FILLER_41_755 ();
 sg13g2_fill_2 FILLER_41_790 ();
 sg13g2_fill_1 FILLER_41_812 ();
 sg13g2_fill_1 FILLER_41_817 ();
 sg13g2_fill_1 FILLER_41_844 ();
 sg13g2_decap_4 FILLER_41_849 ();
 sg13g2_decap_4 FILLER_41_860 ();
 sg13g2_fill_2 FILLER_41_864 ();
 sg13g2_decap_8 FILLER_41_871 ();
 sg13g2_fill_1 FILLER_41_878 ();
 sg13g2_fill_2 FILLER_41_905 ();
 sg13g2_fill_1 FILLER_41_907 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_fill_2 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_974 ();
 sg13g2_decap_8 FILLER_41_981 ();
 sg13g2_decap_8 FILLER_41_988 ();
 sg13g2_fill_2 FILLER_41_1055 ();
 sg13g2_fill_2 FILLER_41_1066 ();
 sg13g2_fill_2 FILLER_41_1079 ();
 sg13g2_fill_1 FILLER_41_1081 ();
 sg13g2_fill_2 FILLER_41_1093 ();
 sg13g2_fill_1 FILLER_41_1103 ();
 sg13g2_fill_1 FILLER_41_1108 ();
 sg13g2_fill_1 FILLER_41_1113 ();
 sg13g2_fill_1 FILLER_41_1124 ();
 sg13g2_fill_2 FILLER_41_1146 ();
 sg13g2_fill_1 FILLER_41_1148 ();
 sg13g2_fill_2 FILLER_41_1219 ();
 sg13g2_fill_1 FILLER_41_1221 ();
 sg13g2_decap_4 FILLER_41_1238 ();
 sg13g2_fill_2 FILLER_41_1258 ();
 sg13g2_fill_1 FILLER_41_1265 ();
 sg13g2_fill_1 FILLER_41_1295 ();
 sg13g2_fill_1 FILLER_41_1350 ();
 sg13g2_fill_1 FILLER_41_1390 ();
 sg13g2_fill_2 FILLER_41_1396 ();
 sg13g2_fill_2 FILLER_41_1409 ();
 sg13g2_fill_1 FILLER_41_1431 ();
 sg13g2_fill_2 FILLER_41_1441 ();
 sg13g2_fill_1 FILLER_41_1443 ();
 sg13g2_fill_2 FILLER_41_1447 ();
 sg13g2_decap_8 FILLER_41_1453 ();
 sg13g2_fill_2 FILLER_41_1460 ();
 sg13g2_fill_1 FILLER_41_1462 ();
 sg13g2_fill_1 FILLER_41_1471 ();
 sg13g2_decap_4 FILLER_41_1481 ();
 sg13g2_fill_1 FILLER_41_1490 ();
 sg13g2_fill_2 FILLER_41_1533 ();
 sg13g2_fill_1 FILLER_41_1540 ();
 sg13g2_decap_4 FILLER_41_1547 ();
 sg13g2_fill_2 FILLER_41_1551 ();
 sg13g2_fill_1 FILLER_41_1561 ();
 sg13g2_fill_2 FILLER_41_1567 ();
 sg13g2_fill_1 FILLER_41_1569 ();
 sg13g2_decap_8 FILLER_41_1630 ();
 sg13g2_decap_8 FILLER_41_1637 ();
 sg13g2_fill_1 FILLER_41_1644 ();
 sg13g2_fill_2 FILLER_41_1650 ();
 sg13g2_fill_2 FILLER_41_1656 ();
 sg13g2_decap_4 FILLER_41_1664 ();
 sg13g2_fill_1 FILLER_41_1668 ();
 sg13g2_fill_2 FILLER_41_1702 ();
 sg13g2_fill_1 FILLER_41_1713 ();
 sg13g2_decap_8 FILLER_41_1753 ();
 sg13g2_decap_4 FILLER_41_1760 ();
 sg13g2_fill_2 FILLER_41_1771 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_fill_1 FILLER_41_1781 ();
 sg13g2_fill_1 FILLER_41_1788 ();
 sg13g2_fill_1 FILLER_41_1800 ();
 sg13g2_fill_2 FILLER_41_1806 ();
 sg13g2_fill_2 FILLER_41_1816 ();
 sg13g2_fill_1 FILLER_41_1818 ();
 sg13g2_fill_1 FILLER_41_1834 ();
 sg13g2_fill_1 FILLER_41_1839 ();
 sg13g2_fill_1 FILLER_41_1845 ();
 sg13g2_fill_2 FILLER_41_1871 ();
 sg13g2_fill_2 FILLER_41_1878 ();
 sg13g2_fill_1 FILLER_41_1880 ();
 sg13g2_fill_2 FILLER_41_1900 ();
 sg13g2_decap_8 FILLER_41_1906 ();
 sg13g2_decap_8 FILLER_41_1913 ();
 sg13g2_decap_8 FILLER_41_1920 ();
 sg13g2_decap_8 FILLER_41_1927 ();
 sg13g2_decap_8 FILLER_41_1934 ();
 sg13g2_decap_8 FILLER_41_1941 ();
 sg13g2_decap_8 FILLER_41_1948 ();
 sg13g2_decap_8 FILLER_41_1955 ();
 sg13g2_decap_8 FILLER_41_1962 ();
 sg13g2_decap_8 FILLER_41_1969 ();
 sg13g2_fill_2 FILLER_41_1976 ();
 sg13g2_decap_8 FILLER_41_1986 ();
 sg13g2_fill_2 FILLER_41_1993 ();
 sg13g2_fill_1 FILLER_41_1995 ();
 sg13g2_decap_8 FILLER_41_2000 ();
 sg13g2_decap_8 FILLER_41_2007 ();
 sg13g2_decap_8 FILLER_41_2014 ();
 sg13g2_decap_8 FILLER_41_2021 ();
 sg13g2_decap_8 FILLER_41_2028 ();
 sg13g2_decap_8 FILLER_41_2035 ();
 sg13g2_decap_8 FILLER_41_2042 ();
 sg13g2_fill_1 FILLER_41_2049 ();
 sg13g2_fill_1 FILLER_41_2080 ();
 sg13g2_fill_1 FILLER_41_2091 ();
 sg13g2_fill_1 FILLER_41_2097 ();
 sg13g2_fill_1 FILLER_41_2102 ();
 sg13g2_decap_4 FILLER_41_2109 ();
 sg13g2_fill_2 FILLER_41_2127 ();
 sg13g2_fill_1 FILLER_41_2134 ();
 sg13g2_fill_1 FILLER_41_2140 ();
 sg13g2_fill_2 FILLER_41_2151 ();
 sg13g2_decap_8 FILLER_41_2167 ();
 sg13g2_fill_1 FILLER_41_2174 ();
 sg13g2_fill_2 FILLER_41_2183 ();
 sg13g2_fill_2 FILLER_41_2193 ();
 sg13g2_fill_1 FILLER_41_2195 ();
 sg13g2_fill_2 FILLER_41_2235 ();
 sg13g2_fill_1 FILLER_41_2243 ();
 sg13g2_fill_1 FILLER_41_2249 ();
 sg13g2_fill_2 FILLER_41_2254 ();
 sg13g2_fill_2 FILLER_41_2308 ();
 sg13g2_fill_1 FILLER_41_2310 ();
 sg13g2_decap_4 FILLER_41_2319 ();
 sg13g2_fill_1 FILLER_41_2345 ();
 sg13g2_decap_4 FILLER_41_2350 ();
 sg13g2_decap_8 FILLER_41_2370 ();
 sg13g2_fill_2 FILLER_41_2377 ();
 sg13g2_decap_8 FILLER_41_2387 ();
 sg13g2_fill_1 FILLER_41_2394 ();
 sg13g2_fill_1 FILLER_41_2409 ();
 sg13g2_fill_2 FILLER_41_2420 ();
 sg13g2_fill_1 FILLER_41_2422 ();
 sg13g2_decap_4 FILLER_41_2427 ();
 sg13g2_fill_2 FILLER_41_2435 ();
 sg13g2_fill_1 FILLER_41_2437 ();
 sg13g2_fill_1 FILLER_41_2443 ();
 sg13g2_fill_2 FILLER_41_2453 ();
 sg13g2_fill_1 FILLER_41_2455 ();
 sg13g2_fill_2 FILLER_41_2475 ();
 sg13g2_fill_1 FILLER_41_2477 ();
 sg13g2_decap_4 FILLER_41_2483 ();
 sg13g2_fill_1 FILLER_41_2501 ();
 sg13g2_fill_2 FILLER_41_2508 ();
 sg13g2_fill_1 FILLER_41_2510 ();
 sg13g2_fill_2 FILLER_41_2522 ();
 sg13g2_fill_1 FILLER_41_2524 ();
 sg13g2_decap_4 FILLER_41_2540 ();
 sg13g2_fill_2 FILLER_41_2544 ();
 sg13g2_fill_1 FILLER_41_2568 ();
 sg13g2_fill_1 FILLER_41_2574 ();
 sg13g2_fill_2 FILLER_41_2579 ();
 sg13g2_fill_1 FILLER_41_2581 ();
 sg13g2_fill_1 FILLER_41_2588 ();
 sg13g2_fill_1 FILLER_41_2601 ();
 sg13g2_decap_8 FILLER_41_2641 ();
 sg13g2_decap_8 FILLER_41_2648 ();
 sg13g2_decap_8 FILLER_41_2655 ();
 sg13g2_decap_8 FILLER_41_2662 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_fill_1 FILLER_42_113 ();
 sg13g2_fill_1 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_160 ();
 sg13g2_fill_1 FILLER_42_187 ();
 sg13g2_fill_1 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_256 ();
 sg13g2_fill_2 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_decap_4 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_fill_2 FILLER_42_460 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_fill_2 FILLER_42_489 ();
 sg13g2_fill_1 FILLER_42_517 ();
 sg13g2_fill_1 FILLER_42_527 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_decap_4 FILLER_42_586 ();
 sg13g2_fill_1 FILLER_42_590 ();
 sg13g2_decap_8 FILLER_42_596 ();
 sg13g2_decap_4 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_646 ();
 sg13g2_fill_1 FILLER_42_653 ();
 sg13g2_fill_2 FILLER_42_659 ();
 sg13g2_fill_1 FILLER_42_661 ();
 sg13g2_fill_1 FILLER_42_688 ();
 sg13g2_fill_2 FILLER_42_782 ();
 sg13g2_fill_2 FILLER_42_809 ();
 sg13g2_decap_4 FILLER_42_860 ();
 sg13g2_fill_2 FILLER_42_864 ();
 sg13g2_decap_8 FILLER_42_910 ();
 sg13g2_fill_1 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_922 ();
 sg13g2_fill_2 FILLER_42_947 ();
 sg13g2_decap_4 FILLER_42_953 ();
 sg13g2_fill_1 FILLER_42_957 ();
 sg13g2_decap_8 FILLER_42_962 ();
 sg13g2_decap_8 FILLER_42_969 ();
 sg13g2_fill_1 FILLER_42_976 ();
 sg13g2_fill_2 FILLER_42_1003 ();
 sg13g2_fill_1 FILLER_42_1005 ();
 sg13g2_decap_4 FILLER_42_1009 ();
 sg13g2_decap_4 FILLER_42_1082 ();
 sg13g2_fill_1 FILLER_42_1086 ();
 sg13g2_fill_1 FILLER_42_1123 ();
 sg13g2_fill_1 FILLER_42_1180 ();
 sg13g2_fill_1 FILLER_42_1193 ();
 sg13g2_fill_2 FILLER_42_1205 ();
 sg13g2_decap_4 FILLER_42_1236 ();
 sg13g2_fill_2 FILLER_42_1271 ();
 sg13g2_fill_1 FILLER_42_1309 ();
 sg13g2_fill_2 FILLER_42_1346 ();
 sg13g2_fill_2 FILLER_42_1354 ();
 sg13g2_fill_1 FILLER_42_1360 ();
 sg13g2_fill_2 FILLER_42_1376 ();
 sg13g2_fill_1 FILLER_42_1388 ();
 sg13g2_fill_2 FILLER_42_1393 ();
 sg13g2_fill_1 FILLER_42_1411 ();
 sg13g2_fill_2 FILLER_42_1432 ();
 sg13g2_fill_1 FILLER_42_1439 ();
 sg13g2_decap_4 FILLER_42_1448 ();
 sg13g2_decap_8 FILLER_42_1469 ();
 sg13g2_decap_8 FILLER_42_1476 ();
 sg13g2_decap_8 FILLER_42_1483 ();
 sg13g2_fill_1 FILLER_42_1490 ();
 sg13g2_fill_2 FILLER_42_1500 ();
 sg13g2_decap_8 FILLER_42_1511 ();
 sg13g2_decap_4 FILLER_42_1518 ();
 sg13g2_fill_2 FILLER_42_1522 ();
 sg13g2_fill_2 FILLER_42_1527 ();
 sg13g2_decap_8 FILLER_42_1532 ();
 sg13g2_decap_8 FILLER_42_1539 ();
 sg13g2_fill_2 FILLER_42_1546 ();
 sg13g2_fill_1 FILLER_42_1548 ();
 sg13g2_decap_4 FILLER_42_1597 ();
 sg13g2_decap_8 FILLER_42_1636 ();
 sg13g2_fill_2 FILLER_42_1643 ();
 sg13g2_fill_1 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1669 ();
 sg13g2_decap_4 FILLER_42_1676 ();
 sg13g2_decap_4 FILLER_42_1710 ();
 sg13g2_decap_4 FILLER_42_1720 ();
 sg13g2_decap_8 FILLER_42_1734 ();
 sg13g2_decap_8 FILLER_42_1741 ();
 sg13g2_fill_2 FILLER_42_1748 ();
 sg13g2_fill_1 FILLER_42_1750 ();
 sg13g2_decap_4 FILLER_42_1760 ();
 sg13g2_fill_2 FILLER_42_1764 ();
 sg13g2_fill_1 FILLER_42_1771 ();
 sg13g2_decap_4 FILLER_42_1797 ();
 sg13g2_fill_1 FILLER_42_1801 ();
 sg13g2_fill_2 FILLER_42_1806 ();
 sg13g2_fill_1 FILLER_42_1829 ();
 sg13g2_fill_1 FILLER_42_1833 ();
 sg13g2_fill_1 FILLER_42_1840 ();
 sg13g2_fill_1 FILLER_42_1858 ();
 sg13g2_decap_4 FILLER_42_1898 ();
 sg13g2_fill_1 FILLER_42_1902 ();
 sg13g2_decap_8 FILLER_42_1907 ();
 sg13g2_decap_8 FILLER_42_1914 ();
 sg13g2_decap_8 FILLER_42_1921 ();
 sg13g2_decap_4 FILLER_42_1928 ();
 sg13g2_fill_1 FILLER_42_1932 ();
 sg13g2_decap_8 FILLER_42_1942 ();
 sg13g2_decap_8 FILLER_42_1949 ();
 sg13g2_decap_8 FILLER_42_1956 ();
 sg13g2_decap_8 FILLER_42_1963 ();
 sg13g2_decap_8 FILLER_42_1970 ();
 sg13g2_decap_8 FILLER_42_1977 ();
 sg13g2_decap_4 FILLER_42_1984 ();
 sg13g2_fill_1 FILLER_42_1988 ();
 sg13g2_decap_4 FILLER_42_1994 ();
 sg13g2_fill_2 FILLER_42_1998 ();
 sg13g2_decap_8 FILLER_42_2008 ();
 sg13g2_decap_8 FILLER_42_2015 ();
 sg13g2_decap_8 FILLER_42_2022 ();
 sg13g2_decap_8 FILLER_42_2029 ();
 sg13g2_decap_8 FILLER_42_2036 ();
 sg13g2_decap_8 FILLER_42_2043 ();
 sg13g2_decap_8 FILLER_42_2050 ();
 sg13g2_decap_8 FILLER_42_2057 ();
 sg13g2_fill_1 FILLER_42_2068 ();
 sg13g2_decap_4 FILLER_42_2152 ();
 sg13g2_decap_8 FILLER_42_2172 ();
 sg13g2_decap_8 FILLER_42_2179 ();
 sg13g2_fill_2 FILLER_42_2186 ();
 sg13g2_decap_8 FILLER_42_2193 ();
 sg13g2_decap_4 FILLER_42_2200 ();
 sg13g2_fill_2 FILLER_42_2204 ();
 sg13g2_decap_8 FILLER_42_2211 ();
 sg13g2_fill_1 FILLER_42_2218 ();
 sg13g2_decap_4 FILLER_42_2232 ();
 sg13g2_fill_1 FILLER_42_2240 ();
 sg13g2_fill_1 FILLER_42_2249 ();
 sg13g2_fill_2 FILLER_42_2279 ();
 sg13g2_fill_1 FILLER_42_2281 ();
 sg13g2_fill_2 FILLER_42_2312 ();
 sg13g2_decap_8 FILLER_42_2370 ();
 sg13g2_decap_8 FILLER_42_2377 ();
 sg13g2_decap_4 FILLER_42_2424 ();
 sg13g2_decap_4 FILLER_42_2464 ();
 sg13g2_decap_4 FILLER_42_2563 ();
 sg13g2_fill_1 FILLER_42_2567 ();
 sg13g2_fill_1 FILLER_42_2617 ();
 sg13g2_decap_8 FILLER_42_2628 ();
 sg13g2_decap_8 FILLER_42_2635 ();
 sg13g2_decap_8 FILLER_42_2642 ();
 sg13g2_decap_8 FILLER_42_2649 ();
 sg13g2_decap_8 FILLER_42_2656 ();
 sg13g2_decap_8 FILLER_42_2663 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_41 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_2 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_156 ();
 sg13g2_decap_4 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_fill_2 FILLER_43_195 ();
 sg13g2_fill_2 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_287 ();
 sg13g2_fill_2 FILLER_43_332 ();
 sg13g2_fill_2 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_fill_2 FILLER_43_394 ();
 sg13g2_fill_1 FILLER_43_396 ();
 sg13g2_fill_1 FILLER_43_435 ();
 sg13g2_fill_1 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_480 ();
 sg13g2_decap_8 FILLER_43_487 ();
 sg13g2_fill_1 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_516 ();
 sg13g2_fill_2 FILLER_43_572 ();
 sg13g2_fill_1 FILLER_43_578 ();
 sg13g2_decap_4 FILLER_43_588 ();
 sg13g2_fill_2 FILLER_43_592 ();
 sg13g2_fill_2 FILLER_43_617 ();
 sg13g2_fill_1 FILLER_43_638 ();
 sg13g2_fill_2 FILLER_43_647 ();
 sg13g2_fill_1 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_fill_2 FILLER_43_669 ();
 sg13g2_fill_1 FILLER_43_671 ();
 sg13g2_decap_8 FILLER_43_681 ();
 sg13g2_fill_1 FILLER_43_688 ();
 sg13g2_decap_4 FILLER_43_692 ();
 sg13g2_fill_2 FILLER_43_733 ();
 sg13g2_fill_1 FILLER_43_793 ();
 sg13g2_fill_2 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_836 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_decap_4 FILLER_43_849 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_4 FILLER_43_868 ();
 sg13g2_fill_2 FILLER_43_877 ();
 sg13g2_decap_4 FILLER_43_905 ();
 sg13g2_decap_8 FILLER_43_913 ();
 sg13g2_fill_2 FILLER_43_954 ();
 sg13g2_fill_1 FILLER_43_956 ();
 sg13g2_decap_8 FILLER_43_963 ();
 sg13g2_fill_2 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_977 ();
 sg13g2_fill_1 FILLER_43_988 ();
 sg13g2_fill_1 FILLER_43_1000 ();
 sg13g2_fill_2 FILLER_43_1040 ();
 sg13g2_decap_4 FILLER_43_1076 ();
 sg13g2_fill_2 FILLER_43_1084 ();
 sg13g2_fill_1 FILLER_43_1086 ();
 sg13g2_decap_8 FILLER_43_1093 ();
 sg13g2_fill_2 FILLER_43_1100 ();
 sg13g2_fill_1 FILLER_43_1102 ();
 sg13g2_fill_2 FILLER_43_1112 ();
 sg13g2_fill_2 FILLER_43_1127 ();
 sg13g2_fill_1 FILLER_43_1129 ();
 sg13g2_fill_2 FILLER_43_1160 ();
 sg13g2_fill_1 FILLER_43_1167 ();
 sg13g2_fill_1 FILLER_43_1172 ();
 sg13g2_fill_2 FILLER_43_1187 ();
 sg13g2_fill_2 FILLER_43_1202 ();
 sg13g2_fill_2 FILLER_43_1211 ();
 sg13g2_decap_4 FILLER_43_1228 ();
 sg13g2_fill_1 FILLER_43_1232 ();
 sg13g2_fill_2 FILLER_43_1242 ();
 sg13g2_fill_1 FILLER_43_1262 ();
 sg13g2_fill_1 FILLER_43_1354 ();
 sg13g2_fill_2 FILLER_43_1387 ();
 sg13g2_fill_1 FILLER_43_1430 ();
 sg13g2_decap_8 FILLER_43_1434 ();
 sg13g2_fill_1 FILLER_43_1441 ();
 sg13g2_decap_4 FILLER_43_1461 ();
 sg13g2_fill_1 FILLER_43_1465 ();
 sg13g2_decap_8 FILLER_43_1471 ();
 sg13g2_fill_2 FILLER_43_1485 ();
 sg13g2_fill_2 FILLER_43_1492 ();
 sg13g2_decap_4 FILLER_43_1498 ();
 sg13g2_fill_1 FILLER_43_1506 ();
 sg13g2_fill_1 FILLER_43_1512 ();
 sg13g2_fill_1 FILLER_43_1590 ();
 sg13g2_fill_2 FILLER_43_1604 ();
 sg13g2_fill_1 FILLER_43_1606 ();
 sg13g2_fill_1 FILLER_43_1615 ();
 sg13g2_fill_1 FILLER_43_1619 ();
 sg13g2_fill_2 FILLER_43_1623 ();
 sg13g2_fill_1 FILLER_43_1625 ();
 sg13g2_fill_2 FILLER_43_1630 ();
 sg13g2_fill_1 FILLER_43_1663 ();
 sg13g2_fill_1 FILLER_43_1683 ();
 sg13g2_fill_1 FILLER_43_1696 ();
 sg13g2_fill_1 FILLER_43_1701 ();
 sg13g2_fill_1 FILLER_43_1709 ();
 sg13g2_fill_2 FILLER_43_1715 ();
 sg13g2_decap_8 FILLER_43_1721 ();
 sg13g2_decap_8 FILLER_43_1738 ();
 sg13g2_decap_8 FILLER_43_1745 ();
 sg13g2_fill_1 FILLER_43_1752 ();
 sg13g2_fill_2 FILLER_43_1805 ();
 sg13g2_decap_8 FILLER_43_1811 ();
 sg13g2_decap_4 FILLER_43_1818 ();
 sg13g2_fill_1 FILLER_43_1822 ();
 sg13g2_fill_1 FILLER_43_1828 ();
 sg13g2_decap_8 FILLER_43_1834 ();
 sg13g2_fill_1 FILLER_43_1841 ();
 sg13g2_fill_2 FILLER_43_1850 ();
 sg13g2_fill_1 FILLER_43_1852 ();
 sg13g2_fill_1 FILLER_43_1858 ();
 sg13g2_decap_4 FILLER_43_1864 ();
 sg13g2_fill_2 FILLER_43_1868 ();
 sg13g2_decap_4 FILLER_43_1875 ();
 sg13g2_fill_2 FILLER_43_1879 ();
 sg13g2_decap_4 FILLER_43_1896 ();
 sg13g2_fill_2 FILLER_43_1900 ();
 sg13g2_decap_8 FILLER_43_1909 ();
 sg13g2_decap_8 FILLER_43_1916 ();
 sg13g2_fill_1 FILLER_43_1923 ();
 sg13g2_fill_1 FILLER_43_1928 ();
 sg13g2_fill_1 FILLER_43_1942 ();
 sg13g2_decap_8 FILLER_43_1960 ();
 sg13g2_decap_8 FILLER_43_1977 ();
 sg13g2_decap_8 FILLER_43_1984 ();
 sg13g2_decap_8 FILLER_43_1991 ();
 sg13g2_decap_8 FILLER_43_1998 ();
 sg13g2_decap_8 FILLER_43_2005 ();
 sg13g2_decap_8 FILLER_43_2012 ();
 sg13g2_decap_8 FILLER_43_2019 ();
 sg13g2_decap_8 FILLER_43_2026 ();
 sg13g2_decap_8 FILLER_43_2033 ();
 sg13g2_decap_8 FILLER_43_2040 ();
 sg13g2_decap_8 FILLER_43_2047 ();
 sg13g2_decap_8 FILLER_43_2054 ();
 sg13g2_decap_8 FILLER_43_2061 ();
 sg13g2_decap_4 FILLER_43_2068 ();
 sg13g2_fill_2 FILLER_43_2072 ();
 sg13g2_fill_2 FILLER_43_2078 ();
 sg13g2_fill_1 FILLER_43_2080 ();
 sg13g2_fill_2 FILLER_43_2094 ();
 sg13g2_decap_8 FILLER_43_2118 ();
 sg13g2_fill_2 FILLER_43_2162 ();
 sg13g2_fill_1 FILLER_43_2164 ();
 sg13g2_fill_1 FILLER_43_2171 ();
 sg13g2_fill_1 FILLER_43_2177 ();
 sg13g2_fill_2 FILLER_43_2182 ();
 sg13g2_decap_4 FILLER_43_2218 ();
 sg13g2_fill_1 FILLER_43_2222 ();
 sg13g2_decap_8 FILLER_43_2228 ();
 sg13g2_decap_8 FILLER_43_2235 ();
 sg13g2_decap_4 FILLER_43_2242 ();
 sg13g2_fill_1 FILLER_43_2246 ();
 sg13g2_fill_2 FILLER_43_2273 ();
 sg13g2_decap_8 FILLER_43_2285 ();
 sg13g2_fill_1 FILLER_43_2292 ();
 sg13g2_fill_1 FILLER_43_2309 ();
 sg13g2_fill_1 FILLER_43_2324 ();
 sg13g2_fill_2 FILLER_43_2335 ();
 sg13g2_fill_1 FILLER_43_2363 ();
 sg13g2_fill_1 FILLER_43_2370 ();
 sg13g2_fill_1 FILLER_43_2381 ();
 sg13g2_fill_1 FILLER_43_2386 ();
 sg13g2_decap_4 FILLER_43_2392 ();
 sg13g2_fill_1 FILLER_43_2396 ();
 sg13g2_decap_4 FILLER_43_2423 ();
 sg13g2_fill_2 FILLER_43_2427 ();
 sg13g2_fill_1 FILLER_43_2499 ();
 sg13g2_fill_1 FILLER_43_2508 ();
 sg13g2_decap_4 FILLER_43_2548 ();
 sg13g2_fill_2 FILLER_43_2552 ();
 sg13g2_fill_2 FILLER_43_2574 ();
 sg13g2_fill_1 FILLER_43_2620 ();
 sg13g2_decap_8 FILLER_43_2651 ();
 sg13g2_decap_8 FILLER_43_2658 ();
 sg13g2_decap_4 FILLER_43_2665 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_36 ();
 sg13g2_fill_1 FILLER_44_43 ();
 sg13g2_fill_2 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_177 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_190 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_1 FILLER_44_271 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_361 ();
 sg13g2_fill_2 FILLER_44_366 ();
 sg13g2_decap_4 FILLER_44_374 ();
 sg13g2_fill_2 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_fill_1 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_405 ();
 sg13g2_fill_2 FILLER_44_411 ();
 sg13g2_fill_1 FILLER_44_413 ();
 sg13g2_fill_2 FILLER_44_432 ();
 sg13g2_decap_8 FILLER_44_470 ();
 sg13g2_decap_4 FILLER_44_477 ();
 sg13g2_fill_1 FILLER_44_481 ();
 sg13g2_decap_4 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_499 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_decap_4 FILLER_44_601 ();
 sg13g2_fill_2 FILLER_44_630 ();
 sg13g2_fill_2 FILLER_44_655 ();
 sg13g2_decap_4 FILLER_44_673 ();
 sg13g2_decap_4 FILLER_44_681 ();
 sg13g2_fill_2 FILLER_44_685 ();
 sg13g2_fill_2 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_713 ();
 sg13g2_decap_8 FILLER_44_720 ();
 sg13g2_decap_4 FILLER_44_727 ();
 sg13g2_fill_2 FILLER_44_731 ();
 sg13g2_fill_2 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_834 ();
 sg13g2_decap_8 FILLER_44_841 ();
 sg13g2_decap_4 FILLER_44_848 ();
 sg13g2_fill_1 FILLER_44_852 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_fill_2 FILLER_44_899 ();
 sg13g2_fill_1 FILLER_44_901 ();
 sg13g2_fill_2 FILLER_44_928 ();
 sg13g2_fill_1 FILLER_44_948 ();
 sg13g2_fill_1 FILLER_44_953 ();
 sg13g2_fill_2 FILLER_44_961 ();
 sg13g2_fill_2 FILLER_44_967 ();
 sg13g2_fill_1 FILLER_44_969 ();
 sg13g2_fill_2 FILLER_44_984 ();
 sg13g2_fill_2 FILLER_44_1008 ();
 sg13g2_fill_2 FILLER_44_1090 ();
 sg13g2_fill_1 FILLER_44_1106 ();
 sg13g2_fill_2 FILLER_44_1110 ();
 sg13g2_fill_1 FILLER_44_1112 ();
 sg13g2_decap_4 FILLER_44_1116 ();
 sg13g2_fill_1 FILLER_44_1120 ();
 sg13g2_decap_8 FILLER_44_1128 ();
 sg13g2_fill_1 FILLER_44_1135 ();
 sg13g2_fill_2 FILLER_44_1152 ();
 sg13g2_decap_4 FILLER_44_1212 ();
 sg13g2_fill_1 FILLER_44_1216 ();
 sg13g2_decap_4 FILLER_44_1222 ();
 sg13g2_fill_2 FILLER_44_1226 ();
 sg13g2_fill_1 FILLER_44_1235 ();
 sg13g2_fill_2 FILLER_44_1250 ();
 sg13g2_fill_2 FILLER_44_1321 ();
 sg13g2_fill_1 FILLER_44_1331 ();
 sg13g2_fill_2 FILLER_44_1359 ();
 sg13g2_fill_1 FILLER_44_1392 ();
 sg13g2_fill_2 FILLER_44_1406 ();
 sg13g2_fill_2 FILLER_44_1424 ();
 sg13g2_fill_2 FILLER_44_1436 ();
 sg13g2_fill_1 FILLER_44_1438 ();
 sg13g2_fill_1 FILLER_44_1460 ();
 sg13g2_fill_2 FILLER_44_1466 ();
 sg13g2_fill_1 FILLER_44_1468 ();
 sg13g2_fill_2 FILLER_44_1474 ();
 sg13g2_fill_2 FILLER_44_1480 ();
 sg13g2_fill_2 FILLER_44_1486 ();
 sg13g2_decap_8 FILLER_44_1497 ();
 sg13g2_decap_4 FILLER_44_1504 ();
 sg13g2_fill_1 FILLER_44_1517 ();
 sg13g2_fill_1 FILLER_44_1543 ();
 sg13g2_fill_2 FILLER_44_1618 ();
 sg13g2_fill_2 FILLER_44_1627 ();
 sg13g2_fill_2 FILLER_44_1633 ();
 sg13g2_fill_1 FILLER_44_1639 ();
 sg13g2_fill_1 FILLER_44_1644 ();
 sg13g2_decap_4 FILLER_44_1648 ();
 sg13g2_decap_4 FILLER_44_1657 ();
 sg13g2_fill_1 FILLER_44_1661 ();
 sg13g2_fill_1 FILLER_44_1667 ();
 sg13g2_fill_2 FILLER_44_1709 ();
 sg13g2_decap_8 FILLER_44_1721 ();
 sg13g2_decap_4 FILLER_44_1728 ();
 sg13g2_fill_1 FILLER_44_1732 ();
 sg13g2_decap_8 FILLER_44_1763 ();
 sg13g2_fill_2 FILLER_44_1770 ();
 sg13g2_fill_1 FILLER_44_1772 ();
 sg13g2_decap_8 FILLER_44_1778 ();
 sg13g2_decap_8 FILLER_44_1785 ();
 sg13g2_decap_8 FILLER_44_1792 ();
 sg13g2_decap_8 FILLER_44_1799 ();
 sg13g2_decap_8 FILLER_44_1806 ();
 sg13g2_decap_8 FILLER_44_1813 ();
 sg13g2_decap_8 FILLER_44_1820 ();
 sg13g2_fill_1 FILLER_44_1827 ();
 sg13g2_decap_8 FILLER_44_1835 ();
 sg13g2_decap_8 FILLER_44_1842 ();
 sg13g2_fill_1 FILLER_44_1849 ();
 sg13g2_decap_8 FILLER_44_1854 ();
 sg13g2_decap_8 FILLER_44_1861 ();
 sg13g2_decap_4 FILLER_44_1868 ();
 sg13g2_fill_1 FILLER_44_1872 ();
 sg13g2_decap_8 FILLER_44_1882 ();
 sg13g2_decap_8 FILLER_44_1889 ();
 sg13g2_decap_8 FILLER_44_1896 ();
 sg13g2_decap_8 FILLER_44_1903 ();
 sg13g2_fill_2 FILLER_44_1910 ();
 sg13g2_decap_8 FILLER_44_1920 ();
 sg13g2_decap_8 FILLER_44_1927 ();
 sg13g2_decap_4 FILLER_44_1934 ();
 sg13g2_fill_1 FILLER_44_1938 ();
 sg13g2_decap_4 FILLER_44_1945 ();
 sg13g2_decap_8 FILLER_44_1953 ();
 sg13g2_decap_4 FILLER_44_1960 ();
 sg13g2_decap_4 FILLER_44_1970 ();
 sg13g2_fill_2 FILLER_44_1974 ();
 sg13g2_decap_8 FILLER_44_1981 ();
 sg13g2_fill_1 FILLER_44_1988 ();
 sg13g2_decap_8 FILLER_44_1993 ();
 sg13g2_fill_2 FILLER_44_2000 ();
 sg13g2_fill_1 FILLER_44_2002 ();
 sg13g2_decap_8 FILLER_44_2008 ();
 sg13g2_decap_8 FILLER_44_2015 ();
 sg13g2_decap_8 FILLER_44_2022 ();
 sg13g2_decap_8 FILLER_44_2029 ();
 sg13g2_decap_8 FILLER_44_2036 ();
 sg13g2_decap_8 FILLER_44_2043 ();
 sg13g2_decap_8 FILLER_44_2050 ();
 sg13g2_decap_8 FILLER_44_2057 ();
 sg13g2_decap_8 FILLER_44_2064 ();
 sg13g2_fill_2 FILLER_44_2071 ();
 sg13g2_decap_8 FILLER_44_2121 ();
 sg13g2_decap_8 FILLER_44_2128 ();
 sg13g2_decap_8 FILLER_44_2135 ();
 sg13g2_fill_1 FILLER_44_2142 ();
 sg13g2_fill_2 FILLER_44_2156 ();
 sg13g2_fill_1 FILLER_44_2158 ();
 sg13g2_fill_1 FILLER_44_2172 ();
 sg13g2_fill_1 FILLER_44_2185 ();
 sg13g2_fill_1 FILLER_44_2192 ();
 sg13g2_fill_1 FILLER_44_2197 ();
 sg13g2_fill_1 FILLER_44_2203 ();
 sg13g2_fill_1 FILLER_44_2208 ();
 sg13g2_fill_1 FILLER_44_2213 ();
 sg13g2_fill_1 FILLER_44_2224 ();
 sg13g2_fill_1 FILLER_44_2240 ();
 sg13g2_decap_8 FILLER_44_2245 ();
 sg13g2_decap_8 FILLER_44_2316 ();
 sg13g2_decap_8 FILLER_44_2323 ();
 sg13g2_fill_2 FILLER_44_2340 ();
 sg13g2_fill_1 FILLER_44_2346 ();
 sg13g2_fill_1 FILLER_44_2357 ();
 sg13g2_fill_2 FILLER_44_2362 ();
 sg13g2_fill_2 FILLER_44_2393 ();
 sg13g2_fill_1 FILLER_44_2409 ();
 sg13g2_fill_2 FILLER_44_2420 ();
 sg13g2_fill_1 FILLER_44_2422 ();
 sg13g2_fill_2 FILLER_44_2453 ();
 sg13g2_fill_1 FILLER_44_2455 ();
 sg13g2_decap_8 FILLER_44_2460 ();
 sg13g2_decap_4 FILLER_44_2467 ();
 sg13g2_fill_1 FILLER_44_2471 ();
 sg13g2_fill_2 FILLER_44_2486 ();
 sg13g2_fill_1 FILLER_44_2488 ();
 sg13g2_fill_1 FILLER_44_2530 ();
 sg13g2_fill_2 FILLER_44_2609 ();
 sg13g2_fill_1 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2622 ();
 sg13g2_fill_1 FILLER_44_2629 ();
 sg13g2_decap_8 FILLER_44_2656 ();
 sg13g2_decap_8 FILLER_44_2663 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_fill_1 FILLER_45_10 ();
 sg13g2_fill_1 FILLER_45_33 ();
 sg13g2_fill_1 FILLER_45_51 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_fill_2 FILLER_45_79 ();
 sg13g2_fill_2 FILLER_45_130 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_fill_2 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_fill_1 FILLER_45_346 ();
 sg13g2_fill_1 FILLER_45_409 ();
 sg13g2_fill_1 FILLER_45_441 ();
 sg13g2_decap_4 FILLER_45_446 ();
 sg13g2_fill_1 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_4 FILLER_45_469 ();
 sg13g2_fill_1 FILLER_45_473 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_fill_1 FILLER_45_522 ();
 sg13g2_fill_1 FILLER_45_536 ();
 sg13g2_fill_1 FILLER_45_606 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_fill_2 FILLER_45_619 ();
 sg13g2_fill_1 FILLER_45_621 ();
 sg13g2_fill_2 FILLER_45_626 ();
 sg13g2_fill_1 FILLER_45_628 ();
 sg13g2_fill_1 FILLER_45_638 ();
 sg13g2_fill_1 FILLER_45_644 ();
 sg13g2_fill_2 FILLER_45_677 ();
 sg13g2_fill_2 FILLER_45_687 ();
 sg13g2_fill_1 FILLER_45_696 ();
 sg13g2_fill_2 FILLER_45_705 ();
 sg13g2_fill_2 FILLER_45_717 ();
 sg13g2_fill_1 FILLER_45_733 ();
 sg13g2_fill_1 FILLER_45_752 ();
 sg13g2_fill_1 FILLER_45_760 ();
 sg13g2_decap_4 FILLER_45_812 ();
 sg13g2_fill_1 FILLER_45_816 ();
 sg13g2_decap_4 FILLER_45_830 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_fill_2 FILLER_45_865 ();
 sg13g2_fill_2 FILLER_45_893 ();
 sg13g2_fill_1 FILLER_45_895 ();
 sg13g2_fill_2 FILLER_45_932 ();
 sg13g2_fill_2 FILLER_45_1023 ();
 sg13g2_fill_2 FILLER_45_1035 ();
 sg13g2_fill_2 FILLER_45_1099 ();
 sg13g2_fill_1 FILLER_45_1101 ();
 sg13g2_fill_2 FILLER_45_1111 ();
 sg13g2_fill_1 FILLER_45_1123 ();
 sg13g2_fill_2 FILLER_45_1135 ();
 sg13g2_decap_4 FILLER_45_1154 ();
 sg13g2_fill_2 FILLER_45_1167 ();
 sg13g2_fill_1 FILLER_45_1169 ();
 sg13g2_fill_2 FILLER_45_1178 ();
 sg13g2_fill_1 FILLER_45_1180 ();
 sg13g2_decap_8 FILLER_45_1185 ();
 sg13g2_decap_8 FILLER_45_1192 ();
 sg13g2_fill_1 FILLER_45_1199 ();
 sg13g2_fill_2 FILLER_45_1204 ();
 sg13g2_fill_2 FILLER_45_1237 ();
 sg13g2_fill_2 FILLER_45_1265 ();
 sg13g2_fill_2 FILLER_45_1289 ();
 sg13g2_fill_2 FILLER_45_1304 ();
 sg13g2_fill_2 FILLER_45_1311 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_fill_1 FILLER_45_1329 ();
 sg13g2_fill_1 FILLER_45_1342 ();
 sg13g2_fill_2 FILLER_45_1360 ();
 sg13g2_fill_1 FILLER_45_1369 ();
 sg13g2_fill_1 FILLER_45_1418 ();
 sg13g2_fill_1 FILLER_45_1442 ();
 sg13g2_fill_1 FILLER_45_1464 ();
 sg13g2_fill_2 FILLER_45_1488 ();
 sg13g2_decap_8 FILLER_45_1494 ();
 sg13g2_fill_2 FILLER_45_1501 ();
 sg13g2_fill_2 FILLER_45_1530 ();
 sg13g2_fill_1 FILLER_45_1546 ();
 sg13g2_fill_1 FILLER_45_1560 ();
 sg13g2_fill_2 FILLER_45_1639 ();
 sg13g2_fill_2 FILLER_45_1648 ();
 sg13g2_fill_2 FILLER_45_1664 ();
 sg13g2_fill_1 FILLER_45_1666 ();
 sg13g2_fill_2 FILLER_45_1696 ();
 sg13g2_decap_8 FILLER_45_1702 ();
 sg13g2_decap_8 FILLER_45_1709 ();
 sg13g2_decap_8 FILLER_45_1716 ();
 sg13g2_decap_4 FILLER_45_1723 ();
 sg13g2_fill_2 FILLER_45_1727 ();
 sg13g2_decap_4 FILLER_45_1746 ();
 sg13g2_decap_8 FILLER_45_1807 ();
 sg13g2_decap_4 FILLER_45_1814 ();
 sg13g2_decap_8 FILLER_45_1825 ();
 sg13g2_decap_8 FILLER_45_1832 ();
 sg13g2_decap_8 FILLER_45_1869 ();
 sg13g2_decap_8 FILLER_45_1876 ();
 sg13g2_decap_8 FILLER_45_1883 ();
 sg13g2_decap_8 FILLER_45_1890 ();
 sg13g2_decap_8 FILLER_45_1897 ();
 sg13g2_decap_8 FILLER_45_1904 ();
 sg13g2_fill_2 FILLER_45_1911 ();
 sg13g2_fill_1 FILLER_45_1913 ();
 sg13g2_decap_4 FILLER_45_1923 ();
 sg13g2_fill_1 FILLER_45_1931 ();
 sg13g2_decap_8 FILLER_45_1937 ();
 sg13g2_decap_4 FILLER_45_1944 ();
 sg13g2_fill_2 FILLER_45_1948 ();
 sg13g2_decap_8 FILLER_45_1955 ();
 sg13g2_decap_8 FILLER_45_1962 ();
 sg13g2_decap_8 FILLER_45_1969 ();
 sg13g2_decap_8 FILLER_45_1976 ();
 sg13g2_decap_8 FILLER_45_1983 ();
 sg13g2_decap_8 FILLER_45_1990 ();
 sg13g2_fill_1 FILLER_45_1997 ();
 sg13g2_decap_8 FILLER_45_2018 ();
 sg13g2_decap_8 FILLER_45_2025 ();
 sg13g2_decap_8 FILLER_45_2032 ();
 sg13g2_decap_8 FILLER_45_2039 ();
 sg13g2_decap_8 FILLER_45_2046 ();
 sg13g2_decap_8 FILLER_45_2053 ();
 sg13g2_fill_2 FILLER_45_2060 ();
 sg13g2_fill_1 FILLER_45_2062 ();
 sg13g2_fill_1 FILLER_45_2089 ();
 sg13g2_fill_1 FILLER_45_2116 ();
 sg13g2_fill_1 FILLER_45_2122 ();
 sg13g2_fill_2 FILLER_45_2127 ();
 sg13g2_fill_1 FILLER_45_2181 ();
 sg13g2_fill_2 FILLER_45_2190 ();
 sg13g2_fill_1 FILLER_45_2192 ();
 sg13g2_fill_2 FILLER_45_2227 ();
 sg13g2_fill_1 FILLER_45_2229 ();
 sg13g2_fill_1 FILLER_45_2297 ();
 sg13g2_fill_2 FILLER_45_2306 ();
 sg13g2_fill_1 FILLER_45_2308 ();
 sg13g2_fill_1 FILLER_45_2313 ();
 sg13g2_fill_1 FILLER_45_2339 ();
 sg13g2_fill_1 FILLER_45_2351 ();
 sg13g2_fill_2 FILLER_45_2382 ();
 sg13g2_decap_4 FILLER_45_2394 ();
 sg13g2_fill_1 FILLER_45_2398 ();
 sg13g2_fill_2 FILLER_45_2416 ();
 sg13g2_fill_1 FILLER_45_2423 ();
 sg13g2_decap_4 FILLER_45_2429 ();
 sg13g2_fill_2 FILLER_45_2433 ();
 sg13g2_fill_1 FILLER_45_2446 ();
 sg13g2_fill_1 FILLER_45_2483 ();
 sg13g2_fill_2 FILLER_45_2514 ();
 sg13g2_fill_1 FILLER_45_2516 ();
 sg13g2_fill_2 FILLER_45_2543 ();
 sg13g2_fill_2 FILLER_45_2561 ();
 sg13g2_fill_2 FILLER_45_2569 ();
 sg13g2_fill_2 FILLER_45_2583 ();
 sg13g2_decap_4 FILLER_45_2607 ();
 sg13g2_fill_2 FILLER_45_2637 ();
 sg13g2_decap_8 FILLER_45_2643 ();
 sg13g2_decap_8 FILLER_45_2650 ();
 sg13g2_decap_8 FILLER_45_2657 ();
 sg13g2_decap_4 FILLER_45_2664 ();
 sg13g2_fill_2 FILLER_45_2668 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_38 ();
 sg13g2_decap_4 FILLER_46_44 ();
 sg13g2_fill_1 FILLER_46_71 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_118 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_293 ();
 sg13g2_fill_1 FILLER_46_305 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_4 FILLER_46_393 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_46_409 ();
 sg13g2_fill_1 FILLER_46_416 ();
 sg13g2_fill_1 FILLER_46_422 ();
 sg13g2_decap_8 FILLER_46_453 ();
 sg13g2_fill_2 FILLER_46_460 ();
 sg13g2_fill_1 FILLER_46_462 ();
 sg13g2_fill_1 FILLER_46_489 ();
 sg13g2_fill_1 FILLER_46_554 ();
 sg13g2_fill_2 FILLER_46_560 ();
 sg13g2_fill_1 FILLER_46_562 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_fill_1 FILLER_46_607 ();
 sg13g2_decap_4 FILLER_46_611 ();
 sg13g2_fill_2 FILLER_46_615 ();
 sg13g2_decap_4 FILLER_46_621 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_1 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_1 FILLER_46_698 ();
 sg13g2_fill_1 FILLER_46_705 ();
 sg13g2_fill_1 FILLER_46_768 ();
 sg13g2_fill_1 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_fill_2 FILLER_46_825 ();
 sg13g2_fill_2 FILLER_46_831 ();
 sg13g2_decap_4 FILLER_46_859 ();
 sg13g2_fill_2 FILLER_46_893 ();
 sg13g2_fill_1 FILLER_46_956 ();
 sg13g2_fill_1 FILLER_46_1023 ();
 sg13g2_fill_1 FILLER_46_1029 ();
 sg13g2_fill_2 FILLER_46_1042 ();
 sg13g2_fill_1 FILLER_46_1048 ();
 sg13g2_fill_2 FILLER_46_1088 ();
 sg13g2_fill_1 FILLER_46_1123 ();
 sg13g2_fill_2 FILLER_46_1156 ();
 sg13g2_fill_1 FILLER_46_1166 ();
 sg13g2_fill_2 FILLER_46_1172 ();
 sg13g2_decap_4 FILLER_46_1194 ();
 sg13g2_fill_1 FILLER_46_1198 ();
 sg13g2_decap_4 FILLER_46_1203 ();
 sg13g2_fill_1 FILLER_46_1207 ();
 sg13g2_fill_1 FILLER_46_1287 ();
 sg13g2_fill_2 FILLER_46_1306 ();
 sg13g2_fill_2 FILLER_46_1333 ();
 sg13g2_fill_2 FILLER_46_1364 ();
 sg13g2_fill_1 FILLER_46_1396 ();
 sg13g2_fill_1 FILLER_46_1442 ();
 sg13g2_fill_2 FILLER_46_1466 ();
 sg13g2_decap_4 FILLER_46_1486 ();
 sg13g2_fill_1 FILLER_46_1490 ();
 sg13g2_fill_1 FILLER_46_1501 ();
 sg13g2_fill_1 FILLER_46_1542 ();
 sg13g2_decap_8 FILLER_46_1655 ();
 sg13g2_decap_8 FILLER_46_1662 ();
 sg13g2_decap_4 FILLER_46_1669 ();
 sg13g2_decap_4 FILLER_46_1699 ();
 sg13g2_decap_8 FILLER_46_1716 ();
 sg13g2_decap_8 FILLER_46_1723 ();
 sg13g2_decap_8 FILLER_46_1730 ();
 sg13g2_decap_8 FILLER_46_1737 ();
 sg13g2_decap_4 FILLER_46_1744 ();
 sg13g2_fill_1 FILLER_46_1748 ();
 sg13g2_fill_2 FILLER_46_1815 ();
 sg13g2_decap_8 FILLER_46_1852 ();
 sg13g2_decap_8 FILLER_46_1859 ();
 sg13g2_fill_1 FILLER_46_1866 ();
 sg13g2_decap_8 FILLER_46_1872 ();
 sg13g2_decap_8 FILLER_46_1879 ();
 sg13g2_decap_8 FILLER_46_1886 ();
 sg13g2_decap_8 FILLER_46_1893 ();
 sg13g2_decap_8 FILLER_46_1900 ();
 sg13g2_decap_8 FILLER_46_1907 ();
 sg13g2_decap_8 FILLER_46_1914 ();
 sg13g2_decap_8 FILLER_46_1921 ();
 sg13g2_decap_8 FILLER_46_1928 ();
 sg13g2_decap_8 FILLER_46_1935 ();
 sg13g2_decap_4 FILLER_46_1942 ();
 sg13g2_fill_2 FILLER_46_1946 ();
 sg13g2_decap_8 FILLER_46_1952 ();
 sg13g2_fill_1 FILLER_46_1959 ();
 sg13g2_fill_2 FILLER_46_1966 ();
 sg13g2_decap_8 FILLER_46_1972 ();
 sg13g2_decap_8 FILLER_46_1979 ();
 sg13g2_decap_4 FILLER_46_1986 ();
 sg13g2_fill_1 FILLER_46_1990 ();
 sg13g2_decap_8 FILLER_46_1999 ();
 sg13g2_decap_8 FILLER_46_2006 ();
 sg13g2_decap_8 FILLER_46_2013 ();
 sg13g2_decap_8 FILLER_46_2020 ();
 sg13g2_decap_4 FILLER_46_2027 ();
 sg13g2_decap_8 FILLER_46_2034 ();
 sg13g2_decap_8 FILLER_46_2041 ();
 sg13g2_decap_8 FILLER_46_2048 ();
 sg13g2_decap_8 FILLER_46_2055 ();
 sg13g2_decap_8 FILLER_46_2062 ();
 sg13g2_decap_4 FILLER_46_2073 ();
 sg13g2_fill_1 FILLER_46_2103 ();
 sg13g2_fill_2 FILLER_46_2107 ();
 sg13g2_fill_1 FILLER_46_2109 ();
 sg13g2_fill_1 FILLER_46_2162 ();
 sg13g2_decap_4 FILLER_46_2167 ();
 sg13g2_fill_1 FILLER_46_2185 ();
 sg13g2_fill_1 FILLER_46_2261 ();
 sg13g2_decap_4 FILLER_46_2274 ();
 sg13g2_fill_1 FILLER_46_2278 ();
 sg13g2_decap_8 FILLER_46_2283 ();
 sg13g2_decap_4 FILLER_46_2290 ();
 sg13g2_fill_1 FILLER_46_2294 ();
 sg13g2_decap_4 FILLER_46_2321 ();
 sg13g2_fill_1 FILLER_46_2325 ();
 sg13g2_decap_8 FILLER_46_2362 ();
 sg13g2_fill_2 FILLER_46_2369 ();
 sg13g2_decap_8 FILLER_46_2443 ();
 sg13g2_decap_4 FILLER_46_2450 ();
 sg13g2_fill_1 FILLER_46_2454 ();
 sg13g2_fill_1 FILLER_46_2464 ();
 sg13g2_decap_4 FILLER_46_2469 ();
 sg13g2_fill_1 FILLER_46_2473 ();
 sg13g2_fill_1 FILLER_46_2484 ();
 sg13g2_fill_1 FILLER_46_2492 ();
 sg13g2_fill_2 FILLER_46_2572 ();
 sg13g2_fill_1 FILLER_46_2574 ();
 sg13g2_decap_8 FILLER_46_2579 ();
 sg13g2_fill_1 FILLER_46_2586 ();
 sg13g2_fill_1 FILLER_46_2612 ();
 sg13g2_fill_1 FILLER_46_2639 ();
 sg13g2_decap_8 FILLER_46_2644 ();
 sg13g2_decap_8 FILLER_46_2651 ();
 sg13g2_decap_8 FILLER_46_2658 ();
 sg13g2_decap_4 FILLER_46_2665 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_55 ();
 sg13g2_fill_1 FILLER_47_66 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_125 ();
 sg13g2_fill_1 FILLER_47_152 ();
 sg13g2_fill_2 FILLER_47_167 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_fill_2 FILLER_47_174 ();
 sg13g2_fill_1 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_198 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_252 ();
 sg13g2_fill_1 FILLER_47_280 ();
 sg13g2_fill_2 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_306 ();
 sg13g2_fill_1 FILLER_47_362 ();
 sg13g2_fill_1 FILLER_47_404 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_419 ();
 sg13g2_fill_1 FILLER_47_426 ();
 sg13g2_fill_1 FILLER_47_431 ();
 sg13g2_decap_8 FILLER_47_443 ();
 sg13g2_decap_8 FILLER_47_450 ();
 sg13g2_decap_4 FILLER_47_457 ();
 sg13g2_fill_1 FILLER_47_461 ();
 sg13g2_fill_2 FILLER_47_466 ();
 sg13g2_fill_1 FILLER_47_468 ();
 sg13g2_decap_8 FILLER_47_473 ();
 sg13g2_fill_1 FILLER_47_480 ();
 sg13g2_fill_2 FILLER_47_512 ();
 sg13g2_fill_1 FILLER_47_539 ();
 sg13g2_fill_1 FILLER_47_545 ();
 sg13g2_fill_2 FILLER_47_555 ();
 sg13g2_decap_4 FILLER_47_562 ();
 sg13g2_fill_1 FILLER_47_581 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_decap_4 FILLER_47_622 ();
 sg13g2_fill_2 FILLER_47_626 ();
 sg13g2_fill_1 FILLER_47_637 ();
 sg13g2_fill_1 FILLER_47_653 ();
 sg13g2_fill_2 FILLER_47_710 ();
 sg13g2_fill_1 FILLER_47_736 ();
 sg13g2_fill_1 FILLER_47_769 ();
 sg13g2_fill_1 FILLER_47_775 ();
 sg13g2_fill_1 FILLER_47_787 ();
 sg13g2_decap_4 FILLER_47_795 ();
 sg13g2_fill_2 FILLER_47_799 ();
 sg13g2_decap_4 FILLER_47_805 ();
 sg13g2_fill_1 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_4 FILLER_47_883 ();
 sg13g2_fill_1 FILLER_47_887 ();
 sg13g2_decap_4 FILLER_47_892 ();
 sg13g2_fill_2 FILLER_47_906 ();
 sg13g2_fill_2 FILLER_47_917 ();
 sg13g2_fill_1 FILLER_47_919 ();
 sg13g2_fill_2 FILLER_47_960 ();
 sg13g2_fill_2 FILLER_47_1002 ();
 sg13g2_fill_1 FILLER_47_1004 ();
 sg13g2_fill_1 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_47_1034 ();
 sg13g2_decap_4 FILLER_47_1041 ();
 sg13g2_fill_1 FILLER_47_1045 ();
 sg13g2_fill_2 FILLER_47_1182 ();
 sg13g2_fill_1 FILLER_47_1184 ();
 sg13g2_fill_1 FILLER_47_1189 ();
 sg13g2_fill_2 FILLER_47_1194 ();
 sg13g2_fill_1 FILLER_47_1196 ();
 sg13g2_fill_2 FILLER_47_1223 ();
 sg13g2_fill_2 FILLER_47_1229 ();
 sg13g2_fill_2 FILLER_47_1267 ();
 sg13g2_fill_2 FILLER_47_1276 ();
 sg13g2_fill_2 FILLER_47_1294 ();
 sg13g2_fill_2 FILLER_47_1303 ();
 sg13g2_fill_1 FILLER_47_1308 ();
 sg13g2_fill_1 FILLER_47_1315 ();
 sg13g2_fill_1 FILLER_47_1321 ();
 sg13g2_fill_2 FILLER_47_1343 ();
 sg13g2_fill_2 FILLER_47_1402 ();
 sg13g2_fill_2 FILLER_47_1410 ();
 sg13g2_fill_2 FILLER_47_1431 ();
 sg13g2_fill_2 FILLER_47_1447 ();
 sg13g2_fill_2 FILLER_47_1494 ();
 sg13g2_fill_1 FILLER_47_1496 ();
 sg13g2_fill_2 FILLER_47_1540 ();
 sg13g2_fill_1 FILLER_47_1554 ();
 sg13g2_fill_1 FILLER_47_1572 ();
 sg13g2_fill_2 FILLER_47_1578 ();
 sg13g2_fill_2 FILLER_47_1626 ();
 sg13g2_fill_1 FILLER_47_1670 ();
 sg13g2_fill_2 FILLER_47_1675 ();
 sg13g2_decap_8 FILLER_47_1682 ();
 sg13g2_fill_2 FILLER_47_1689 ();
 sg13g2_decap_8 FILLER_47_1702 ();
 sg13g2_decap_8 FILLER_47_1714 ();
 sg13g2_fill_2 FILLER_47_1721 ();
 sg13g2_fill_1 FILLER_47_1723 ();
 sg13g2_decap_8 FILLER_47_1728 ();
 sg13g2_decap_8 FILLER_47_1735 ();
 sg13g2_decap_8 FILLER_47_1742 ();
 sg13g2_decap_4 FILLER_47_1749 ();
 sg13g2_fill_2 FILLER_47_1757 ();
 sg13g2_fill_1 FILLER_47_1759 ();
 sg13g2_decap_4 FILLER_47_1816 ();
 sg13g2_fill_2 FILLER_47_1825 ();
 sg13g2_decap_8 FILLER_47_1835 ();
 sg13g2_decap_4 FILLER_47_1842 ();
 sg13g2_fill_1 FILLER_47_1846 ();
 sg13g2_decap_4 FILLER_47_1852 ();
 sg13g2_fill_1 FILLER_47_1856 ();
 sg13g2_decap_8 FILLER_47_1861 ();
 sg13g2_decap_8 FILLER_47_1868 ();
 sg13g2_decap_8 FILLER_47_1875 ();
 sg13g2_decap_8 FILLER_47_1882 ();
 sg13g2_decap_4 FILLER_47_1889 ();
 sg13g2_fill_2 FILLER_47_1893 ();
 sg13g2_decap_8 FILLER_47_1899 ();
 sg13g2_decap_8 FILLER_47_1906 ();
 sg13g2_decap_8 FILLER_47_1913 ();
 sg13g2_decap_8 FILLER_47_1920 ();
 sg13g2_decap_4 FILLER_47_1927 ();
 sg13g2_decap_8 FILLER_47_1935 ();
 sg13g2_decap_8 FILLER_47_1942 ();
 sg13g2_decap_8 FILLER_47_1949 ();
 sg13g2_decap_8 FILLER_47_1956 ();
 sg13g2_decap_8 FILLER_47_1963 ();
 sg13g2_decap_8 FILLER_47_1970 ();
 sg13g2_decap_8 FILLER_47_1977 ();
 sg13g2_decap_8 FILLER_47_1984 ();
 sg13g2_decap_8 FILLER_47_1991 ();
 sg13g2_decap_8 FILLER_47_1998 ();
 sg13g2_decap_8 FILLER_47_2005 ();
 sg13g2_decap_8 FILLER_47_2012 ();
 sg13g2_decap_8 FILLER_47_2019 ();
 sg13g2_decap_4 FILLER_47_2026 ();
 sg13g2_fill_1 FILLER_47_2030 ();
 sg13g2_decap_8 FILLER_47_2034 ();
 sg13g2_decap_8 FILLER_47_2041 ();
 sg13g2_decap_8 FILLER_47_2048 ();
 sg13g2_decap_8 FILLER_47_2055 ();
 sg13g2_decap_8 FILLER_47_2062 ();
 sg13g2_decap_8 FILLER_47_2069 ();
 sg13g2_fill_2 FILLER_47_2076 ();
 sg13g2_fill_2 FILLER_47_2087 ();
 sg13g2_fill_2 FILLER_47_2098 ();
 sg13g2_fill_1 FILLER_47_2100 ();
 sg13g2_decap_4 FILLER_47_2133 ();
 sg13g2_fill_1 FILLER_47_2137 ();
 sg13g2_fill_2 FILLER_47_2142 ();
 sg13g2_fill_1 FILLER_47_2162 ();
 sg13g2_fill_1 FILLER_47_2168 ();
 sg13g2_fill_2 FILLER_47_2173 ();
 sg13g2_fill_1 FILLER_47_2175 ();
 sg13g2_decap_8 FILLER_47_2185 ();
 sg13g2_decap_4 FILLER_47_2192 ();
 sg13g2_fill_1 FILLER_47_2196 ();
 sg13g2_fill_1 FILLER_47_2240 ();
 sg13g2_fill_1 FILLER_47_2246 ();
 sg13g2_fill_1 FILLER_47_2252 ();
 sg13g2_decap_4 FILLER_47_2292 ();
 sg13g2_fill_1 FILLER_47_2296 ();
 sg13g2_decap_4 FILLER_47_2301 ();
 sg13g2_fill_2 FILLER_47_2305 ();
 sg13g2_fill_1 FILLER_47_2342 ();
 sg13g2_decap_8 FILLER_47_2347 ();
 sg13g2_decap_8 FILLER_47_2354 ();
 sg13g2_decap_4 FILLER_47_2361 ();
 sg13g2_fill_2 FILLER_47_2365 ();
 sg13g2_fill_1 FILLER_47_2370 ();
 sg13g2_fill_1 FILLER_47_2381 ();
 sg13g2_fill_2 FILLER_47_2448 ();
 sg13g2_fill_2 FILLER_47_2460 ();
 sg13g2_decap_4 FILLER_47_2472 ();
 sg13g2_fill_1 FILLER_47_2495 ();
 sg13g2_fill_1 FILLER_47_2506 ();
 sg13g2_fill_1 FILLER_47_2517 ();
 sg13g2_fill_1 FILLER_47_2524 ();
 sg13g2_decap_4 FILLER_47_2545 ();
 sg13g2_fill_2 FILLER_47_2553 ();
 sg13g2_fill_1 FILLER_47_2555 ();
 sg13g2_fill_2 FILLER_47_2565 ();
 sg13g2_fill_1 FILLER_47_2567 ();
 sg13g2_decap_4 FILLER_47_2577 ();
 sg13g2_fill_2 FILLER_47_2581 ();
 sg13g2_decap_4 FILLER_47_2588 ();
 sg13g2_decap_4 FILLER_47_2601 ();
 sg13g2_fill_1 FILLER_47_2605 ();
 sg13g2_fill_1 FILLER_47_2616 ();
 sg13g2_decap_8 FILLER_47_2643 ();
 sg13g2_decap_8 FILLER_47_2650 ();
 sg13g2_decap_8 FILLER_47_2657 ();
 sg13g2_decap_4 FILLER_47_2664 ();
 sg13g2_fill_2 FILLER_47_2668 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_76 ();
 sg13g2_fill_2 FILLER_48_88 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_decap_8 FILLER_48_118 ();
 sg13g2_fill_2 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_decap_8 FILLER_48_181 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_decap_8 FILLER_48_195 ();
 sg13g2_decap_8 FILLER_48_202 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_252 ();
 sg13g2_fill_1 FILLER_48_374 ();
 sg13g2_fill_2 FILLER_48_400 ();
 sg13g2_decap_4 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_411 ();
 sg13g2_decap_8 FILLER_48_443 ();
 sg13g2_fill_2 FILLER_48_481 ();
 sg13g2_fill_1 FILLER_48_483 ();
 sg13g2_decap_4 FILLER_48_509 ();
 sg13g2_fill_2 FILLER_48_513 ();
 sg13g2_fill_2 FILLER_48_520 ();
 sg13g2_fill_1 FILLER_48_522 ();
 sg13g2_fill_1 FILLER_48_549 ();
 sg13g2_fill_1 FILLER_48_555 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_fill_2 FILLER_48_567 ();
 sg13g2_decap_4 FILLER_48_578 ();
 sg13g2_fill_1 FILLER_48_582 ();
 sg13g2_decap_4 FILLER_48_588 ();
 sg13g2_fill_1 FILLER_48_597 ();
 sg13g2_fill_1 FILLER_48_602 ();
 sg13g2_fill_1 FILLER_48_613 ();
 sg13g2_fill_2 FILLER_48_619 ();
 sg13g2_fill_2 FILLER_48_626 ();
 sg13g2_decap_4 FILLER_48_632 ();
 sg13g2_fill_2 FILLER_48_636 ();
 sg13g2_fill_2 FILLER_48_666 ();
 sg13g2_fill_1 FILLER_48_687 ();
 sg13g2_fill_2 FILLER_48_701 ();
 sg13g2_fill_2 FILLER_48_708 ();
 sg13g2_fill_1 FILLER_48_714 ();
 sg13g2_fill_1 FILLER_48_754 ();
 sg13g2_fill_1 FILLER_48_766 ();
 sg13g2_fill_1 FILLER_48_787 ();
 sg13g2_fill_1 FILLER_48_797 ();
 sg13g2_decap_4 FILLER_48_802 ();
 sg13g2_decap_4 FILLER_48_814 ();
 sg13g2_decap_4 FILLER_48_823 ();
 sg13g2_fill_1 FILLER_48_827 ();
 sg13g2_decap_4 FILLER_48_838 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_fill_2 FILLER_48_849 ();
 sg13g2_fill_1 FILLER_48_881 ();
 sg13g2_decap_4 FILLER_48_887 ();
 sg13g2_decap_8 FILLER_48_909 ();
 sg13g2_fill_2 FILLER_48_916 ();
 sg13g2_fill_1 FILLER_48_918 ();
 sg13g2_decap_4 FILLER_48_923 ();
 sg13g2_fill_1 FILLER_48_927 ();
 sg13g2_fill_2 FILLER_48_937 ();
 sg13g2_fill_1 FILLER_48_942 ();
 sg13g2_decap_4 FILLER_48_948 ();
 sg13g2_fill_2 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_fill_2 FILLER_48_974 ();
 sg13g2_decap_4 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_1004 ();
 sg13g2_decap_8 FILLER_48_1020 ();
 sg13g2_decap_4 FILLER_48_1027 ();
 sg13g2_fill_2 FILLER_48_1031 ();
 sg13g2_fill_1 FILLER_48_1083 ();
 sg13g2_fill_2 FILLER_48_1103 ();
 sg13g2_fill_2 FILLER_48_1119 ();
 sg13g2_fill_2 FILLER_48_1131 ();
 sg13g2_fill_2 FILLER_48_1164 ();
 sg13g2_fill_2 FILLER_48_1172 ();
 sg13g2_fill_1 FILLER_48_1174 ();
 sg13g2_fill_1 FILLER_48_1179 ();
 sg13g2_fill_1 FILLER_48_1195 ();
 sg13g2_fill_2 FILLER_48_1248 ();
 sg13g2_fill_1 FILLER_48_1280 ();
 sg13g2_fill_1 FILLER_48_1299 ();
 sg13g2_fill_1 FILLER_48_1331 ();
 sg13g2_fill_2 FILLER_48_1355 ();
 sg13g2_fill_1 FILLER_48_1375 ();
 sg13g2_fill_2 FILLER_48_1387 ();
 sg13g2_fill_1 FILLER_48_1410 ();
 sg13g2_fill_1 FILLER_48_1415 ();
 sg13g2_fill_1 FILLER_48_1421 ();
 sg13g2_fill_1 FILLER_48_1429 ();
 sg13g2_fill_1 FILLER_48_1435 ();
 sg13g2_fill_2 FILLER_48_1446 ();
 sg13g2_fill_2 FILLER_48_1472 ();
 sg13g2_fill_1 FILLER_48_1474 ();
 sg13g2_fill_1 FILLER_48_1520 ();
 sg13g2_fill_2 FILLER_48_1525 ();
 sg13g2_fill_2 FILLER_48_1554 ();
 sg13g2_fill_2 FILLER_48_1577 ();
 sg13g2_fill_1 FILLER_48_1584 ();
 sg13g2_decap_8 FILLER_48_1605 ();
 sg13g2_decap_4 FILLER_48_1612 ();
 sg13g2_fill_1 FILLER_48_1616 ();
 sg13g2_fill_1 FILLER_48_1626 ();
 sg13g2_decap_4 FILLER_48_1667 ();
 sg13g2_fill_2 FILLER_48_1710 ();
 sg13g2_fill_2 FILLER_48_1719 ();
 sg13g2_fill_1 FILLER_48_1721 ();
 sg13g2_fill_1 FILLER_48_1727 ();
 sg13g2_decap_4 FILLER_48_1733 ();
 sg13g2_fill_2 FILLER_48_1737 ();
 sg13g2_fill_1 FILLER_48_1750 ();
 sg13g2_decap_8 FILLER_48_1758 ();
 sg13g2_decap_8 FILLER_48_1769 ();
 sg13g2_fill_2 FILLER_48_1776 ();
 sg13g2_fill_1 FILLER_48_1778 ();
 sg13g2_fill_1 FILLER_48_1783 ();
 sg13g2_fill_2 FILLER_48_1788 ();
 sg13g2_fill_1 FILLER_48_1790 ();
 sg13g2_decap_8 FILLER_48_1803 ();
 sg13g2_fill_2 FILLER_48_1810 ();
 sg13g2_fill_1 FILLER_48_1812 ();
 sg13g2_decap_4 FILLER_48_1817 ();
 sg13g2_decap_8 FILLER_48_1873 ();
 sg13g2_decap_8 FILLER_48_1880 ();
 sg13g2_decap_8 FILLER_48_1887 ();
 sg13g2_decap_8 FILLER_48_1894 ();
 sg13g2_fill_2 FILLER_48_1901 ();
 sg13g2_fill_1 FILLER_48_1903 ();
 sg13g2_decap_4 FILLER_48_1908 ();
 sg13g2_fill_2 FILLER_48_1912 ();
 sg13g2_fill_1 FILLER_48_1918 ();
 sg13g2_decap_8 FILLER_48_1938 ();
 sg13g2_decap_8 FILLER_48_1945 ();
 sg13g2_fill_2 FILLER_48_1952 ();
 sg13g2_fill_1 FILLER_48_1954 ();
 sg13g2_decap_8 FILLER_48_1959 ();
 sg13g2_decap_8 FILLER_48_1966 ();
 sg13g2_decap_8 FILLER_48_1973 ();
 sg13g2_decap_8 FILLER_48_1980 ();
 sg13g2_decap_8 FILLER_48_1987 ();
 sg13g2_fill_2 FILLER_48_1994 ();
 sg13g2_fill_1 FILLER_48_1996 ();
 sg13g2_decap_8 FILLER_48_2002 ();
 sg13g2_fill_1 FILLER_48_2009 ();
 sg13g2_decap_8 FILLER_48_2022 ();
 sg13g2_decap_8 FILLER_48_2029 ();
 sg13g2_decap_8 FILLER_48_2036 ();
 sg13g2_decap_8 FILLER_48_2043 ();
 sg13g2_decap_8 FILLER_48_2050 ();
 sg13g2_decap_8 FILLER_48_2057 ();
 sg13g2_decap_8 FILLER_48_2064 ();
 sg13g2_decap_8 FILLER_48_2071 ();
 sg13g2_decap_8 FILLER_48_2078 ();
 sg13g2_decap_4 FILLER_48_2085 ();
 sg13g2_fill_1 FILLER_48_2089 ();
 sg13g2_decap_4 FILLER_48_2125 ();
 sg13g2_fill_1 FILLER_48_2129 ();
 sg13g2_fill_1 FILLER_48_2135 ();
 sg13g2_fill_2 FILLER_48_2183 ();
 sg13g2_fill_2 FILLER_48_2195 ();
 sg13g2_decap_4 FILLER_48_2206 ();
 sg13g2_fill_1 FILLER_48_2210 ();
 sg13g2_fill_2 FILLER_48_2229 ();
 sg13g2_fill_1 FILLER_48_2249 ();
 sg13g2_fill_2 FILLER_48_2263 ();
 sg13g2_decap_8 FILLER_48_2270 ();
 sg13g2_decap_8 FILLER_48_2281 ();
 sg13g2_decap_8 FILLER_48_2288 ();
 sg13g2_fill_2 FILLER_48_2295 ();
 sg13g2_fill_1 FILLER_48_2297 ();
 sg13g2_fill_2 FILLER_48_2302 ();
 sg13g2_fill_1 FILLER_48_2332 ();
 sg13g2_fill_1 FILLER_48_2371 ();
 sg13g2_fill_2 FILLER_48_2395 ();
 sg13g2_decap_4 FILLER_48_2418 ();
 sg13g2_decap_4 FILLER_48_2426 ();
 sg13g2_fill_1 FILLER_48_2474 ();
 sg13g2_decap_4 FILLER_48_2481 ();
 sg13g2_fill_1 FILLER_48_2485 ();
 sg13g2_fill_1 FILLER_48_2534 ();
 sg13g2_decap_8 FILLER_48_2569 ();
 sg13g2_decap_8 FILLER_48_2576 ();
 sg13g2_fill_1 FILLER_48_2583 ();
 sg13g2_decap_4 FILLER_48_2613 ();
 sg13g2_fill_1 FILLER_48_2617 ();
 sg13g2_decap_8 FILLER_48_2644 ();
 sg13g2_decap_8 FILLER_48_2651 ();
 sg13g2_decap_8 FILLER_48_2658 ();
 sg13g2_decap_4 FILLER_48_2665 ();
 sg13g2_fill_1 FILLER_48_2669 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_92 ();
 sg13g2_fill_2 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_121 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_decap_8 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_153 ();
 sg13g2_decap_4 FILLER_49_160 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_8 FILLER_49_178 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_decap_4 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_229 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_fill_2 FILLER_49_424 ();
 sg13g2_fill_1 FILLER_49_426 ();
 sg13g2_fill_2 FILLER_49_453 ();
 sg13g2_fill_1 FILLER_49_460 ();
 sg13g2_fill_2 FILLER_49_487 ();
 sg13g2_fill_1 FILLER_49_511 ();
 sg13g2_fill_2 FILLER_49_517 ();
 sg13g2_decap_4 FILLER_49_568 ();
 sg13g2_decap_8 FILLER_49_576 ();
 sg13g2_decap_4 FILLER_49_583 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_654 ();
 sg13g2_fill_2 FILLER_49_664 ();
 sg13g2_fill_1 FILLER_49_712 ();
 sg13g2_fill_1 FILLER_49_722 ();
 sg13g2_fill_1 FILLER_49_732 ();
 sg13g2_fill_1 FILLER_49_762 ();
 sg13g2_fill_2 FILLER_49_786 ();
 sg13g2_fill_2 FILLER_49_793 ();
 sg13g2_fill_2 FILLER_49_823 ();
 sg13g2_fill_1 FILLER_49_829 ();
 sg13g2_fill_2 FILLER_49_844 ();
 sg13g2_fill_1 FILLER_49_846 ();
 sg13g2_fill_1 FILLER_49_865 ();
 sg13g2_fill_1 FILLER_49_892 ();
 sg13g2_fill_1 FILLER_49_898 ();
 sg13g2_fill_1 FILLER_49_904 ();
 sg13g2_fill_1 FILLER_49_909 ();
 sg13g2_fill_1 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_921 ();
 sg13g2_decap_8 FILLER_49_932 ();
 sg13g2_decap_8 FILLER_49_939 ();
 sg13g2_decap_8 FILLER_49_946 ();
 sg13g2_decap_8 FILLER_49_953 ();
 sg13g2_decap_4 FILLER_49_960 ();
 sg13g2_fill_2 FILLER_49_973 ();
 sg13g2_fill_1 FILLER_49_975 ();
 sg13g2_decap_8 FILLER_49_981 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_fill_1 FILLER_49_1067 ();
 sg13g2_decap_8 FILLER_49_1072 ();
 sg13g2_decap_4 FILLER_49_1079 ();
 sg13g2_fill_2 FILLER_49_1096 ();
 sg13g2_fill_2 FILLER_49_1108 ();
 sg13g2_fill_1 FILLER_49_1180 ();
 sg13g2_fill_2 FILLER_49_1219 ();
 sg13g2_fill_1 FILLER_49_1326 ();
 sg13g2_fill_1 FILLER_49_1331 ();
 sg13g2_fill_1 FILLER_49_1432 ();
 sg13g2_fill_1 FILLER_49_1443 ();
 sg13g2_fill_2 FILLER_49_1448 ();
 sg13g2_fill_2 FILLER_49_1494 ();
 sg13g2_fill_1 FILLER_49_1513 ();
 sg13g2_fill_1 FILLER_49_1519 ();
 sg13g2_fill_1 FILLER_49_1527 ();
 sg13g2_fill_1 FILLER_49_1531 ();
 sg13g2_fill_1 FILLER_49_1559 ();
 sg13g2_fill_1 FILLER_49_1601 ();
 sg13g2_decap_8 FILLER_49_1612 ();
 sg13g2_decap_8 FILLER_49_1619 ();
 sg13g2_decap_4 FILLER_49_1626 ();
 sg13g2_fill_2 FILLER_49_1630 ();
 sg13g2_fill_2 FILLER_49_1681 ();
 sg13g2_fill_2 FILLER_49_1708 ();
 sg13g2_fill_1 FILLER_49_1710 ();
 sg13g2_decap_4 FILLER_49_1720 ();
 sg13g2_fill_2 FILLER_49_1728 ();
 sg13g2_fill_2 FILLER_49_1735 ();
 sg13g2_fill_1 FILLER_49_1741 ();
 sg13g2_fill_1 FILLER_49_1746 ();
 sg13g2_fill_1 FILLER_49_1755 ();
 sg13g2_decap_4 FILLER_49_1764 ();
 sg13g2_fill_2 FILLER_49_1768 ();
 sg13g2_decap_8 FILLER_49_1775 ();
 sg13g2_decap_4 FILLER_49_1787 ();
 sg13g2_fill_1 FILLER_49_1791 ();
 sg13g2_decap_4 FILLER_49_1796 ();
 sg13g2_fill_2 FILLER_49_1800 ();
 sg13g2_decap_4 FILLER_49_1806 ();
 sg13g2_fill_2 FILLER_49_1810 ();
 sg13g2_fill_1 FILLER_49_1817 ();
 sg13g2_decap_8 FILLER_49_1821 ();
 sg13g2_decap_8 FILLER_49_1832 ();
 sg13g2_decap_8 FILLER_49_1839 ();
 sg13g2_decap_8 FILLER_49_1846 ();
 sg13g2_fill_2 FILLER_49_1853 ();
 sg13g2_fill_1 FILLER_49_1855 ();
 sg13g2_decap_4 FILLER_49_1860 ();
 sg13g2_fill_1 FILLER_49_1864 ();
 sg13g2_decap_8 FILLER_49_1870 ();
 sg13g2_decap_4 FILLER_49_1877 ();
 sg13g2_decap_8 FILLER_49_1887 ();
 sg13g2_fill_1 FILLER_49_1900 ();
 sg13g2_decap_4 FILLER_49_1909 ();
 sg13g2_fill_2 FILLER_49_1913 ();
 sg13g2_decap_8 FILLER_49_1919 ();
 sg13g2_fill_2 FILLER_49_1926 ();
 sg13g2_decap_4 FILLER_49_1934 ();
 sg13g2_fill_1 FILLER_49_1938 ();
 sg13g2_decap_8 FILLER_49_1945 ();
 sg13g2_decap_8 FILLER_49_1952 ();
 sg13g2_fill_2 FILLER_49_1959 ();
 sg13g2_decap_8 FILLER_49_1966 ();
 sg13g2_decap_8 FILLER_49_1973 ();
 sg13g2_decap_8 FILLER_49_1980 ();
 sg13g2_decap_8 FILLER_49_1987 ();
 sg13g2_decap_8 FILLER_49_1994 ();
 sg13g2_decap_8 FILLER_49_2001 ();
 sg13g2_decap_8 FILLER_49_2008 ();
 sg13g2_decap_8 FILLER_49_2015 ();
 sg13g2_decap_8 FILLER_49_2022 ();
 sg13g2_decap_8 FILLER_49_2029 ();
 sg13g2_decap_8 FILLER_49_2036 ();
 sg13g2_decap_8 FILLER_49_2043 ();
 sg13g2_decap_8 FILLER_49_2050 ();
 sg13g2_decap_8 FILLER_49_2057 ();
 sg13g2_decap_8 FILLER_49_2064 ();
 sg13g2_decap_8 FILLER_49_2071 ();
 sg13g2_fill_1 FILLER_49_2078 ();
 sg13g2_fill_2 FILLER_49_2088 ();
 sg13g2_fill_1 FILLER_49_2090 ();
 sg13g2_fill_1 FILLER_49_2117 ();
 sg13g2_decap_4 FILLER_49_2148 ();
 sg13g2_fill_1 FILLER_49_2202 ();
 sg13g2_fill_2 FILLER_49_2229 ();
 sg13g2_decap_4 FILLER_49_2241 ();
 sg13g2_fill_1 FILLER_49_2261 ();
 sg13g2_fill_1 FILLER_49_2267 ();
 sg13g2_fill_1 FILLER_49_2274 ();
 sg13g2_fill_1 FILLER_49_2301 ();
 sg13g2_fill_1 FILLER_49_2307 ();
 sg13g2_fill_1 FILLER_49_2338 ();
 sg13g2_fill_1 FILLER_49_2349 ();
 sg13g2_fill_2 FILLER_49_2366 ();
 sg13g2_fill_1 FILLER_49_2368 ();
 sg13g2_fill_1 FILLER_49_2373 ();
 sg13g2_fill_1 FILLER_49_2410 ();
 sg13g2_decap_8 FILLER_49_2441 ();
 sg13g2_fill_2 FILLER_49_2474 ();
 sg13g2_fill_2 FILLER_49_2486 ();
 sg13g2_fill_2 FILLER_49_2498 ();
 sg13g2_fill_1 FILLER_49_2552 ();
 sg13g2_decap_4 FILLER_49_2603 ();
 sg13g2_fill_1 FILLER_49_2607 ();
 sg13g2_decap_8 FILLER_49_2640 ();
 sg13g2_decap_8 FILLER_49_2647 ();
 sg13g2_decap_8 FILLER_49_2654 ();
 sg13g2_decap_8 FILLER_49_2661 ();
 sg13g2_fill_2 FILLER_49_2668 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_11 ();
 sg13g2_fill_1 FILLER_50_16 ();
 sg13g2_fill_1 FILLER_50_22 ();
 sg13g2_fill_2 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_29 ();
 sg13g2_fill_1 FILLER_50_40 ();
 sg13g2_decap_8 FILLER_50_48 ();
 sg13g2_fill_1 FILLER_50_59 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_4 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_130 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_decap_4 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_152 ();
 sg13g2_fill_2 FILLER_50_168 ();
 sg13g2_decap_4 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_189 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_fill_1 FILLER_50_404 ();
 sg13g2_fill_2 FILLER_50_410 ();
 sg13g2_fill_2 FILLER_50_420 ();
 sg13g2_fill_2 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_434 ();
 sg13g2_fill_2 FILLER_50_439 ();
 sg13g2_fill_1 FILLER_50_441 ();
 sg13g2_fill_1 FILLER_50_446 ();
 sg13g2_fill_1 FILLER_50_487 ();
 sg13g2_fill_2 FILLER_50_493 ();
 sg13g2_fill_1 FILLER_50_495 ();
 sg13g2_fill_1 FILLER_50_506 ();
 sg13g2_fill_1 FILLER_50_517 ();
 sg13g2_fill_2 FILLER_50_531 ();
 sg13g2_fill_2 FILLER_50_538 ();
 sg13g2_fill_1 FILLER_50_545 ();
 sg13g2_fill_2 FILLER_50_551 ();
 sg13g2_fill_1 FILLER_50_571 ();
 sg13g2_fill_1 FILLER_50_626 ();
 sg13g2_fill_1 FILLER_50_637 ();
 sg13g2_fill_1 FILLER_50_650 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_694 ();
 sg13g2_fill_2 FILLER_50_706 ();
 sg13g2_fill_2 FILLER_50_748 ();
 sg13g2_fill_2 FILLER_50_760 ();
 sg13g2_fill_1 FILLER_50_762 ();
 sg13g2_fill_1 FILLER_50_774 ();
 sg13g2_decap_4 FILLER_50_824 ();
 sg13g2_fill_2 FILLER_50_828 ();
 sg13g2_fill_2 FILLER_50_836 ();
 sg13g2_fill_2 FILLER_50_843 ();
 sg13g2_fill_1 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_923 ();
 sg13g2_decap_4 FILLER_50_944 ();
 sg13g2_fill_1 FILLER_50_948 ();
 sg13g2_fill_1 FILLER_50_1010 ();
 sg13g2_fill_2 FILLER_50_1015 ();
 sg13g2_decap_4 FILLER_50_1027 ();
 sg13g2_fill_1 FILLER_50_1035 ();
 sg13g2_decap_8 FILLER_50_1067 ();
 sg13g2_fill_1 FILLER_50_1080 ();
 sg13g2_fill_1 FILLER_50_1086 ();
 sg13g2_fill_2 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1102 ();
 sg13g2_fill_2 FILLER_50_1115 ();
 sg13g2_fill_1 FILLER_50_1117 ();
 sg13g2_fill_2 FILLER_50_1162 ();
 sg13g2_fill_1 FILLER_50_1211 ();
 sg13g2_fill_1 FILLER_50_1230 ();
 sg13g2_fill_1 FILLER_50_1236 ();
 sg13g2_fill_2 FILLER_50_1242 ();
 sg13g2_fill_1 FILLER_50_1336 ();
 sg13g2_fill_2 FILLER_50_1343 ();
 sg13g2_fill_1 FILLER_50_1427 ();
 sg13g2_fill_2 FILLER_50_1472 ();
 sg13g2_fill_1 FILLER_50_1474 ();
 sg13g2_fill_2 FILLER_50_1481 ();
 sg13g2_fill_1 FILLER_50_1483 ();
 sg13g2_fill_1 FILLER_50_1497 ();
 sg13g2_fill_2 FILLER_50_1510 ();
 sg13g2_fill_1 FILLER_50_1529 ();
 sg13g2_fill_2 FILLER_50_1622 ();
 sg13g2_fill_1 FILLER_50_1643 ();
 sg13g2_fill_1 FILLER_50_1652 ();
 sg13g2_fill_1 FILLER_50_1658 ();
 sg13g2_fill_1 FILLER_50_1665 ();
 sg13g2_fill_2 FILLER_50_1679 ();
 sg13g2_fill_2 FILLER_50_1686 ();
 sg13g2_fill_1 FILLER_50_1688 ();
 sg13g2_fill_2 FILLER_50_1696 ();
 sg13g2_fill_2 FILLER_50_1703 ();
 sg13g2_fill_1 FILLER_50_1718 ();
 sg13g2_fill_1 FILLER_50_1723 ();
 sg13g2_fill_2 FILLER_50_1729 ();
 sg13g2_fill_2 FILLER_50_1739 ();
 sg13g2_fill_2 FILLER_50_1764 ();
 sg13g2_fill_2 FILLER_50_1770 ();
 sg13g2_fill_2 FILLER_50_1776 ();
 sg13g2_fill_2 FILLER_50_1786 ();
 sg13g2_fill_2 FILLER_50_1793 ();
 sg13g2_fill_1 FILLER_50_1799 ();
 sg13g2_fill_2 FILLER_50_1808 ();
 sg13g2_decap_8 FILLER_50_1826 ();
 sg13g2_decap_8 FILLER_50_1833 ();
 sg13g2_fill_1 FILLER_50_1840 ();
 sg13g2_decap_4 FILLER_50_1845 ();
 sg13g2_fill_1 FILLER_50_1849 ();
 sg13g2_decap_8 FILLER_50_1854 ();
 sg13g2_decap_8 FILLER_50_1861 ();
 sg13g2_decap_4 FILLER_50_1868 ();
 sg13g2_decap_8 FILLER_50_1876 ();
 sg13g2_decap_8 FILLER_50_1883 ();
 sg13g2_decap_8 FILLER_50_1890 ();
 sg13g2_decap_4 FILLER_50_1897 ();
 sg13g2_decap_4 FILLER_50_1906 ();
 sg13g2_fill_1 FILLER_50_1910 ();
 sg13g2_fill_2 FILLER_50_1916 ();
 sg13g2_decap_8 FILLER_50_1931 ();
 sg13g2_decap_8 FILLER_50_1938 ();
 sg13g2_decap_8 FILLER_50_1950 ();
 sg13g2_fill_2 FILLER_50_1967 ();
 sg13g2_fill_1 FILLER_50_1969 ();
 sg13g2_decap_8 FILLER_50_1974 ();
 sg13g2_decap_8 FILLER_50_1981 ();
 sg13g2_decap_4 FILLER_50_1988 ();
 sg13g2_fill_1 FILLER_50_1992 ();
 sg13g2_fill_1 FILLER_50_2011 ();
 sg13g2_decap_8 FILLER_50_2018 ();
 sg13g2_decap_8 FILLER_50_2025 ();
 sg13g2_decap_8 FILLER_50_2032 ();
 sg13g2_decap_8 FILLER_50_2039 ();
 sg13g2_decap_8 FILLER_50_2046 ();
 sg13g2_decap_8 FILLER_50_2053 ();
 sg13g2_decap_8 FILLER_50_2060 ();
 sg13g2_decap_4 FILLER_50_2067 ();
 sg13g2_fill_2 FILLER_50_2127 ();
 sg13g2_decap_8 FILLER_50_2133 ();
 sg13g2_decap_8 FILLER_50_2140 ();
 sg13g2_decap_4 FILLER_50_2147 ();
 sg13g2_fill_1 FILLER_50_2151 ();
 sg13g2_fill_2 FILLER_50_2161 ();
 sg13g2_fill_1 FILLER_50_2197 ();
 sg13g2_decap_4 FILLER_50_2224 ();
 sg13g2_fill_1 FILLER_50_2228 ();
 sg13g2_fill_2 FILLER_50_2279 ();
 sg13g2_fill_1 FILLER_50_2311 ();
 sg13g2_fill_2 FILLER_50_2317 ();
 sg13g2_fill_2 FILLER_50_2354 ();
 sg13g2_fill_2 FILLER_50_2377 ();
 sg13g2_fill_2 FILLER_50_2393 ();
 sg13g2_fill_1 FILLER_50_2395 ();
 sg13g2_decap_4 FILLER_50_2449 ();
 sg13g2_fill_1 FILLER_50_2453 ();
 sg13g2_fill_1 FILLER_50_2502 ();
 sg13g2_fill_2 FILLER_50_2513 ();
 sg13g2_fill_2 FILLER_50_2519 ();
 sg13g2_fill_1 FILLER_50_2526 ();
 sg13g2_fill_1 FILLER_50_2531 ();
 sg13g2_fill_2 FILLER_50_2575 ();
 sg13g2_fill_1 FILLER_50_2577 ();
 sg13g2_decap_4 FILLER_50_2630 ();
 sg13g2_fill_1 FILLER_50_2634 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_decap_8 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2660 ();
 sg13g2_fill_2 FILLER_50_2667 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_decap_4 FILLER_51_37 ();
 sg13g2_fill_1 FILLER_51_75 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_decap_4 FILLER_51_92 ();
 sg13g2_decap_4 FILLER_51_100 ();
 sg13g2_fill_2 FILLER_51_104 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_fill_1 FILLER_51_207 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_2 FILLER_51_381 ();
 sg13g2_fill_1 FILLER_51_414 ();
 sg13g2_decap_8 FILLER_51_419 ();
 sg13g2_decap_8 FILLER_51_426 ();
 sg13g2_decap_8 FILLER_51_433 ();
 sg13g2_decap_8 FILLER_51_440 ();
 sg13g2_decap_8 FILLER_51_447 ();
 sg13g2_fill_2 FILLER_51_454 ();
 sg13g2_decap_4 FILLER_51_465 ();
 sg13g2_fill_2 FILLER_51_473 ();
 sg13g2_fill_1 FILLER_51_541 ();
 sg13g2_fill_2 FILLER_51_546 ();
 sg13g2_fill_1 FILLER_51_574 ();
 sg13g2_fill_1 FILLER_51_605 ();
 sg13g2_decap_8 FILLER_51_618 ();
 sg13g2_fill_1 FILLER_51_681 ();
 sg13g2_fill_1 FILLER_51_692 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_fill_2 FILLER_51_743 ();
 sg13g2_fill_2 FILLER_51_750 ();
 sg13g2_decap_4 FILLER_51_756 ();
 sg13g2_fill_1 FILLER_51_760 ();
 sg13g2_decap_4 FILLER_51_770 ();
 sg13g2_fill_1 FILLER_51_774 ();
 sg13g2_fill_2 FILLER_51_794 ();
 sg13g2_fill_1 FILLER_51_824 ();
 sg13g2_fill_1 FILLER_51_842 ();
 sg13g2_fill_1 FILLER_51_853 ();
 sg13g2_fill_1 FILLER_51_867 ();
 sg13g2_decap_4 FILLER_51_883 ();
 sg13g2_fill_1 FILLER_51_887 ();
 sg13g2_fill_1 FILLER_51_893 ();
 sg13g2_fill_1 FILLER_51_898 ();
 sg13g2_fill_2 FILLER_51_903 ();
 sg13g2_fill_1 FILLER_51_909 ();
 sg13g2_fill_1 FILLER_51_936 ();
 sg13g2_fill_1 FILLER_51_941 ();
 sg13g2_fill_2 FILLER_51_952 ();
 sg13g2_fill_1 FILLER_51_954 ();
 sg13g2_fill_1 FILLER_51_964 ();
 sg13g2_fill_2 FILLER_51_969 ();
 sg13g2_fill_1 FILLER_51_984 ();
 sg13g2_decap_8 FILLER_51_1015 ();
 sg13g2_fill_2 FILLER_51_1022 ();
 sg13g2_fill_2 FILLER_51_1050 ();
 sg13g2_fill_2 FILLER_51_1057 ();
 sg13g2_fill_1 FILLER_51_1085 ();
 sg13g2_fill_1 FILLER_51_1109 ();
 sg13g2_fill_1 FILLER_51_1124 ();
 sg13g2_decap_8 FILLER_51_1133 ();
 sg13g2_fill_2 FILLER_51_1229 ();
 sg13g2_fill_1 FILLER_51_1304 ();
 sg13g2_fill_2 FILLER_51_1344 ();
 sg13g2_fill_2 FILLER_51_1350 ();
 sg13g2_fill_1 FILLER_51_1358 ();
 sg13g2_fill_1 FILLER_51_1373 ();
 sg13g2_fill_1 FILLER_51_1383 ();
 sg13g2_fill_2 FILLER_51_1451 ();
 sg13g2_fill_1 FILLER_51_1453 ();
 sg13g2_fill_1 FILLER_51_1462 ();
 sg13g2_fill_2 FILLER_51_1500 ();
 sg13g2_fill_2 FILLER_51_1559 ();
 sg13g2_fill_2 FILLER_51_1574 ();
 sg13g2_fill_1 FILLER_51_1594 ();
 sg13g2_decap_4 FILLER_51_1621 ();
 sg13g2_fill_1 FILLER_51_1625 ();
 sg13g2_fill_1 FILLER_51_1630 ();
 sg13g2_fill_1 FILLER_51_1644 ();
 sg13g2_fill_1 FILLER_51_1649 ();
 sg13g2_decap_8 FILLER_51_1670 ();
 sg13g2_decap_4 FILLER_51_1677 ();
 sg13g2_fill_2 FILLER_51_1681 ();
 sg13g2_fill_2 FILLER_51_1690 ();
 sg13g2_fill_1 FILLER_51_1692 ();
 sg13g2_fill_2 FILLER_51_1714 ();
 sg13g2_fill_1 FILLER_51_1716 ();
 sg13g2_fill_1 FILLER_51_1726 ();
 sg13g2_fill_2 FILLER_51_1732 ();
 sg13g2_fill_1 FILLER_51_1772 ();
 sg13g2_fill_2 FILLER_51_1800 ();
 sg13g2_decap_8 FILLER_51_1806 ();
 sg13g2_decap_8 FILLER_51_1813 ();
 sg13g2_decap_4 FILLER_51_1820 ();
 sg13g2_decap_8 FILLER_51_1829 ();
 sg13g2_decap_8 FILLER_51_1836 ();
 sg13g2_decap_4 FILLER_51_1843 ();
 sg13g2_fill_2 FILLER_51_1847 ();
 sg13g2_decap_8 FILLER_51_1854 ();
 sg13g2_decap_8 FILLER_51_1861 ();
 sg13g2_decap_8 FILLER_51_1868 ();
 sg13g2_decap_8 FILLER_51_1875 ();
 sg13g2_decap_8 FILLER_51_1882 ();
 sg13g2_decap_4 FILLER_51_1889 ();
 sg13g2_decap_8 FILLER_51_1901 ();
 sg13g2_decap_8 FILLER_51_1908 ();
 sg13g2_decap_8 FILLER_51_1915 ();
 sg13g2_fill_1 FILLER_51_1922 ();
 sg13g2_decap_4 FILLER_51_1927 ();
 sg13g2_decap_8 FILLER_51_1935 ();
 sg13g2_decap_8 FILLER_51_1942 ();
 sg13g2_decap_4 FILLER_51_1949 ();
 sg13g2_fill_2 FILLER_51_1953 ();
 sg13g2_decap_8 FILLER_51_1959 ();
 sg13g2_decap_8 FILLER_51_1966 ();
 sg13g2_decap_8 FILLER_51_1973 ();
 sg13g2_decap_4 FILLER_51_1980 ();
 sg13g2_fill_1 FILLER_51_1984 ();
 sg13g2_decap_8 FILLER_51_1989 ();
 sg13g2_fill_1 FILLER_51_1996 ();
 sg13g2_fill_2 FILLER_51_2006 ();
 sg13g2_decap_4 FILLER_51_2013 ();
 sg13g2_fill_2 FILLER_51_2017 ();
 sg13g2_fill_2 FILLER_51_2025 ();
 sg13g2_decap_8 FILLER_51_2032 ();
 sg13g2_decap_8 FILLER_51_2039 ();
 sg13g2_decap_8 FILLER_51_2046 ();
 sg13g2_decap_8 FILLER_51_2053 ();
 sg13g2_decap_8 FILLER_51_2060 ();
 sg13g2_decap_8 FILLER_51_2067 ();
 sg13g2_fill_2 FILLER_51_2078 ();
 sg13g2_fill_1 FILLER_51_2119 ();
 sg13g2_fill_2 FILLER_51_2154 ();
 sg13g2_decap_4 FILLER_51_2162 ();
 sg13g2_fill_1 FILLER_51_2166 ();
 sg13g2_fill_2 FILLER_51_2176 ();
 sg13g2_fill_1 FILLER_51_2178 ();
 sg13g2_fill_1 FILLER_51_2183 ();
 sg13g2_fill_1 FILLER_51_2188 ();
 sg13g2_decap_4 FILLER_51_2193 ();
 sg13g2_fill_2 FILLER_51_2197 ();
 sg13g2_fill_1 FILLER_51_2208 ();
 sg13g2_fill_2 FILLER_51_2213 ();
 sg13g2_decap_8 FILLER_51_2222 ();
 sg13g2_fill_2 FILLER_51_2229 ();
 sg13g2_fill_1 FILLER_51_2231 ();
 sg13g2_fill_1 FILLER_51_2236 ();
 sg13g2_decap_8 FILLER_51_2247 ();
 sg13g2_decap_4 FILLER_51_2280 ();
 sg13g2_fill_1 FILLER_51_2284 ();
 sg13g2_fill_2 FILLER_51_2288 ();
 sg13g2_fill_2 FILLER_51_2311 ();
 sg13g2_fill_2 FILLER_51_2316 ();
 sg13g2_fill_2 FILLER_51_2344 ();
 sg13g2_fill_2 FILLER_51_2372 ();
 sg13g2_fill_1 FILLER_51_2374 ();
 sg13g2_fill_2 FILLER_51_2423 ();
 sg13g2_fill_1 FILLER_51_2425 ();
 sg13g2_decap_8 FILLER_51_2452 ();
 sg13g2_decap_4 FILLER_51_2459 ();
 sg13g2_fill_2 FILLER_51_2463 ();
 sg13g2_decap_8 FILLER_51_2469 ();
 sg13g2_fill_1 FILLER_51_2476 ();
 sg13g2_fill_2 FILLER_51_2493 ();
 sg13g2_fill_1 FILLER_51_2534 ();
 sg13g2_fill_2 FILLER_51_2539 ();
 sg13g2_fill_1 FILLER_51_2541 ();
 sg13g2_fill_2 FILLER_51_2547 ();
 sg13g2_fill_1 FILLER_51_2556 ();
 sg13g2_fill_1 FILLER_51_2566 ();
 sg13g2_fill_2 FILLER_51_2610 ();
 sg13g2_decap_8 FILLER_51_2652 ();
 sg13g2_decap_8 FILLER_51_2659 ();
 sg13g2_decap_4 FILLER_51_2666 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_52_186 ();
 sg13g2_fill_2 FILLER_52_210 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_389 ();
 sg13g2_decap_8 FILLER_52_424 ();
 sg13g2_fill_1 FILLER_52_431 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_4 FILLER_52_469 ();
 sg13g2_fill_1 FILLER_52_473 ();
 sg13g2_fill_2 FILLER_52_483 ();
 sg13g2_fill_1 FILLER_52_485 ();
 sg13g2_fill_2 FILLER_52_500 ();
 sg13g2_fill_1 FILLER_52_502 ();
 sg13g2_fill_2 FILLER_52_516 ();
 sg13g2_fill_2 FILLER_52_531 ();
 sg13g2_fill_2 FILLER_52_538 ();
 sg13g2_fill_2 FILLER_52_544 ();
 sg13g2_fill_2 FILLER_52_551 ();
 sg13g2_fill_1 FILLER_52_553 ();
 sg13g2_fill_2 FILLER_52_558 ();
 sg13g2_fill_1 FILLER_52_560 ();
 sg13g2_fill_2 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_568 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_decap_4 FILLER_52_629 ();
 sg13g2_fill_1 FILLER_52_683 ();
 sg13g2_fill_2 FILLER_52_689 ();
 sg13g2_fill_2 FILLER_52_695 ();
 sg13g2_fill_2 FILLER_52_702 ();
 sg13g2_fill_2 FILLER_52_725 ();
 sg13g2_fill_1 FILLER_52_727 ();
 sg13g2_fill_1 FILLER_52_741 ();
 sg13g2_fill_2 FILLER_52_750 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_fill_1 FILLER_52_828 ();
 sg13g2_fill_2 FILLER_52_863 ();
 sg13g2_fill_1 FILLER_52_865 ();
 sg13g2_fill_1 FILLER_52_870 ();
 sg13g2_decap_4 FILLER_52_879 ();
 sg13g2_fill_2 FILLER_52_883 ();
 sg13g2_decap_4 FILLER_52_890 ();
 sg13g2_fill_1 FILLER_52_894 ();
 sg13g2_decap_8 FILLER_52_905 ();
 sg13g2_fill_1 FILLER_52_965 ();
 sg13g2_decap_8 FILLER_52_1009 ();
 sg13g2_fill_2 FILLER_52_1016 ();
 sg13g2_fill_1 FILLER_52_1018 ();
 sg13g2_decap_4 FILLER_52_1027 ();
 sg13g2_fill_1 FILLER_52_1031 ();
 sg13g2_fill_2 FILLER_52_1046 ();
 sg13g2_fill_1 FILLER_52_1048 ();
 sg13g2_decap_4 FILLER_52_1054 ();
 sg13g2_fill_1 FILLER_52_1099 ();
 sg13g2_decap_4 FILLER_52_1173 ();
 sg13g2_fill_1 FILLER_52_1177 ();
 sg13g2_fill_1 FILLER_52_1181 ();
 sg13g2_fill_1 FILLER_52_1255 ();
 sg13g2_fill_1 FILLER_52_1276 ();
 sg13g2_fill_2 FILLER_52_1306 ();
 sg13g2_fill_1 FILLER_52_1312 ();
 sg13g2_fill_2 FILLER_52_1376 ();
 sg13g2_fill_1 FILLER_52_1378 ();
 sg13g2_fill_2 FILLER_52_1387 ();
 sg13g2_fill_2 FILLER_52_1415 ();
 sg13g2_fill_2 FILLER_52_1422 ();
 sg13g2_fill_2 FILLER_52_1428 ();
 sg13g2_fill_1 FILLER_52_1430 ();
 sg13g2_decap_8 FILLER_52_1441 ();
 sg13g2_fill_2 FILLER_52_1448 ();
 sg13g2_fill_1 FILLER_52_1450 ();
 sg13g2_fill_1 FILLER_52_1468 ();
 sg13g2_fill_1 FILLER_52_1474 ();
 sg13g2_fill_1 FILLER_52_1480 ();
 sg13g2_fill_2 FILLER_52_1489 ();
 sg13g2_fill_1 FILLER_52_1505 ();
 sg13g2_fill_1 FILLER_52_1511 ();
 sg13g2_fill_1 FILLER_52_1516 ();
 sg13g2_fill_1 FILLER_52_1522 ();
 sg13g2_fill_1 FILLER_52_1532 ();
 sg13g2_fill_2 FILLER_52_1546 ();
 sg13g2_fill_2 FILLER_52_1554 ();
 sg13g2_fill_2 FILLER_52_1587 ();
 sg13g2_fill_2 FILLER_52_1598 ();
 sg13g2_decap_8 FILLER_52_1687 ();
 sg13g2_decap_4 FILLER_52_1694 ();
 sg13g2_fill_1 FILLER_52_1698 ();
 sg13g2_decap_4 FILLER_52_1718 ();
 sg13g2_fill_2 FILLER_52_1722 ();
 sg13g2_decap_4 FILLER_52_1728 ();
 sg13g2_fill_1 FILLER_52_1761 ();
 sg13g2_fill_2 FILLER_52_1767 ();
 sg13g2_fill_2 FILLER_52_1779 ();
 sg13g2_fill_1 FILLER_52_1792 ();
 sg13g2_fill_2 FILLER_52_1797 ();
 sg13g2_fill_2 FILLER_52_1804 ();
 sg13g2_fill_1 FILLER_52_1816 ();
 sg13g2_fill_2 FILLER_52_1822 ();
 sg13g2_fill_1 FILLER_52_1824 ();
 sg13g2_decap_8 FILLER_52_1828 ();
 sg13g2_decap_8 FILLER_52_1835 ();
 sg13g2_fill_2 FILLER_52_1842 ();
 sg13g2_decap_8 FILLER_52_1850 ();
 sg13g2_decap_8 FILLER_52_1857 ();
 sg13g2_decap_8 FILLER_52_1864 ();
 sg13g2_decap_8 FILLER_52_1871 ();
 sg13g2_fill_2 FILLER_52_1878 ();
 sg13g2_fill_1 FILLER_52_1880 ();
 sg13g2_decap_8 FILLER_52_1886 ();
 sg13g2_decap_4 FILLER_52_1893 ();
 sg13g2_fill_2 FILLER_52_1897 ();
 sg13g2_decap_8 FILLER_52_1909 ();
 sg13g2_decap_8 FILLER_52_1916 ();
 sg13g2_decap_8 FILLER_52_1923 ();
 sg13g2_decap_8 FILLER_52_1930 ();
 sg13g2_fill_1 FILLER_52_1937 ();
 sg13g2_decap_8 FILLER_52_1942 ();
 sg13g2_decap_8 FILLER_52_1949 ();
 sg13g2_decap_8 FILLER_52_1956 ();
 sg13g2_decap_8 FILLER_52_1963 ();
 sg13g2_decap_8 FILLER_52_1970 ();
 sg13g2_decap_8 FILLER_52_1977 ();
 sg13g2_decap_8 FILLER_52_1984 ();
 sg13g2_decap_8 FILLER_52_1991 ();
 sg13g2_decap_8 FILLER_52_1998 ();
 sg13g2_decap_4 FILLER_52_2005 ();
 sg13g2_fill_2 FILLER_52_2009 ();
 sg13g2_decap_8 FILLER_52_2015 ();
 sg13g2_decap_8 FILLER_52_2022 ();
 sg13g2_decap_8 FILLER_52_2029 ();
 sg13g2_decap_8 FILLER_52_2036 ();
 sg13g2_decap_8 FILLER_52_2043 ();
 sg13g2_decap_8 FILLER_52_2070 ();
 sg13g2_decap_8 FILLER_52_2077 ();
 sg13g2_decap_8 FILLER_52_2084 ();
 sg13g2_fill_2 FILLER_52_2091 ();
 sg13g2_fill_1 FILLER_52_2105 ();
 sg13g2_fill_1 FILLER_52_2111 ();
 sg13g2_fill_1 FILLER_52_2116 ();
 sg13g2_fill_2 FILLER_52_2166 ();
 sg13g2_fill_1 FILLER_52_2168 ();
 sg13g2_fill_1 FILLER_52_2175 ();
 sg13g2_fill_1 FILLER_52_2216 ();
 sg13g2_fill_1 FILLER_52_2271 ();
 sg13g2_fill_2 FILLER_52_2298 ();
 sg13g2_fill_2 FILLER_52_2343 ();
 sg13g2_fill_2 FILLER_52_2376 ();
 sg13g2_fill_1 FILLER_52_2378 ();
 sg13g2_fill_2 FILLER_52_2397 ();
 sg13g2_fill_1 FILLER_52_2399 ();
 sg13g2_fill_1 FILLER_52_2412 ();
 sg13g2_decap_4 FILLER_52_2457 ();
 sg13g2_fill_2 FILLER_52_2461 ();
 sg13g2_fill_1 FILLER_52_2467 ();
 sg13g2_fill_2 FILLER_52_2474 ();
 sg13g2_fill_2 FILLER_52_2482 ();
 sg13g2_fill_2 FILLER_52_2489 ();
 sg13g2_fill_1 FILLER_52_2491 ();
 sg13g2_fill_2 FILLER_52_2510 ();
 sg13g2_fill_1 FILLER_52_2512 ();
 sg13g2_fill_2 FILLER_52_2536 ();
 sg13g2_fill_1 FILLER_52_2538 ();
 sg13g2_fill_2 FILLER_52_2553 ();
 sg13g2_fill_1 FILLER_52_2561 ();
 sg13g2_decap_4 FILLER_52_2573 ();
 sg13g2_fill_2 FILLER_52_2577 ();
 sg13g2_fill_1 FILLER_52_2583 ();
 sg13g2_decap_4 FILLER_52_2588 ();
 sg13g2_fill_2 FILLER_52_2592 ();
 sg13g2_decap_8 FILLER_52_2630 ();
 sg13g2_decap_8 FILLER_52_2637 ();
 sg13g2_decap_8 FILLER_52_2644 ();
 sg13g2_decap_8 FILLER_52_2651 ();
 sg13g2_decap_8 FILLER_52_2658 ();
 sg13g2_decap_4 FILLER_52_2665 ();
 sg13g2_fill_1 FILLER_52_2669 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_13 ();
 sg13g2_decap_4 FILLER_53_22 ();
 sg13g2_fill_1 FILLER_53_60 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_73 ();
 sg13g2_decap_4 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_97 ();
 sg13g2_decap_4 FILLER_53_102 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_fill_1 FILLER_53_136 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_decap_4 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_188 ();
 sg13g2_decap_8 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_212 ();
 sg13g2_decap_4 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_fill_2 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_285 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_362 ();
 sg13g2_fill_1 FILLER_53_392 ();
 sg13g2_fill_1 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_457 ();
 sg13g2_fill_2 FILLER_53_494 ();
 sg13g2_fill_1 FILLER_53_496 ();
 sg13g2_fill_1 FILLER_53_507 ();
 sg13g2_fill_2 FILLER_53_513 ();
 sg13g2_fill_1 FILLER_53_515 ();
 sg13g2_fill_1 FILLER_53_521 ();
 sg13g2_fill_1 FILLER_53_545 ();
 sg13g2_fill_2 FILLER_53_550 ();
 sg13g2_fill_1 FILLER_53_566 ();
 sg13g2_fill_2 FILLER_53_593 ();
 sg13g2_fill_2 FILLER_53_600 ();
 sg13g2_decap_4 FILLER_53_611 ();
 sg13g2_fill_2 FILLER_53_619 ();
 sg13g2_fill_1 FILLER_53_630 ();
 sg13g2_fill_1 FILLER_53_636 ();
 sg13g2_decap_4 FILLER_53_642 ();
 sg13g2_fill_1 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_fill_2 FILLER_53_663 ();
 sg13g2_fill_1 FILLER_53_665 ();
 sg13g2_decap_4 FILLER_53_671 ();
 sg13g2_decap_4 FILLER_53_679 ();
 sg13g2_decap_4 FILLER_53_687 ();
 sg13g2_fill_2 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_707 ();
 sg13g2_fill_1 FILLER_53_721 ();
 sg13g2_fill_1 FILLER_53_761 ();
 sg13g2_fill_2 FILLER_53_772 ();
 sg13g2_fill_2 FILLER_53_809 ();
 sg13g2_decap_4 FILLER_53_815 ();
 sg13g2_fill_2 FILLER_53_819 ();
 sg13g2_fill_2 FILLER_53_835 ();
 sg13g2_fill_2 FILLER_53_869 ();
 sg13g2_fill_1 FILLER_53_875 ();
 sg13g2_fill_1 FILLER_53_884 ();
 sg13g2_fill_2 FILLER_53_894 ();
 sg13g2_fill_1 FILLER_53_905 ();
 sg13g2_decap_4 FILLER_53_910 ();
 sg13g2_decap_4 FILLER_53_922 ();
 sg13g2_decap_8 FILLER_53_931 ();
 sg13g2_fill_1 FILLER_53_938 ();
 sg13g2_fill_2 FILLER_53_943 ();
 sg13g2_fill_1 FILLER_53_945 ();
 sg13g2_fill_2 FILLER_53_960 ();
 sg13g2_fill_2 FILLER_53_1009 ();
 sg13g2_decap_8 FILLER_53_1037 ();
 sg13g2_decap_8 FILLER_53_1044 ();
 sg13g2_decap_4 FILLER_53_1051 ();
 sg13g2_fill_1 FILLER_53_1078 ();
 sg13g2_fill_1 FILLER_53_1083 ();
 sg13g2_decap_4 FILLER_53_1132 ();
 sg13g2_fill_1 FILLER_53_1136 ();
 sg13g2_fill_2 FILLER_53_1141 ();
 sg13g2_fill_2 FILLER_53_1162 ();
 sg13g2_fill_1 FILLER_53_1172 ();
 sg13g2_decap_8 FILLER_53_1187 ();
 sg13g2_decap_8 FILLER_53_1194 ();
 sg13g2_fill_2 FILLER_53_1201 ();
 sg13g2_fill_1 FILLER_53_1203 ();
 sg13g2_fill_2 FILLER_53_1208 ();
 sg13g2_fill_2 FILLER_53_1239 ();
 sg13g2_fill_1 FILLER_53_1246 ();
 sg13g2_fill_2 FILLER_53_1253 ();
 sg13g2_fill_2 FILLER_53_1312 ();
 sg13g2_fill_2 FILLER_53_1326 ();
 sg13g2_decap_8 FILLER_53_1370 ();
 sg13g2_decap_8 FILLER_53_1377 ();
 sg13g2_decap_8 FILLER_53_1384 ();
 sg13g2_decap_4 FILLER_53_1391 ();
 sg13g2_fill_2 FILLER_53_1399 ();
 sg13g2_decap_8 FILLER_53_1414 ();
 sg13g2_fill_2 FILLER_53_1421 ();
 sg13g2_decap_8 FILLER_53_1431 ();
 sg13g2_decap_8 FILLER_53_1438 ();
 sg13g2_decap_4 FILLER_53_1445 ();
 sg13g2_fill_1 FILLER_53_1449 ();
 sg13g2_fill_1 FILLER_53_1458 ();
 sg13g2_fill_2 FILLER_53_1466 ();
 sg13g2_fill_1 FILLER_53_1468 ();
 sg13g2_fill_2 FILLER_53_1474 ();
 sg13g2_fill_2 FILLER_53_1499 ();
 sg13g2_fill_1 FILLER_53_1535 ();
 sg13g2_decap_8 FILLER_53_1583 ();
 sg13g2_decap_8 FILLER_53_1590 ();
 sg13g2_decap_8 FILLER_53_1597 ();
 sg13g2_fill_2 FILLER_53_1604 ();
 sg13g2_decap_4 FILLER_53_1610 ();
 sg13g2_fill_2 FILLER_53_1614 ();
 sg13g2_fill_2 FILLER_53_1619 ();
 sg13g2_fill_1 FILLER_53_1632 ();
 sg13g2_fill_1 FILLER_53_1638 ();
 sg13g2_fill_1 FILLER_53_1657 ();
 sg13g2_fill_1 FILLER_53_1676 ();
 sg13g2_fill_2 FILLER_53_1690 ();
 sg13g2_fill_1 FILLER_53_1692 ();
 sg13g2_fill_2 FILLER_53_1697 ();
 sg13g2_fill_1 FILLER_53_1699 ();
 sg13g2_decap_8 FILLER_53_1706 ();
 sg13g2_decap_8 FILLER_53_1713 ();
 sg13g2_decap_8 FILLER_53_1720 ();
 sg13g2_decap_4 FILLER_53_1727 ();
 sg13g2_fill_1 FILLER_53_1731 ();
 sg13g2_decap_4 FILLER_53_1740 ();
 sg13g2_fill_2 FILLER_53_1796 ();
 sg13g2_fill_2 FILLER_53_1803 ();
 sg13g2_fill_1 FILLER_53_1805 ();
 sg13g2_fill_1 FILLER_53_1809 ();
 sg13g2_fill_2 FILLER_53_1815 ();
 sg13g2_decap_8 FILLER_53_1826 ();
 sg13g2_decap_8 FILLER_53_1833 ();
 sg13g2_decap_8 FILLER_53_1840 ();
 sg13g2_decap_8 FILLER_53_1847 ();
 sg13g2_decap_4 FILLER_53_1854 ();
 sg13g2_fill_2 FILLER_53_1858 ();
 sg13g2_decap_4 FILLER_53_1869 ();
 sg13g2_fill_2 FILLER_53_1873 ();
 sg13g2_fill_1 FILLER_53_1892 ();
 sg13g2_decap_8 FILLER_53_1898 ();
 sg13g2_decap_8 FILLER_53_1905 ();
 sg13g2_decap_8 FILLER_53_1912 ();
 sg13g2_decap_8 FILLER_53_1919 ();
 sg13g2_decap_8 FILLER_53_1926 ();
 sg13g2_fill_2 FILLER_53_1933 ();
 sg13g2_fill_1 FILLER_53_1935 ();
 sg13g2_fill_2 FILLER_53_1948 ();
 sg13g2_decap_8 FILLER_53_1960 ();
 sg13g2_decap_4 FILLER_53_1967 ();
 sg13g2_fill_2 FILLER_53_1971 ();
 sg13g2_decap_8 FILLER_53_1977 ();
 sg13g2_decap_8 FILLER_53_1984 ();
 sg13g2_decap_8 FILLER_53_1991 ();
 sg13g2_decap_8 FILLER_53_1998 ();
 sg13g2_decap_8 FILLER_53_2005 ();
 sg13g2_decap_8 FILLER_53_2012 ();
 sg13g2_decap_8 FILLER_53_2019 ();
 sg13g2_decap_8 FILLER_53_2026 ();
 sg13g2_decap_8 FILLER_53_2033 ();
 sg13g2_decap_8 FILLER_53_2040 ();
 sg13g2_decap_8 FILLER_53_2047 ();
 sg13g2_decap_8 FILLER_53_2054 ();
 sg13g2_decap_8 FILLER_53_2061 ();
 sg13g2_decap_8 FILLER_53_2068 ();
 sg13g2_decap_8 FILLER_53_2075 ();
 sg13g2_decap_8 FILLER_53_2082 ();
 sg13g2_decap_8 FILLER_53_2089 ();
 sg13g2_decap_8 FILLER_53_2096 ();
 sg13g2_fill_2 FILLER_53_2103 ();
 sg13g2_decap_4 FILLER_53_2110 ();
 sg13g2_fill_1 FILLER_53_2114 ();
 sg13g2_fill_1 FILLER_53_2119 ();
 sg13g2_fill_2 FILLER_53_2128 ();
 sg13g2_decap_4 FILLER_53_2138 ();
 sg13g2_decap_4 FILLER_53_2155 ();
 sg13g2_fill_1 FILLER_53_2159 ();
 sg13g2_fill_1 FILLER_53_2168 ();
 sg13g2_fill_2 FILLER_53_2195 ();
 sg13g2_fill_2 FILLER_53_2202 ();
 sg13g2_fill_1 FILLER_53_2216 ();
 sg13g2_fill_2 FILLER_53_2229 ();
 sg13g2_fill_1 FILLER_53_2244 ();
 sg13g2_fill_1 FILLER_53_2250 ();
 sg13g2_decap_4 FILLER_53_2256 ();
 sg13g2_fill_1 FILLER_53_2269 ();
 sg13g2_fill_1 FILLER_53_2274 ();
 sg13g2_fill_1 FILLER_53_2370 ();
 sg13g2_decap_4 FILLER_53_2378 ();
 sg13g2_fill_2 FILLER_53_2392 ();
 sg13g2_fill_1 FILLER_53_2398 ();
 sg13g2_fill_1 FILLER_53_2411 ();
 sg13g2_fill_1 FILLER_53_2422 ();
 sg13g2_fill_1 FILLER_53_2449 ();
 sg13g2_fill_2 FILLER_53_2460 ();
 sg13g2_fill_2 FILLER_53_2467 ();
 sg13g2_fill_1 FILLER_53_2475 ();
 sg13g2_fill_1 FILLER_53_2502 ();
 sg13g2_fill_1 FILLER_53_2513 ();
 sg13g2_fill_1 FILLER_53_2540 ();
 sg13g2_fill_2 FILLER_53_2567 ();
 sg13g2_fill_2 FILLER_53_2579 ();
 sg13g2_fill_1 FILLER_53_2581 ();
 sg13g2_decap_8 FILLER_53_2588 ();
 sg13g2_decap_8 FILLER_53_2595 ();
 sg13g2_fill_1 FILLER_53_2602 ();
 sg13g2_fill_1 FILLER_53_2626 ();
 sg13g2_decap_8 FILLER_53_2653 ();
 sg13g2_decap_8 FILLER_53_2660 ();
 sg13g2_fill_2 FILLER_53_2667 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_decap_4 FILLER_54_31 ();
 sg13g2_fill_2 FILLER_54_96 ();
 sg13g2_fill_1 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_174 ();
 sg13g2_decap_8 FILLER_54_214 ();
 sg13g2_fill_2 FILLER_54_233 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_280 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_307 ();
 sg13g2_fill_2 FILLER_54_338 ();
 sg13g2_fill_2 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_403 ();
 sg13g2_fill_2 FILLER_54_408 ();
 sg13g2_fill_1 FILLER_54_462 ();
 sg13g2_fill_2 FILLER_54_468 ();
 sg13g2_fill_2 FILLER_54_485 ();
 sg13g2_decap_8 FILLER_54_617 ();
 sg13g2_fill_1 FILLER_54_624 ();
 sg13g2_decap_4 FILLER_54_658 ();
 sg13g2_fill_1 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_671 ();
 sg13g2_fill_1 FILLER_54_678 ();
 sg13g2_fill_1 FILLER_54_724 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_fill_2 FILLER_54_760 ();
 sg13g2_fill_1 FILLER_54_762 ();
 sg13g2_fill_1 FILLER_54_793 ();
 sg13g2_fill_2 FILLER_54_803 ();
 sg13g2_fill_1 FILLER_54_831 ();
 sg13g2_fill_1 FILLER_54_863 ();
 sg13g2_fill_1 FILLER_54_869 ();
 sg13g2_fill_1 FILLER_54_875 ();
 sg13g2_fill_2 FILLER_54_881 ();
 sg13g2_fill_1 FILLER_54_888 ();
 sg13g2_fill_2 FILLER_54_894 ();
 sg13g2_fill_2 FILLER_54_922 ();
 sg13g2_decap_8 FILLER_54_960 ();
 sg13g2_decap_8 FILLER_54_967 ();
 sg13g2_fill_1 FILLER_54_980 ();
 sg13g2_fill_2 FILLER_54_997 ();
 sg13g2_fill_1 FILLER_54_999 ();
 sg13g2_fill_1 FILLER_54_1005 ();
 sg13g2_decap_8 FILLER_54_1051 ();
 sg13g2_fill_1 FILLER_54_1058 ();
 sg13g2_fill_2 FILLER_54_1112 ();
 sg13g2_fill_1 FILLER_54_1118 ();
 sg13g2_decap_8 FILLER_54_1127 ();
 sg13g2_decap_8 FILLER_54_1134 ();
 sg13g2_fill_2 FILLER_54_1141 ();
 sg13g2_decap_8 FILLER_54_1146 ();
 sg13g2_fill_2 FILLER_54_1153 ();
 sg13g2_fill_1 FILLER_54_1155 ();
 sg13g2_fill_2 FILLER_54_1166 ();
 sg13g2_decap_4 FILLER_54_1180 ();
 sg13g2_fill_2 FILLER_54_1184 ();
 sg13g2_decap_8 FILLER_54_1201 ();
 sg13g2_fill_2 FILLER_54_1208 ();
 sg13g2_fill_2 FILLER_54_1224 ();
 sg13g2_fill_2 FILLER_54_1258 ();
 sg13g2_fill_1 FILLER_54_1285 ();
 sg13g2_fill_1 FILLER_54_1310 ();
 sg13g2_fill_1 FILLER_54_1342 ();
 sg13g2_fill_2 FILLER_54_1373 ();
 sg13g2_fill_1 FILLER_54_1375 ();
 sg13g2_decap_8 FILLER_54_1420 ();
 sg13g2_fill_2 FILLER_54_1427 ();
 sg13g2_decap_8 FILLER_54_1443 ();
 sg13g2_fill_2 FILLER_54_1450 ();
 sg13g2_fill_1 FILLER_54_1452 ();
 sg13g2_fill_2 FILLER_54_1457 ();
 sg13g2_fill_1 FILLER_54_1464 ();
 sg13g2_decap_4 FILLER_54_1473 ();
 sg13g2_fill_1 FILLER_54_1477 ();
 sg13g2_fill_1 FILLER_54_1492 ();
 sg13g2_fill_2 FILLER_54_1498 ();
 sg13g2_fill_2 FILLER_54_1505 ();
 sg13g2_fill_1 FILLER_54_1507 ();
 sg13g2_decap_8 FILLER_54_1516 ();
 sg13g2_fill_2 FILLER_54_1523 ();
 sg13g2_decap_8 FILLER_54_1543 ();
 sg13g2_decap_4 FILLER_54_1550 ();
 sg13g2_fill_2 FILLER_54_1554 ();
 sg13g2_decap_8 FILLER_54_1567 ();
 sg13g2_fill_2 FILLER_54_1574 ();
 sg13g2_fill_2 FILLER_54_1580 ();
 sg13g2_decap_8 FILLER_54_1586 ();
 sg13g2_decap_8 FILLER_54_1593 ();
 sg13g2_decap_4 FILLER_54_1600 ();
 sg13g2_fill_2 FILLER_54_1604 ();
 sg13g2_fill_1 FILLER_54_1637 ();
 sg13g2_fill_2 FILLER_54_1659 ();
 sg13g2_fill_1 FILLER_54_1694 ();
 sg13g2_decap_4 FILLER_54_1701 ();
 sg13g2_fill_1 FILLER_54_1705 ();
 sg13g2_decap_8 FILLER_54_1711 ();
 sg13g2_fill_2 FILLER_54_1718 ();
 sg13g2_decap_4 FILLER_54_1729 ();
 sg13g2_fill_2 FILLER_54_1737 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_fill_1 FILLER_54_1750 ();
 sg13g2_fill_1 FILLER_54_1770 ();
 sg13g2_fill_1 FILLER_54_1785 ();
 sg13g2_fill_1 FILLER_54_1792 ();
 sg13g2_fill_1 FILLER_54_1801 ();
 sg13g2_fill_2 FILLER_54_1841 ();
 sg13g2_fill_1 FILLER_54_1843 ();
 sg13g2_fill_1 FILLER_54_1848 ();
 sg13g2_fill_2 FILLER_54_1853 ();
 sg13g2_fill_1 FILLER_54_1855 ();
 sg13g2_fill_2 FILLER_54_1870 ();
 sg13g2_fill_1 FILLER_54_1878 ();
 sg13g2_decap_4 FILLER_54_1883 ();
 sg13g2_fill_2 FILLER_54_1902 ();
 sg13g2_fill_1 FILLER_54_1904 ();
 sg13g2_decap_4 FILLER_54_1919 ();
 sg13g2_decap_4 FILLER_54_1928 ();
 sg13g2_fill_2 FILLER_54_1932 ();
 sg13g2_decap_8 FILLER_54_1940 ();
 sg13g2_fill_1 FILLER_54_1947 ();
 sg13g2_fill_1 FILLER_54_1953 ();
 sg13g2_decap_8 FILLER_54_1959 ();
 sg13g2_fill_2 FILLER_54_1966 ();
 sg13g2_fill_1 FILLER_54_1968 ();
 sg13g2_fill_2 FILLER_54_1978 ();
 sg13g2_fill_1 FILLER_54_1980 ();
 sg13g2_decap_8 FILLER_54_1986 ();
 sg13g2_fill_2 FILLER_54_1993 ();
 sg13g2_decap_8 FILLER_54_2000 ();
 sg13g2_decap_8 FILLER_54_2007 ();
 sg13g2_decap_4 FILLER_54_2014 ();
 sg13g2_fill_2 FILLER_54_2018 ();
 sg13g2_fill_1 FILLER_54_2026 ();
 sg13g2_decap_8 FILLER_54_2033 ();
 sg13g2_decap_8 FILLER_54_2040 ();
 sg13g2_decap_8 FILLER_54_2047 ();
 sg13g2_decap_8 FILLER_54_2054 ();
 sg13g2_decap_8 FILLER_54_2061 ();
 sg13g2_decap_8 FILLER_54_2068 ();
 sg13g2_decap_8 FILLER_54_2075 ();
 sg13g2_decap_4 FILLER_54_2082 ();
 sg13g2_fill_1 FILLER_54_2086 ();
 sg13g2_fill_2 FILLER_54_2092 ();
 sg13g2_fill_2 FILLER_54_2128 ();
 sg13g2_fill_2 FILLER_54_2135 ();
 sg13g2_fill_1 FILLER_54_2137 ();
 sg13g2_fill_2 FILLER_54_2142 ();
 sg13g2_fill_1 FILLER_54_2144 ();
 sg13g2_fill_2 FILLER_54_2151 ();
 sg13g2_fill_1 FILLER_54_2153 ();
 sg13g2_fill_1 FILLER_54_2164 ();
 sg13g2_fill_1 FILLER_54_2170 ();
 sg13g2_fill_2 FILLER_54_2176 ();
 sg13g2_fill_2 FILLER_54_2189 ();
 sg13g2_fill_1 FILLER_54_2225 ();
 sg13g2_fill_1 FILLER_54_2274 ();
 sg13g2_fill_2 FILLER_54_2283 ();
 sg13g2_fill_1 FILLER_54_2304 ();
 sg13g2_fill_1 FILLER_54_2310 ();
 sg13g2_fill_1 FILLER_54_2361 ();
 sg13g2_fill_2 FILLER_54_2391 ();
 sg13g2_fill_1 FILLER_54_2393 ();
 sg13g2_fill_1 FILLER_54_2451 ();
 sg13g2_fill_1 FILLER_54_2478 ();
 sg13g2_fill_2 FILLER_54_2484 ();
 sg13g2_fill_2 FILLER_54_2490 ();
 sg13g2_fill_2 FILLER_54_2498 ();
 sg13g2_fill_1 FILLER_54_2530 ();
 sg13g2_fill_2 FILLER_54_2578 ();
 sg13g2_decap_8 FILLER_54_2606 ();
 sg13g2_fill_2 FILLER_54_2613 ();
 sg13g2_decap_8 FILLER_54_2625 ();
 sg13g2_fill_2 FILLER_54_2632 ();
 sg13g2_decap_8 FILLER_54_2642 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_49 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_decap_4 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_2 FILLER_55_74 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_fill_2 FILLER_55_114 ();
 sg13g2_decap_8 FILLER_55_120 ();
 sg13g2_decap_4 FILLER_55_127 ();
 sg13g2_fill_1 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_decap_4 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_163 ();
 sg13g2_decap_8 FILLER_55_169 ();
 sg13g2_decap_8 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_193 ();
 sg13g2_fill_1 FILLER_55_195 ();
 sg13g2_fill_2 FILLER_55_259 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_367 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_decap_4 FILLER_55_411 ();
 sg13g2_fill_1 FILLER_55_434 ();
 sg13g2_decap_4 FILLER_55_548 ();
 sg13g2_fill_2 FILLER_55_596 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_fill_2 FILLER_55_613 ();
 sg13g2_decap_8 FILLER_55_620 ();
 sg13g2_decap_8 FILLER_55_635 ();
 sg13g2_fill_1 FILLER_55_642 ();
 sg13g2_decap_8 FILLER_55_647 ();
 sg13g2_fill_2 FILLER_55_654 ();
 sg13g2_decap_8 FILLER_55_659 ();
 sg13g2_decap_8 FILLER_55_666 ();
 sg13g2_decap_8 FILLER_55_673 ();
 sg13g2_decap_8 FILLER_55_680 ();
 sg13g2_fill_1 FILLER_55_687 ();
 sg13g2_fill_2 FILLER_55_728 ();
 sg13g2_fill_2 FILLER_55_747 ();
 sg13g2_fill_2 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_769 ();
 sg13g2_decap_4 FILLER_55_784 ();
 sg13g2_fill_1 FILLER_55_788 ();
 sg13g2_fill_2 FILLER_55_800 ();
 sg13g2_fill_2 FILLER_55_807 ();
 sg13g2_fill_1 FILLER_55_814 ();
 sg13g2_fill_2 FILLER_55_819 ();
 sg13g2_decap_4 FILLER_55_826 ();
 sg13g2_fill_1 FILLER_55_830 ();
 sg13g2_fill_1 FILLER_55_915 ();
 sg13g2_fill_2 FILLER_55_994 ();
 sg13g2_fill_2 FILLER_55_1022 ();
 sg13g2_fill_1 FILLER_55_1038 ();
 sg13g2_fill_2 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1047 ();
 sg13g2_fill_1 FILLER_55_1052 ();
 sg13g2_fill_2 FILLER_55_1064 ();
 sg13g2_fill_1 FILLER_55_1109 ();
 sg13g2_fill_2 FILLER_55_1119 ();
 sg13g2_fill_1 FILLER_55_1136 ();
 sg13g2_fill_2 FILLER_55_1142 ();
 sg13g2_fill_2 FILLER_55_1177 ();
 sg13g2_fill_1 FILLER_55_1179 ();
 sg13g2_fill_1 FILLER_55_1188 ();
 sg13g2_fill_2 FILLER_55_1197 ();
 sg13g2_fill_1 FILLER_55_1199 ();
 sg13g2_fill_2 FILLER_55_1214 ();
 sg13g2_fill_1 FILLER_55_1233 ();
 sg13g2_fill_1 FILLER_55_1238 ();
 sg13g2_decap_8 FILLER_55_1246 ();
 sg13g2_decap_8 FILLER_55_1253 ();
 sg13g2_decap_8 FILLER_55_1260 ();
 sg13g2_decap_4 FILLER_55_1267 ();
 sg13g2_fill_2 FILLER_55_1278 ();
 sg13g2_fill_1 FILLER_55_1329 ();
 sg13g2_decap_8 FILLER_55_1416 ();
 sg13g2_decap_8 FILLER_55_1423 ();
 sg13g2_decap_4 FILLER_55_1430 ();
 sg13g2_fill_2 FILLER_55_1456 ();
 sg13g2_fill_1 FILLER_55_1465 ();
 sg13g2_decap_4 FILLER_55_1475 ();
 sg13g2_fill_1 FILLER_55_1479 ();
 sg13g2_decap_8 FILLER_55_1492 ();
 sg13g2_fill_2 FILLER_55_1499 ();
 sg13g2_fill_1 FILLER_55_1501 ();
 sg13g2_fill_2 FILLER_55_1528 ();
 sg13g2_fill_1 FILLER_55_1530 ();
 sg13g2_fill_1 FILLER_55_1535 ();
 sg13g2_decap_8 FILLER_55_1540 ();
 sg13g2_decap_8 FILLER_55_1547 ();
 sg13g2_decap_8 FILLER_55_1554 ();
 sg13g2_fill_2 FILLER_55_1561 ();
 sg13g2_fill_1 FILLER_55_1563 ();
 sg13g2_fill_1 FILLER_55_1597 ();
 sg13g2_decap_8 FILLER_55_1608 ();
 sg13g2_decap_8 FILLER_55_1615 ();
 sg13g2_fill_1 FILLER_55_1622 ();
 sg13g2_fill_2 FILLER_55_1658 ();
 sg13g2_fill_1 FILLER_55_1660 ();
 sg13g2_decap_8 FILLER_55_1680 ();
 sg13g2_decap_8 FILLER_55_1687 ();
 sg13g2_fill_2 FILLER_55_1694 ();
 sg13g2_decap_8 FILLER_55_1714 ();
 sg13g2_decap_8 FILLER_55_1721 ();
 sg13g2_fill_2 FILLER_55_1733 ();
 sg13g2_fill_1 FILLER_55_1746 ();
 sg13g2_decap_4 FILLER_55_1770 ();
 sg13g2_fill_1 FILLER_55_1774 ();
 sg13g2_decap_8 FILLER_55_1780 ();
 sg13g2_fill_2 FILLER_55_1787 ();
 sg13g2_fill_1 FILLER_55_1789 ();
 sg13g2_fill_1 FILLER_55_1799 ();
 sg13g2_fill_1 FILLER_55_1809 ();
 sg13g2_fill_1 FILLER_55_1818 ();
 sg13g2_fill_1 FILLER_55_1836 ();
 sg13g2_decap_8 FILLER_55_1846 ();
 sg13g2_decap_4 FILLER_55_1853 ();
 sg13g2_fill_2 FILLER_55_1857 ();
 sg13g2_decap_4 FILLER_55_1865 ();
 sg13g2_fill_2 FILLER_55_1869 ();
 sg13g2_decap_8 FILLER_55_1879 ();
 sg13g2_fill_2 FILLER_55_1886 ();
 sg13g2_fill_1 FILLER_55_1894 ();
 sg13g2_fill_2 FILLER_55_1900 ();
 sg13g2_fill_1 FILLER_55_1916 ();
 sg13g2_fill_2 FILLER_55_1921 ();
 sg13g2_decap_8 FILLER_55_1928 ();
 sg13g2_decap_8 FILLER_55_1935 ();
 sg13g2_decap_8 FILLER_55_1942 ();
 sg13g2_decap_8 FILLER_55_1949 ();
 sg13g2_fill_2 FILLER_55_1956 ();
 sg13g2_fill_1 FILLER_55_1958 ();
 sg13g2_decap_8 FILLER_55_1969 ();
 sg13g2_fill_2 FILLER_55_1976 ();
 sg13g2_fill_1 FILLER_55_1978 ();
 sg13g2_decap_4 FILLER_55_1984 ();
 sg13g2_fill_1 FILLER_55_1988 ();
 sg13g2_fill_1 FILLER_55_1994 ();
 sg13g2_decap_8 FILLER_55_1999 ();
 sg13g2_decap_8 FILLER_55_2006 ();
 sg13g2_decap_4 FILLER_55_2013 ();
 sg13g2_decap_8 FILLER_55_2053 ();
 sg13g2_decap_8 FILLER_55_2060 ();
 sg13g2_decap_8 FILLER_55_2067 ();
 sg13g2_decap_8 FILLER_55_2074 ();
 sg13g2_decap_8 FILLER_55_2081 ();
 sg13g2_fill_2 FILLER_55_2088 ();
 sg13g2_fill_1 FILLER_55_2116 ();
 sg13g2_fill_2 FILLER_55_2147 ();
 sg13g2_fill_1 FILLER_55_2149 ();
 sg13g2_fill_1 FILLER_55_2176 ();
 sg13g2_fill_1 FILLER_55_2185 ();
 sg13g2_fill_1 FILLER_55_2202 ();
 sg13g2_fill_2 FILLER_55_2234 ();
 sg13g2_fill_2 FILLER_55_2275 ();
 sg13g2_fill_1 FILLER_55_2331 ();
 sg13g2_fill_1 FILLER_55_2337 ();
 sg13g2_fill_1 FILLER_55_2369 ();
 sg13g2_fill_1 FILLER_55_2450 ();
 sg13g2_fill_2 FILLER_55_2461 ();
 sg13g2_decap_8 FILLER_55_2492 ();
 sg13g2_fill_1 FILLER_55_2499 ();
 sg13g2_fill_2 FILLER_55_2520 ();
 sg13g2_fill_2 FILLER_55_2526 ();
 sg13g2_fill_1 FILLER_55_2528 ();
 sg13g2_fill_2 FILLER_55_2535 ();
 sg13g2_fill_2 FILLER_55_2563 ();
 sg13g2_fill_1 FILLER_55_2571 ();
 sg13g2_fill_1 FILLER_55_2577 ();
 sg13g2_decap_8 FILLER_55_2653 ();
 sg13g2_decap_8 FILLER_55_2660 ();
 sg13g2_fill_2 FILLER_55_2667 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_1 FILLER_56_44 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_2 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_134 ();
 sg13g2_fill_2 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_143 ();
 sg13g2_decap_4 FILLER_56_152 ();
 sg13g2_decap_8 FILLER_56_166 ();
 sg13g2_fill_2 FILLER_56_173 ();
 sg13g2_decap_4 FILLER_56_179 ();
 sg13g2_fill_1 FILLER_56_223 ();
 sg13g2_fill_1 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_377 ();
 sg13g2_fill_2 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_fill_1 FILLER_56_404 ();
 sg13g2_fill_2 FILLER_56_428 ();
 sg13g2_fill_1 FILLER_56_430 ();
 sg13g2_fill_2 FILLER_56_456 ();
 sg13g2_fill_2 FILLER_56_462 ();
 sg13g2_fill_2 FILLER_56_499 ();
 sg13g2_decap_8 FILLER_56_546 ();
 sg13g2_decap_4 FILLER_56_553 ();
 sg13g2_fill_2 FILLER_56_557 ();
 sg13g2_fill_2 FILLER_56_569 ();
 sg13g2_fill_1 FILLER_56_571 ();
 sg13g2_fill_2 FILLER_56_591 ();
 sg13g2_fill_2 FILLER_56_615 ();
 sg13g2_decap_4 FILLER_56_652 ();
 sg13g2_fill_2 FILLER_56_670 ();
 sg13g2_decap_8 FILLER_56_681 ();
 sg13g2_decap_8 FILLER_56_688 ();
 sg13g2_decap_4 FILLER_56_695 ();
 sg13g2_fill_2 FILLER_56_699 ();
 sg13g2_fill_2 FILLER_56_705 ();
 sg13g2_fill_1 FILLER_56_763 ();
 sg13g2_decap_4 FILLER_56_767 ();
 sg13g2_fill_2 FILLER_56_771 ();
 sg13g2_fill_2 FILLER_56_805 ();
 sg13g2_fill_1 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_813 ();
 sg13g2_fill_2 FILLER_56_820 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_870 ();
 sg13g2_fill_2 FILLER_56_885 ();
 sg13g2_fill_1 FILLER_56_887 ();
 sg13g2_fill_1 FILLER_56_893 ();
 sg13g2_fill_1 FILLER_56_924 ();
 sg13g2_fill_1 FILLER_56_934 ();
 sg13g2_fill_1 FILLER_56_952 ();
 sg13g2_fill_2 FILLER_56_1002 ();
 sg13g2_fill_1 FILLER_56_1090 ();
 sg13g2_fill_2 FILLER_56_1100 ();
 sg13g2_fill_2 FILLER_56_1119 ();
 sg13g2_fill_1 FILLER_56_1126 ();
 sg13g2_fill_1 FILLER_56_1135 ();
 sg13g2_fill_1 FILLER_56_1149 ();
 sg13g2_fill_1 FILLER_56_1159 ();
 sg13g2_fill_1 FILLER_56_1165 ();
 sg13g2_fill_1 FILLER_56_1172 ();
 sg13g2_fill_1 FILLER_56_1196 ();
 sg13g2_decap_8 FILLER_56_1207 ();
 sg13g2_decap_8 FILLER_56_1265 ();
 sg13g2_decap_4 FILLER_56_1272 ();
 sg13g2_fill_2 FILLER_56_1276 ();
 sg13g2_fill_1 FILLER_56_1304 ();
 sg13g2_fill_2 FILLER_56_1308 ();
 sg13g2_fill_1 FILLER_56_1335 ();
 sg13g2_fill_1 FILLER_56_1356 ();
 sg13g2_fill_2 FILLER_56_1361 ();
 sg13g2_fill_1 FILLER_56_1381 ();
 sg13g2_fill_2 FILLER_56_1409 ();
 sg13g2_decap_8 FILLER_56_1415 ();
 sg13g2_fill_1 FILLER_56_1422 ();
 sg13g2_fill_2 FILLER_56_1427 ();
 sg13g2_fill_1 FILLER_56_1429 ();
 sg13g2_fill_1 FILLER_56_1448 ();
 sg13g2_fill_1 FILLER_56_1471 ();
 sg13g2_fill_1 FILLER_56_1477 ();
 sg13g2_fill_1 FILLER_56_1484 ();
 sg13g2_fill_1 FILLER_56_1489 ();
 sg13g2_fill_2 FILLER_56_1516 ();
 sg13g2_decap_8 FILLER_56_1523 ();
 sg13g2_fill_2 FILLER_56_1530 ();
 sg13g2_fill_1 FILLER_56_1532 ();
 sg13g2_fill_1 FILLER_56_1547 ();
 sg13g2_fill_2 FILLER_56_1561 ();
 sg13g2_fill_1 FILLER_56_1568 ();
 sg13g2_fill_2 FILLER_56_1591 ();
 sg13g2_decap_8 FILLER_56_1598 ();
 sg13g2_decap_4 FILLER_56_1605 ();
 sg13g2_fill_1 FILLER_56_1609 ();
 sg13g2_decap_8 FILLER_56_1614 ();
 sg13g2_decap_8 FILLER_56_1621 ();
 sg13g2_fill_2 FILLER_56_1628 ();
 sg13g2_fill_1 FILLER_56_1630 ();
 sg13g2_decap_8 FILLER_56_1635 ();
 sg13g2_decap_8 FILLER_56_1642 ();
 sg13g2_fill_2 FILLER_56_1665 ();
 sg13g2_fill_1 FILLER_56_1667 ();
 sg13g2_fill_1 FILLER_56_1673 ();
 sg13g2_decap_4 FILLER_56_1679 ();
 sg13g2_fill_2 FILLER_56_1683 ();
 sg13g2_decap_4 FILLER_56_1689 ();
 sg13g2_decap_4 FILLER_56_1698 ();
 sg13g2_fill_1 FILLER_56_1702 ();
 sg13g2_decap_4 FILLER_56_1708 ();
 sg13g2_fill_1 FILLER_56_1712 ();
 sg13g2_decap_4 FILLER_56_1718 ();
 sg13g2_fill_2 FILLER_56_1722 ();
 sg13g2_decap_8 FILLER_56_1750 ();
 sg13g2_fill_2 FILLER_56_1757 ();
 sg13g2_decap_8 FILLER_56_1770 ();
 sg13g2_decap_8 FILLER_56_1777 ();
 sg13g2_fill_1 FILLER_56_1784 ();
 sg13g2_fill_1 FILLER_56_1804 ();
 sg13g2_decap_8 FILLER_56_1810 ();
 sg13g2_decap_4 FILLER_56_1817 ();
 sg13g2_fill_2 FILLER_56_1821 ();
 sg13g2_fill_2 FILLER_56_1833 ();
 sg13g2_decap_8 FILLER_56_1839 ();
 sg13g2_decap_4 FILLER_56_1846 ();
 sg13g2_fill_1 FILLER_56_1856 ();
 sg13g2_decap_4 FILLER_56_1862 ();
 sg13g2_decap_8 FILLER_56_1870 ();
 sg13g2_fill_2 FILLER_56_1882 ();
 sg13g2_fill_1 FILLER_56_1884 ();
 sg13g2_fill_2 FILLER_56_1894 ();
 sg13g2_fill_1 FILLER_56_1901 ();
 sg13g2_fill_1 FILLER_56_1912 ();
 sg13g2_fill_1 FILLER_56_1917 ();
 sg13g2_decap_4 FILLER_56_1922 ();
 sg13g2_decap_8 FILLER_56_1930 ();
 sg13g2_decap_8 FILLER_56_1937 ();
 sg13g2_decap_8 FILLER_56_1944 ();
 sg13g2_decap_8 FILLER_56_1951 ();
 sg13g2_decap_8 FILLER_56_1958 ();
 sg13g2_decap_8 FILLER_56_1965 ();
 sg13g2_decap_8 FILLER_56_1972 ();
 sg13g2_decap_8 FILLER_56_1979 ();
 sg13g2_fill_2 FILLER_56_1986 ();
 sg13g2_fill_1 FILLER_56_1988 ();
 sg13g2_decap_8 FILLER_56_1993 ();
 sg13g2_decap_8 FILLER_56_2000 ();
 sg13g2_decap_8 FILLER_56_2007 ();
 sg13g2_decap_4 FILLER_56_2014 ();
 sg13g2_decap_4 FILLER_56_2023 ();
 sg13g2_fill_1 FILLER_56_2027 ();
 sg13g2_decap_8 FILLER_56_2052 ();
 sg13g2_decap_8 FILLER_56_2059 ();
 sg13g2_decap_8 FILLER_56_2066 ();
 sg13g2_decap_8 FILLER_56_2073 ();
 sg13g2_decap_8 FILLER_56_2080 ();
 sg13g2_fill_2 FILLER_56_2117 ();
 sg13g2_fill_1 FILLER_56_2119 ();
 sg13g2_fill_1 FILLER_56_2146 ();
 sg13g2_fill_2 FILLER_56_2153 ();
 sg13g2_fill_1 FILLER_56_2159 ();
 sg13g2_decap_4 FILLER_56_2174 ();
 sg13g2_fill_2 FILLER_56_2229 ();
 sg13g2_fill_2 FILLER_56_2244 ();
 sg13g2_decap_8 FILLER_56_2266 ();
 sg13g2_fill_2 FILLER_56_2273 ();
 sg13g2_fill_1 FILLER_56_2326 ();
 sg13g2_fill_1 FILLER_56_2334 ();
 sg13g2_fill_2 FILLER_56_2361 ();
 sg13g2_fill_1 FILLER_56_2377 ();
 sg13g2_fill_2 FILLER_56_2439 ();
 sg13g2_fill_1 FILLER_56_2481 ();
 sg13g2_fill_1 FILLER_56_2486 ();
 sg13g2_fill_1 FILLER_56_2522 ();
 sg13g2_fill_2 FILLER_56_2529 ();
 sg13g2_fill_2 FILLER_56_2541 ();
 sg13g2_fill_2 FILLER_56_2547 ();
 sg13g2_fill_1 FILLER_56_2549 ();
 sg13g2_fill_1 FILLER_56_2554 ();
 sg13g2_fill_1 FILLER_56_2581 ();
 sg13g2_fill_1 FILLER_56_2587 ();
 sg13g2_decap_8 FILLER_56_2650 ();
 sg13g2_decap_8 FILLER_56_2657 ();
 sg13g2_decap_4 FILLER_56_2664 ();
 sg13g2_fill_2 FILLER_56_2668 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_fill_1 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_208 ();
 sg13g2_fill_1 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_218 ();
 sg13g2_fill_2 FILLER_57_224 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_fill_1 FILLER_57_337 ();
 sg13g2_fill_2 FILLER_57_342 ();
 sg13g2_fill_2 FILLER_57_392 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_2 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_467 ();
 sg13g2_fill_1 FILLER_57_493 ();
 sg13g2_fill_2 FILLER_57_508 ();
 sg13g2_fill_2 FILLER_57_521 ();
 sg13g2_decap_8 FILLER_57_558 ();
 sg13g2_decap_4 FILLER_57_565 ();
 sg13g2_fill_1 FILLER_57_569 ();
 sg13g2_fill_1 FILLER_57_574 ();
 sg13g2_fill_2 FILLER_57_588 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_fill_2 FILLER_57_650 ();
 sg13g2_fill_1 FILLER_57_687 ();
 sg13g2_fill_2 FILLER_57_737 ();
 sg13g2_fill_1 FILLER_57_739 ();
 sg13g2_fill_1 FILLER_57_745 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_fill_1 FILLER_57_772 ();
 sg13g2_fill_1 FILLER_57_823 ();
 sg13g2_fill_1 FILLER_57_889 ();
 sg13g2_decap_4 FILLER_57_898 ();
 sg13g2_fill_1 FILLER_57_915 ();
 sg13g2_fill_1 FILLER_57_930 ();
 sg13g2_fill_1 FILLER_57_970 ();
 sg13g2_fill_1 FILLER_57_1103 ();
 sg13g2_fill_2 FILLER_57_1114 ();
 sg13g2_fill_1 FILLER_57_1125 ();
 sg13g2_fill_1 FILLER_57_1131 ();
 sg13g2_fill_1 FILLER_57_1138 ();
 sg13g2_decap_4 FILLER_57_1196 ();
 sg13g2_fill_1 FILLER_57_1200 ();
 sg13g2_decap_8 FILLER_57_1207 ();
 sg13g2_decap_8 FILLER_57_1214 ();
 sg13g2_fill_2 FILLER_57_1221 ();
 sg13g2_fill_2 FILLER_57_1290 ();
 sg13g2_fill_2 FILLER_57_1331 ();
 sg13g2_fill_1 FILLER_57_1333 ();
 sg13g2_decap_8 FILLER_57_1342 ();
 sg13g2_fill_2 FILLER_57_1356 ();
 sg13g2_fill_1 FILLER_57_1358 ();
 sg13g2_fill_2 FILLER_57_1388 ();
 sg13g2_fill_1 FILLER_57_1390 ();
 sg13g2_fill_2 FILLER_57_1397 ();
 sg13g2_fill_2 FILLER_57_1407 ();
 sg13g2_fill_2 FILLER_57_1413 ();
 sg13g2_decap_4 FILLER_57_1418 ();
 sg13g2_fill_2 FILLER_57_1422 ();
 sg13g2_fill_1 FILLER_57_1428 ();
 sg13g2_fill_2 FILLER_57_1434 ();
 sg13g2_fill_1 FILLER_57_1442 ();
 sg13g2_fill_1 FILLER_57_1455 ();
 sg13g2_fill_1 FILLER_57_1470 ();
 sg13g2_decap_8 FILLER_57_1483 ();
 sg13g2_fill_1 FILLER_57_1510 ();
 sg13g2_decap_8 FILLER_57_1520 ();
 sg13g2_fill_1 FILLER_57_1527 ();
 sg13g2_decap_4 FILLER_57_1532 ();
 sg13g2_fill_2 FILLER_57_1571 ();
 sg13g2_decap_8 FILLER_57_1603 ();
 sg13g2_decap_8 FILLER_57_1610 ();
 sg13g2_decap_4 FILLER_57_1625 ();
 sg13g2_decap_8 FILLER_57_1633 ();
 sg13g2_decap_8 FILLER_57_1647 ();
 sg13g2_decap_8 FILLER_57_1669 ();
 sg13g2_fill_2 FILLER_57_1676 ();
 sg13g2_fill_1 FILLER_57_1678 ();
 sg13g2_fill_1 FILLER_57_1694 ();
 sg13g2_decap_8 FILLER_57_1699 ();
 sg13g2_decap_8 FILLER_57_1710 ();
 sg13g2_fill_2 FILLER_57_1717 ();
 sg13g2_decap_8 FILLER_57_1763 ();
 sg13g2_decap_8 FILLER_57_1770 ();
 sg13g2_fill_2 FILLER_57_1777 ();
 sg13g2_fill_1 FILLER_57_1779 ();
 sg13g2_decap_8 FILLER_57_1785 ();
 sg13g2_decap_8 FILLER_57_1792 ();
 sg13g2_decap_8 FILLER_57_1799 ();
 sg13g2_fill_2 FILLER_57_1806 ();
 sg13g2_fill_1 FILLER_57_1808 ();
 sg13g2_fill_1 FILLER_57_1813 ();
 sg13g2_decap_8 FILLER_57_1822 ();
 sg13g2_fill_2 FILLER_57_1829 ();
 sg13g2_decap_8 FILLER_57_1836 ();
 sg13g2_decap_8 FILLER_57_1843 ();
 sg13g2_decap_8 FILLER_57_1850 ();
 sg13g2_fill_1 FILLER_57_1857 ();
 sg13g2_decap_4 FILLER_57_1863 ();
 sg13g2_fill_1 FILLER_57_1875 ();
 sg13g2_fill_1 FILLER_57_1881 ();
 sg13g2_fill_2 FILLER_57_1896 ();
 sg13g2_fill_2 FILLER_57_1902 ();
 sg13g2_fill_1 FILLER_57_1913 ();
 sg13g2_decap_8 FILLER_57_1929 ();
 sg13g2_fill_1 FILLER_57_1936 ();
 sg13g2_decap_4 FILLER_57_1942 ();
 sg13g2_decap_8 FILLER_57_1950 ();
 sg13g2_decap_8 FILLER_57_1965 ();
 sg13g2_decap_8 FILLER_57_1972 ();
 sg13g2_decap_8 FILLER_57_1979 ();
 sg13g2_decap_8 FILLER_57_1986 ();
 sg13g2_fill_1 FILLER_57_1993 ();
 sg13g2_decap_8 FILLER_57_2002 ();
 sg13g2_decap_8 FILLER_57_2009 ();
 sg13g2_fill_2 FILLER_57_2016 ();
 sg13g2_decap_8 FILLER_57_2031 ();
 sg13g2_fill_1 FILLER_57_2038 ();
 sg13g2_decap_8 FILLER_57_2044 ();
 sg13g2_decap_8 FILLER_57_2051 ();
 sg13g2_decap_8 FILLER_57_2058 ();
 sg13g2_decap_8 FILLER_57_2065 ();
 sg13g2_decap_8 FILLER_57_2072 ();
 sg13g2_decap_4 FILLER_57_2079 ();
 sg13g2_fill_2 FILLER_57_2083 ();
 sg13g2_fill_2 FILLER_57_2102 ();
 sg13g2_fill_2 FILLER_57_2113 ();
 sg13g2_fill_1 FILLER_57_2121 ();
 sg13g2_fill_1 FILLER_57_2156 ();
 sg13g2_fill_1 FILLER_57_2206 ();
 sg13g2_fill_2 FILLER_57_2220 ();
 sg13g2_fill_1 FILLER_57_2227 ();
 sg13g2_fill_2 FILLER_57_2307 ();
 sg13g2_fill_2 FILLER_57_2312 ();
 sg13g2_decap_8 FILLER_57_2432 ();
 sg13g2_decap_8 FILLER_57_2439 ();
 sg13g2_fill_2 FILLER_57_2446 ();
 sg13g2_decap_8 FILLER_57_2461 ();
 sg13g2_fill_1 FILLER_57_2468 ();
 sg13g2_decap_8 FILLER_57_2474 ();
 sg13g2_decap_4 FILLER_57_2481 ();
 sg13g2_fill_2 FILLER_57_2485 ();
 sg13g2_decap_8 FILLER_57_2514 ();
 sg13g2_decap_8 FILLER_57_2521 ();
 sg13g2_fill_1 FILLER_57_2528 ();
 sg13g2_decap_8 FILLER_57_2533 ();
 sg13g2_decap_4 FILLER_57_2540 ();
 sg13g2_fill_1 FILLER_57_2572 ();
 sg13g2_fill_2 FILLER_57_2577 ();
 sg13g2_fill_1 FILLER_57_2579 ();
 sg13g2_fill_2 FILLER_57_2585 ();
 sg13g2_fill_1 FILLER_57_2591 ();
 sg13g2_decap_8 FILLER_57_2598 ();
 sg13g2_fill_1 FILLER_57_2605 ();
 sg13g2_decap_8 FILLER_57_2624 ();
 sg13g2_fill_1 FILLER_57_2631 ();
 sg13g2_decap_8 FILLER_57_2636 ();
 sg13g2_decap_8 FILLER_57_2643 ();
 sg13g2_decap_8 FILLER_57_2650 ();
 sg13g2_decap_8 FILLER_57_2657 ();
 sg13g2_decap_4 FILLER_57_2664 ();
 sg13g2_fill_2 FILLER_57_2668 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_fill_2 FILLER_58_136 ();
 sg13g2_fill_2 FILLER_58_143 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_fill_1 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_fill_1 FILLER_58_387 ();
 sg13g2_fill_1 FILLER_58_414 ();
 sg13g2_fill_1 FILLER_58_474 ();
 sg13g2_fill_2 FILLER_58_485 ();
 sg13g2_fill_2 FILLER_58_510 ();
 sg13g2_fill_2 FILLER_58_542 ();
 sg13g2_fill_2 FILLER_58_550 ();
 sg13g2_fill_1 FILLER_58_558 ();
 sg13g2_decap_4 FILLER_58_565 ();
 sg13g2_fill_1 FILLER_58_595 ();
 sg13g2_fill_2 FILLER_58_609 ();
 sg13g2_fill_1 FILLER_58_626 ();
 sg13g2_fill_1 FILLER_58_681 ();
 sg13g2_fill_1 FILLER_58_687 ();
 sg13g2_fill_1 FILLER_58_693 ();
 sg13g2_fill_1 FILLER_58_698 ();
 sg13g2_fill_2 FILLER_58_730 ();
 sg13g2_fill_2 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_769 ();
 sg13g2_fill_1 FILLER_58_775 ();
 sg13g2_fill_2 FILLER_58_826 ();
 sg13g2_fill_1 FILLER_58_828 ();
 sg13g2_fill_1 FILLER_58_834 ();
 sg13g2_decap_8 FILLER_58_839 ();
 sg13g2_fill_2 FILLER_58_861 ();
 sg13g2_fill_2 FILLER_58_868 ();
 sg13g2_fill_1 FILLER_58_870 ();
 sg13g2_fill_2 FILLER_58_903 ();
 sg13g2_fill_1 FILLER_58_905 ();
 sg13g2_decap_8 FILLER_58_910 ();
 sg13g2_decap_4 FILLER_58_925 ();
 sg13g2_fill_1 FILLER_58_929 ();
 sg13g2_fill_1 FILLER_58_960 ();
 sg13g2_fill_2 FILLER_58_974 ();
 sg13g2_fill_2 FILLER_58_992 ();
 sg13g2_fill_1 FILLER_58_1013 ();
 sg13g2_fill_1 FILLER_58_1040 ();
 sg13g2_fill_2 FILLER_58_1076 ();
 sg13g2_fill_1 FILLER_58_1078 ();
 sg13g2_fill_1 FILLER_58_1110 ();
 sg13g2_fill_1 FILLER_58_1116 ();
 sg13g2_fill_1 FILLER_58_1151 ();
 sg13g2_fill_2 FILLER_58_1235 ();
 sg13g2_decap_8 FILLER_58_1291 ();
 sg13g2_fill_1 FILLER_58_1298 ();
 sg13g2_fill_1 FILLER_58_1328 ();
 sg13g2_fill_1 FILLER_58_1352 ();
 sg13g2_decap_4 FILLER_58_1374 ();
 sg13g2_fill_2 FILLER_58_1378 ();
 sg13g2_fill_1 FILLER_58_1393 ();
 sg13g2_fill_2 FILLER_58_1403 ();
 sg13g2_fill_1 FILLER_58_1405 ();
 sg13g2_fill_2 FILLER_58_1455 ();
 sg13g2_fill_1 FILLER_58_1467 ();
 sg13g2_fill_2 FILLER_58_1474 ();
 sg13g2_decap_8 FILLER_58_1486 ();
 sg13g2_decap_8 FILLER_58_1493 ();
 sg13g2_decap_8 FILLER_58_1500 ();
 sg13g2_decap_4 FILLER_58_1507 ();
 sg13g2_fill_1 FILLER_58_1511 ();
 sg13g2_fill_2 FILLER_58_1530 ();
 sg13g2_fill_1 FILLER_58_1547 ();
 sg13g2_fill_1 FILLER_58_1562 ();
 sg13g2_fill_1 FILLER_58_1567 ();
 sg13g2_fill_2 FILLER_58_1621 ();
 sg13g2_fill_1 FILLER_58_1623 ();
 sg13g2_decap_4 FILLER_58_1640 ();
 sg13g2_fill_2 FILLER_58_1644 ();
 sg13g2_fill_1 FILLER_58_1653 ();
 sg13g2_fill_1 FILLER_58_1659 ();
 sg13g2_fill_2 FILLER_58_1665 ();
 sg13g2_fill_2 FILLER_58_1672 ();
 sg13g2_fill_1 FILLER_58_1691 ();
 sg13g2_decap_8 FILLER_58_1695 ();
 sg13g2_decap_8 FILLER_58_1702 ();
 sg13g2_fill_2 FILLER_58_1709 ();
 sg13g2_fill_1 FILLER_58_1711 ();
 sg13g2_decap_4 FILLER_58_1738 ();
 sg13g2_decap_8 FILLER_58_1746 ();
 sg13g2_decap_4 FILLER_58_1765 ();
 sg13g2_fill_1 FILLER_58_1773 ();
 sg13g2_decap_8 FILLER_58_1789 ();
 sg13g2_decap_8 FILLER_58_1796 ();
 sg13g2_decap_4 FILLER_58_1811 ();
 sg13g2_fill_2 FILLER_58_1815 ();
 sg13g2_decap_4 FILLER_58_1821 ();
 sg13g2_fill_2 FILLER_58_1825 ();
 sg13g2_decap_8 FILLER_58_1832 ();
 sg13g2_fill_1 FILLER_58_1839 ();
 sg13g2_decap_8 FILLER_58_1851 ();
 sg13g2_decap_8 FILLER_58_1858 ();
 sg13g2_fill_2 FILLER_58_1869 ();
 sg13g2_fill_1 FILLER_58_1871 ();
 sg13g2_decap_4 FILLER_58_1881 ();
 sg13g2_fill_1 FILLER_58_1885 ();
 sg13g2_fill_2 FILLER_58_1908 ();
 sg13g2_decap_8 FILLER_58_1931 ();
 sg13g2_decap_8 FILLER_58_1938 ();
 sg13g2_decap_4 FILLER_58_1945 ();
 sg13g2_fill_1 FILLER_58_1949 ();
 sg13g2_decap_8 FILLER_58_1955 ();
 sg13g2_fill_2 FILLER_58_1962 ();
 sg13g2_decap_8 FILLER_58_1969 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_decap_8 FILLER_58_1988 ();
 sg13g2_decap_8 FILLER_58_1995 ();
 sg13g2_decap_8 FILLER_58_2002 ();
 sg13g2_decap_8 FILLER_58_2009 ();
 sg13g2_decap_8 FILLER_58_2016 ();
 sg13g2_fill_1 FILLER_58_2023 ();
 sg13g2_decap_8 FILLER_58_2032 ();
 sg13g2_decap_8 FILLER_58_2039 ();
 sg13g2_decap_8 FILLER_58_2046 ();
 sg13g2_decap_8 FILLER_58_2053 ();
 sg13g2_decap_8 FILLER_58_2060 ();
 sg13g2_decap_8 FILLER_58_2067 ();
 sg13g2_decap_8 FILLER_58_2074 ();
 sg13g2_decap_4 FILLER_58_2081 ();
 sg13g2_fill_2 FILLER_58_2085 ();
 sg13g2_decap_8 FILLER_58_2092 ();
 sg13g2_decap_8 FILLER_58_2099 ();
 sg13g2_decap_8 FILLER_58_2106 ();
 sg13g2_fill_2 FILLER_58_2113 ();
 sg13g2_fill_1 FILLER_58_2130 ();
 sg13g2_fill_2 FILLER_58_2160 ();
 sg13g2_fill_2 FILLER_58_2269 ();
 sg13g2_fill_2 FILLER_58_2315 ();
 sg13g2_fill_2 FILLER_58_2460 ();
 sg13g2_fill_2 FILLER_58_2476 ();
 sg13g2_fill_1 FILLER_58_2478 ();
 sg13g2_fill_1 FILLER_58_2496 ();
 sg13g2_decap_4 FILLER_58_2525 ();
 sg13g2_fill_1 FILLER_58_2529 ();
 sg13g2_decap_8 FILLER_58_2534 ();
 sg13g2_decap_8 FILLER_58_2571 ();
 sg13g2_fill_2 FILLER_58_2578 ();
 sg13g2_fill_1 FILLER_58_2580 ();
 sg13g2_fill_2 FILLER_58_2587 ();
 sg13g2_decap_4 FILLER_58_2593 ();
 sg13g2_fill_1 FILLER_58_2597 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_decap_8 FILLER_58_2622 ();
 sg13g2_decap_8 FILLER_58_2629 ();
 sg13g2_decap_8 FILLER_58_2636 ();
 sg13g2_decap_8 FILLER_58_2643 ();
 sg13g2_decap_8 FILLER_58_2650 ();
 sg13g2_decap_8 FILLER_58_2657 ();
 sg13g2_decap_4 FILLER_58_2664 ();
 sg13g2_fill_2 FILLER_58_2668 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_38 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_fill_1 FILLER_59_52 ();
 sg13g2_fill_1 FILLER_59_75 ();
 sg13g2_fill_2 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_fill_1 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_decap_8 FILLER_59_250 ();
 sg13g2_decap_4 FILLER_59_257 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_decap_8 FILLER_59_270 ();
 sg13g2_fill_2 FILLER_59_277 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_317 ();
 sg13g2_fill_2 FILLER_59_345 ();
 sg13g2_decap_4 FILLER_59_374 ();
 sg13g2_decap_4 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_480 ();
 sg13g2_fill_1 FILLER_59_497 ();
 sg13g2_fill_1 FILLER_59_547 ();
 sg13g2_decap_8 FILLER_59_564 ();
 sg13g2_fill_2 FILLER_59_606 ();
 sg13g2_decap_8 FILLER_59_639 ();
 sg13g2_fill_2 FILLER_59_646 ();
 sg13g2_fill_1 FILLER_59_648 ();
 sg13g2_fill_2 FILLER_59_659 ();
 sg13g2_fill_1 FILLER_59_661 ();
 sg13g2_decap_4 FILLER_59_670 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_fill_2 FILLER_59_684 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_fill_2 FILLER_59_710 ();
 sg13g2_fill_2 FILLER_59_736 ();
 sg13g2_fill_1 FILLER_59_738 ();
 sg13g2_fill_1 FILLER_59_744 ();
 sg13g2_fill_2 FILLER_59_773 ();
 sg13g2_fill_1 FILLER_59_775 ();
 sg13g2_fill_2 FILLER_59_784 ();
 sg13g2_fill_1 FILLER_59_815 ();
 sg13g2_decap_8 FILLER_59_842 ();
 sg13g2_fill_2 FILLER_59_891 ();
 sg13g2_fill_1 FILLER_59_908 ();
 sg13g2_fill_1 FILLER_59_913 ();
 sg13g2_fill_1 FILLER_59_920 ();
 sg13g2_fill_1 FILLER_59_927 ();
 sg13g2_fill_1 FILLER_59_936 ();
 sg13g2_fill_2 FILLER_59_946 ();
 sg13g2_fill_1 FILLER_59_948 ();
 sg13g2_fill_1 FILLER_59_975 ();
 sg13g2_fill_1 FILLER_59_1019 ();
 sg13g2_fill_2 FILLER_59_1064 ();
 sg13g2_fill_1 FILLER_59_1066 ();
 sg13g2_fill_2 FILLER_59_1085 ();
 sg13g2_fill_2 FILLER_59_1142 ();
 sg13g2_decap_4 FILLER_59_1174 ();
 sg13g2_fill_1 FILLER_59_1178 ();
 sg13g2_fill_2 FILLER_59_1188 ();
 sg13g2_fill_1 FILLER_59_1190 ();
 sg13g2_decap_4 FILLER_59_1199 ();
 sg13g2_fill_1 FILLER_59_1203 ();
 sg13g2_fill_2 FILLER_59_1214 ();
 sg13g2_decap_8 FILLER_59_1242 ();
 sg13g2_fill_2 FILLER_59_1249 ();
 sg13g2_decap_8 FILLER_59_1289 ();
 sg13g2_decap_8 FILLER_59_1296 ();
 sg13g2_fill_1 FILLER_59_1303 ();
 sg13g2_fill_1 FILLER_59_1312 ();
 sg13g2_decap_4 FILLER_59_1338 ();
 sg13g2_fill_1 FILLER_59_1342 ();
 sg13g2_fill_1 FILLER_59_1348 ();
 sg13g2_fill_1 FILLER_59_1354 ();
 sg13g2_fill_1 FILLER_59_1360 ();
 sg13g2_fill_2 FILLER_59_1377 ();
 sg13g2_fill_2 FILLER_59_1384 ();
 sg13g2_fill_1 FILLER_59_1386 ();
 sg13g2_fill_2 FILLER_59_1397 ();
 sg13g2_fill_2 FILLER_59_1408 ();
 sg13g2_fill_1 FILLER_59_1410 ();
 sg13g2_decap_8 FILLER_59_1423 ();
 sg13g2_fill_2 FILLER_59_1444 ();
 sg13g2_fill_1 FILLER_59_1466 ();
 sg13g2_decap_4 FILLER_59_1476 ();
 sg13g2_fill_1 FILLER_59_1480 ();
 sg13g2_decap_4 FILLER_59_1486 ();
 sg13g2_fill_2 FILLER_59_1513 ();
 sg13g2_fill_1 FILLER_59_1535 ();
 sg13g2_fill_1 FILLER_59_1542 ();
 sg13g2_decap_4 FILLER_59_1561 ();
 sg13g2_fill_1 FILLER_59_1565 ();
 sg13g2_fill_2 FILLER_59_1610 ();
 sg13g2_decap_8 FILLER_59_1651 ();
 sg13g2_decap_4 FILLER_59_1689 ();
 sg13g2_fill_1 FILLER_59_1693 ();
 sg13g2_decap_8 FILLER_59_1698 ();
 sg13g2_decap_4 FILLER_59_1705 ();
 sg13g2_fill_1 FILLER_59_1709 ();
 sg13g2_fill_2 FILLER_59_1714 ();
 sg13g2_fill_1 FILLER_59_1716 ();
 sg13g2_fill_1 FILLER_59_1763 ();
 sg13g2_fill_1 FILLER_59_1778 ();
 sg13g2_fill_1 FILLER_59_1792 ();
 sg13g2_decap_4 FILLER_59_1797 ();
 sg13g2_fill_2 FILLER_59_1801 ();
 sg13g2_decap_4 FILLER_59_1828 ();
 sg13g2_fill_1 FILLER_59_1832 ();
 sg13g2_decap_4 FILLER_59_1838 ();
 sg13g2_fill_2 FILLER_59_1842 ();
 sg13g2_fill_1 FILLER_59_1849 ();
 sg13g2_decap_8 FILLER_59_1853 ();
 sg13g2_decap_4 FILLER_59_1860 ();
 sg13g2_fill_1 FILLER_59_1864 ();
 sg13g2_fill_1 FILLER_59_1870 ();
 sg13g2_fill_2 FILLER_59_1886 ();
 sg13g2_fill_1 FILLER_59_1888 ();
 sg13g2_fill_2 FILLER_59_1894 ();
 sg13g2_decap_8 FILLER_59_1901 ();
 sg13g2_decap_8 FILLER_59_1908 ();
 sg13g2_decap_8 FILLER_59_1915 ();
 sg13g2_decap_8 FILLER_59_1927 ();
 sg13g2_decap_8 FILLER_59_1934 ();
 sg13g2_fill_2 FILLER_59_1941 ();
 sg13g2_fill_1 FILLER_59_1943 ();
 sg13g2_decap_8 FILLER_59_1948 ();
 sg13g2_decap_8 FILLER_59_1955 ();
 sg13g2_decap_8 FILLER_59_1962 ();
 sg13g2_decap_8 FILLER_59_1969 ();
 sg13g2_fill_1 FILLER_59_1976 ();
 sg13g2_decap_8 FILLER_59_1982 ();
 sg13g2_decap_8 FILLER_59_1989 ();
 sg13g2_decap_8 FILLER_59_1996 ();
 sg13g2_decap_8 FILLER_59_2003 ();
 sg13g2_decap_8 FILLER_59_2010 ();
 sg13g2_decap_8 FILLER_59_2017 ();
 sg13g2_decap_8 FILLER_59_2024 ();
 sg13g2_decap_8 FILLER_59_2037 ();
 sg13g2_decap_8 FILLER_59_2044 ();
 sg13g2_decap_8 FILLER_59_2051 ();
 sg13g2_decap_8 FILLER_59_2058 ();
 sg13g2_decap_8 FILLER_59_2065 ();
 sg13g2_decap_8 FILLER_59_2072 ();
 sg13g2_decap_8 FILLER_59_2079 ();
 sg13g2_decap_8 FILLER_59_2086 ();
 sg13g2_decap_4 FILLER_59_2093 ();
 sg13g2_fill_1 FILLER_59_2097 ();
 sg13g2_fill_2 FILLER_59_2107 ();
 sg13g2_fill_1 FILLER_59_2109 ();
 sg13g2_fill_2 FILLER_59_2114 ();
 sg13g2_decap_4 FILLER_59_2122 ();
 sg13g2_fill_2 FILLER_59_2139 ();
 sg13g2_fill_1 FILLER_59_2141 ();
 sg13g2_fill_2 FILLER_59_2152 ();
 sg13g2_fill_1 FILLER_59_2154 ();
 sg13g2_fill_2 FILLER_59_2180 ();
 sg13g2_fill_1 FILLER_59_2188 ();
 sg13g2_fill_2 FILLER_59_2193 ();
 sg13g2_fill_2 FILLER_59_2199 ();
 sg13g2_fill_2 FILLER_59_2209 ();
 sg13g2_fill_2 FILLER_59_2216 ();
 sg13g2_fill_2 FILLER_59_2226 ();
 sg13g2_fill_1 FILLER_59_2280 ();
 sg13g2_fill_2 FILLER_59_2285 ();
 sg13g2_fill_2 FILLER_59_2313 ();
 sg13g2_fill_1 FILLER_59_2328 ();
 sg13g2_fill_2 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2426 ();
 sg13g2_decap_4 FILLER_59_2433 ();
 sg13g2_fill_1 FILLER_59_2499 ();
 sg13g2_decap_8 FILLER_59_2530 ();
 sg13g2_fill_1 FILLER_59_2537 ();
 sg13g2_fill_2 FILLER_59_2570 ();
 sg13g2_decap_8 FILLER_59_2637 ();
 sg13g2_decap_8 FILLER_59_2644 ();
 sg13g2_decap_8 FILLER_59_2651 ();
 sg13g2_decap_8 FILLER_59_2658 ();
 sg13g2_decap_4 FILLER_59_2665 ();
 sg13g2_fill_1 FILLER_59_2669 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_24 ();
 sg13g2_fill_1 FILLER_60_33 ();
 sg13g2_fill_1 FILLER_60_39 ();
 sg13g2_decap_8 FILLER_60_44 ();
 sg13g2_decap_4 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_55 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_99 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_130 ();
 sg13g2_decap_4 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_145 ();
 sg13g2_decap_8 FILLER_60_152 ();
 sg13g2_fill_2 FILLER_60_159 ();
 sg13g2_fill_2 FILLER_60_221 ();
 sg13g2_fill_1 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_228 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_fill_2 FILLER_60_266 ();
 sg13g2_decap_4 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_276 ();
 sg13g2_decap_4 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_306 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_decap_8 FILLER_60_370 ();
 sg13g2_decap_8 FILLER_60_377 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_decap_4 FILLER_60_395 ();
 sg13g2_fill_1 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_414 ();
 sg13g2_fill_1 FILLER_60_416 ();
 sg13g2_fill_2 FILLER_60_421 ();
 sg13g2_fill_2 FILLER_60_522 ();
 sg13g2_fill_1 FILLER_60_529 ();
 sg13g2_fill_1 FILLER_60_556 ();
 sg13g2_fill_2 FILLER_60_561 ();
 sg13g2_fill_1 FILLER_60_563 ();
 sg13g2_fill_1 FILLER_60_568 ();
 sg13g2_fill_2 FILLER_60_582 ();
 sg13g2_fill_1 FILLER_60_584 ();
 sg13g2_decap_8 FILLER_60_629 ();
 sg13g2_fill_1 FILLER_60_636 ();
 sg13g2_fill_1 FILLER_60_641 ();
 sg13g2_decap_4 FILLER_60_648 ();
 sg13g2_decap_8 FILLER_60_656 ();
 sg13g2_decap_4 FILLER_60_663 ();
 sg13g2_decap_8 FILLER_60_683 ();
 sg13g2_decap_8 FILLER_60_690 ();
 sg13g2_fill_1 FILLER_60_697 ();
 sg13g2_fill_1 FILLER_60_702 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_fill_2 FILLER_60_714 ();
 sg13g2_fill_1 FILLER_60_716 ();
 sg13g2_fill_1 FILLER_60_722 ();
 sg13g2_fill_2 FILLER_60_732 ();
 sg13g2_fill_1 FILLER_60_734 ();
 sg13g2_fill_2 FILLER_60_781 ();
 sg13g2_fill_2 FILLER_60_808 ();
 sg13g2_fill_1 FILLER_60_825 ();
 sg13g2_fill_2 FILLER_60_831 ();
 sg13g2_fill_1 FILLER_60_930 ();
 sg13g2_fill_1 FILLER_60_975 ();
 sg13g2_fill_2 FILLER_60_1005 ();
 sg13g2_fill_1 FILLER_60_1057 ();
 sg13g2_fill_2 FILLER_60_1062 ();
 sg13g2_fill_1 FILLER_60_1064 ();
 sg13g2_fill_2 FILLER_60_1105 ();
 sg13g2_fill_1 FILLER_60_1115 ();
 sg13g2_fill_2 FILLER_60_1121 ();
 sg13g2_decap_8 FILLER_60_1134 ();
 sg13g2_fill_1 FILLER_60_1141 ();
 sg13g2_fill_1 FILLER_60_1155 ();
 sg13g2_fill_2 FILLER_60_1168 ();
 sg13g2_fill_2 FILLER_60_1173 ();
 sg13g2_fill_1 FILLER_60_1175 ();
 sg13g2_decap_4 FILLER_60_1186 ();
 sg13g2_fill_2 FILLER_60_1190 ();
 sg13g2_fill_2 FILLER_60_1196 ();
 sg13g2_decap_4 FILLER_60_1206 ();
 sg13g2_fill_1 FILLER_60_1228 ();
 sg13g2_fill_2 FILLER_60_1239 ();
 sg13g2_decap_8 FILLER_60_1267 ();
 sg13g2_decap_8 FILLER_60_1274 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_fill_2 FILLER_60_1288 ();
 sg13g2_fill_1 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_4 FILLER_60_1302 ();
 sg13g2_fill_1 FILLER_60_1306 ();
 sg13g2_fill_1 FILLER_60_1312 ();
 sg13g2_fill_1 FILLER_60_1319 ();
 sg13g2_fill_2 FILLER_60_1330 ();
 sg13g2_fill_1 FILLER_60_1332 ();
 sg13g2_fill_1 FILLER_60_1345 ();
 sg13g2_fill_1 FILLER_60_1351 ();
 sg13g2_fill_1 FILLER_60_1356 ();
 sg13g2_decap_4 FILLER_60_1362 ();
 sg13g2_fill_1 FILLER_60_1366 ();
 sg13g2_fill_1 FILLER_60_1371 ();
 sg13g2_fill_1 FILLER_60_1376 ();
 sg13g2_fill_1 FILLER_60_1382 ();
 sg13g2_fill_1 FILLER_60_1395 ();
 sg13g2_decap_4 FILLER_60_1405 ();
 sg13g2_fill_1 FILLER_60_1414 ();
 sg13g2_decap_4 FILLER_60_1420 ();
 sg13g2_fill_1 FILLER_60_1424 ();
 sg13g2_fill_1 FILLER_60_1433 ();
 sg13g2_fill_2 FILLER_60_1438 ();
 sg13g2_fill_1 FILLER_60_1450 ();
 sg13g2_fill_1 FILLER_60_1470 ();
 sg13g2_fill_2 FILLER_60_1476 ();
 sg13g2_fill_1 FILLER_60_1482 ();
 sg13g2_fill_1 FILLER_60_1513 ();
 sg13g2_fill_1 FILLER_60_1528 ();
 sg13g2_fill_2 FILLER_60_1537 ();
 sg13g2_fill_1 FILLER_60_1548 ();
 sg13g2_fill_1 FILLER_60_1554 ();
 sg13g2_fill_2 FILLER_60_1585 ();
 sg13g2_fill_2 FILLER_60_1591 ();
 sg13g2_fill_1 FILLER_60_1597 ();
 sg13g2_fill_1 FILLER_60_1624 ();
 sg13g2_fill_2 FILLER_60_1639 ();
 sg13g2_fill_1 FILLER_60_1641 ();
 sg13g2_fill_2 FILLER_60_1647 ();
 sg13g2_decap_4 FILLER_60_1653 ();
 sg13g2_fill_2 FILLER_60_1657 ();
 sg13g2_fill_1 FILLER_60_1670 ();
 sg13g2_decap_4 FILLER_60_1689 ();
 sg13g2_fill_1 FILLER_60_1693 ();
 sg13g2_fill_1 FILLER_60_1698 ();
 sg13g2_fill_1 FILLER_60_1703 ();
 sg13g2_decap_4 FILLER_60_1709 ();
 sg13g2_fill_1 FILLER_60_1713 ();
 sg13g2_fill_2 FILLER_60_1723 ();
 sg13g2_fill_1 FILLER_60_1725 ();
 sg13g2_decap_8 FILLER_60_1733 ();
 sg13g2_fill_2 FILLER_60_1758 ();
 sg13g2_fill_2 FILLER_60_1764 ();
 sg13g2_fill_2 FILLER_60_1771 ();
 sg13g2_decap_4 FILLER_60_1785 ();
 sg13g2_decap_8 FILLER_60_1803 ();
 sg13g2_decap_4 FILLER_60_1810 ();
 sg13g2_fill_2 FILLER_60_1814 ();
 sg13g2_decap_8 FILLER_60_1821 ();
 sg13g2_fill_2 FILLER_60_1828 ();
 sg13g2_fill_1 FILLER_60_1830 ();
 sg13g2_decap_4 FILLER_60_1836 ();
 sg13g2_fill_1 FILLER_60_1840 ();
 sg13g2_decap_8 FILLER_60_1845 ();
 sg13g2_decap_8 FILLER_60_1852 ();
 sg13g2_decap_8 FILLER_60_1859 ();
 sg13g2_decap_8 FILLER_60_1870 ();
 sg13g2_fill_2 FILLER_60_1891 ();
 sg13g2_fill_2 FILLER_60_1897 ();
 sg13g2_fill_2 FILLER_60_1909 ();
 sg13g2_fill_1 FILLER_60_1911 ();
 sg13g2_fill_1 FILLER_60_1925 ();
 sg13g2_decap_8 FILLER_60_1932 ();
 sg13g2_decap_8 FILLER_60_1939 ();
 sg13g2_decap_8 FILLER_60_1946 ();
 sg13g2_decap_8 FILLER_60_1953 ();
 sg13g2_decap_4 FILLER_60_1960 ();
 sg13g2_fill_2 FILLER_60_1964 ();
 sg13g2_decap_8 FILLER_60_1972 ();
 sg13g2_decap_8 FILLER_60_1979 ();
 sg13g2_decap_8 FILLER_60_1986 ();
 sg13g2_decap_8 FILLER_60_1993 ();
 sg13g2_decap_8 FILLER_60_2000 ();
 sg13g2_decap_4 FILLER_60_2007 ();
 sg13g2_fill_2 FILLER_60_2011 ();
 sg13g2_decap_8 FILLER_60_2017 ();
 sg13g2_decap_8 FILLER_60_2024 ();
 sg13g2_decap_8 FILLER_60_2031 ();
 sg13g2_decap_8 FILLER_60_2038 ();
 sg13g2_decap_8 FILLER_60_2045 ();
 sg13g2_decap_8 FILLER_60_2052 ();
 sg13g2_decap_8 FILLER_60_2059 ();
 sg13g2_decap_8 FILLER_60_2066 ();
 sg13g2_decap_8 FILLER_60_2073 ();
 sg13g2_decap_8 FILLER_60_2080 ();
 sg13g2_decap_4 FILLER_60_2087 ();
 sg13g2_fill_1 FILLER_60_2091 ();
 sg13g2_fill_2 FILLER_60_2144 ();
 sg13g2_fill_1 FILLER_60_2146 ();
 sg13g2_fill_2 FILLER_60_2158 ();
 sg13g2_fill_1 FILLER_60_2160 ();
 sg13g2_fill_2 FILLER_60_2196 ();
 sg13g2_fill_2 FILLER_60_2202 ();
 sg13g2_fill_1 FILLER_60_2241 ();
 sg13g2_fill_2 FILLER_60_2287 ();
 sg13g2_fill_1 FILLER_60_2289 ();
 sg13g2_fill_1 FILLER_60_2332 ();
 sg13g2_decap_4 FILLER_60_2415 ();
 sg13g2_fill_2 FILLER_60_2419 ();
 sg13g2_fill_2 FILLER_60_2455 ();
 sg13g2_decap_4 FILLER_60_2461 ();
 sg13g2_fill_1 FILLER_60_2465 ();
 sg13g2_fill_1 FILLER_60_2548 ();
 sg13g2_fill_1 FILLER_60_2565 ();
 sg13g2_fill_1 FILLER_60_2618 ();
 sg13g2_decap_8 FILLER_60_2645 ();
 sg13g2_decap_8 FILLER_60_2652 ();
 sg13g2_decap_8 FILLER_60_2659 ();
 sg13g2_decap_4 FILLER_60_2666 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_11 ();
 sg13g2_decap_8 FILLER_61_17 ();
 sg13g2_decap_8 FILLER_61_24 ();
 sg13g2_decap_8 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_38 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_120 ();
 sg13g2_fill_1 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_131 ();
 sg13g2_fill_1 FILLER_61_144 ();
 sg13g2_decap_8 FILLER_61_158 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_fill_1 FILLER_61_167 ();
 sg13g2_fill_2 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_decap_4 FILLER_61_234 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_fill_2 FILLER_61_249 ();
 sg13g2_fill_2 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_290 ();
 sg13g2_decap_8 FILLER_61_300 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_decap_4 FILLER_61_355 ();
 sg13g2_fill_2 FILLER_61_359 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_8 FILLER_61_405 ();
 sg13g2_fill_2 FILLER_61_412 ();
 sg13g2_fill_1 FILLER_61_414 ();
 sg13g2_fill_1 FILLER_61_435 ();
 sg13g2_fill_1 FILLER_61_469 ();
 sg13g2_fill_1 FILLER_61_474 ();
 sg13g2_fill_1 FILLER_61_480 ();
 sg13g2_fill_1 FILLER_61_487 ();
 sg13g2_fill_1 FILLER_61_493 ();
 sg13g2_fill_1 FILLER_61_508 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_fill_1 FILLER_61_526 ();
 sg13g2_fill_1 FILLER_61_532 ();
 sg13g2_fill_1 FILLER_61_545 ();
 sg13g2_decap_4 FILLER_61_572 ();
 sg13g2_fill_2 FILLER_61_592 ();
 sg13g2_fill_1 FILLER_61_594 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_610 ();
 sg13g2_decap_4 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_639 ();
 sg13g2_fill_2 FILLER_61_722 ();
 sg13g2_fill_1 FILLER_61_724 ();
 sg13g2_fill_1 FILLER_61_760 ();
 sg13g2_fill_2 FILLER_61_770 ();
 sg13g2_fill_2 FILLER_61_776 ();
 sg13g2_fill_2 FILLER_61_804 ();
 sg13g2_fill_2 FILLER_61_837 ();
 sg13g2_fill_1 FILLER_61_839 ();
 sg13g2_fill_2 FILLER_61_858 ();
 sg13g2_fill_1 FILLER_61_930 ();
 sg13g2_fill_1 FILLER_61_941 ();
 sg13g2_fill_1 FILLER_61_947 ();
 sg13g2_fill_1 FILLER_61_952 ();
 sg13g2_fill_1 FILLER_61_1001 ();
 sg13g2_fill_2 FILLER_61_1007 ();
 sg13g2_fill_1 FILLER_61_1009 ();
 sg13g2_decap_8 FILLER_61_1042 ();
 sg13g2_decap_8 FILLER_61_1049 ();
 sg13g2_decap_8 FILLER_61_1056 ();
 sg13g2_decap_8 FILLER_61_1063 ();
 sg13g2_decap_4 FILLER_61_1070 ();
 sg13g2_fill_2 FILLER_61_1074 ();
 sg13g2_fill_1 FILLER_61_1122 ();
 sg13g2_decap_8 FILLER_61_1130 ();
 sg13g2_fill_2 FILLER_61_1147 ();
 sg13g2_fill_1 FILLER_61_1149 ();
 sg13g2_fill_1 FILLER_61_1154 ();
 sg13g2_decap_8 FILLER_61_1159 ();
 sg13g2_decap_4 FILLER_61_1166 ();
 sg13g2_fill_1 FILLER_61_1170 ();
 sg13g2_decap_8 FILLER_61_1176 ();
 sg13g2_decap_8 FILLER_61_1209 ();
 sg13g2_decap_8 FILLER_61_1216 ();
 sg13g2_decap_8 FILLER_61_1223 ();
 sg13g2_fill_2 FILLER_61_1240 ();
 sg13g2_fill_1 FILLER_61_1242 ();
 sg13g2_decap_8 FILLER_61_1296 ();
 sg13g2_decap_8 FILLER_61_1303 ();
 sg13g2_fill_2 FILLER_61_1310 ();
 sg13g2_fill_1 FILLER_61_1317 ();
 sg13g2_decap_4 FILLER_61_1332 ();
 sg13g2_fill_2 FILLER_61_1336 ();
 sg13g2_decap_8 FILLER_61_1347 ();
 sg13g2_fill_1 FILLER_61_1354 ();
 sg13g2_fill_1 FILLER_61_1386 ();
 sg13g2_fill_1 FILLER_61_1390 ();
 sg13g2_fill_1 FILLER_61_1460 ();
 sg13g2_decap_4 FILLER_61_1470 ();
 sg13g2_fill_2 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1490 ();
 sg13g2_fill_1 FILLER_61_1502 ();
 sg13g2_decap_4 FILLER_61_1509 ();
 sg13g2_fill_1 FILLER_61_1540 ();
 sg13g2_decap_4 FILLER_61_1546 ();
 sg13g2_fill_1 FILLER_61_1550 ();
 sg13g2_fill_2 FILLER_61_1598 ();
 sg13g2_fill_1 FILLER_61_1600 ();
 sg13g2_decap_8 FILLER_61_1609 ();
 sg13g2_decap_8 FILLER_61_1616 ();
 sg13g2_decap_8 FILLER_61_1623 ();
 sg13g2_decap_8 FILLER_61_1635 ();
 sg13g2_decap_8 FILLER_61_1642 ();
 sg13g2_decap_8 FILLER_61_1649 ();
 sg13g2_decap_8 FILLER_61_1656 ();
 sg13g2_fill_1 FILLER_61_1663 ();
 sg13g2_fill_2 FILLER_61_1668 ();
 sg13g2_decap_8 FILLER_61_1674 ();
 sg13g2_fill_2 FILLER_61_1681 ();
 sg13g2_fill_1 FILLER_61_1683 ();
 sg13g2_fill_2 FILLER_61_1688 ();
 sg13g2_fill_1 FILLER_61_1698 ();
 sg13g2_decap_8 FILLER_61_1703 ();
 sg13g2_fill_1 FILLER_61_1710 ();
 sg13g2_decap_8 FILLER_61_1719 ();
 sg13g2_decap_8 FILLER_61_1726 ();
 sg13g2_decap_8 FILLER_61_1733 ();
 sg13g2_decap_8 FILLER_61_1740 ();
 sg13g2_decap_8 FILLER_61_1747 ();
 sg13g2_decap_8 FILLER_61_1754 ();
 sg13g2_decap_4 FILLER_61_1761 ();
 sg13g2_fill_1 FILLER_61_1765 ();
 sg13g2_decap_8 FILLER_61_1778 ();
 sg13g2_decap_8 FILLER_61_1785 ();
 sg13g2_decap_4 FILLER_61_1792 ();
 sg13g2_fill_1 FILLER_61_1796 ();
 sg13g2_decap_8 FILLER_61_1802 ();
 sg13g2_decap_8 FILLER_61_1809 ();
 sg13g2_decap_8 FILLER_61_1816 ();
 sg13g2_decap_8 FILLER_61_1823 ();
 sg13g2_decap_8 FILLER_61_1830 ();
 sg13g2_decap_8 FILLER_61_1837 ();
 sg13g2_decap_8 FILLER_61_1844 ();
 sg13g2_decap_8 FILLER_61_1851 ();
 sg13g2_decap_8 FILLER_61_1858 ();
 sg13g2_fill_1 FILLER_61_1865 ();
 sg13g2_decap_8 FILLER_61_1876 ();
 sg13g2_decap_8 FILLER_61_1883 ();
 sg13g2_fill_2 FILLER_61_1890 ();
 sg13g2_fill_1 FILLER_61_1892 ();
 sg13g2_decap_4 FILLER_61_1898 ();
 sg13g2_fill_1 FILLER_61_1902 ();
 sg13g2_decap_8 FILLER_61_1907 ();
 sg13g2_decap_8 FILLER_61_1914 ();
 sg13g2_decap_8 FILLER_61_1926 ();
 sg13g2_decap_8 FILLER_61_1933 ();
 sg13g2_decap_8 FILLER_61_1940 ();
 sg13g2_fill_2 FILLER_61_1947 ();
 sg13g2_fill_1 FILLER_61_1949 ();
 sg13g2_decap_8 FILLER_61_1956 ();
 sg13g2_decap_4 FILLER_61_1969 ();
 sg13g2_fill_1 FILLER_61_1973 ();
 sg13g2_decap_8 FILLER_61_1985 ();
 sg13g2_decap_4 FILLER_61_1997 ();
 sg13g2_fill_1 FILLER_61_2001 ();
 sg13g2_decap_8 FILLER_61_2006 ();
 sg13g2_fill_1 FILLER_61_2013 ();
 sg13g2_decap_8 FILLER_61_2037 ();
 sg13g2_decap_8 FILLER_61_2044 ();
 sg13g2_decap_8 FILLER_61_2051 ();
 sg13g2_decap_8 FILLER_61_2058 ();
 sg13g2_decap_8 FILLER_61_2065 ();
 sg13g2_decap_8 FILLER_61_2072 ();
 sg13g2_decap_8 FILLER_61_2079 ();
 sg13g2_fill_1 FILLER_61_2086 ();
 sg13g2_fill_2 FILLER_61_2191 ();
 sg13g2_fill_1 FILLER_61_2228 ();
 sg13g2_fill_1 FILLER_61_2239 ();
 sg13g2_fill_2 FILLER_61_2266 ();
 sg13g2_fill_1 FILLER_61_2279 ();
 sg13g2_fill_1 FILLER_61_2333 ();
 sg13g2_fill_2 FILLER_61_2373 ();
 sg13g2_fill_1 FILLER_61_2426 ();
 sg13g2_fill_1 FILLER_61_2437 ();
 sg13g2_fill_1 FILLER_61_2444 ();
 sg13g2_fill_2 FILLER_61_2451 ();
 sg13g2_fill_2 FILLER_61_2463 ();
 sg13g2_fill_1 FILLER_61_2465 ();
 sg13g2_decap_4 FILLER_61_2474 ();
 sg13g2_decap_8 FILLER_61_2492 ();
 sg13g2_decap_4 FILLER_61_2499 ();
 sg13g2_fill_1 FILLER_61_2503 ();
 sg13g2_fill_1 FILLER_61_2529 ();
 sg13g2_fill_2 FILLER_61_2551 ();
 sg13g2_fill_1 FILLER_61_2553 ();
 sg13g2_fill_2 FILLER_61_2557 ();
 sg13g2_fill_1 FILLER_61_2567 ();
 sg13g2_fill_1 FILLER_61_2578 ();
 sg13g2_decap_8 FILLER_61_2650 ();
 sg13g2_decap_8 FILLER_61_2657 ();
 sg13g2_decap_4 FILLER_61_2664 ();
 sg13g2_fill_2 FILLER_61_2668 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_94 ();
 sg13g2_decap_4 FILLER_62_101 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_151 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_decap_8 FILLER_62_207 ();
 sg13g2_decap_8 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_221 ();
 sg13g2_decap_8 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_decap_4 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_313 ();
 sg13g2_decap_4 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_decap_4 FILLER_62_327 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_decap_4 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_decap_4 FILLER_62_356 ();
 sg13g2_fill_1 FILLER_62_360 ();
 sg13g2_decap_4 FILLER_62_366 ();
 sg13g2_fill_2 FILLER_62_370 ();
 sg13g2_fill_2 FILLER_62_398 ();
 sg13g2_fill_2 FILLER_62_432 ();
 sg13g2_fill_2 FILLER_62_490 ();
 sg13g2_fill_1 FILLER_62_534 ();
 sg13g2_fill_1 FILLER_62_539 ();
 sg13g2_decap_4 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_585 ();
 sg13g2_decap_8 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_607 ();
 sg13g2_fill_1 FILLER_62_613 ();
 sg13g2_fill_1 FILLER_62_662 ();
 sg13g2_fill_2 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_699 ();
 sg13g2_decap_4 FILLER_62_739 ();
 sg13g2_fill_2 FILLER_62_760 ();
 sg13g2_fill_1 FILLER_62_762 ();
 sg13g2_fill_2 FILLER_62_768 ();
 sg13g2_fill_1 FILLER_62_770 ();
 sg13g2_fill_2 FILLER_62_776 ();
 sg13g2_fill_1 FILLER_62_778 ();
 sg13g2_fill_2 FILLER_62_784 ();
 sg13g2_fill_2 FILLER_62_831 ();
 sg13g2_fill_2 FILLER_62_839 ();
 sg13g2_decap_4 FILLER_62_874 ();
 sg13g2_decap_4 FILLER_62_882 ();
 sg13g2_fill_2 FILLER_62_886 ();
 sg13g2_fill_2 FILLER_62_893 ();
 sg13g2_fill_1 FILLER_62_895 ();
 sg13g2_fill_2 FILLER_62_927 ();
 sg13g2_fill_1 FILLER_62_953 ();
 sg13g2_fill_1 FILLER_62_1009 ();
 sg13g2_decap_8 FILLER_62_1018 ();
 sg13g2_decap_4 FILLER_62_1025 ();
 sg13g2_fill_2 FILLER_62_1029 ();
 sg13g2_decap_4 FILLER_62_1049 ();
 sg13g2_fill_2 FILLER_62_1053 ();
 sg13g2_decap_4 FILLER_62_1059 ();
 sg13g2_fill_1 FILLER_62_1063 ();
 sg13g2_decap_8 FILLER_62_1070 ();
 sg13g2_fill_1 FILLER_62_1077 ();
 sg13g2_decap_8 FILLER_62_1083 ();
 sg13g2_fill_2 FILLER_62_1090 ();
 sg13g2_fill_2 FILLER_62_1096 ();
 sg13g2_fill_1 FILLER_62_1132 ();
 sg13g2_decap_8 FILLER_62_1203 ();
 sg13g2_fill_2 FILLER_62_1210 ();
 sg13g2_fill_1 FILLER_62_1212 ();
 sg13g2_decap_4 FILLER_62_1295 ();
 sg13g2_fill_2 FILLER_62_1299 ();
 sg13g2_fill_2 FILLER_62_1340 ();
 sg13g2_decap_8 FILLER_62_1349 ();
 sg13g2_fill_2 FILLER_62_1356 ();
 sg13g2_fill_2 FILLER_62_1361 ();
 sg13g2_fill_1 FILLER_62_1363 ();
 sg13g2_fill_2 FILLER_62_1382 ();
 sg13g2_fill_1 FILLER_62_1398 ();
 sg13g2_fill_1 FILLER_62_1444 ();
 sg13g2_fill_1 FILLER_62_1454 ();
 sg13g2_fill_2 FILLER_62_1460 ();
 sg13g2_decap_8 FILLER_62_1478 ();
 sg13g2_decap_8 FILLER_62_1485 ();
 sg13g2_decap_8 FILLER_62_1492 ();
 sg13g2_fill_1 FILLER_62_1499 ();
 sg13g2_fill_1 FILLER_62_1566 ();
 sg13g2_fill_2 FILLER_62_1576 ();
 sg13g2_decap_4 FILLER_62_1591 ();
 sg13g2_fill_1 FILLER_62_1595 ();
 sg13g2_decap_8 FILLER_62_1612 ();
 sg13g2_decap_8 FILLER_62_1619 ();
 sg13g2_decap_8 FILLER_62_1626 ();
 sg13g2_decap_8 FILLER_62_1633 ();
 sg13g2_decap_8 FILLER_62_1640 ();
 sg13g2_decap_8 FILLER_62_1647 ();
 sg13g2_decap_8 FILLER_62_1654 ();
 sg13g2_decap_8 FILLER_62_1661 ();
 sg13g2_decap_8 FILLER_62_1668 ();
 sg13g2_decap_4 FILLER_62_1675 ();
 sg13g2_fill_2 FILLER_62_1679 ();
 sg13g2_decap_4 FILLER_62_1685 ();
 sg13g2_fill_2 FILLER_62_1689 ();
 sg13g2_decap_8 FILLER_62_1709 ();
 sg13g2_decap_8 FILLER_62_1716 ();
 sg13g2_decap_4 FILLER_62_1723 ();
 sg13g2_decap_8 FILLER_62_1732 ();
 sg13g2_decap_8 FILLER_62_1739 ();
 sg13g2_decap_8 FILLER_62_1746 ();
 sg13g2_decap_8 FILLER_62_1753 ();
 sg13g2_decap_8 FILLER_62_1760 ();
 sg13g2_decap_8 FILLER_62_1767 ();
 sg13g2_decap_8 FILLER_62_1778 ();
 sg13g2_decap_8 FILLER_62_1785 ();
 sg13g2_fill_2 FILLER_62_1792 ();
 sg13g2_decap_4 FILLER_62_1802 ();
 sg13g2_fill_2 FILLER_62_1806 ();
 sg13g2_decap_8 FILLER_62_1813 ();
 sg13g2_decap_8 FILLER_62_1820 ();
 sg13g2_decap_8 FILLER_62_1827 ();
 sg13g2_decap_8 FILLER_62_1834 ();
 sg13g2_decap_8 FILLER_62_1841 ();
 sg13g2_decap_8 FILLER_62_1848 ();
 sg13g2_decap_8 FILLER_62_1855 ();
 sg13g2_decap_8 FILLER_62_1862 ();
 sg13g2_fill_2 FILLER_62_1875 ();
 sg13g2_fill_1 FILLER_62_1877 ();
 sg13g2_decap_8 FILLER_62_1883 ();
 sg13g2_decap_8 FILLER_62_1890 ();
 sg13g2_fill_1 FILLER_62_1897 ();
 sg13g2_decap_8 FILLER_62_1910 ();
 sg13g2_decap_8 FILLER_62_1917 ();
 sg13g2_decap_8 FILLER_62_1924 ();
 sg13g2_decap_8 FILLER_62_1931 ();
 sg13g2_decap_4 FILLER_62_1938 ();
 sg13g2_fill_1 FILLER_62_1942 ();
 sg13g2_decap_8 FILLER_62_1948 ();
 sg13g2_decap_4 FILLER_62_1955 ();
 sg13g2_decap_8 FILLER_62_1968 ();
 sg13g2_decap_8 FILLER_62_1975 ();
 sg13g2_decap_8 FILLER_62_1982 ();
 sg13g2_decap_8 FILLER_62_1989 ();
 sg13g2_decap_8 FILLER_62_1996 ();
 sg13g2_decap_8 FILLER_62_2003 ();
 sg13g2_decap_8 FILLER_62_2010 ();
 sg13g2_fill_2 FILLER_62_2017 ();
 sg13g2_fill_1 FILLER_62_2019 ();
 sg13g2_fill_2 FILLER_62_2026 ();
 sg13g2_decap_8 FILLER_62_2036 ();
 sg13g2_decap_8 FILLER_62_2043 ();
 sg13g2_decap_8 FILLER_62_2050 ();
 sg13g2_decap_8 FILLER_62_2057 ();
 sg13g2_decap_8 FILLER_62_2064 ();
 sg13g2_decap_8 FILLER_62_2071 ();
 sg13g2_decap_8 FILLER_62_2078 ();
 sg13g2_decap_8 FILLER_62_2085 ();
 sg13g2_decap_8 FILLER_62_2096 ();
 sg13g2_fill_1 FILLER_62_2108 ();
 sg13g2_fill_2 FILLER_62_2113 ();
 sg13g2_decap_4 FILLER_62_2129 ();
 sg13g2_fill_1 FILLER_62_2157 ();
 sg13g2_fill_1 FILLER_62_2162 ();
 sg13g2_fill_2 FILLER_62_2192 ();
 sg13g2_fill_1 FILLER_62_2199 ();
 sg13g2_fill_1 FILLER_62_2238 ();
 sg13g2_fill_1 FILLER_62_2248 ();
 sg13g2_fill_1 FILLER_62_2259 ();
 sg13g2_fill_1 FILLER_62_2273 ();
 sg13g2_fill_2 FILLER_62_2284 ();
 sg13g2_fill_1 FILLER_62_2286 ();
 sg13g2_fill_1 FILLER_62_2291 ();
 sg13g2_fill_2 FILLER_62_2301 ();
 sg13g2_fill_1 FILLER_62_2376 ();
 sg13g2_fill_1 FILLER_62_2399 ();
 sg13g2_fill_1 FILLER_62_2550 ();
 sg13g2_fill_1 FILLER_62_2564 ();
 sg13g2_fill_2 FILLER_62_2575 ();
 sg13g2_fill_1 FILLER_62_2630 ();
 sg13g2_decap_8 FILLER_62_2659 ();
 sg13g2_decap_4 FILLER_62_2666 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_24 ();
 sg13g2_fill_1 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_103 ();
 sg13g2_fill_1 FILLER_63_138 ();
 sg13g2_fill_1 FILLER_63_144 ();
 sg13g2_decap_8 FILLER_63_193 ();
 sg13g2_decap_8 FILLER_63_200 ();
 sg13g2_decap_8 FILLER_63_207 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_226 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_fill_1 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_332 ();
 sg13g2_decap_8 FILLER_63_368 ();
 sg13g2_decap_4 FILLER_63_375 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_decap_4 FILLER_63_384 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_fill_2 FILLER_63_487 ();
 sg13g2_fill_1 FILLER_63_499 ();
 sg13g2_fill_2 FILLER_63_509 ();
 sg13g2_fill_1 FILLER_63_520 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_537 ();
 sg13g2_fill_1 FILLER_63_545 ();
 sg13g2_fill_2 FILLER_63_550 ();
 sg13g2_fill_1 FILLER_63_562 ();
 sg13g2_fill_2 FILLER_63_572 ();
 sg13g2_fill_2 FILLER_63_597 ();
 sg13g2_fill_1 FILLER_63_599 ();
 sg13g2_fill_2 FILLER_63_643 ();
 sg13g2_fill_1 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_720 ();
 sg13g2_fill_2 FILLER_63_732 ();
 sg13g2_fill_1 FILLER_63_734 ();
 sg13g2_decap_4 FILLER_63_761 ();
 sg13g2_decap_8 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_776 ();
 sg13g2_fill_2 FILLER_63_783 ();
 sg13g2_fill_1 FILLER_63_785 ();
 sg13g2_decap_4 FILLER_63_815 ();
 sg13g2_fill_2 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_decap_8 FILLER_63_837 ();
 sg13g2_fill_2 FILLER_63_844 ();
 sg13g2_fill_1 FILLER_63_846 ();
 sg13g2_fill_1 FILLER_63_856 ();
 sg13g2_fill_1 FILLER_63_893 ();
 sg13g2_decap_8 FILLER_63_898 ();
 sg13g2_fill_1 FILLER_63_905 ();
 sg13g2_fill_2 FILLER_63_912 ();
 sg13g2_fill_1 FILLER_63_914 ();
 sg13g2_fill_1 FILLER_63_924 ();
 sg13g2_fill_2 FILLER_63_930 ();
 sg13g2_fill_1 FILLER_63_947 ();
 sg13g2_fill_1 FILLER_63_977 ();
 sg13g2_fill_1 FILLER_63_1020 ();
 sg13g2_fill_1 FILLER_63_1035 ();
 sg13g2_fill_2 FILLER_63_1046 ();
 sg13g2_fill_1 FILLER_63_1074 ();
 sg13g2_fill_2 FILLER_63_1101 ();
 sg13g2_fill_2 FILLER_63_1107 ();
 sg13g2_decap_4 FILLER_63_1123 ();
 sg13g2_decap_8 FILLER_63_1134 ();
 sg13g2_decap_4 FILLER_63_1141 ();
 sg13g2_fill_1 FILLER_63_1187 ();
 sg13g2_fill_2 FILLER_63_1196 ();
 sg13g2_fill_1 FILLER_63_1198 ();
 sg13g2_fill_2 FILLER_63_1235 ();
 sg13g2_fill_1 FILLER_63_1237 ();
 sg13g2_decap_8 FILLER_63_1291 ();
 sg13g2_decap_8 FILLER_63_1298 ();
 sg13g2_fill_1 FILLER_63_1305 ();
 sg13g2_fill_1 FILLER_63_1324 ();
 sg13g2_decap_8 FILLER_63_1373 ();
 sg13g2_fill_1 FILLER_63_1380 ();
 sg13g2_fill_1 FILLER_63_1399 ();
 sg13g2_fill_1 FILLER_63_1414 ();
 sg13g2_fill_1 FILLER_63_1441 ();
 sg13g2_fill_1 FILLER_63_1447 ();
 sg13g2_decap_4 FILLER_63_1456 ();
 sg13g2_fill_2 FILLER_63_1460 ();
 sg13g2_decap_8 FILLER_63_1466 ();
 sg13g2_decap_8 FILLER_63_1473 ();
 sg13g2_decap_8 FILLER_63_1532 ();
 sg13g2_fill_1 FILLER_63_1539 ();
 sg13g2_decap_8 FILLER_63_1544 ();
 sg13g2_decap_4 FILLER_63_1561 ();
 sg13g2_fill_1 FILLER_63_1565 ();
 sg13g2_decap_8 FILLER_63_1581 ();
 sg13g2_decap_4 FILLER_63_1599 ();
 sg13g2_decap_8 FILLER_63_1607 ();
 sg13g2_decap_8 FILLER_63_1614 ();
 sg13g2_decap_8 FILLER_63_1621 ();
 sg13g2_decap_8 FILLER_63_1628 ();
 sg13g2_decap_8 FILLER_63_1635 ();
 sg13g2_decap_8 FILLER_63_1642 ();
 sg13g2_decap_8 FILLER_63_1649 ();
 sg13g2_decap_8 FILLER_63_1656 ();
 sg13g2_decap_8 FILLER_63_1663 ();
 sg13g2_decap_8 FILLER_63_1670 ();
 sg13g2_decap_8 FILLER_63_1677 ();
 sg13g2_fill_1 FILLER_63_1693 ();
 sg13g2_fill_1 FILLER_63_1699 ();
 sg13g2_fill_2 FILLER_63_1713 ();
 sg13g2_fill_2 FILLER_63_1727 ();
 sg13g2_fill_2 FILLER_63_1750 ();
 sg13g2_fill_1 FILLER_63_1752 ();
 sg13g2_decap_8 FILLER_63_1758 ();
 sg13g2_decap_8 FILLER_63_1765 ();
 sg13g2_decap_4 FILLER_63_1772 ();
 sg13g2_fill_1 FILLER_63_1776 ();
 sg13g2_fill_1 FILLER_63_1782 ();
 sg13g2_fill_2 FILLER_63_1790 ();
 sg13g2_fill_1 FILLER_63_1792 ();
 sg13g2_fill_2 FILLER_63_1805 ();
 sg13g2_decap_8 FILLER_63_1812 ();
 sg13g2_fill_1 FILLER_63_1819 ();
 sg13g2_decap_8 FILLER_63_1829 ();
 sg13g2_decap_8 FILLER_63_1836 ();
 sg13g2_decap_4 FILLER_63_1843 ();
 sg13g2_fill_2 FILLER_63_1847 ();
 sg13g2_decap_8 FILLER_63_1854 ();
 sg13g2_decap_8 FILLER_63_1861 ();
 sg13g2_decap_8 FILLER_63_1868 ();
 sg13g2_decap_8 FILLER_63_1875 ();
 sg13g2_decap_8 FILLER_63_1882 ();
 sg13g2_fill_1 FILLER_63_1889 ();
 sg13g2_fill_1 FILLER_63_1895 ();
 sg13g2_decap_4 FILLER_63_1900 ();
 sg13g2_decap_8 FILLER_63_1912 ();
 sg13g2_decap_4 FILLER_63_1919 ();
 sg13g2_fill_2 FILLER_63_1923 ();
 sg13g2_decap_8 FILLER_63_1931 ();
 sg13g2_decap_8 FILLER_63_1938 ();
 sg13g2_decap_8 FILLER_63_1945 ();
 sg13g2_decap_8 FILLER_63_1952 ();
 sg13g2_decap_8 FILLER_63_1959 ();
 sg13g2_decap_8 FILLER_63_1966 ();
 sg13g2_decap_8 FILLER_63_1973 ();
 sg13g2_decap_8 FILLER_63_1980 ();
 sg13g2_decap_8 FILLER_63_1991 ();
 sg13g2_decap_8 FILLER_63_1998 ();
 sg13g2_decap_4 FILLER_63_2005 ();
 sg13g2_fill_1 FILLER_63_2009 ();
 sg13g2_decap_8 FILLER_63_2018 ();
 sg13g2_decap_8 FILLER_63_2025 ();
 sg13g2_decap_8 FILLER_63_2032 ();
 sg13g2_decap_8 FILLER_63_2039 ();
 sg13g2_decap_8 FILLER_63_2046 ();
 sg13g2_decap_8 FILLER_63_2053 ();
 sg13g2_decap_8 FILLER_63_2060 ();
 sg13g2_decap_8 FILLER_63_2067 ();
 sg13g2_decap_8 FILLER_63_2074 ();
 sg13g2_decap_8 FILLER_63_2081 ();
 sg13g2_decap_4 FILLER_63_2088 ();
 sg13g2_fill_2 FILLER_63_2092 ();
 sg13g2_fill_1 FILLER_63_2138 ();
 sg13g2_fill_2 FILLER_63_2147 ();
 sg13g2_fill_1 FILLER_63_2149 ();
 sg13g2_fill_1 FILLER_63_2177 ();
 sg13g2_fill_2 FILLER_63_2200 ();
 sg13g2_decap_4 FILLER_63_2206 ();
 sg13g2_fill_2 FILLER_63_2210 ();
 sg13g2_decap_8 FILLER_63_2220 ();
 sg13g2_decap_8 FILLER_63_2227 ();
 sg13g2_decap_4 FILLER_63_2264 ();
 sg13g2_fill_2 FILLER_63_2268 ();
 sg13g2_decap_8 FILLER_63_2274 ();
 sg13g2_decap_4 FILLER_63_2281 ();
 sg13g2_fill_2 FILLER_63_2285 ();
 sg13g2_fill_1 FILLER_63_2292 ();
 sg13g2_fill_1 FILLER_63_2374 ();
 sg13g2_fill_1 FILLER_63_2417 ();
 sg13g2_fill_1 FILLER_63_2460 ();
 sg13g2_fill_1 FILLER_63_2467 ();
 sg13g2_decap_8 FILLER_63_2472 ();
 sg13g2_decap_8 FILLER_63_2479 ();
 sg13g2_decap_8 FILLER_63_2486 ();
 sg13g2_fill_2 FILLER_63_2493 ();
 sg13g2_fill_1 FILLER_63_2495 ();
 sg13g2_fill_2 FILLER_63_2511 ();
 sg13g2_decap_4 FILLER_63_2617 ();
 sg13g2_decap_8 FILLER_63_2647 ();
 sg13g2_decap_8 FILLER_63_2654 ();
 sg13g2_decap_8 FILLER_63_2661 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_64 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_decap_4 FILLER_64_180 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_fill_2 FILLER_64_225 ();
 sg13g2_fill_1 FILLER_64_227 ();
 sg13g2_fill_1 FILLER_64_262 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_270 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_286 ();
 sg13g2_fill_1 FILLER_64_291 ();
 sg13g2_fill_2 FILLER_64_300 ();
 sg13g2_decap_8 FILLER_64_310 ();
 sg13g2_fill_2 FILLER_64_341 ();
 sg13g2_fill_2 FILLER_64_356 ();
 sg13g2_fill_1 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_390 ();
 sg13g2_fill_1 FILLER_64_460 ();
 sg13g2_fill_1 FILLER_64_465 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_fill_1 FILLER_64_481 ();
 sg13g2_fill_1 FILLER_64_496 ();
 sg13g2_fill_1 FILLER_64_505 ();
 sg13g2_fill_2 FILLER_64_539 ();
 sg13g2_fill_1 FILLER_64_541 ();
 sg13g2_fill_1 FILLER_64_551 ();
 sg13g2_fill_2 FILLER_64_556 ();
 sg13g2_fill_1 FILLER_64_558 ();
 sg13g2_fill_2 FILLER_64_564 ();
 sg13g2_fill_1 FILLER_64_571 ();
 sg13g2_fill_1 FILLER_64_577 ();
 sg13g2_fill_2 FILLER_64_604 ();
 sg13g2_fill_1 FILLER_64_610 ();
 sg13g2_fill_1 FILLER_64_620 ();
 sg13g2_fill_1 FILLER_64_626 ();
 sg13g2_fill_2 FILLER_64_632 ();
 sg13g2_fill_1 FILLER_64_663 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_4 FILLER_64_689 ();
 sg13g2_fill_2 FILLER_64_693 ();
 sg13g2_fill_1 FILLER_64_699 ();
 sg13g2_fill_2 FILLER_64_711 ();
 sg13g2_fill_1 FILLER_64_713 ();
 sg13g2_decap_8 FILLER_64_762 ();
 sg13g2_decap_8 FILLER_64_769 ();
 sg13g2_decap_8 FILLER_64_776 ();
 sg13g2_decap_8 FILLER_64_783 ();
 sg13g2_decap_8 FILLER_64_835 ();
 sg13g2_decap_4 FILLER_64_842 ();
 sg13g2_fill_2 FILLER_64_846 ();
 sg13g2_fill_1 FILLER_64_851 ();
 sg13g2_fill_1 FILLER_64_858 ();
 sg13g2_fill_2 FILLER_64_868 ();
 sg13g2_fill_2 FILLER_64_880 ();
 sg13g2_fill_1 FILLER_64_882 ();
 sg13g2_decap_8 FILLER_64_893 ();
 sg13g2_fill_2 FILLER_64_905 ();
 sg13g2_fill_1 FILLER_64_907 ();
 sg13g2_fill_1 FILLER_64_925 ();
 sg13g2_fill_2 FILLER_64_949 ();
 sg13g2_fill_2 FILLER_64_956 ();
 sg13g2_fill_1 FILLER_64_970 ();
 sg13g2_fill_1 FILLER_64_1017 ();
 sg13g2_decap_4 FILLER_64_1049 ();
 sg13g2_fill_1 FILLER_64_1081 ();
 sg13g2_fill_2 FILLER_64_1108 ();
 sg13g2_fill_1 FILLER_64_1110 ();
 sg13g2_decap_8 FILLER_64_1145 ();
 sg13g2_decap_4 FILLER_64_1156 ();
 sg13g2_fill_1 FILLER_64_1160 ();
 sg13g2_decap_4 FILLER_64_1220 ();
 sg13g2_decap_8 FILLER_64_1281 ();
 sg13g2_decap_8 FILLER_64_1288 ();
 sg13g2_decap_8 FILLER_64_1295 ();
 sg13g2_decap_8 FILLER_64_1306 ();
 sg13g2_decap_4 FILLER_64_1313 ();
 sg13g2_fill_1 FILLER_64_1317 ();
 sg13g2_fill_1 FILLER_64_1323 ();
 sg13g2_fill_1 FILLER_64_1329 ();
 sg13g2_fill_2 FILLER_64_1338 ();
 sg13g2_fill_2 FILLER_64_1344 ();
 sg13g2_fill_2 FILLER_64_1350 ();
 sg13g2_fill_1 FILLER_64_1352 ();
 sg13g2_fill_1 FILLER_64_1371 ();
 sg13g2_fill_1 FILLER_64_1376 ();
 sg13g2_fill_1 FILLER_64_1383 ();
 sg13g2_decap_8 FILLER_64_1403 ();
 sg13g2_fill_1 FILLER_64_1410 ();
 sg13g2_decap_8 FILLER_64_1453 ();
 sg13g2_decap_4 FILLER_64_1460 ();
 sg13g2_fill_2 FILLER_64_1464 ();
 sg13g2_fill_2 FILLER_64_1479 ();
 sg13g2_decap_4 FILLER_64_1517 ();
 sg13g2_fill_1 FILLER_64_1521 ();
 sg13g2_fill_2 FILLER_64_1533 ();
 sg13g2_fill_1 FILLER_64_1535 ();
 sg13g2_fill_2 FILLER_64_1546 ();
 sg13g2_fill_2 FILLER_64_1553 ();
 sg13g2_fill_1 FILLER_64_1555 ();
 sg13g2_decap_4 FILLER_64_1561 ();
 sg13g2_fill_1 FILLER_64_1565 ();
 sg13g2_fill_1 FILLER_64_1574 ();
 sg13g2_fill_2 FILLER_64_1603 ();
 sg13g2_fill_1 FILLER_64_1605 ();
 sg13g2_decap_8 FILLER_64_1610 ();
 sg13g2_fill_2 FILLER_64_1617 ();
 sg13g2_fill_1 FILLER_64_1619 ();
 sg13g2_decap_8 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1633 ();
 sg13g2_decap_8 FILLER_64_1640 ();
 sg13g2_decap_4 FILLER_64_1647 ();
 sg13g2_fill_2 FILLER_64_1651 ();
 sg13g2_decap_4 FILLER_64_1681 ();
 sg13g2_fill_1 FILLER_64_1685 ();
 sg13g2_decap_8 FILLER_64_1690 ();
 sg13g2_decap_8 FILLER_64_1697 ();
 sg13g2_fill_1 FILLER_64_1712 ();
 sg13g2_fill_2 FILLER_64_1749 ();
 sg13g2_fill_1 FILLER_64_1751 ();
 sg13g2_decap_8 FILLER_64_1757 ();
 sg13g2_decap_8 FILLER_64_1764 ();
 sg13g2_decap_4 FILLER_64_1771 ();
 sg13g2_fill_1 FILLER_64_1775 ();
 sg13g2_decap_8 FILLER_64_1784 ();
 sg13g2_decap_8 FILLER_64_1791 ();
 sg13g2_decap_8 FILLER_64_1798 ();
 sg13g2_decap_4 FILLER_64_1805 ();
 sg13g2_fill_1 FILLER_64_1809 ();
 sg13g2_decap_4 FILLER_64_1815 ();
 sg13g2_fill_2 FILLER_64_1819 ();
 sg13g2_decap_8 FILLER_64_1834 ();
 sg13g2_decap_4 FILLER_64_1841 ();
 sg13g2_decap_8 FILLER_64_1853 ();
 sg13g2_decap_8 FILLER_64_1860 ();
 sg13g2_decap_8 FILLER_64_1867 ();
 sg13g2_decap_8 FILLER_64_1874 ();
 sg13g2_decap_4 FILLER_64_1881 ();
 sg13g2_decap_8 FILLER_64_1891 ();
 sg13g2_decap_8 FILLER_64_1898 ();
 sg13g2_decap_8 FILLER_64_1905 ();
 sg13g2_decap_8 FILLER_64_1912 ();
 sg13g2_decap_8 FILLER_64_1919 ();
 sg13g2_decap_8 FILLER_64_1926 ();
 sg13g2_decap_8 FILLER_64_1933 ();
 sg13g2_decap_8 FILLER_64_1940 ();
 sg13g2_decap_8 FILLER_64_1947 ();
 sg13g2_decap_8 FILLER_64_1954 ();
 sg13g2_decap_8 FILLER_64_1961 ();
 sg13g2_decap_8 FILLER_64_1968 ();
 sg13g2_decap_8 FILLER_64_1975 ();
 sg13g2_decap_8 FILLER_64_1982 ();
 sg13g2_decap_8 FILLER_64_1995 ();
 sg13g2_decap_8 FILLER_64_2002 ();
 sg13g2_decap_8 FILLER_64_2009 ();
 sg13g2_decap_8 FILLER_64_2016 ();
 sg13g2_decap_4 FILLER_64_2023 ();
 sg13g2_fill_2 FILLER_64_2027 ();
 sg13g2_decap_8 FILLER_64_2035 ();
 sg13g2_decap_8 FILLER_64_2042 ();
 sg13g2_decap_8 FILLER_64_2049 ();
 sg13g2_decap_8 FILLER_64_2056 ();
 sg13g2_decap_8 FILLER_64_2063 ();
 sg13g2_decap_8 FILLER_64_2070 ();
 sg13g2_decap_8 FILLER_64_2077 ();
 sg13g2_fill_2 FILLER_64_2084 ();
 sg13g2_fill_1 FILLER_64_2086 ();
 sg13g2_fill_1 FILLER_64_2118 ();
 sg13g2_fill_1 FILLER_64_2139 ();
 sg13g2_fill_1 FILLER_64_2224 ();
 sg13g2_fill_1 FILLER_64_2238 ();
 sg13g2_fill_1 FILLER_64_2270 ();
 sg13g2_fill_2 FILLER_64_2320 ();
 sg13g2_fill_2 FILLER_64_2334 ();
 sg13g2_fill_1 FILLER_64_2379 ();
 sg13g2_fill_2 FILLER_64_2410 ();
 sg13g2_fill_1 FILLER_64_2418 ();
 sg13g2_decap_8 FILLER_64_2424 ();
 sg13g2_fill_1 FILLER_64_2457 ();
 sg13g2_fill_1 FILLER_64_2470 ();
 sg13g2_fill_1 FILLER_64_2481 ();
 sg13g2_fill_1 FILLER_64_2508 ();
 sg13g2_fill_2 FILLER_64_2561 ();
 sg13g2_decap_4 FILLER_64_2610 ();
 sg13g2_decap_4 FILLER_64_2624 ();
 sg13g2_decap_8 FILLER_64_2632 ();
 sg13g2_decap_8 FILLER_64_2639 ();
 sg13g2_decap_8 FILLER_64_2646 ();
 sg13g2_decap_8 FILLER_64_2653 ();
 sg13g2_decap_8 FILLER_64_2660 ();
 sg13g2_fill_2 FILLER_64_2667 ();
 sg13g2_fill_1 FILLER_64_2669 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_38 ();
 sg13g2_fill_1 FILLER_65_45 ();
 sg13g2_fill_2 FILLER_65_82 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_fill_1 FILLER_65_124 ();
 sg13g2_fill_1 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_182 ();
 sg13g2_fill_2 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_215 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_291 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_decap_4 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_314 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_2 FILLER_65_374 ();
 sg13g2_decap_8 FILLER_65_380 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_decap_4 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_424 ();
 sg13g2_fill_2 FILLER_65_463 ();
 sg13g2_fill_1 FILLER_65_469 ();
 sg13g2_decap_4 FILLER_65_474 ();
 sg13g2_fill_2 FILLER_65_478 ();
 sg13g2_fill_1 FILLER_65_484 ();
 sg13g2_fill_2 FILLER_65_539 ();
 sg13g2_fill_1 FILLER_65_541 ();
 sg13g2_fill_2 FILLER_65_591 ();
 sg13g2_fill_1 FILLER_65_607 ();
 sg13g2_fill_2 FILLER_65_613 ();
 sg13g2_fill_2 FILLER_65_665 ();
 sg13g2_fill_1 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_fill_2 FILLER_65_718 ();
 sg13g2_fill_1 FILLER_65_720 ();
 sg13g2_fill_2 FILLER_65_733 ();
 sg13g2_fill_1 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_773 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_4 FILLER_65_791 ();
 sg13g2_fill_1 FILLER_65_820 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_4 FILLER_65_885 ();
 sg13g2_fill_1 FILLER_65_920 ();
 sg13g2_fill_2 FILLER_65_942 ();
 sg13g2_fill_2 FILLER_65_1010 ();
 sg13g2_decap_8 FILLER_65_1041 ();
 sg13g2_decap_4 FILLER_65_1068 ();
 sg13g2_decap_4 FILLER_65_1076 ();
 sg13g2_fill_1 FILLER_65_1089 ();
 sg13g2_fill_2 FILLER_65_1114 ();
 sg13g2_decap_8 FILLER_65_1152 ();
 sg13g2_decap_4 FILLER_65_1159 ();
 sg13g2_fill_1 FILLER_65_1163 ();
 sg13g2_decap_4 FILLER_65_1169 ();
 sg13g2_fill_1 FILLER_65_1173 ();
 sg13g2_fill_1 FILLER_65_1184 ();
 sg13g2_fill_2 FILLER_65_1219 ();
 sg13g2_fill_1 FILLER_65_1221 ();
 sg13g2_fill_2 FILLER_65_1232 ();
 sg13g2_fill_1 FILLER_65_1234 ();
 sg13g2_fill_2 FILLER_65_1247 ();
 sg13g2_decap_8 FILLER_65_1259 ();
 sg13g2_decap_8 FILLER_65_1270 ();
 sg13g2_decap_8 FILLER_65_1277 ();
 sg13g2_decap_8 FILLER_65_1284 ();
 sg13g2_decap_4 FILLER_65_1291 ();
 sg13g2_decap_8 FILLER_65_1329 ();
 sg13g2_decap_8 FILLER_65_1340 ();
 sg13g2_fill_1 FILLER_65_1347 ();
 sg13g2_decap_4 FILLER_65_1353 ();
 sg13g2_fill_1 FILLER_65_1357 ();
 sg13g2_fill_2 FILLER_65_1364 ();
 sg13g2_fill_2 FILLER_65_1372 ();
 sg13g2_fill_1 FILLER_65_1382 ();
 sg13g2_fill_1 FILLER_65_1406 ();
 sg13g2_decap_8 FILLER_65_1412 ();
 sg13g2_fill_1 FILLER_65_1429 ();
 sg13g2_fill_1 FILLER_65_1435 ();
 sg13g2_fill_1 FILLER_65_1442 ();
 sg13g2_fill_2 FILLER_65_1448 ();
 sg13g2_fill_1 FILLER_65_1454 ();
 sg13g2_fill_2 FILLER_65_1462 ();
 sg13g2_fill_1 FILLER_65_1473 ();
 sg13g2_fill_2 FILLER_65_1487 ();
 sg13g2_decap_4 FILLER_65_1493 ();
 sg13g2_fill_2 FILLER_65_1502 ();
 sg13g2_fill_2 FILLER_65_1508 ();
 sg13g2_fill_1 FILLER_65_1510 ();
 sg13g2_fill_1 FILLER_65_1515 ();
 sg13g2_fill_2 FILLER_65_1546 ();
 sg13g2_fill_1 FILLER_65_1548 ();
 sg13g2_decap_8 FILLER_65_1553 ();
 sg13g2_fill_2 FILLER_65_1560 ();
 sg13g2_decap_8 FILLER_65_1566 ();
 sg13g2_decap_4 FILLER_65_1573 ();
 sg13g2_fill_2 FILLER_65_1577 ();
 sg13g2_fill_1 FILLER_65_1598 ();
 sg13g2_decap_8 FILLER_65_1629 ();
 sg13g2_decap_8 FILLER_65_1636 ();
 sg13g2_decap_8 FILLER_65_1643 ();
 sg13g2_decap_8 FILLER_65_1650 ();
 sg13g2_fill_2 FILLER_65_1657 ();
 sg13g2_fill_1 FILLER_65_1673 ();
 sg13g2_decap_4 FILLER_65_1683 ();
 sg13g2_fill_1 FILLER_65_1691 ();
 sg13g2_decap_8 FILLER_65_1701 ();
 sg13g2_decap_8 FILLER_65_1708 ();
 sg13g2_decap_4 FILLER_65_1715 ();
 sg13g2_fill_1 FILLER_65_1719 ();
 sg13g2_decap_4 FILLER_65_1729 ();
 sg13g2_fill_1 FILLER_65_1756 ();
 sg13g2_fill_2 FILLER_65_1767 ();
 sg13g2_fill_1 FILLER_65_1773 ();
 sg13g2_decap_8 FILLER_65_1784 ();
 sg13g2_decap_8 FILLER_65_1791 ();
 sg13g2_decap_8 FILLER_65_1798 ();
 sg13g2_decap_4 FILLER_65_1805 ();
 sg13g2_fill_1 FILLER_65_1809 ();
 sg13g2_decap_8 FILLER_65_1815 ();
 sg13g2_decap_8 FILLER_65_1822 ();
 sg13g2_decap_8 FILLER_65_1829 ();
 sg13g2_decap_8 FILLER_65_1836 ();
 sg13g2_decap_8 FILLER_65_1843 ();
 sg13g2_decap_8 FILLER_65_1850 ();
 sg13g2_decap_8 FILLER_65_1857 ();
 sg13g2_decap_8 FILLER_65_1864 ();
 sg13g2_decap_8 FILLER_65_1871 ();
 sg13g2_decap_8 FILLER_65_1878 ();
 sg13g2_fill_1 FILLER_65_1885 ();
 sg13g2_decap_8 FILLER_65_1890 ();
 sg13g2_decap_8 FILLER_65_1897 ();
 sg13g2_decap_8 FILLER_65_1904 ();
 sg13g2_decap_8 FILLER_65_1911 ();
 sg13g2_decap_8 FILLER_65_1918 ();
 sg13g2_fill_1 FILLER_65_1925 ();
 sg13g2_decap_8 FILLER_65_1931 ();
 sg13g2_decap_8 FILLER_65_1938 ();
 sg13g2_decap_8 FILLER_65_1945 ();
 sg13g2_decap_4 FILLER_65_1952 ();
 sg13g2_decap_8 FILLER_65_1962 ();
 sg13g2_decap_8 FILLER_65_1969 ();
 sg13g2_decap_8 FILLER_65_1976 ();
 sg13g2_decap_8 FILLER_65_1983 ();
 sg13g2_decap_4 FILLER_65_1990 ();
 sg13g2_fill_2 FILLER_65_1994 ();
 sg13g2_decap_8 FILLER_65_2002 ();
 sg13g2_decap_8 FILLER_65_2009 ();
 sg13g2_decap_8 FILLER_65_2016 ();
 sg13g2_fill_2 FILLER_65_2023 ();
 sg13g2_decap_8 FILLER_65_2039 ();
 sg13g2_decap_8 FILLER_65_2046 ();
 sg13g2_decap_8 FILLER_65_2053 ();
 sg13g2_decap_8 FILLER_65_2060 ();
 sg13g2_decap_8 FILLER_65_2067 ();
 sg13g2_decap_8 FILLER_65_2074 ();
 sg13g2_decap_8 FILLER_65_2081 ();
 sg13g2_fill_1 FILLER_65_2088 ();
 sg13g2_decap_8 FILLER_65_2094 ();
 sg13g2_fill_1 FILLER_65_2101 ();
 sg13g2_decap_8 FILLER_65_2106 ();
 sg13g2_decap_8 FILLER_65_2113 ();
 sg13g2_fill_2 FILLER_65_2130 ();
 sg13g2_fill_1 FILLER_65_2132 ();
 sg13g2_fill_2 FILLER_65_2206 ();
 sg13g2_fill_1 FILLER_65_2222 ();
 sg13g2_fill_2 FILLER_65_2257 ();
 sg13g2_fill_1 FILLER_65_2332 ();
 sg13g2_fill_2 FILLER_65_2341 ();
 sg13g2_fill_1 FILLER_65_2379 ();
 sg13g2_fill_1 FILLER_65_2390 ();
 sg13g2_decap_4 FILLER_65_2460 ();
 sg13g2_fill_2 FILLER_65_2523 ();
 sg13g2_fill_1 FILLER_65_2562 ();
 sg13g2_fill_1 FILLER_65_2569 ();
 sg13g2_fill_1 FILLER_65_2580 ();
 sg13g2_fill_1 FILLER_65_2607 ();
 sg13g2_decap_8 FILLER_65_2644 ();
 sg13g2_decap_8 FILLER_65_2651 ();
 sg13g2_decap_8 FILLER_65_2658 ();
 sg13g2_decap_4 FILLER_65_2665 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_17 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_fill_2 FILLER_66_63 ();
 sg13g2_fill_1 FILLER_66_95 ();
 sg13g2_fill_1 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_148 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_fill_2 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_183 ();
 sg13g2_fill_1 FILLER_66_185 ();
 sg13g2_fill_2 FILLER_66_190 ();
 sg13g2_fill_1 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_283 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_decap_4 FILLER_66_302 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_348 ();
 sg13g2_fill_2 FILLER_66_363 ();
 sg13g2_decap_8 FILLER_66_391 ();
 sg13g2_fill_1 FILLER_66_496 ();
 sg13g2_fill_2 FILLER_66_519 ();
 sg13g2_fill_2 FILLER_66_526 ();
 sg13g2_decap_8 FILLER_66_542 ();
 sg13g2_decap_4 FILLER_66_549 ();
 sg13g2_fill_2 FILLER_66_553 ();
 sg13g2_decap_4 FILLER_66_559 ();
 sg13g2_fill_1 FILLER_66_563 ();
 sg13g2_fill_2 FILLER_66_568 ();
 sg13g2_fill_1 FILLER_66_570 ();
 sg13g2_fill_2 FILLER_66_575 ();
 sg13g2_fill_1 FILLER_66_577 ();
 sg13g2_fill_2 FILLER_66_584 ();
 sg13g2_fill_2 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_619 ();
 sg13g2_fill_1 FILLER_66_630 ();
 sg13g2_fill_1 FILLER_66_715 ();
 sg13g2_fill_1 FILLER_66_747 ();
 sg13g2_fill_2 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_890 ();
 sg13g2_fill_2 FILLER_66_999 ();
 sg13g2_fill_1 FILLER_66_1060 ();
 sg13g2_decap_4 FILLER_66_1071 ();
 sg13g2_fill_2 FILLER_66_1075 ();
 sg13g2_fill_2 FILLER_66_1088 ();
 sg13g2_fill_1 FILLER_66_1103 ();
 sg13g2_fill_2 FILLER_66_1145 ();
 sg13g2_fill_1 FILLER_66_1193 ();
 sg13g2_fill_1 FILLER_66_1204 ();
 sg13g2_decap_8 FILLER_66_1209 ();
 sg13g2_decap_8 FILLER_66_1216 ();
 sg13g2_decap_8 FILLER_66_1223 ();
 sg13g2_decap_8 FILLER_66_1242 ();
 sg13g2_fill_2 FILLER_66_1285 ();
 sg13g2_fill_2 FILLER_66_1328 ();
 sg13g2_fill_1 FILLER_66_1338 ();
 sg13g2_fill_1 FILLER_66_1364 ();
 sg13g2_fill_1 FILLER_66_1375 ();
 sg13g2_decap_4 FILLER_66_1419 ();
 sg13g2_fill_1 FILLER_66_1423 ();
 sg13g2_fill_1 FILLER_66_1429 ();
 sg13g2_fill_2 FILLER_66_1446 ();
 sg13g2_fill_1 FILLER_66_1448 ();
 sg13g2_decap_4 FILLER_66_1453 ();
 sg13g2_fill_2 FILLER_66_1482 ();
 sg13g2_decap_4 FILLER_66_1495 ();
 sg13g2_fill_1 FILLER_66_1499 ();
 sg13g2_decap_8 FILLER_66_1504 ();
 sg13g2_fill_1 FILLER_66_1515 ();
 sg13g2_fill_2 FILLER_66_1526 ();
 sg13g2_decap_4 FILLER_66_1533 ();
 sg13g2_fill_1 FILLER_66_1537 ();
 sg13g2_decap_8 FILLER_66_1543 ();
 sg13g2_decap_4 FILLER_66_1550 ();
 sg13g2_decap_8 FILLER_66_1559 ();
 sg13g2_fill_1 FILLER_66_1566 ();
 sg13g2_decap_8 FILLER_66_1577 ();
 sg13g2_fill_1 FILLER_66_1589 ();
 sg13g2_decap_8 FILLER_66_1620 ();
 sg13g2_decap_8 FILLER_66_1627 ();
 sg13g2_decap_8 FILLER_66_1634 ();
 sg13g2_decap_8 FILLER_66_1641 ();
 sg13g2_fill_2 FILLER_66_1653 ();
 sg13g2_fill_1 FILLER_66_1664 ();
 sg13g2_fill_2 FILLER_66_1687 ();
 sg13g2_decap_8 FILLER_66_1693 ();
 sg13g2_decap_8 FILLER_66_1700 ();
 sg13g2_decap_8 FILLER_66_1707 ();
 sg13g2_decap_8 FILLER_66_1714 ();
 sg13g2_decap_4 FILLER_66_1721 ();
 sg13g2_fill_2 FILLER_66_1725 ();
 sg13g2_decap_4 FILLER_66_1758 ();
 sg13g2_fill_2 FILLER_66_1762 ();
 sg13g2_fill_2 FILLER_66_1774 ();
 sg13g2_fill_1 FILLER_66_1781 ();
 sg13g2_decap_8 FILLER_66_1792 ();
 sg13g2_decap_8 FILLER_66_1799 ();
 sg13g2_decap_8 FILLER_66_1806 ();
 sg13g2_decap_8 FILLER_66_1813 ();
 sg13g2_decap_8 FILLER_66_1820 ();
 sg13g2_decap_8 FILLER_66_1827 ();
 sg13g2_decap_4 FILLER_66_1834 ();
 sg13g2_fill_2 FILLER_66_1838 ();
 sg13g2_decap_8 FILLER_66_1843 ();
 sg13g2_fill_2 FILLER_66_1850 ();
 sg13g2_decap_8 FILLER_66_1857 ();
 sg13g2_fill_2 FILLER_66_1864 ();
 sg13g2_fill_1 FILLER_66_1866 ();
 sg13g2_decap_8 FILLER_66_1872 ();
 sg13g2_fill_1 FILLER_66_1879 ();
 sg13g2_decap_8 FILLER_66_1892 ();
 sg13g2_decap_8 FILLER_66_1899 ();
 sg13g2_fill_1 FILLER_66_1906 ();
 sg13g2_decap_8 FILLER_66_1911 ();
 sg13g2_decap_8 FILLER_66_1918 ();
 sg13g2_decap_8 FILLER_66_1925 ();
 sg13g2_decap_8 FILLER_66_1932 ();
 sg13g2_decap_8 FILLER_66_1939 ();
 sg13g2_decap_4 FILLER_66_1946 ();
 sg13g2_fill_2 FILLER_66_1950 ();
 sg13g2_decap_8 FILLER_66_1958 ();
 sg13g2_decap_8 FILLER_66_1965 ();
 sg13g2_decap_8 FILLER_66_1972 ();
 sg13g2_decap_8 FILLER_66_1979 ();
 sg13g2_fill_2 FILLER_66_1986 ();
 sg13g2_fill_1 FILLER_66_1988 ();
 sg13g2_decap_8 FILLER_66_2001 ();
 sg13g2_decap_8 FILLER_66_2008 ();
 sg13g2_decap_4 FILLER_66_2015 ();
 sg13g2_fill_2 FILLER_66_2019 ();
 sg13g2_decap_8 FILLER_66_2027 ();
 sg13g2_decap_8 FILLER_66_2034 ();
 sg13g2_decap_8 FILLER_66_2041 ();
 sg13g2_decap_8 FILLER_66_2048 ();
 sg13g2_decap_8 FILLER_66_2055 ();
 sg13g2_decap_8 FILLER_66_2062 ();
 sg13g2_decap_8 FILLER_66_2069 ();
 sg13g2_decap_8 FILLER_66_2076 ();
 sg13g2_decap_8 FILLER_66_2083 ();
 sg13g2_decap_4 FILLER_66_2090 ();
 sg13g2_fill_1 FILLER_66_2094 ();
 sg13g2_decap_4 FILLER_66_2103 ();
 sg13g2_fill_2 FILLER_66_2107 ();
 sg13g2_fill_1 FILLER_66_2149 ();
 sg13g2_decap_8 FILLER_66_2164 ();
 sg13g2_fill_1 FILLER_66_2171 ();
 sg13g2_fill_1 FILLER_66_2177 ();
 sg13g2_fill_2 FILLER_66_2182 ();
 sg13g2_fill_1 FILLER_66_2184 ();
 sg13g2_fill_2 FILLER_66_2194 ();
 sg13g2_fill_2 FILLER_66_2248 ();
 sg13g2_fill_2 FILLER_66_2284 ();
 sg13g2_fill_2 FILLER_66_2328 ();
 sg13g2_fill_1 FILLER_66_2362 ();
 sg13g2_fill_2 FILLER_66_2374 ();
 sg13g2_fill_1 FILLER_66_2380 ();
 sg13g2_fill_1 FILLER_66_2407 ();
 sg13g2_fill_1 FILLER_66_2413 ();
 sg13g2_fill_1 FILLER_66_2418 ();
 sg13g2_fill_1 FILLER_66_2439 ();
 sg13g2_fill_2 FILLER_66_2482 ();
 sg13g2_decap_8 FILLER_66_2544 ();
 sg13g2_decap_8 FILLER_66_2551 ();
 sg13g2_fill_1 FILLER_66_2565 ();
 sg13g2_fill_1 FILLER_66_2586 ();
 sg13g2_decap_8 FILLER_66_2617 ();
 sg13g2_fill_1 FILLER_66_2624 ();
 sg13g2_decap_8 FILLER_66_2629 ();
 sg13g2_decap_8 FILLER_66_2636 ();
 sg13g2_decap_8 FILLER_66_2643 ();
 sg13g2_decap_8 FILLER_66_2650 ();
 sg13g2_decap_8 FILLER_66_2657 ();
 sg13g2_decap_4 FILLER_66_2664 ();
 sg13g2_fill_2 FILLER_66_2668 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_12 ();
 sg13g2_fill_1 FILLER_67_39 ();
 sg13g2_fill_1 FILLER_67_54 ();
 sg13g2_fill_1 FILLER_67_117 ();
 sg13g2_fill_1 FILLER_67_122 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_2 FILLER_67_216 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_decap_4 FILLER_67_231 ();
 sg13g2_fill_2 FILLER_67_253 ();
 sg13g2_fill_1 FILLER_67_296 ();
 sg13g2_fill_1 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_decap_8 FILLER_67_317 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_fill_2 FILLER_67_336 ();
 sg13g2_fill_1 FILLER_67_338 ();
 sg13g2_fill_2 FILLER_67_348 ();
 sg13g2_fill_1 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_384 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_409 ();
 sg13g2_fill_2 FILLER_67_415 ();
 sg13g2_decap_4 FILLER_67_445 ();
 sg13g2_fill_1 FILLER_67_449 ();
 sg13g2_decap_4 FILLER_67_490 ();
 sg13g2_fill_1 FILLER_67_499 ();
 sg13g2_decap_8 FILLER_67_510 ();
 sg13g2_fill_2 FILLER_67_522 ();
 sg13g2_fill_2 FILLER_67_550 ();
 sg13g2_fill_1 FILLER_67_557 ();
 sg13g2_fill_2 FILLER_67_563 ();
 sg13g2_fill_2 FILLER_67_570 ();
 sg13g2_fill_1 FILLER_67_598 ();
 sg13g2_fill_2 FILLER_67_604 ();
 sg13g2_fill_1 FILLER_67_615 ();
 sg13g2_fill_1 FILLER_67_700 ();
 sg13g2_fill_2 FILLER_67_711 ();
 sg13g2_fill_2 FILLER_67_739 ();
 sg13g2_fill_1 FILLER_67_741 ();
 sg13g2_fill_1 FILLER_67_747 ();
 sg13g2_fill_1 FILLER_67_759 ();
 sg13g2_fill_2 FILLER_67_771 ();
 sg13g2_fill_2 FILLER_67_777 ();
 sg13g2_fill_1 FILLER_67_779 ();
 sg13g2_fill_1 FILLER_67_816 ();
 sg13g2_fill_1 FILLER_67_821 ();
 sg13g2_fill_1 FILLER_67_865 ();
 sg13g2_fill_2 FILLER_67_885 ();
 sg13g2_fill_2 FILLER_67_937 ();
 sg13g2_fill_2 FILLER_67_973 ();
 sg13g2_fill_2 FILLER_67_998 ();
 sg13g2_fill_1 FILLER_67_1021 ();
 sg13g2_fill_1 FILLER_67_1034 ();
 sg13g2_fill_2 FILLER_67_1091 ();
 sg13g2_fill_1 FILLER_67_1093 ();
 sg13g2_fill_2 FILLER_67_1120 ();
 sg13g2_decap_4 FILLER_67_1173 ();
 sg13g2_fill_1 FILLER_67_1177 ();
 sg13g2_fill_2 FILLER_67_1191 ();
 sg13g2_fill_1 FILLER_67_1193 ();
 sg13g2_fill_1 FILLER_67_1220 ();
 sg13g2_decap_4 FILLER_67_1231 ();
 sg13g2_fill_1 FILLER_67_1235 ();
 sg13g2_fill_2 FILLER_67_1248 ();
 sg13g2_decap_8 FILLER_67_1286 ();
 sg13g2_fill_2 FILLER_67_1293 ();
 sg13g2_fill_1 FILLER_67_1295 ();
 sg13g2_fill_1 FILLER_67_1333 ();
 sg13g2_fill_2 FILLER_67_1349 ();
 sg13g2_fill_1 FILLER_67_1351 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_decap_8 FILLER_67_1420 ();
 sg13g2_decap_4 FILLER_67_1427 ();
 sg13g2_fill_1 FILLER_67_1431 ();
 sg13g2_decap_8 FILLER_67_1443 ();
 sg13g2_fill_2 FILLER_67_1450 ();
 sg13g2_decap_8 FILLER_67_1457 ();
 sg13g2_decap_8 FILLER_67_1464 ();
 sg13g2_decap_8 FILLER_67_1471 ();
 sg13g2_decap_4 FILLER_67_1478 ();
 sg13g2_fill_2 FILLER_67_1486 ();
 sg13g2_fill_1 FILLER_67_1488 ();
 sg13g2_fill_2 FILLER_67_1522 ();
 sg13g2_fill_1 FILLER_67_1524 ();
 sg13g2_fill_2 FILLER_67_1543 ();
 sg13g2_fill_2 FILLER_67_1554 ();
 sg13g2_fill_1 FILLER_67_1561 ();
 sg13g2_decap_4 FILLER_67_1587 ();
 sg13g2_fill_2 FILLER_67_1591 ();
 sg13g2_fill_2 FILLER_67_1613 ();
 sg13g2_fill_1 FILLER_67_1615 ();
 sg13g2_decap_8 FILLER_67_1621 ();
 sg13g2_decap_8 FILLER_67_1628 ();
 sg13g2_decap_8 FILLER_67_1635 ();
 sg13g2_decap_8 FILLER_67_1642 ();
 sg13g2_decap_8 FILLER_67_1659 ();
 sg13g2_decap_8 FILLER_67_1666 ();
 sg13g2_decap_8 FILLER_67_1673 ();
 sg13g2_decap_8 FILLER_67_1680 ();
 sg13g2_decap_8 FILLER_67_1687 ();
 sg13g2_decap_4 FILLER_67_1694 ();
 sg13g2_fill_1 FILLER_67_1698 ();
 sg13g2_fill_1 FILLER_67_1715 ();
 sg13g2_fill_1 FILLER_67_1747 ();
 sg13g2_decap_4 FILLER_67_1798 ();
 sg13g2_decap_4 FILLER_67_1814 ();
 sg13g2_fill_2 FILLER_67_1818 ();
 sg13g2_decap_8 FILLER_67_1823 ();
 sg13g2_fill_2 FILLER_67_1830 ();
 sg13g2_fill_1 FILLER_67_1832 ();
 sg13g2_fill_2 FILLER_67_1838 ();
 sg13g2_decap_8 FILLER_67_1844 ();
 sg13g2_decap_8 FILLER_67_1851 ();
 sg13g2_decap_8 FILLER_67_1858 ();
 sg13g2_decap_8 FILLER_67_1865 ();
 sg13g2_decap_8 FILLER_67_1872 ();
 sg13g2_decap_4 FILLER_67_1879 ();
 sg13g2_fill_1 FILLER_67_1883 ();
 sg13g2_decap_8 FILLER_67_1890 ();
 sg13g2_decap_8 FILLER_67_1897 ();
 sg13g2_fill_2 FILLER_67_1913 ();
 sg13g2_fill_2 FILLER_67_1920 ();
 sg13g2_fill_2 FILLER_67_1928 ();
 sg13g2_decap_8 FILLER_67_1934 ();
 sg13g2_decap_8 FILLER_67_1941 ();
 sg13g2_decap_4 FILLER_67_1948 ();
 sg13g2_decap_8 FILLER_67_1958 ();
 sg13g2_decap_8 FILLER_67_1965 ();
 sg13g2_decap_8 FILLER_67_1972 ();
 sg13g2_decap_8 FILLER_67_1979 ();
 sg13g2_decap_4 FILLER_67_1986 ();
 sg13g2_fill_1 FILLER_67_1990 ();
 sg13g2_decap_8 FILLER_67_2002 ();
 sg13g2_decap_8 FILLER_67_2009 ();
 sg13g2_decap_8 FILLER_67_2016 ();
 sg13g2_decap_8 FILLER_67_2029 ();
 sg13g2_decap_8 FILLER_67_2036 ();
 sg13g2_decap_8 FILLER_67_2043 ();
 sg13g2_decap_8 FILLER_67_2050 ();
 sg13g2_decap_8 FILLER_67_2057 ();
 sg13g2_decap_8 FILLER_67_2064 ();
 sg13g2_decap_8 FILLER_67_2071 ();
 sg13g2_fill_2 FILLER_67_2078 ();
 sg13g2_decap_8 FILLER_67_2154 ();
 sg13g2_decap_8 FILLER_67_2161 ();
 sg13g2_decap_8 FILLER_67_2168 ();
 sg13g2_fill_1 FILLER_67_2175 ();
 sg13g2_fill_1 FILLER_67_2211 ();
 sg13g2_fill_1 FILLER_67_2242 ();
 sg13g2_fill_1 FILLER_67_2253 ();
 sg13g2_fill_2 FILLER_67_2267 ();
 sg13g2_fill_2 FILLER_67_2283 ();
 sg13g2_fill_1 FILLER_67_2367 ();
 sg13g2_fill_2 FILLER_67_2430 ();
 sg13g2_fill_2 FILLER_67_2436 ();
 sg13g2_fill_1 FILLER_67_2449 ();
 sg13g2_fill_1 FILLER_67_2456 ();
 sg13g2_fill_1 FILLER_67_2489 ();
 sg13g2_fill_2 FILLER_67_2494 ();
 sg13g2_fill_2 FILLER_67_2500 ();
 sg13g2_decap_4 FILLER_67_2535 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_1 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_188 ();
 sg13g2_decap_4 FILLER_68_198 ();
 sg13g2_fill_1 FILLER_68_202 ();
 sg13g2_decap_4 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_224 ();
 sg13g2_fill_1 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_283 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_fill_2 FILLER_68_375 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_68_388 ();
 sg13g2_fill_2 FILLER_68_410 ();
 sg13g2_fill_1 FILLER_68_412 ();
 sg13g2_fill_1 FILLER_68_433 ();
 sg13g2_fill_2 FILLER_68_438 ();
 sg13g2_fill_2 FILLER_68_460 ();
 sg13g2_fill_1 FILLER_68_508 ();
 sg13g2_fill_1 FILLER_68_517 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_fill_1 FILLER_68_571 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_fill_1 FILLER_68_660 ();
 sg13g2_fill_1 FILLER_68_679 ();
 sg13g2_fill_2 FILLER_68_714 ();
 sg13g2_fill_1 FILLER_68_716 ();
 sg13g2_fill_1 FILLER_68_728 ();
 sg13g2_fill_2 FILLER_68_774 ();
 sg13g2_fill_2 FILLER_68_780 ();
 sg13g2_fill_2 FILLER_68_852 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_68_896 ();
 sg13g2_decap_8 FILLER_68_903 ();
 sg13g2_fill_1 FILLER_68_910 ();
 sg13g2_fill_1 FILLER_68_948 ();
 sg13g2_fill_2 FILLER_68_995 ();
 sg13g2_fill_1 FILLER_68_1008 ();
 sg13g2_fill_2 FILLER_68_1012 ();
 sg13g2_fill_2 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1080 ();
 sg13g2_fill_1 FILLER_68_1087 ();
 sg13g2_fill_1 FILLER_68_1110 ();
 sg13g2_decap_4 FILLER_68_1167 ();
 sg13g2_fill_2 FILLER_68_1171 ();
 sg13g2_decap_4 FILLER_68_1213 ();
 sg13g2_fill_1 FILLER_68_1217 ();
 sg13g2_fill_1 FILLER_68_1255 ();
 sg13g2_fill_2 FILLER_68_1270 ();
 sg13g2_fill_1 FILLER_68_1272 ();
 sg13g2_fill_2 FILLER_68_1299 ();
 sg13g2_fill_1 FILLER_68_1301 ();
 sg13g2_fill_1 FILLER_68_1306 ();
 sg13g2_fill_1 FILLER_68_1319 ();
 sg13g2_fill_2 FILLER_68_1330 ();
 sg13g2_fill_1 FILLER_68_1371 ();
 sg13g2_fill_2 FILLER_68_1383 ();
 sg13g2_decap_4 FILLER_68_1390 ();
 sg13g2_decap_4 FILLER_68_1403 ();
 sg13g2_fill_2 FILLER_68_1411 ();
 sg13g2_fill_1 FILLER_68_1413 ();
 sg13g2_fill_1 FILLER_68_1432 ();
 sg13g2_fill_2 FILLER_68_1437 ();
 sg13g2_fill_1 FILLER_68_1444 ();
 sg13g2_fill_2 FILLER_68_1450 ();
 sg13g2_fill_2 FILLER_68_1464 ();
 sg13g2_decap_8 FILLER_68_1490 ();
 sg13g2_decap_4 FILLER_68_1504 ();
 sg13g2_fill_1 FILLER_68_1512 ();
 sg13g2_fill_2 FILLER_68_1547 ();
 sg13g2_fill_2 FILLER_68_1554 ();
 sg13g2_fill_2 FILLER_68_1559 ();
 sg13g2_decap_8 FILLER_68_1567 ();
 sg13g2_fill_2 FILLER_68_1574 ();
 sg13g2_fill_1 FILLER_68_1592 ();
 sg13g2_decap_8 FILLER_68_1627 ();
 sg13g2_decap_8 FILLER_68_1634 ();
 sg13g2_decap_8 FILLER_68_1641 ();
 sg13g2_decap_4 FILLER_68_1648 ();
 sg13g2_fill_2 FILLER_68_1660 ();
 sg13g2_fill_2 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1680 ();
 sg13g2_decap_8 FILLER_68_1687 ();
 sg13g2_fill_1 FILLER_68_1702 ();
 sg13g2_decap_8 FILLER_68_1711 ();
 sg13g2_decap_8 FILLER_68_1718 ();
 sg13g2_fill_2 FILLER_68_1769 ();
 sg13g2_decap_8 FILLER_68_1781 ();
 sg13g2_fill_1 FILLER_68_1788 ();
 sg13g2_decap_4 FILLER_68_1806 ();
 sg13g2_fill_1 FILLER_68_1810 ();
 sg13g2_decap_4 FILLER_68_1816 ();
 sg13g2_fill_1 FILLER_68_1820 ();
 sg13g2_decap_8 FILLER_68_1835 ();
 sg13g2_decap_8 FILLER_68_1842 ();
 sg13g2_decap_8 FILLER_68_1849 ();
 sg13g2_decap_8 FILLER_68_1856 ();
 sg13g2_fill_2 FILLER_68_1863 ();
 sg13g2_decap_8 FILLER_68_1870 ();
 sg13g2_decap_8 FILLER_68_1877 ();
 sg13g2_decap_8 FILLER_68_1884 ();
 sg13g2_decap_8 FILLER_68_1891 ();
 sg13g2_decap_8 FILLER_68_1898 ();
 sg13g2_decap_4 FILLER_68_1905 ();
 sg13g2_decap_8 FILLER_68_1918 ();
 sg13g2_decap_8 FILLER_68_1925 ();
 sg13g2_decap_8 FILLER_68_1932 ();
 sg13g2_decap_8 FILLER_68_1957 ();
 sg13g2_decap_8 FILLER_68_1964 ();
 sg13g2_decap_8 FILLER_68_1971 ();
 sg13g2_fill_2 FILLER_68_1978 ();
 sg13g2_fill_1 FILLER_68_1980 ();
 sg13g2_decap_8 FILLER_68_1986 ();
 sg13g2_decap_8 FILLER_68_1998 ();
 sg13g2_decap_8 FILLER_68_2005 ();
 sg13g2_decap_8 FILLER_68_2012 ();
 sg13g2_decap_8 FILLER_68_2019 ();
 sg13g2_decap_4 FILLER_68_2026 ();
 sg13g2_decap_8 FILLER_68_2036 ();
 sg13g2_decap_8 FILLER_68_2043 ();
 sg13g2_decap_8 FILLER_68_2050 ();
 sg13g2_decap_8 FILLER_68_2057 ();
 sg13g2_decap_8 FILLER_68_2064 ();
 sg13g2_decap_8 FILLER_68_2071 ();
 sg13g2_decap_4 FILLER_68_2078 ();
 sg13g2_fill_2 FILLER_68_2082 ();
 sg13g2_fill_1 FILLER_68_2100 ();
 sg13g2_fill_2 FILLER_68_2105 ();
 sg13g2_fill_1 FILLER_68_2107 ();
 sg13g2_fill_2 FILLER_68_2131 ();
 sg13g2_fill_1 FILLER_68_2133 ();
 sg13g2_fill_2 FILLER_68_2148 ();
 sg13g2_fill_1 FILLER_68_2150 ();
 sg13g2_decap_8 FILLER_68_2161 ();
 sg13g2_decap_8 FILLER_68_2168 ();
 sg13g2_decap_8 FILLER_68_2175 ();
 sg13g2_decap_4 FILLER_68_2187 ();
 sg13g2_fill_2 FILLER_68_2195 ();
 sg13g2_fill_2 FILLER_68_2209 ();
 sg13g2_fill_2 FILLER_68_2219 ();
 sg13g2_fill_2 FILLER_68_2247 ();
 sg13g2_fill_2 FILLER_68_2291 ();
 sg13g2_fill_1 FILLER_68_2333 ();
 sg13g2_fill_1 FILLER_68_2344 ();
 sg13g2_fill_2 FILLER_68_2421 ();
 sg13g2_decap_8 FILLER_68_2470 ();
 sg13g2_decap_8 FILLER_68_2477 ();
 sg13g2_fill_2 FILLER_68_2484 ();
 sg13g2_decap_4 FILLER_68_2490 ();
 sg13g2_fill_2 FILLER_68_2494 ();
 sg13g2_fill_2 FILLER_68_2506 ();
 sg13g2_fill_1 FILLER_68_2518 ();
 sg13g2_fill_1 FILLER_68_2525 ();
 sg13g2_fill_2 FILLER_68_2596 ();
 sg13g2_decap_8 FILLER_68_2638 ();
 sg13g2_decap_8 FILLER_68_2645 ();
 sg13g2_decap_8 FILLER_68_2652 ();
 sg13g2_decap_8 FILLER_68_2659 ();
 sg13g2_decap_4 FILLER_68_2666 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_4 ();
 sg13g2_fill_2 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_43 ();
 sg13g2_fill_2 FILLER_69_58 ();
 sg13g2_fill_2 FILLER_69_65 ();
 sg13g2_fill_2 FILLER_69_82 ();
 sg13g2_fill_2 FILLER_69_139 ();
 sg13g2_decap_4 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_decap_4 FILLER_69_215 ();
 sg13g2_fill_2 FILLER_69_219 ();
 sg13g2_fill_2 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_decap_4 FILLER_69_336 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_2 FILLER_69_419 ();
 sg13g2_fill_2 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_504 ();
 sg13g2_fill_2 FILLER_69_538 ();
 sg13g2_fill_1 FILLER_69_540 ();
 sg13g2_fill_2 FILLER_69_551 ();
 sg13g2_fill_2 FILLER_69_557 ();
 sg13g2_fill_1 FILLER_69_559 ();
 sg13g2_fill_1 FILLER_69_586 ();
 sg13g2_fill_2 FILLER_69_597 ();
 sg13g2_fill_1 FILLER_69_599 ();
 sg13g2_fill_1 FILLER_69_611 ();
 sg13g2_fill_1 FILLER_69_666 ();
 sg13g2_decap_4 FILLER_69_673 ();
 sg13g2_decap_8 FILLER_69_684 ();
 sg13g2_fill_2 FILLER_69_691 ();
 sg13g2_fill_1 FILLER_69_693 ();
 sg13g2_fill_2 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_714 ();
 sg13g2_fill_1 FILLER_69_725 ();
 sg13g2_fill_1 FILLER_69_738 ();
 sg13g2_decap_4 FILLER_69_743 ();
 sg13g2_fill_1 FILLER_69_747 ();
 sg13g2_fill_1 FILLER_69_771 ();
 sg13g2_fill_1 FILLER_69_786 ();
 sg13g2_fill_2 FILLER_69_883 ();
 sg13g2_decap_4 FILLER_69_914 ();
 sg13g2_fill_1 FILLER_69_918 ();
 sg13g2_fill_2 FILLER_69_923 ();
 sg13g2_fill_1 FILLER_69_939 ();
 sg13g2_fill_1 FILLER_69_945 ();
 sg13g2_fill_1 FILLER_69_973 ();
 sg13g2_fill_2 FILLER_69_1003 ();
 sg13g2_fill_2 FILLER_69_1010 ();
 sg13g2_decap_8 FILLER_69_1038 ();
 sg13g2_decap_4 FILLER_69_1045 ();
 sg13g2_fill_1 FILLER_69_1085 ();
 sg13g2_fill_1 FILLER_69_1107 ();
 sg13g2_fill_2 FILLER_69_1144 ();
 sg13g2_decap_4 FILLER_69_1150 ();
 sg13g2_fill_1 FILLER_69_1154 ();
 sg13g2_decap_8 FILLER_69_1159 ();
 sg13g2_decap_8 FILLER_69_1166 ();
 sg13g2_decap_8 FILLER_69_1173 ();
 sg13g2_decap_8 FILLER_69_1180 ();
 sg13g2_decap_8 FILLER_69_1197 ();
 sg13g2_decap_4 FILLER_69_1204 ();
 sg13g2_decap_8 FILLER_69_1253 ();
 sg13g2_fill_2 FILLER_69_1260 ();
 sg13g2_fill_1 FILLER_69_1262 ();
 sg13g2_decap_4 FILLER_69_1268 ();
 sg13g2_fill_1 FILLER_69_1282 ();
 sg13g2_fill_2 FILLER_69_1300 ();
 sg13g2_fill_1 FILLER_69_1302 ();
 sg13g2_decap_8 FILLER_69_1307 ();
 sg13g2_fill_2 FILLER_69_1314 ();
 sg13g2_decap_4 FILLER_69_1326 ();
 sg13g2_fill_1 FILLER_69_1350 ();
 sg13g2_decap_8 FILLER_69_1379 ();
 sg13g2_decap_4 FILLER_69_1386 ();
 sg13g2_fill_1 FILLER_69_1390 ();
 sg13g2_decap_8 FILLER_69_1404 ();
 sg13g2_decap_4 FILLER_69_1411 ();
 sg13g2_fill_2 FILLER_69_1415 ();
 sg13g2_decap_4 FILLER_69_1430 ();
 sg13g2_fill_2 FILLER_69_1434 ();
 sg13g2_fill_2 FILLER_69_1448 ();
 sg13g2_fill_1 FILLER_69_1450 ();
 sg13g2_fill_1 FILLER_69_1458 ();
 sg13g2_decap_8 FILLER_69_1466 ();
 sg13g2_fill_2 FILLER_69_1499 ();
 sg13g2_fill_1 FILLER_69_1523 ();
 sg13g2_decap_4 FILLER_69_1575 ();
 sg13g2_fill_1 FILLER_69_1586 ();
 sg13g2_fill_2 FILLER_69_1591 ();
 sg13g2_fill_2 FILLER_69_1609 ();
 sg13g2_fill_2 FILLER_69_1615 ();
 sg13g2_decap_8 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1635 ();
 sg13g2_decap_8 FILLER_69_1642 ();
 sg13g2_decap_4 FILLER_69_1649 ();
 sg13g2_decap_8 FILLER_69_1663 ();
 sg13g2_decap_8 FILLER_69_1670 ();
 sg13g2_fill_2 FILLER_69_1677 ();
 sg13g2_fill_1 FILLER_69_1679 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_decap_8 FILLER_69_1692 ();
 sg13g2_decap_8 FILLER_69_1699 ();
 sg13g2_decap_8 FILLER_69_1706 ();
 sg13g2_decap_8 FILLER_69_1713 ();
 sg13g2_decap_4 FILLER_69_1720 ();
 sg13g2_decap_4 FILLER_69_1733 ();
 sg13g2_fill_2 FILLER_69_1737 ();
 sg13g2_fill_1 FILLER_69_1754 ();
 sg13g2_decap_8 FILLER_69_1765 ();
 sg13g2_decap_4 FILLER_69_1772 ();
 sg13g2_fill_1 FILLER_69_1776 ();
 sg13g2_fill_2 FILLER_69_1782 ();
 sg13g2_fill_1 FILLER_69_1784 ();
 sg13g2_decap_4 FILLER_69_1791 ();
 sg13g2_fill_1 FILLER_69_1795 ();
 sg13g2_decap_8 FILLER_69_1804 ();
 sg13g2_decap_8 FILLER_69_1811 ();
 sg13g2_decap_8 FILLER_69_1827 ();
 sg13g2_decap_8 FILLER_69_1834 ();
 sg13g2_fill_2 FILLER_69_1841 ();
 sg13g2_fill_2 FILLER_69_1847 ();
 sg13g2_decap_8 FILLER_69_1853 ();
 sg13g2_decap_8 FILLER_69_1860 ();
 sg13g2_decap_8 FILLER_69_1867 ();
 sg13g2_decap_8 FILLER_69_1874 ();
 sg13g2_decap_8 FILLER_69_1881 ();
 sg13g2_decap_8 FILLER_69_1888 ();
 sg13g2_decap_8 FILLER_69_1895 ();
 sg13g2_decap_8 FILLER_69_1902 ();
 sg13g2_decap_8 FILLER_69_1909 ();
 sg13g2_decap_8 FILLER_69_1916 ();
 sg13g2_decap_8 FILLER_69_1923 ();
 sg13g2_decap_4 FILLER_69_1930 ();
 sg13g2_fill_2 FILLER_69_1934 ();
 sg13g2_fill_2 FILLER_69_1941 ();
 sg13g2_decap_8 FILLER_69_1953 ();
 sg13g2_decap_8 FILLER_69_1960 ();
 sg13g2_decap_8 FILLER_69_1967 ();
 sg13g2_decap_4 FILLER_69_1974 ();
 sg13g2_fill_1 FILLER_69_1978 ();
 sg13g2_decap_4 FILLER_69_1985 ();
 sg13g2_fill_2 FILLER_69_1989 ();
 sg13g2_decap_8 FILLER_69_1995 ();
 sg13g2_decap_8 FILLER_69_2002 ();
 sg13g2_decap_8 FILLER_69_2009 ();
 sg13g2_decap_8 FILLER_69_2016 ();
 sg13g2_decap_8 FILLER_69_2023 ();
 sg13g2_decap_8 FILLER_69_2030 ();
 sg13g2_decap_8 FILLER_69_2037 ();
 sg13g2_decap_8 FILLER_69_2044 ();
 sg13g2_decap_8 FILLER_69_2051 ();
 sg13g2_decap_8 FILLER_69_2058 ();
 sg13g2_decap_8 FILLER_69_2065 ();
 sg13g2_decap_8 FILLER_69_2072 ();
 sg13g2_decap_8 FILLER_69_2079 ();
 sg13g2_fill_1 FILLER_69_2114 ();
 sg13g2_fill_2 FILLER_69_2141 ();
 sg13g2_fill_2 FILLER_69_2169 ();
 sg13g2_fill_2 FILLER_69_2197 ();
 sg13g2_fill_1 FILLER_69_2242 ();
 sg13g2_fill_2 FILLER_69_2252 ();
 sg13g2_fill_1 FILLER_69_2335 ();
 sg13g2_fill_1 FILLER_69_2346 ();
 sg13g2_fill_2 FILLER_69_2383 ();
 sg13g2_fill_2 FILLER_69_2415 ();
 sg13g2_fill_1 FILLER_69_2443 ();
 sg13g2_fill_2 FILLER_69_2483 ();
 sg13g2_fill_1 FILLER_69_2558 ();
 sg13g2_fill_2 FILLER_69_2578 ();
 sg13g2_decap_8 FILLER_69_2606 ();
 sg13g2_decap_4 FILLER_69_2613 ();
 sg13g2_fill_2 FILLER_69_2617 ();
 sg13g2_decap_8 FILLER_69_2623 ();
 sg13g2_decap_8 FILLER_69_2630 ();
 sg13g2_decap_8 FILLER_69_2637 ();
 sg13g2_decap_8 FILLER_69_2644 ();
 sg13g2_decap_8 FILLER_69_2651 ();
 sg13g2_decap_8 FILLER_69_2658 ();
 sg13g2_decap_4 FILLER_69_2665 ();
 sg13g2_fill_1 FILLER_69_2669 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_18 ();
 sg13g2_decap_8 FILLER_70_25 ();
 sg13g2_fill_1 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_87 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_decap_4 FILLER_70_98 ();
 sg13g2_decap_4 FILLER_70_112 ();
 sg13g2_decap_4 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_124 ();
 sg13g2_fill_1 FILLER_70_169 ();
 sg13g2_fill_1 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_1 FILLER_70_249 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_269 ();
 sg13g2_decap_4 FILLER_70_302 ();
 sg13g2_fill_2 FILLER_70_317 ();
 sg13g2_decap_4 FILLER_70_324 ();
 sg13g2_decap_4 FILLER_70_359 ();
 sg13g2_fill_2 FILLER_70_363 ();
 sg13g2_decap_8 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_decap_4 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_397 ();
 sg13g2_fill_1 FILLER_70_399 ();
 sg13g2_fill_2 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_416 ();
 sg13g2_fill_2 FILLER_70_455 ();
 sg13g2_fill_1 FILLER_70_457 ();
 sg13g2_fill_1 FILLER_70_471 ();
 sg13g2_fill_2 FILLER_70_485 ();
 sg13g2_fill_1 FILLER_70_487 ();
 sg13g2_fill_1 FILLER_70_529 ();
 sg13g2_fill_1 FILLER_70_543 ();
 sg13g2_fill_2 FILLER_70_554 ();
 sg13g2_decap_8 FILLER_70_560 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_fill_1 FILLER_70_596 ();
 sg13g2_fill_1 FILLER_70_620 ();
 sg13g2_fill_1 FILLER_70_646 ();
 sg13g2_fill_1 FILLER_70_651 ();
 sg13g2_decap_8 FILLER_70_682 ();
 sg13g2_fill_1 FILLER_70_689 ();
 sg13g2_fill_2 FILLER_70_733 ();
 sg13g2_decap_4 FILLER_70_745 ();
 sg13g2_fill_1 FILLER_70_836 ();
 sg13g2_fill_2 FILLER_70_851 ();
 sg13g2_fill_1 FILLER_70_857 ();
 sg13g2_fill_2 FILLER_70_893 ();
 sg13g2_decap_4 FILLER_70_926 ();
 sg13g2_fill_2 FILLER_70_942 ();
 sg13g2_fill_2 FILLER_70_959 ();
 sg13g2_fill_1 FILLER_70_999 ();
 sg13g2_decap_8 FILLER_70_1033 ();
 sg13g2_decap_8 FILLER_70_1048 ();
 sg13g2_decap_4 FILLER_70_1055 ();
 sg13g2_fill_2 FILLER_70_1063 ();
 sg13g2_fill_2 FILLER_70_1083 ();
 sg13g2_fill_1 FILLER_70_1085 ();
 sg13g2_fill_2 FILLER_70_1100 ();
 sg13g2_fill_1 FILLER_70_1102 ();
 sg13g2_fill_1 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1148 ();
 sg13g2_fill_2 FILLER_70_1155 ();
 sg13g2_decap_8 FILLER_70_1189 ();
 sg13g2_decap_4 FILLER_70_1200 ();
 sg13g2_fill_1 FILLER_70_1204 ();
 sg13g2_fill_1 FILLER_70_1210 ();
 sg13g2_fill_1 FILLER_70_1247 ();
 sg13g2_decap_4 FILLER_70_1252 ();
 sg13g2_decap_4 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1322 ();
 sg13g2_fill_2 FILLER_70_1329 ();
 sg13g2_decap_8 FILLER_70_1337 ();
 sg13g2_decap_8 FILLER_70_1377 ();
 sg13g2_decap_8 FILLER_70_1384 ();
 sg13g2_decap_8 FILLER_70_1391 ();
 sg13g2_decap_8 FILLER_70_1398 ();
 sg13g2_decap_4 FILLER_70_1441 ();
 sg13g2_fill_1 FILLER_70_1465 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_fill_2 FILLER_70_1481 ();
 sg13g2_fill_1 FILLER_70_1483 ();
 sg13g2_fill_1 FILLER_70_1488 ();
 sg13g2_fill_1 FILLER_70_1497 ();
 sg13g2_fill_1 FILLER_70_1502 ();
 sg13g2_fill_1 FILLER_70_1516 ();
 sg13g2_fill_2 FILLER_70_1527 ();
 sg13g2_fill_2 FILLER_70_1533 ();
 sg13g2_fill_1 FILLER_70_1535 ();
 sg13g2_fill_1 FILLER_70_1541 ();
 sg13g2_fill_2 FILLER_70_1555 ();
 sg13g2_decap_8 FILLER_70_1562 ();
 sg13g2_decap_4 FILLER_70_1578 ();
 sg13g2_fill_2 FILLER_70_1587 ();
 sg13g2_fill_1 FILLER_70_1589 ();
 sg13g2_fill_1 FILLER_70_1594 ();
 sg13g2_decap_4 FILLER_70_1603 ();
 sg13g2_fill_1 FILLER_70_1607 ();
 sg13g2_decap_8 FILLER_70_1611 ();
 sg13g2_decap_8 FILLER_70_1618 ();
 sg13g2_decap_8 FILLER_70_1625 ();
 sg13g2_decap_8 FILLER_70_1632 ();
 sg13g2_decap_8 FILLER_70_1639 ();
 sg13g2_fill_2 FILLER_70_1646 ();
 sg13g2_fill_1 FILLER_70_1648 ();
 sg13g2_decap_8 FILLER_70_1662 ();
 sg13g2_decap_8 FILLER_70_1669 ();
 sg13g2_decap_8 FILLER_70_1681 ();
 sg13g2_decap_8 FILLER_70_1688 ();
 sg13g2_decap_8 FILLER_70_1695 ();
 sg13g2_decap_4 FILLER_70_1708 ();
 sg13g2_decap_4 FILLER_70_1717 ();
 sg13g2_fill_2 FILLER_70_1721 ();
 sg13g2_decap_8 FILLER_70_1727 ();
 sg13g2_decap_8 FILLER_70_1734 ();
 sg13g2_decap_8 FILLER_70_1741 ();
 sg13g2_decap_8 FILLER_70_1748 ();
 sg13g2_decap_4 FILLER_70_1755 ();
 sg13g2_fill_2 FILLER_70_1764 ();
 sg13g2_fill_1 FILLER_70_1766 ();
 sg13g2_decap_8 FILLER_70_1771 ();
 sg13g2_decap_8 FILLER_70_1778 ();
 sg13g2_fill_1 FILLER_70_1785 ();
 sg13g2_decap_8 FILLER_70_1796 ();
 sg13g2_decap_4 FILLER_70_1803 ();
 sg13g2_fill_2 FILLER_70_1807 ();
 sg13g2_decap_8 FILLER_70_1814 ();
 sg13g2_decap_8 FILLER_70_1821 ();
 sg13g2_fill_1 FILLER_70_1828 ();
 sg13g2_decap_8 FILLER_70_1834 ();
 sg13g2_decap_8 FILLER_70_1849 ();
 sg13g2_decap_8 FILLER_70_1856 ();
 sg13g2_decap_8 FILLER_70_1863 ();
 sg13g2_decap_8 FILLER_70_1870 ();
 sg13g2_decap_8 FILLER_70_1877 ();
 sg13g2_decap_8 FILLER_70_1884 ();
 sg13g2_decap_4 FILLER_70_1891 ();
 sg13g2_fill_2 FILLER_70_1895 ();
 sg13g2_decap_8 FILLER_70_1902 ();
 sg13g2_decap_8 FILLER_70_1909 ();
 sg13g2_decap_8 FILLER_70_1916 ();
 sg13g2_decap_8 FILLER_70_1923 ();
 sg13g2_decap_8 FILLER_70_1930 ();
 sg13g2_decap_8 FILLER_70_1937 ();
 sg13g2_decap_8 FILLER_70_1944 ();
 sg13g2_decap_8 FILLER_70_1951 ();
 sg13g2_decap_8 FILLER_70_1958 ();
 sg13g2_decap_8 FILLER_70_1965 ();
 sg13g2_decap_8 FILLER_70_1972 ();
 sg13g2_decap_8 FILLER_70_1979 ();
 sg13g2_decap_8 FILLER_70_1990 ();
 sg13g2_decap_8 FILLER_70_1997 ();
 sg13g2_decap_8 FILLER_70_2004 ();
 sg13g2_decap_8 FILLER_70_2011 ();
 sg13g2_fill_2 FILLER_70_2018 ();
 sg13g2_decap_8 FILLER_70_2026 ();
 sg13g2_decap_8 FILLER_70_2033 ();
 sg13g2_decap_8 FILLER_70_2040 ();
 sg13g2_decap_8 FILLER_70_2047 ();
 sg13g2_decap_8 FILLER_70_2054 ();
 sg13g2_decap_8 FILLER_70_2061 ();
 sg13g2_decap_8 FILLER_70_2068 ();
 sg13g2_decap_8 FILLER_70_2075 ();
 sg13g2_decap_8 FILLER_70_2082 ();
 sg13g2_decap_8 FILLER_70_2089 ();
 sg13g2_fill_1 FILLER_70_2096 ();
 sg13g2_decap_8 FILLER_70_2132 ();
 sg13g2_fill_2 FILLER_70_2139 ();
 sg13g2_fill_2 FILLER_70_2206 ();
 sg13g2_fill_1 FILLER_70_2208 ();
 sg13g2_fill_1 FILLER_70_2244 ();
 sg13g2_fill_2 FILLER_70_2271 ();
 sg13g2_fill_1 FILLER_70_2277 ();
 sg13g2_fill_1 FILLER_70_2282 ();
 sg13g2_fill_1 FILLER_70_2287 ();
 sg13g2_fill_2 FILLER_70_2296 ();
 sg13g2_fill_1 FILLER_70_2328 ();
 sg13g2_fill_2 FILLER_70_2416 ();
 sg13g2_fill_1 FILLER_70_2518 ();
 sg13g2_fill_1 FILLER_70_2523 ();
 sg13g2_fill_1 FILLER_70_2534 ();
 sg13g2_fill_2 FILLER_70_2553 ();
 sg13g2_fill_1 FILLER_70_2575 ();
 sg13g2_decap_8 FILLER_70_2614 ();
 sg13g2_decap_8 FILLER_70_2621 ();
 sg13g2_decap_8 FILLER_70_2628 ();
 sg13g2_decap_8 FILLER_70_2635 ();
 sg13g2_decap_8 FILLER_70_2642 ();
 sg13g2_decap_8 FILLER_70_2649 ();
 sg13g2_decap_8 FILLER_70_2656 ();
 sg13g2_decap_8 FILLER_70_2663 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_39 ();
 sg13g2_fill_1 FILLER_71_67 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_2 FILLER_71_92 ();
 sg13g2_fill_2 FILLER_71_99 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_205 ();
 sg13g2_decap_4 FILLER_71_212 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_decap_4 FILLER_71_226 ();
 sg13g2_fill_2 FILLER_71_230 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_fill_2 FILLER_71_257 ();
 sg13g2_fill_1 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_284 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_decap_8 FILLER_71_316 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_4 FILLER_71_330 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_4 FILLER_71_371 ();
 sg13g2_fill_1 FILLER_71_375 ();
 sg13g2_decap_4 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_decap_4 FILLER_71_475 ();
 sg13g2_fill_2 FILLER_71_479 ();
 sg13g2_fill_1 FILLER_71_516 ();
 sg13g2_decap_8 FILLER_71_521 ();
 sg13g2_fill_1 FILLER_71_528 ();
 sg13g2_fill_1 FILLER_71_533 ();
 sg13g2_fill_2 FILLER_71_561 ();
 sg13g2_fill_1 FILLER_71_577 ();
 sg13g2_fill_1 FILLER_71_582 ();
 sg13g2_decap_8 FILLER_71_592 ();
 sg13g2_decap_4 FILLER_71_599 ();
 sg13g2_fill_2 FILLER_71_645 ();
 sg13g2_fill_1 FILLER_71_666 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_fill_2 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_685 ();
 sg13g2_fill_2 FILLER_71_723 ();
 sg13g2_fill_1 FILLER_71_780 ();
 sg13g2_fill_2 FILLER_71_789 ();
 sg13g2_fill_2 FILLER_71_796 ();
 sg13g2_fill_1 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_873 ();
 sg13g2_fill_2 FILLER_71_882 ();
 sg13g2_fill_1 FILLER_71_893 ();
 sg13g2_fill_2 FILLER_71_985 ();
 sg13g2_decap_8 FILLER_71_1022 ();
 sg13g2_decap_8 FILLER_71_1029 ();
 sg13g2_decap_8 FILLER_71_1036 ();
 sg13g2_decap_8 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_fill_1 FILLER_71_1057 ();
 sg13g2_fill_2 FILLER_71_1062 ();
 sg13g2_fill_1 FILLER_71_1064 ();
 sg13g2_fill_2 FILLER_71_1073 ();
 sg13g2_fill_1 FILLER_71_1075 ();
 sg13g2_fill_2 FILLER_71_1105 ();
 sg13g2_fill_1 FILLER_71_1107 ();
 sg13g2_decap_4 FILLER_71_1143 ();
 sg13g2_fill_2 FILLER_71_1147 ();
 sg13g2_fill_2 FILLER_71_1173 ();
 sg13g2_fill_1 FILLER_71_1175 ();
 sg13g2_decap_8 FILLER_71_1241 ();
 sg13g2_decap_4 FILLER_71_1248 ();
 sg13g2_fill_1 FILLER_71_1252 ();
 sg13g2_fill_1 FILLER_71_1269 ();
 sg13g2_fill_1 FILLER_71_1296 ();
 sg13g2_decap_8 FILLER_71_1301 ();
 sg13g2_decap_8 FILLER_71_1308 ();
 sg13g2_decap_8 FILLER_71_1319 ();
 sg13g2_fill_2 FILLER_71_1326 ();
 sg13g2_decap_8 FILLER_71_1336 ();
 sg13g2_fill_2 FILLER_71_1343 ();
 sg13g2_fill_1 FILLER_71_1345 ();
 sg13g2_decap_8 FILLER_71_1358 ();
 sg13g2_decap_8 FILLER_71_1365 ();
 sg13g2_fill_2 FILLER_71_1385 ();
 sg13g2_fill_1 FILLER_71_1387 ();
 sg13g2_fill_1 FILLER_71_1413 ();
 sg13g2_decap_8 FILLER_71_1421 ();
 sg13g2_fill_2 FILLER_71_1428 ();
 sg13g2_fill_1 FILLER_71_1442 ();
 sg13g2_fill_1 FILLER_71_1461 ();
 sg13g2_fill_1 FILLER_71_1475 ();
 sg13g2_fill_1 FILLER_71_1481 ();
 sg13g2_fill_1 FILLER_71_1513 ();
 sg13g2_fill_1 FILLER_71_1518 ();
 sg13g2_decap_4 FILLER_71_1532 ();
 sg13g2_fill_1 FILLER_71_1540 ();
 sg13g2_decap_8 FILLER_71_1546 ();
 sg13g2_decap_8 FILLER_71_1553 ();
 sg13g2_decap_4 FILLER_71_1560 ();
 sg13g2_fill_2 FILLER_71_1564 ();
 sg13g2_fill_2 FILLER_71_1580 ();
 sg13g2_decap_8 FILLER_71_1620 ();
 sg13g2_decap_8 FILLER_71_1627 ();
 sg13g2_decap_8 FILLER_71_1634 ();
 sg13g2_decap_4 FILLER_71_1641 ();
 sg13g2_fill_1 FILLER_71_1645 ();
 sg13g2_decap_4 FILLER_71_1654 ();
 sg13g2_fill_2 FILLER_71_1658 ();
 sg13g2_decap_8 FILLER_71_1664 ();
 sg13g2_decap_8 FILLER_71_1671 ();
 sg13g2_decap_8 FILLER_71_1682 ();
 sg13g2_decap_8 FILLER_71_1689 ();
 sg13g2_fill_2 FILLER_71_1696 ();
 sg13g2_fill_1 FILLER_71_1698 ();
 sg13g2_fill_2 FILLER_71_1709 ();
 sg13g2_decap_8 FILLER_71_1715 ();
 sg13g2_decap_8 FILLER_71_1722 ();
 sg13g2_fill_1 FILLER_71_1729 ();
 sg13g2_decap_8 FILLER_71_1734 ();
 sg13g2_decap_8 FILLER_71_1741 ();
 sg13g2_decap_8 FILLER_71_1748 ();
 sg13g2_decap_8 FILLER_71_1755 ();
 sg13g2_fill_1 FILLER_71_1766 ();
 sg13g2_fill_2 FILLER_71_1773 ();
 sg13g2_decap_4 FILLER_71_1785 ();
 sg13g2_fill_2 FILLER_71_1789 ();
 sg13g2_decap_8 FILLER_71_1795 ();
 sg13g2_decap_8 FILLER_71_1802 ();
 sg13g2_decap_8 FILLER_71_1809 ();
 sg13g2_decap_8 FILLER_71_1816 ();
 sg13g2_decap_8 FILLER_71_1823 ();
 sg13g2_decap_8 FILLER_71_1830 ();
 sg13g2_decap_8 FILLER_71_1837 ();
 sg13g2_decap_8 FILLER_71_1844 ();
 sg13g2_decap_8 FILLER_71_1851 ();
 sg13g2_decap_4 FILLER_71_1858 ();
 sg13g2_fill_1 FILLER_71_1862 ();
 sg13g2_decap_8 FILLER_71_1868 ();
 sg13g2_decap_8 FILLER_71_1875 ();
 sg13g2_fill_2 FILLER_71_1882 ();
 sg13g2_fill_1 FILLER_71_1884 ();
 sg13g2_fill_1 FILLER_71_1899 ();
 sg13g2_fill_1 FILLER_71_1905 ();
 sg13g2_decap_8 FILLER_71_1910 ();
 sg13g2_decap_8 FILLER_71_1917 ();
 sg13g2_decap_8 FILLER_71_1924 ();
 sg13g2_decap_8 FILLER_71_1931 ();
 sg13g2_decap_8 FILLER_71_1938 ();
 sg13g2_fill_1 FILLER_71_1945 ();
 sg13g2_decap_8 FILLER_71_1952 ();
 sg13g2_decap_8 FILLER_71_1959 ();
 sg13g2_decap_8 FILLER_71_1966 ();
 sg13g2_decap_8 FILLER_71_1973 ();
 sg13g2_fill_2 FILLER_71_1980 ();
 sg13g2_decap_8 FILLER_71_1992 ();
 sg13g2_decap_8 FILLER_71_1999 ();
 sg13g2_decap_8 FILLER_71_2006 ();
 sg13g2_fill_1 FILLER_71_2013 ();
 sg13g2_decap_4 FILLER_71_2025 ();
 sg13g2_fill_1 FILLER_71_2029 ();
 sg13g2_decap_8 FILLER_71_2036 ();
 sg13g2_decap_8 FILLER_71_2043 ();
 sg13g2_decap_8 FILLER_71_2050 ();
 sg13g2_decap_8 FILLER_71_2057 ();
 sg13g2_decap_8 FILLER_71_2064 ();
 sg13g2_decap_8 FILLER_71_2071 ();
 sg13g2_decap_8 FILLER_71_2078 ();
 sg13g2_fill_2 FILLER_71_2155 ();
 sg13g2_fill_1 FILLER_71_2163 ();
 sg13g2_fill_1 FILLER_71_2200 ();
 sg13g2_fill_1 FILLER_71_2206 ();
 sg13g2_fill_2 FILLER_71_2380 ();
 sg13g2_fill_2 FILLER_71_2392 ();
 sg13g2_fill_1 FILLER_71_2445 ();
 sg13g2_fill_1 FILLER_71_2529 ();
 sg13g2_fill_2 FILLER_71_2572 ();
 sg13g2_decap_8 FILLER_71_2603 ();
 sg13g2_decap_8 FILLER_71_2610 ();
 sg13g2_decap_8 FILLER_71_2617 ();
 sg13g2_decap_8 FILLER_71_2624 ();
 sg13g2_decap_8 FILLER_71_2631 ();
 sg13g2_decap_8 FILLER_71_2638 ();
 sg13g2_decap_8 FILLER_71_2645 ();
 sg13g2_decap_8 FILLER_71_2652 ();
 sg13g2_decap_8 FILLER_71_2659 ();
 sg13g2_decap_4 FILLER_71_2666 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_41 ();
 sg13g2_fill_2 FILLER_72_76 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_1 FILLER_72_109 ();
 sg13g2_fill_1 FILLER_72_152 ();
 sg13g2_fill_1 FILLER_72_168 ();
 sg13g2_fill_1 FILLER_72_178 ();
 sg13g2_decap_4 FILLER_72_183 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_fill_2 FILLER_72_193 ();
 sg13g2_fill_1 FILLER_72_195 ();
 sg13g2_fill_2 FILLER_72_201 ();
 sg13g2_fill_1 FILLER_72_203 ();
 sg13g2_decap_4 FILLER_72_230 ();
 sg13g2_decap_4 FILLER_72_239 ();
 sg13g2_fill_2 FILLER_72_243 ();
 sg13g2_decap_8 FILLER_72_253 ();
 sg13g2_fill_1 FILLER_72_260 ();
 sg13g2_fill_2 FILLER_72_275 ();
 sg13g2_fill_2 FILLER_72_292 ();
 sg13g2_fill_1 FILLER_72_299 ();
 sg13g2_decap_4 FILLER_72_312 ();
 sg13g2_fill_1 FILLER_72_316 ();
 sg13g2_decap_8 FILLER_72_347 ();
 sg13g2_decap_8 FILLER_72_354 ();
 sg13g2_decap_8 FILLER_72_361 ();
 sg13g2_decap_4 FILLER_72_368 ();
 sg13g2_fill_1 FILLER_72_392 ();
 sg13g2_fill_2 FILLER_72_419 ();
 sg13g2_fill_1 FILLER_72_421 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_492 ();
 sg13g2_fill_2 FILLER_72_515 ();
 sg13g2_fill_1 FILLER_72_517 ();
 sg13g2_fill_1 FILLER_72_544 ();
 sg13g2_fill_1 FILLER_72_582 ();
 sg13g2_fill_1 FILLER_72_589 ();
 sg13g2_fill_1 FILLER_72_600 ();
 sg13g2_fill_1 FILLER_72_627 ();
 sg13g2_fill_1 FILLER_72_634 ();
 sg13g2_fill_1 FILLER_72_641 ();
 sg13g2_fill_1 FILLER_72_650 ();
 sg13g2_fill_1 FILLER_72_697 ();
 sg13g2_fill_2 FILLER_72_717 ();
 sg13g2_fill_1 FILLER_72_729 ();
 sg13g2_fill_2 FILLER_72_740 ();
 sg13g2_fill_1 FILLER_72_746 ();
 sg13g2_fill_1 FILLER_72_796 ();
 sg13g2_fill_1 FILLER_72_805 ();
 sg13g2_fill_2 FILLER_72_813 ();
 sg13g2_fill_2 FILLER_72_872 ();
 sg13g2_fill_2 FILLER_72_884 ();
 sg13g2_fill_1 FILLER_72_904 ();
 sg13g2_fill_1 FILLER_72_931 ();
 sg13g2_fill_1 FILLER_72_945 ();
 sg13g2_fill_1 FILLER_72_955 ();
 sg13g2_fill_2 FILLER_72_978 ();
 sg13g2_fill_2 FILLER_72_1011 ();
 sg13g2_fill_2 FILLER_72_1026 ();
 sg13g2_fill_1 FILLER_72_1028 ();
 sg13g2_fill_1 FILLER_72_1069 ();
 sg13g2_fill_2 FILLER_72_1080 ();
 sg13g2_fill_1 FILLER_72_1092 ();
 sg13g2_decap_8 FILLER_72_1132 ();
 sg13g2_decap_8 FILLER_72_1139 ();
 sg13g2_decap_8 FILLER_72_1146 ();
 sg13g2_fill_1 FILLER_72_1153 ();
 sg13g2_decap_4 FILLER_72_1238 ();
 sg13g2_fill_2 FILLER_72_1242 ();
 sg13g2_fill_2 FILLER_72_1248 ();
 sg13g2_fill_2 FILLER_72_1256 ();
 sg13g2_fill_2 FILLER_72_1279 ();
 sg13g2_fill_2 FILLER_72_1285 ();
 sg13g2_fill_1 FILLER_72_1287 ();
 sg13g2_decap_4 FILLER_72_1327 ();
 sg13g2_decap_8 FILLER_72_1343 ();
 sg13g2_fill_2 FILLER_72_1376 ();
 sg13g2_fill_1 FILLER_72_1378 ();
 sg13g2_fill_1 FILLER_72_1399 ();
 sg13g2_fill_2 FILLER_72_1406 ();
 sg13g2_fill_1 FILLER_72_1413 ();
 sg13g2_fill_1 FILLER_72_1421 ();
 sg13g2_fill_1 FILLER_72_1427 ();
 sg13g2_decap_4 FILLER_72_1438 ();
 sg13g2_fill_1 FILLER_72_1450 ();
 sg13g2_fill_1 FILLER_72_1456 ();
 sg13g2_fill_1 FILLER_72_1462 ();
 sg13g2_fill_1 FILLER_72_1477 ();
 sg13g2_fill_1 FILLER_72_1526 ();
 sg13g2_decap_8 FILLER_72_1534 ();
 sg13g2_decap_8 FILLER_72_1544 ();
 sg13g2_decap_8 FILLER_72_1551 ();
 sg13g2_fill_2 FILLER_72_1558 ();
 sg13g2_fill_1 FILLER_72_1583 ();
 sg13g2_fill_1 FILLER_72_1599 ();
 sg13g2_fill_1 FILLER_72_1605 ();
 sg13g2_fill_1 FILLER_72_1611 ();
 sg13g2_decap_8 FILLER_72_1616 ();
 sg13g2_decap_8 FILLER_72_1623 ();
 sg13g2_decap_8 FILLER_72_1630 ();
 sg13g2_decap_8 FILLER_72_1637 ();
 sg13g2_decap_8 FILLER_72_1644 ();
 sg13g2_decap_4 FILLER_72_1651 ();
 sg13g2_fill_2 FILLER_72_1655 ();
 sg13g2_decap_8 FILLER_72_1665 ();
 sg13g2_decap_8 FILLER_72_1672 ();
 sg13g2_decap_8 FILLER_72_1683 ();
 sg13g2_decap_8 FILLER_72_1690 ();
 sg13g2_fill_2 FILLER_72_1697 ();
 sg13g2_fill_1 FILLER_72_1699 ();
 sg13g2_decap_8 FILLER_72_1704 ();
 sg13g2_decap_8 FILLER_72_1711 ();
 sg13g2_decap_8 FILLER_72_1718 ();
 sg13g2_decap_8 FILLER_72_1725 ();
 sg13g2_decap_8 FILLER_72_1732 ();
 sg13g2_decap_8 FILLER_72_1739 ();
 sg13g2_decap_8 FILLER_72_1746 ();
 sg13g2_decap_8 FILLER_72_1753 ();
 sg13g2_fill_1 FILLER_72_1760 ();
 sg13g2_decap_8 FILLER_72_1766 ();
 sg13g2_decap_8 FILLER_72_1773 ();
 sg13g2_decap_8 FILLER_72_1784 ();
 sg13g2_decap_8 FILLER_72_1791 ();
 sg13g2_decap_8 FILLER_72_1798 ();
 sg13g2_decap_8 FILLER_72_1805 ();
 sg13g2_decap_8 FILLER_72_1812 ();
 sg13g2_decap_8 FILLER_72_1819 ();
 sg13g2_decap_4 FILLER_72_1826 ();
 sg13g2_decap_8 FILLER_72_1835 ();
 sg13g2_decap_4 FILLER_72_1842 ();
 sg13g2_fill_2 FILLER_72_1846 ();
 sg13g2_fill_2 FILLER_72_1854 ();
 sg13g2_decap_8 FILLER_72_1863 ();
 sg13g2_decap_8 FILLER_72_1870 ();
 sg13g2_decap_8 FILLER_72_1877 ();
 sg13g2_decap_8 FILLER_72_1889 ();
 sg13g2_decap_8 FILLER_72_1896 ();
 sg13g2_decap_8 FILLER_72_1903 ();
 sg13g2_decap_8 FILLER_72_1910 ();
 sg13g2_decap_8 FILLER_72_1917 ();
 sg13g2_decap_8 FILLER_72_1924 ();
 sg13g2_decap_8 FILLER_72_1931 ();
 sg13g2_fill_2 FILLER_72_1938 ();
 sg13g2_decap_8 FILLER_72_1957 ();
 sg13g2_decap_8 FILLER_72_1964 ();
 sg13g2_decap_8 FILLER_72_1971 ();
 sg13g2_decap_4 FILLER_72_1978 ();
 sg13g2_fill_1 FILLER_72_1982 ();
 sg13g2_decap_8 FILLER_72_1989 ();
 sg13g2_decap_8 FILLER_72_1996 ();
 sg13g2_decap_8 FILLER_72_2003 ();
 sg13g2_decap_8 FILLER_72_2010 ();
 sg13g2_decap_8 FILLER_72_2017 ();
 sg13g2_decap_8 FILLER_72_2024 ();
 sg13g2_decap_8 FILLER_72_2031 ();
 sg13g2_fill_1 FILLER_72_2038 ();
 sg13g2_decap_8 FILLER_72_2045 ();
 sg13g2_decap_8 FILLER_72_2052 ();
 sg13g2_decap_8 FILLER_72_2059 ();
 sg13g2_decap_8 FILLER_72_2066 ();
 sg13g2_decap_8 FILLER_72_2073 ();
 sg13g2_decap_8 FILLER_72_2080 ();
 sg13g2_fill_2 FILLER_72_2169 ();
 sg13g2_fill_1 FILLER_72_2175 ();
 sg13g2_fill_2 FILLER_72_2208 ();
 sg13g2_fill_1 FILLER_72_2210 ();
 sg13g2_fill_1 FILLER_72_2241 ();
 sg13g2_fill_2 FILLER_72_2246 ();
 sg13g2_fill_1 FILLER_72_2248 ();
 sg13g2_fill_1 FILLER_72_2284 ();
 sg13g2_fill_1 FILLER_72_2333 ();
 sg13g2_fill_1 FILLER_72_2406 ();
 sg13g2_fill_1 FILLER_72_2449 ();
 sg13g2_fill_1 FILLER_72_2500 ();
 sg13g2_fill_1 FILLER_72_2518 ();
 sg13g2_fill_2 FILLER_72_2525 ();
 sg13g2_fill_1 FILLER_72_2576 ();
 sg13g2_decap_8 FILLER_72_2629 ();
 sg13g2_decap_8 FILLER_72_2636 ();
 sg13g2_decap_8 FILLER_72_2643 ();
 sg13g2_decap_8 FILLER_72_2650 ();
 sg13g2_decap_8 FILLER_72_2657 ();
 sg13g2_decap_4 FILLER_72_2664 ();
 sg13g2_fill_2 FILLER_72_2668 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_27 ();
 sg13g2_fill_2 FILLER_73_34 ();
 sg13g2_fill_2 FILLER_73_40 ();
 sg13g2_fill_1 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_79 ();
 sg13g2_fill_1 FILLER_73_120 ();
 sg13g2_fill_1 FILLER_73_126 ();
 sg13g2_fill_1 FILLER_73_148 ();
 sg13g2_fill_2 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_164 ();
 sg13g2_fill_1 FILLER_73_166 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_decap_4 FILLER_73_203 ();
 sg13g2_fill_2 FILLER_73_207 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_decap_4 FILLER_73_251 ();
 sg13g2_fill_1 FILLER_73_255 ();
 sg13g2_fill_2 FILLER_73_264 ();
 sg13g2_decap_4 FILLER_73_271 ();
 sg13g2_fill_1 FILLER_73_275 ();
 sg13g2_fill_1 FILLER_73_316 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_368 ();
 sg13g2_fill_1 FILLER_73_390 ();
 sg13g2_decap_4 FILLER_73_476 ();
 sg13g2_decap_8 FILLER_73_506 ();
 sg13g2_fill_1 FILLER_73_521 ();
 sg13g2_fill_2 FILLER_73_553 ();
 sg13g2_fill_1 FILLER_73_559 ();
 sg13g2_fill_1 FILLER_73_586 ();
 sg13g2_fill_1 FILLER_73_593 ();
 sg13g2_fill_1 FILLER_73_599 ();
 sg13g2_fill_1 FILLER_73_626 ();
 sg13g2_fill_1 FILLER_73_643 ();
 sg13g2_fill_2 FILLER_73_651 ();
 sg13g2_fill_2 FILLER_73_661 ();
 sg13g2_fill_1 FILLER_73_667 ();
 sg13g2_fill_2 FILLER_73_700 ();
 sg13g2_fill_1 FILLER_73_770 ();
 sg13g2_fill_2 FILLER_73_775 ();
 sg13g2_fill_1 FILLER_73_840 ();
 sg13g2_fill_1 FILLER_73_844 ();
 sg13g2_fill_1 FILLER_73_865 ();
 sg13g2_fill_1 FILLER_73_874 ();
 sg13g2_fill_1 FILLER_73_886 ();
 sg13g2_fill_2 FILLER_73_926 ();
 sg13g2_fill_2 FILLER_73_932 ();
 sg13g2_fill_1 FILLER_73_938 ();
 sg13g2_fill_2 FILLER_73_967 ();
 sg13g2_fill_1 FILLER_73_1025 ();
 sg13g2_fill_2 FILLER_73_1146 ();
 sg13g2_decap_8 FILLER_73_1153 ();
 sg13g2_decap_4 FILLER_73_1160 ();
 sg13g2_fill_2 FILLER_73_1164 ();
 sg13g2_fill_1 FILLER_73_1185 ();
 sg13g2_fill_2 FILLER_73_1196 ();
 sg13g2_fill_1 FILLER_73_1198 ();
 sg13g2_decap_4 FILLER_73_1216 ();
 sg13g2_decap_8 FILLER_73_1308 ();
 sg13g2_decap_8 FILLER_73_1315 ();
 sg13g2_fill_2 FILLER_73_1322 ();
 sg13g2_fill_1 FILLER_73_1328 ();
 sg13g2_fill_2 FILLER_73_1334 ();
 sg13g2_fill_2 FILLER_73_1351 ();
 sg13g2_fill_1 FILLER_73_1353 ();
 sg13g2_fill_1 FILLER_73_1366 ();
 sg13g2_fill_1 FILLER_73_1380 ();
 sg13g2_fill_1 FILLER_73_1392 ();
 sg13g2_fill_2 FILLER_73_1398 ();
 sg13g2_fill_1 FILLER_73_1400 ();
 sg13g2_fill_2 FILLER_73_1409 ();
 sg13g2_decap_4 FILLER_73_1420 ();
 sg13g2_fill_2 FILLER_73_1424 ();
 sg13g2_fill_2 FILLER_73_1439 ();
 sg13g2_fill_1 FILLER_73_1446 ();
 sg13g2_fill_1 FILLER_73_1452 ();
 sg13g2_fill_1 FILLER_73_1457 ();
 sg13g2_fill_2 FILLER_73_1463 ();
 sg13g2_fill_1 FILLER_73_1469 ();
 sg13g2_fill_1 FILLER_73_1533 ();
 sg13g2_fill_1 FILLER_73_1546 ();
 sg13g2_fill_2 FILLER_73_1577 ();
 sg13g2_fill_1 FILLER_73_1579 ();
 sg13g2_fill_1 FILLER_73_1586 ();
 sg13g2_fill_1 FILLER_73_1598 ();
 sg13g2_decap_4 FILLER_73_1604 ();
 sg13g2_fill_2 FILLER_73_1608 ();
 sg13g2_decap_8 FILLER_73_1615 ();
 sg13g2_decap_8 FILLER_73_1622 ();
 sg13g2_decap_8 FILLER_73_1629 ();
 sg13g2_decap_8 FILLER_73_1636 ();
 sg13g2_decap_8 FILLER_73_1643 ();
 sg13g2_decap_8 FILLER_73_1650 ();
 sg13g2_decap_8 FILLER_73_1657 ();
 sg13g2_decap_8 FILLER_73_1664 ();
 sg13g2_decap_8 FILLER_73_1675 ();
 sg13g2_decap_8 FILLER_73_1682 ();
 sg13g2_decap_8 FILLER_73_1689 ();
 sg13g2_fill_2 FILLER_73_1696 ();
 sg13g2_decap_8 FILLER_73_1714 ();
 sg13g2_decap_4 FILLER_73_1721 ();
 sg13g2_decap_8 FILLER_73_1733 ();
 sg13g2_fill_2 FILLER_73_1740 ();
 sg13g2_fill_1 FILLER_73_1742 ();
 sg13g2_decap_8 FILLER_73_1748 ();
 sg13g2_decap_8 FILLER_73_1767 ();
 sg13g2_decap_8 FILLER_73_1774 ();
 sg13g2_decap_8 FILLER_73_1785 ();
 sg13g2_decap_8 FILLER_73_1792 ();
 sg13g2_decap_8 FILLER_73_1799 ();
 sg13g2_decap_8 FILLER_73_1806 ();
 sg13g2_fill_2 FILLER_73_1813 ();
 sg13g2_fill_1 FILLER_73_1815 ();
 sg13g2_fill_2 FILLER_73_1824 ();
 sg13g2_fill_1 FILLER_73_1826 ();
 sg13g2_decap_8 FILLER_73_1847 ();
 sg13g2_decap_8 FILLER_73_1854 ();
 sg13g2_fill_2 FILLER_73_1861 ();
 sg13g2_fill_1 FILLER_73_1863 ();
 sg13g2_decap_8 FILLER_73_1868 ();
 sg13g2_decap_8 FILLER_73_1875 ();
 sg13g2_decap_4 FILLER_73_1882 ();
 sg13g2_fill_1 FILLER_73_1886 ();
 sg13g2_decap_8 FILLER_73_1895 ();
 sg13g2_decap_8 FILLER_73_1902 ();
 sg13g2_fill_2 FILLER_73_1909 ();
 sg13g2_fill_1 FILLER_73_1911 ();
 sg13g2_decap_8 FILLER_73_1916 ();
 sg13g2_decap_8 FILLER_73_1923 ();
 sg13g2_decap_8 FILLER_73_1930 ();
 sg13g2_decap_8 FILLER_73_1937 ();
 sg13g2_fill_2 FILLER_73_1944 ();
 sg13g2_fill_2 FILLER_73_1950 ();
 sg13g2_fill_1 FILLER_73_1952 ();
 sg13g2_decap_8 FILLER_73_1957 ();
 sg13g2_decap_8 FILLER_73_1964 ();
 sg13g2_decap_8 FILLER_73_1971 ();
 sg13g2_fill_2 FILLER_73_1978 ();
 sg13g2_fill_1 FILLER_73_1980 ();
 sg13g2_decap_8 FILLER_73_1989 ();
 sg13g2_decap_8 FILLER_73_1996 ();
 sg13g2_decap_8 FILLER_73_2003 ();
 sg13g2_decap_8 FILLER_73_2010 ();
 sg13g2_decap_8 FILLER_73_2017 ();
 sg13g2_fill_1 FILLER_73_2024 ();
 sg13g2_fill_2 FILLER_73_2035 ();
 sg13g2_decap_8 FILLER_73_2042 ();
 sg13g2_decap_8 FILLER_73_2049 ();
 sg13g2_decap_8 FILLER_73_2056 ();
 sg13g2_decap_8 FILLER_73_2063 ();
 sg13g2_decap_8 FILLER_73_2070 ();
 sg13g2_decap_8 FILLER_73_2077 ();
 sg13g2_decap_8 FILLER_73_2084 ();
 sg13g2_fill_1 FILLER_73_2103 ();
 sg13g2_fill_1 FILLER_73_2110 ();
 sg13g2_fill_1 FILLER_73_2125 ();
 sg13g2_decap_8 FILLER_73_2129 ();
 sg13g2_decap_8 FILLER_73_2136 ();
 sg13g2_fill_1 FILLER_73_2143 ();
 sg13g2_fill_2 FILLER_73_2161 ();
 sg13g2_decap_8 FILLER_73_2193 ();
 sg13g2_decap_4 FILLER_73_2200 ();
 sg13g2_fill_2 FILLER_73_2204 ();
 sg13g2_decap_8 FILLER_73_2209 ();
 sg13g2_fill_1 FILLER_73_2216 ();
 sg13g2_fill_2 FILLER_73_2221 ();
 sg13g2_fill_1 FILLER_73_2223 ();
 sg13g2_fill_1 FILLER_73_2237 ();
 sg13g2_decap_8 FILLER_73_2244 ();
 sg13g2_decap_8 FILLER_73_2251 ();
 sg13g2_fill_2 FILLER_73_2258 ();
 sg13g2_fill_1 FILLER_73_2286 ();
 sg13g2_fill_2 FILLER_73_2317 ();
 sg13g2_fill_2 FILLER_73_2353 ();
 sg13g2_fill_2 FILLER_73_2424 ();
 sg13g2_fill_1 FILLER_73_2460 ();
 sg13g2_fill_1 FILLER_73_2492 ();
 sg13g2_fill_2 FILLER_73_2565 ();
 sg13g2_fill_1 FILLER_73_2593 ();
 sg13g2_decap_8 FILLER_73_2620 ();
 sg13g2_decap_8 FILLER_73_2627 ();
 sg13g2_decap_8 FILLER_73_2634 ();
 sg13g2_decap_8 FILLER_73_2641 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_90 ();
 sg13g2_fill_2 FILLER_74_96 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_fill_1 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_160 ();
 sg13g2_fill_1 FILLER_74_162 ();
 sg13g2_fill_2 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_fill_1 FILLER_74_220 ();
 sg13g2_decap_4 FILLER_74_234 ();
 sg13g2_fill_1 FILLER_74_238 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_decap_8 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_2 FILLER_74_350 ();
 sg13g2_fill_1 FILLER_74_441 ();
 sg13g2_fill_2 FILLER_74_468 ();
 sg13g2_fill_1 FILLER_74_478 ();
 sg13g2_fill_2 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_511 ();
 sg13g2_fill_1 FILLER_74_516 ();
 sg13g2_decap_4 FILLER_74_522 ();
 sg13g2_fill_1 FILLER_74_526 ();
 sg13g2_fill_2 FILLER_74_531 ();
 sg13g2_fill_1 FILLER_74_533 ();
 sg13g2_fill_2 FILLER_74_538 ();
 sg13g2_decap_4 FILLER_74_562 ();
 sg13g2_fill_1 FILLER_74_592 ();
 sg13g2_fill_1 FILLER_74_690 ();
 sg13g2_fill_1 FILLER_74_695 ();
 sg13g2_fill_2 FILLER_74_704 ();
 sg13g2_fill_1 FILLER_74_732 ();
 sg13g2_fill_2 FILLER_74_738 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_fill_2 FILLER_74_792 ();
 sg13g2_fill_1 FILLER_74_799 ();
 sg13g2_fill_2 FILLER_74_805 ();
 sg13g2_fill_2 FILLER_74_812 ();
 sg13g2_fill_2 FILLER_74_818 ();
 sg13g2_fill_1 FILLER_74_885 ();
 sg13g2_fill_1 FILLER_74_903 ();
 sg13g2_fill_2 FILLER_74_917 ();
 sg13g2_fill_1 FILLER_74_1029 ();
 sg13g2_fill_2 FILLER_74_1050 ();
 sg13g2_fill_1 FILLER_74_1052 ();
 sg13g2_fill_2 FILLER_74_1079 ();
 sg13g2_fill_1 FILLER_74_1081 ();
 sg13g2_fill_1 FILLER_74_1110 ();
 sg13g2_decap_4 FILLER_74_1115 ();
 sg13g2_decap_4 FILLER_74_1124 ();
 sg13g2_fill_1 FILLER_74_1173 ();
 sg13g2_fill_2 FILLER_74_1180 ();
 sg13g2_fill_1 FILLER_74_1182 ();
 sg13g2_fill_1 FILLER_74_1197 ();
 sg13g2_fill_1 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1282 ();
 sg13g2_decap_8 FILLER_74_1289 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_4 FILLER_74_1309 ();
 sg13g2_fill_2 FILLER_74_1326 ();
 sg13g2_fill_2 FILLER_74_1334 ();
 sg13g2_fill_1 FILLER_74_1354 ();
 sg13g2_fill_1 FILLER_74_1372 ();
 sg13g2_decap_8 FILLER_74_1404 ();
 sg13g2_decap_8 FILLER_74_1411 ();
 sg13g2_decap_8 FILLER_74_1418 ();
 sg13g2_fill_2 FILLER_74_1425 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_decap_8 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1449 ();
 sg13g2_fill_1 FILLER_74_1456 ();
 sg13g2_fill_1 FILLER_74_1491 ();
 sg13g2_decap_8 FILLER_74_1498 ();
 sg13g2_decap_4 FILLER_74_1505 ();
 sg13g2_fill_1 FILLER_74_1509 ();
 sg13g2_fill_1 FILLER_74_1528 ();
 sg13g2_fill_1 FILLER_74_1533 ();
 sg13g2_fill_2 FILLER_74_1554 ();
 sg13g2_fill_2 FILLER_74_1560 ();
 sg13g2_fill_1 FILLER_74_1562 ();
 sg13g2_fill_2 FILLER_74_1567 ();
 sg13g2_fill_1 FILLER_74_1569 ();
 sg13g2_decap_4 FILLER_74_1575 ();
 sg13g2_fill_2 FILLER_74_1583 ();
 sg13g2_fill_1 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1626 ();
 sg13g2_decap_8 FILLER_74_1633 ();
 sg13g2_decap_8 FILLER_74_1640 ();
 sg13g2_decap_8 FILLER_74_1647 ();
 sg13g2_fill_2 FILLER_74_1654 ();
 sg13g2_fill_1 FILLER_74_1656 ();
 sg13g2_decap_8 FILLER_74_1661 ();
 sg13g2_decap_8 FILLER_74_1668 ();
 sg13g2_decap_8 FILLER_74_1675 ();
 sg13g2_decap_8 FILLER_74_1682 ();
 sg13g2_decap_8 FILLER_74_1689 ();
 sg13g2_decap_8 FILLER_74_1696 ();
 sg13g2_fill_1 FILLER_74_1703 ();
 sg13g2_decap_4 FILLER_74_1710 ();
 sg13g2_fill_1 FILLER_74_1714 ();
 sg13g2_fill_2 FILLER_74_1721 ();
 sg13g2_fill_2 FILLER_74_1736 ();
 sg13g2_fill_2 FILLER_74_1746 ();
 sg13g2_decap_8 FILLER_74_1756 ();
 sg13g2_decap_8 FILLER_74_1763 ();
 sg13g2_decap_8 FILLER_74_1770 ();
 sg13g2_decap_8 FILLER_74_1777 ();
 sg13g2_decap_8 FILLER_74_1784 ();
 sg13g2_decap_8 FILLER_74_1791 ();
 sg13g2_decap_8 FILLER_74_1798 ();
 sg13g2_decap_8 FILLER_74_1829 ();
 sg13g2_decap_8 FILLER_74_1836 ();
 sg13g2_decap_8 FILLER_74_1843 ();
 sg13g2_decap_8 FILLER_74_1850 ();
 sg13g2_decap_8 FILLER_74_1857 ();
 sg13g2_decap_8 FILLER_74_1864 ();
 sg13g2_decap_8 FILLER_74_1871 ();
 sg13g2_decap_8 FILLER_74_1878 ();
 sg13g2_decap_8 FILLER_74_1885 ();
 sg13g2_decap_8 FILLER_74_1892 ();
 sg13g2_decap_8 FILLER_74_1899 ();
 sg13g2_decap_8 FILLER_74_1906 ();
 sg13g2_decap_8 FILLER_74_1913 ();
 sg13g2_decap_8 FILLER_74_1920 ();
 sg13g2_decap_8 FILLER_74_1927 ();
 sg13g2_decap_8 FILLER_74_1934 ();
 sg13g2_decap_8 FILLER_74_1941 ();
 sg13g2_fill_1 FILLER_74_1948 ();
 sg13g2_decap_8 FILLER_74_1954 ();
 sg13g2_decap_8 FILLER_74_1961 ();
 sg13g2_decap_8 FILLER_74_1968 ();
 sg13g2_decap_8 FILLER_74_1975 ();
 sg13g2_decap_8 FILLER_74_1982 ();
 sg13g2_decap_8 FILLER_74_1989 ();
 sg13g2_decap_8 FILLER_74_1996 ();
 sg13g2_decap_8 FILLER_74_2003 ();
 sg13g2_decap_8 FILLER_74_2010 ();
 sg13g2_decap_8 FILLER_74_2017 ();
 sg13g2_decap_8 FILLER_74_2024 ();
 sg13g2_decap_8 FILLER_74_2031 ();
 sg13g2_decap_8 FILLER_74_2038 ();
 sg13g2_decap_8 FILLER_74_2045 ();
 sg13g2_decap_8 FILLER_74_2052 ();
 sg13g2_decap_8 FILLER_74_2059 ();
 sg13g2_decap_8 FILLER_74_2066 ();
 sg13g2_decap_8 FILLER_74_2073 ();
 sg13g2_decap_8 FILLER_74_2080 ();
 sg13g2_decap_8 FILLER_74_2087 ();
 sg13g2_fill_2 FILLER_74_2094 ();
 sg13g2_fill_1 FILLER_74_2096 ();
 sg13g2_decap_4 FILLER_74_2100 ();
 sg13g2_decap_4 FILLER_74_2132 ();
 sg13g2_decap_8 FILLER_74_2172 ();
 sg13g2_fill_1 FILLER_74_2179 ();
 sg13g2_fill_1 FILLER_74_2189 ();
 sg13g2_fill_1 FILLER_74_2196 ();
 sg13g2_decap_4 FILLER_74_2201 ();
 sg13g2_fill_1 FILLER_74_2205 ();
 sg13g2_fill_1 FILLER_74_2246 ();
 sg13g2_fill_1 FILLER_74_2256 ();
 sg13g2_fill_1 FILLER_74_2398 ();
 sg13g2_fill_2 FILLER_74_2409 ();
 sg13g2_fill_2 FILLER_74_2416 ();
 sg13g2_fill_2 FILLER_74_2422 ();
 sg13g2_fill_2 FILLER_74_2432 ();
 sg13g2_fill_2 FILLER_74_2469 ();
 sg13g2_fill_1 FILLER_74_2496 ();
 sg13g2_decap_8 FILLER_74_2614 ();
 sg13g2_decap_8 FILLER_74_2621 ();
 sg13g2_decap_8 FILLER_74_2628 ();
 sg13g2_decap_8 FILLER_74_2635 ();
 sg13g2_decap_8 FILLER_74_2642 ();
 sg13g2_decap_8 FILLER_74_2649 ();
 sg13g2_decap_8 FILLER_74_2656 ();
 sg13g2_decap_8 FILLER_74_2663 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_4 ();
 sg13g2_decap_8 FILLER_75_48 ();
 sg13g2_decap_4 FILLER_75_55 ();
 sg13g2_fill_1 FILLER_75_59 ();
 sg13g2_decap_4 FILLER_75_64 ();
 sg13g2_fill_1 FILLER_75_73 ();
 sg13g2_decap_4 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_104 ();
 sg13g2_decap_8 FILLER_75_111 ();
 sg13g2_decap_8 FILLER_75_118 ();
 sg13g2_fill_2 FILLER_75_125 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_1 FILLER_75_139 ();
 sg13g2_decap_4 FILLER_75_158 ();
 sg13g2_fill_1 FILLER_75_162 ();
 sg13g2_decap_4 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_230 ();
 sg13g2_decap_4 FILLER_75_242 ();
 sg13g2_fill_1 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_decap_4 FILLER_75_312 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_2 FILLER_75_409 ();
 sg13g2_fill_1 FILLER_75_460 ();
 sg13g2_fill_1 FILLER_75_468 ();
 sg13g2_fill_2 FILLER_75_478 ();
 sg13g2_fill_1 FILLER_75_485 ();
 sg13g2_fill_1 FILLER_75_491 ();
 sg13g2_fill_2 FILLER_75_496 ();
 sg13g2_fill_2 FILLER_75_503 ();
 sg13g2_decap_4 FILLER_75_510 ();
 sg13g2_fill_1 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_530 ();
 sg13g2_fill_2 FILLER_75_540 ();
 sg13g2_fill_1 FILLER_75_542 ();
 sg13g2_decap_8 FILLER_75_548 ();
 sg13g2_decap_8 FILLER_75_555 ();
 sg13g2_fill_2 FILLER_75_562 ();
 sg13g2_fill_1 FILLER_75_568 ();
 sg13g2_fill_2 FILLER_75_574 ();
 sg13g2_fill_1 FILLER_75_576 ();
 sg13g2_decap_4 FILLER_75_585 ();
 sg13g2_fill_2 FILLER_75_593 ();
 sg13g2_fill_1 FILLER_75_595 ();
 sg13g2_fill_1 FILLER_75_612 ();
 sg13g2_fill_1 FILLER_75_617 ();
 sg13g2_fill_1 FILLER_75_627 ();
 sg13g2_fill_2 FILLER_75_658 ();
 sg13g2_fill_2 FILLER_75_700 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_fill_1 FILLER_75_708 ();
 sg13g2_fill_2 FILLER_75_735 ();
 sg13g2_fill_1 FILLER_75_781 ();
 sg13g2_fill_1 FILLER_75_867 ();
 sg13g2_fill_2 FILLER_75_880 ();
 sg13g2_fill_1 FILLER_75_886 ();
 sg13g2_fill_2 FILLER_75_922 ();
 sg13g2_fill_1 FILLER_75_924 ();
 sg13g2_fill_2 FILLER_75_977 ();
 sg13g2_fill_1 FILLER_75_1034 ();
 sg13g2_fill_1 FILLER_75_1047 ();
 sg13g2_fill_1 FILLER_75_1054 ();
 sg13g2_fill_1 FILLER_75_1085 ();
 sg13g2_decap_8 FILLER_75_1112 ();
 sg13g2_fill_2 FILLER_75_1119 ();
 sg13g2_fill_1 FILLER_75_1121 ();
 sg13g2_fill_2 FILLER_75_1130 ();
 sg13g2_fill_1 FILLER_75_1137 ();
 sg13g2_fill_2 FILLER_75_1142 ();
 sg13g2_fill_1 FILLER_75_1144 ();
 sg13g2_fill_2 FILLER_75_1155 ();
 sg13g2_fill_1 FILLER_75_1157 ();
 sg13g2_fill_1 FILLER_75_1194 ();
 sg13g2_fill_1 FILLER_75_1251 ();
 sg13g2_decap_4 FILLER_75_1278 ();
 sg13g2_fill_2 FILLER_75_1285 ();
 sg13g2_decap_8 FILLER_75_1304 ();
 sg13g2_decap_8 FILLER_75_1311 ();
 sg13g2_decap_8 FILLER_75_1318 ();
 sg13g2_fill_2 FILLER_75_1325 ();
 sg13g2_fill_1 FILLER_75_1332 ();
 sg13g2_fill_2 FILLER_75_1356 ();
 sg13g2_fill_2 FILLER_75_1374 ();
 sg13g2_fill_1 FILLER_75_1382 ();
 sg13g2_decap_8 FILLER_75_1408 ();
 sg13g2_fill_2 FILLER_75_1415 ();
 sg13g2_decap_4 FILLER_75_1426 ();
 sg13g2_fill_2 FILLER_75_1439 ();
 sg13g2_fill_1 FILLER_75_1441 ();
 sg13g2_decap_8 FILLER_75_1447 ();
 sg13g2_decap_8 FILLER_75_1454 ();
 sg13g2_fill_1 FILLER_75_1466 ();
 sg13g2_fill_1 FILLER_75_1473 ();
 sg13g2_fill_1 FILLER_75_1478 ();
 sg13g2_decap_4 FILLER_75_1483 ();
 sg13g2_fill_1 FILLER_75_1487 ();
 sg13g2_decap_4 FILLER_75_1491 ();
 sg13g2_fill_1 FILLER_75_1495 ();
 sg13g2_fill_2 FILLER_75_1504 ();
 sg13g2_fill_1 FILLER_75_1506 ();
 sg13g2_fill_2 FILLER_75_1516 ();
 sg13g2_fill_1 FILLER_75_1524 ();
 sg13g2_fill_1 FILLER_75_1530 ();
 sg13g2_fill_2 FILLER_75_1535 ();
 sg13g2_fill_1 FILLER_75_1541 ();
 sg13g2_fill_1 FILLER_75_1552 ();
 sg13g2_decap_8 FILLER_75_1557 ();
 sg13g2_fill_1 FILLER_75_1564 ();
 sg13g2_fill_2 FILLER_75_1570 ();
 sg13g2_fill_2 FILLER_75_1591 ();
 sg13g2_decap_4 FILLER_75_1601 ();
 sg13g2_fill_2 FILLER_75_1605 ();
 sg13g2_decap_8 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1618 ();
 sg13g2_decap_8 FILLER_75_1625 ();
 sg13g2_decap_8 FILLER_75_1632 ();
 sg13g2_decap_8 FILLER_75_1639 ();
 sg13g2_decap_4 FILLER_75_1646 ();
 sg13g2_fill_2 FILLER_75_1650 ();
 sg13g2_decap_8 FILLER_75_1657 ();
 sg13g2_decap_8 FILLER_75_1664 ();
 sg13g2_decap_8 FILLER_75_1671 ();
 sg13g2_decap_8 FILLER_75_1678 ();
 sg13g2_decap_8 FILLER_75_1685 ();
 sg13g2_decap_8 FILLER_75_1692 ();
 sg13g2_decap_8 FILLER_75_1699 ();
 sg13g2_decap_8 FILLER_75_1706 ();
 sg13g2_fill_1 FILLER_75_1713 ();
 sg13g2_decap_8 FILLER_75_1719 ();
 sg13g2_decap_8 FILLER_75_1726 ();
 sg13g2_decap_8 FILLER_75_1733 ();
 sg13g2_decap_8 FILLER_75_1740 ();
 sg13g2_decap_8 FILLER_75_1747 ();
 sg13g2_decap_8 FILLER_75_1754 ();
 sg13g2_decap_8 FILLER_75_1761 ();
 sg13g2_decap_8 FILLER_75_1768 ();
 sg13g2_decap_8 FILLER_75_1775 ();
 sg13g2_decap_8 FILLER_75_1782 ();
 sg13g2_decap_8 FILLER_75_1789 ();
 sg13g2_decap_8 FILLER_75_1796 ();
 sg13g2_decap_8 FILLER_75_1807 ();
 sg13g2_fill_2 FILLER_75_1814 ();
 sg13g2_fill_1 FILLER_75_1816 ();
 sg13g2_decap_8 FILLER_75_1827 ();
 sg13g2_decap_4 FILLER_75_1834 ();
 sg13g2_decap_8 FILLER_75_1847 ();
 sg13g2_decap_8 FILLER_75_1854 ();
 sg13g2_decap_8 FILLER_75_1861 ();
 sg13g2_decap_8 FILLER_75_1868 ();
 sg13g2_decap_8 FILLER_75_1875 ();
 sg13g2_decap_8 FILLER_75_1882 ();
 sg13g2_decap_8 FILLER_75_1889 ();
 sg13g2_decap_8 FILLER_75_1896 ();
 sg13g2_decap_8 FILLER_75_1903 ();
 sg13g2_decap_8 FILLER_75_1910 ();
 sg13g2_decap_8 FILLER_75_1917 ();
 sg13g2_decap_8 FILLER_75_1924 ();
 sg13g2_decap_8 FILLER_75_1931 ();
 sg13g2_decap_8 FILLER_75_1938 ();
 sg13g2_fill_2 FILLER_75_1945 ();
 sg13g2_fill_1 FILLER_75_1947 ();
 sg13g2_decap_8 FILLER_75_1953 ();
 sg13g2_decap_8 FILLER_75_1960 ();
 sg13g2_decap_8 FILLER_75_1967 ();
 sg13g2_decap_8 FILLER_75_1974 ();
 sg13g2_decap_8 FILLER_75_1981 ();
 sg13g2_decap_8 FILLER_75_1988 ();
 sg13g2_decap_8 FILLER_75_1995 ();
 sg13g2_decap_8 FILLER_75_2002 ();
 sg13g2_decap_4 FILLER_75_2009 ();
 sg13g2_fill_2 FILLER_75_2019 ();
 sg13g2_decap_8 FILLER_75_2027 ();
 sg13g2_decap_8 FILLER_75_2034 ();
 sg13g2_decap_8 FILLER_75_2041 ();
 sg13g2_decap_8 FILLER_75_2048 ();
 sg13g2_decap_8 FILLER_75_2055 ();
 sg13g2_decap_8 FILLER_75_2062 ();
 sg13g2_decap_8 FILLER_75_2069 ();
 sg13g2_decap_8 FILLER_75_2076 ();
 sg13g2_decap_8 FILLER_75_2083 ();
 sg13g2_decap_8 FILLER_75_2090 ();
 sg13g2_decap_4 FILLER_75_2097 ();
 sg13g2_fill_1 FILLER_75_2101 ();
 sg13g2_decap_4 FILLER_75_2148 ();
 sg13g2_fill_2 FILLER_75_2152 ();
 sg13g2_fill_2 FILLER_75_2160 ();
 sg13g2_fill_1 FILLER_75_2162 ();
 sg13g2_decap_8 FILLER_75_2169 ();
 sg13g2_fill_1 FILLER_75_2176 ();
 sg13g2_fill_1 FILLER_75_2182 ();
 sg13g2_fill_2 FILLER_75_2187 ();
 sg13g2_fill_2 FILLER_75_2223 ();
 sg13g2_fill_1 FILLER_75_2269 ();
 sg13g2_fill_1 FILLER_75_2283 ();
 sg13g2_fill_1 FILLER_75_2366 ();
 sg13g2_fill_1 FILLER_75_2408 ();
 sg13g2_fill_1 FILLER_75_2418 ();
 sg13g2_fill_1 FILLER_75_2429 ();
 sg13g2_fill_2 FILLER_75_2438 ();
 sg13g2_fill_1 FILLER_75_2449 ();
 sg13g2_fill_1 FILLER_75_2454 ();
 sg13g2_fill_1 FILLER_75_2501 ();
 sg13g2_fill_1 FILLER_75_2525 ();
 sg13g2_decap_8 FILLER_75_2610 ();
 sg13g2_decap_8 FILLER_75_2617 ();
 sg13g2_decap_8 FILLER_75_2624 ();
 sg13g2_decap_8 FILLER_75_2631 ();
 sg13g2_decap_8 FILLER_75_2638 ();
 sg13g2_decap_8 FILLER_75_2645 ();
 sg13g2_decap_8 FILLER_75_2652 ();
 sg13g2_decap_8 FILLER_75_2659 ();
 sg13g2_decap_4 FILLER_75_2666 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_decap_4 FILLER_76_66 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_fill_2 FILLER_76_76 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_decap_8 FILLER_76_110 ();
 sg13g2_fill_2 FILLER_76_117 ();
 sg13g2_decap_4 FILLER_76_122 ();
 sg13g2_fill_1 FILLER_76_126 ();
 sg13g2_fill_2 FILLER_76_190 ();
 sg13g2_decap_8 FILLER_76_237 ();
 sg13g2_decap_8 FILLER_76_244 ();
 sg13g2_decap_8 FILLER_76_251 ();
 sg13g2_fill_1 FILLER_76_313 ();
 sg13g2_fill_2 FILLER_76_324 ();
 sg13g2_fill_1 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_342 ();
 sg13g2_fill_2 FILLER_76_401 ();
 sg13g2_fill_2 FILLER_76_445 ();
 sg13g2_fill_1 FILLER_76_455 ();
 sg13g2_fill_1 FILLER_76_461 ();
 sg13g2_fill_2 FILLER_76_484 ();
 sg13g2_decap_4 FILLER_76_491 ();
 sg13g2_fill_2 FILLER_76_495 ();
 sg13g2_fill_1 FILLER_76_502 ();
 sg13g2_fill_2 FILLER_76_535 ();
 sg13g2_fill_1 FILLER_76_537 ();
 sg13g2_fill_2 FILLER_76_543 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_fill_1 FILLER_76_553 ();
 sg13g2_decap_4 FILLER_76_563 ();
 sg13g2_fill_2 FILLER_76_586 ();
 sg13g2_decap_4 FILLER_76_598 ();
 sg13g2_fill_2 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_612 ();
 sg13g2_fill_1 FILLER_76_619 ();
 sg13g2_fill_1 FILLER_76_630 ();
 sg13g2_fill_1 FILLER_76_651 ();
 sg13g2_fill_1 FILLER_76_657 ();
 sg13g2_fill_2 FILLER_76_689 ();
 sg13g2_fill_2 FILLER_76_696 ();
 sg13g2_fill_2 FILLER_76_729 ();
 sg13g2_fill_2 FILLER_76_770 ();
 sg13g2_fill_2 FILLER_76_796 ();
 sg13g2_fill_2 FILLER_76_838 ();
 sg13g2_fill_1 FILLER_76_844 ();
 sg13g2_fill_2 FILLER_76_871 ();
 sg13g2_fill_1 FILLER_76_911 ();
 sg13g2_fill_1 FILLER_76_917 ();
 sg13g2_fill_1 FILLER_76_959 ();
 sg13g2_fill_1 FILLER_76_1040 ();
 sg13g2_fill_2 FILLER_76_1091 ();
 sg13g2_fill_1 FILLER_76_1141 ();
 sg13g2_fill_2 FILLER_76_1152 ();
 sg13g2_fill_1 FILLER_76_1158 ();
 sg13g2_decap_8 FILLER_76_1195 ();
 sg13g2_fill_2 FILLER_76_1202 ();
 sg13g2_fill_1 FILLER_76_1204 ();
 sg13g2_fill_1 FILLER_76_1209 ();
 sg13g2_fill_1 FILLER_76_1216 ();
 sg13g2_fill_2 FILLER_76_1254 ();
 sg13g2_fill_2 FILLER_76_1270 ();
 sg13g2_fill_1 FILLER_76_1272 ();
 sg13g2_fill_2 FILLER_76_1312 ();
 sg13g2_fill_1 FILLER_76_1314 ();
 sg13g2_fill_2 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1323 ();
 sg13g2_decap_8 FILLER_76_1330 ();
 sg13g2_decap_4 FILLER_76_1337 ();
 sg13g2_fill_1 FILLER_76_1369 ();
 sg13g2_fill_2 FILLER_76_1374 ();
 sg13g2_fill_1 FILLER_76_1411 ();
 sg13g2_fill_1 FILLER_76_1426 ();
 sg13g2_fill_2 FILLER_76_1432 ();
 sg13g2_fill_1 FILLER_76_1461 ();
 sg13g2_fill_1 FILLER_76_1479 ();
 sg13g2_fill_2 FILLER_76_1545 ();
 sg13g2_fill_1 FILLER_76_1552 ();
 sg13g2_decap_8 FILLER_76_1603 ();
 sg13g2_decap_8 FILLER_76_1610 ();
 sg13g2_decap_8 FILLER_76_1617 ();
 sg13g2_decap_8 FILLER_76_1624 ();
 sg13g2_decap_8 FILLER_76_1631 ();
 sg13g2_decap_8 FILLER_76_1638 ();
 sg13g2_fill_2 FILLER_76_1645 ();
 sg13g2_decap_8 FILLER_76_1651 ();
 sg13g2_decap_8 FILLER_76_1658 ();
 sg13g2_fill_2 FILLER_76_1674 ();
 sg13g2_decap_8 FILLER_76_1682 ();
 sg13g2_decap_8 FILLER_76_1689 ();
 sg13g2_decap_8 FILLER_76_1696 ();
 sg13g2_decap_8 FILLER_76_1703 ();
 sg13g2_decap_8 FILLER_76_1710 ();
 sg13g2_decap_4 FILLER_76_1717 ();
 sg13g2_fill_2 FILLER_76_1721 ();
 sg13g2_fill_1 FILLER_76_1727 ();
 sg13g2_fill_1 FILLER_76_1733 ();
 sg13g2_fill_2 FILLER_76_1742 ();
 sg13g2_fill_1 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1753 ();
 sg13g2_decap_8 FILLER_76_1765 ();
 sg13g2_decap_4 FILLER_76_1772 ();
 sg13g2_fill_1 FILLER_76_1776 ();
 sg13g2_decap_8 FILLER_76_1782 ();
 sg13g2_decap_8 FILLER_76_1789 ();
 sg13g2_fill_2 FILLER_76_1796 ();
 sg13g2_fill_2 FILLER_76_1803 ();
 sg13g2_fill_1 FILLER_76_1805 ();
 sg13g2_fill_2 FILLER_76_1815 ();
 sg13g2_decap_4 FILLER_76_1822 ();
 sg13g2_fill_2 FILLER_76_1826 ();
 sg13g2_decap_8 FILLER_76_1832 ();
 sg13g2_decap_8 FILLER_76_1839 ();
 sg13g2_decap_8 FILLER_76_1846 ();
 sg13g2_decap_8 FILLER_76_1853 ();
 sg13g2_decap_8 FILLER_76_1860 ();
 sg13g2_decap_8 FILLER_76_1867 ();
 sg13g2_decap_8 FILLER_76_1874 ();
 sg13g2_decap_8 FILLER_76_1881 ();
 sg13g2_decap_8 FILLER_76_1904 ();
 sg13g2_decap_8 FILLER_76_1911 ();
 sg13g2_decap_8 FILLER_76_1918 ();
 sg13g2_decap_8 FILLER_76_1925 ();
 sg13g2_decap_8 FILLER_76_1932 ();
 sg13g2_decap_8 FILLER_76_1950 ();
 sg13g2_decap_8 FILLER_76_1957 ();
 sg13g2_decap_8 FILLER_76_1964 ();
 sg13g2_decap_4 FILLER_76_1971 ();
 sg13g2_fill_2 FILLER_76_1975 ();
 sg13g2_fill_1 FILLER_76_1982 ();
 sg13g2_decap_8 FILLER_76_1993 ();
 sg13g2_decap_8 FILLER_76_2000 ();
 sg13g2_decap_8 FILLER_76_2007 ();
 sg13g2_decap_8 FILLER_76_2020 ();
 sg13g2_decap_8 FILLER_76_2027 ();
 sg13g2_decap_8 FILLER_76_2034 ();
 sg13g2_decap_8 FILLER_76_2041 ();
 sg13g2_decap_8 FILLER_76_2048 ();
 sg13g2_decap_8 FILLER_76_2055 ();
 sg13g2_decap_8 FILLER_76_2062 ();
 sg13g2_decap_8 FILLER_76_2069 ();
 sg13g2_decap_8 FILLER_76_2076 ();
 sg13g2_fill_2 FILLER_76_2083 ();
 sg13g2_fill_2 FILLER_76_2145 ();
 sg13g2_decap_4 FILLER_76_2173 ();
 sg13g2_fill_2 FILLER_76_2203 ();
 sg13g2_fill_2 FILLER_76_2210 ();
 sg13g2_fill_1 FILLER_76_2212 ();
 sg13g2_fill_1 FILLER_76_2217 ();
 sg13g2_fill_1 FILLER_76_2222 ();
 sg13g2_fill_1 FILLER_76_2228 ();
 sg13g2_fill_2 FILLER_76_2242 ();
 sg13g2_fill_1 FILLER_76_2291 ();
 sg13g2_fill_1 FILLER_76_2296 ();
 sg13g2_fill_1 FILLER_76_2393 ();
 sg13g2_fill_1 FILLER_76_2418 ();
 sg13g2_fill_1 FILLER_76_2461 ();
 sg13g2_fill_1 FILLER_76_2476 ();
 sg13g2_fill_2 FILLER_76_2487 ();
 sg13g2_fill_1 FILLER_76_2521 ();
 sg13g2_decap_8 FILLER_76_2604 ();
 sg13g2_decap_8 FILLER_76_2611 ();
 sg13g2_decap_8 FILLER_76_2618 ();
 sg13g2_decap_8 FILLER_76_2625 ();
 sg13g2_decap_8 FILLER_76_2632 ();
 sg13g2_decap_8 FILLER_76_2639 ();
 sg13g2_decap_8 FILLER_76_2646 ();
 sg13g2_decap_8 FILLER_76_2653 ();
 sg13g2_decap_8 FILLER_76_2660 ();
 sg13g2_fill_2 FILLER_76_2667 ();
 sg13g2_fill_1 FILLER_76_2669 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_4 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_25 ();
 sg13g2_fill_2 FILLER_77_100 ();
 sg13g2_fill_1 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_fill_1 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_167 ();
 sg13g2_decap_8 FILLER_77_174 ();
 sg13g2_decap_4 FILLER_77_181 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_2 FILLER_77_235 ();
 sg13g2_decap_4 FILLER_77_303 ();
 sg13g2_decap_4 FILLER_77_312 ();
 sg13g2_fill_1 FILLER_77_316 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_fill_2 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_fill_2 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_421 ();
 sg13g2_fill_1 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_468 ();
 sg13g2_fill_1 FILLER_77_496 ();
 sg13g2_fill_1 FILLER_77_574 ();
 sg13g2_decap_4 FILLER_77_595 ();
 sg13g2_fill_1 FILLER_77_599 ();
 sg13g2_fill_2 FILLER_77_604 ();
 sg13g2_fill_1 FILLER_77_622 ();
 sg13g2_fill_1 FILLER_77_636 ();
 sg13g2_fill_2 FILLER_77_651 ();
 sg13g2_fill_2 FILLER_77_659 ();
 sg13g2_fill_2 FILLER_77_667 ();
 sg13g2_fill_2 FILLER_77_673 ();
 sg13g2_fill_1 FILLER_77_675 ();
 sg13g2_fill_1 FILLER_77_681 ();
 sg13g2_fill_1 FILLER_77_716 ();
 sg13g2_fill_2 FILLER_77_815 ();
 sg13g2_fill_2 FILLER_77_910 ();
 sg13g2_fill_1 FILLER_77_912 ();
 sg13g2_fill_2 FILLER_77_934 ();
 sg13g2_fill_1 FILLER_77_936 ();
 sg13g2_fill_2 FILLER_77_963 ();
 sg13g2_fill_2 FILLER_77_970 ();
 sg13g2_fill_2 FILLER_77_1005 ();
 sg13g2_fill_1 FILLER_77_1071 ();
 sg13g2_fill_1 FILLER_77_1082 ();
 sg13g2_fill_1 FILLER_77_1109 ();
 sg13g2_fill_1 FILLER_77_1116 ();
 sg13g2_fill_1 FILLER_77_1121 ();
 sg13g2_fill_2 FILLER_77_1132 ();
 sg13g2_decap_4 FILLER_77_1140 ();
 sg13g2_fill_2 FILLER_77_1144 ();
 sg13g2_fill_1 FILLER_77_1180 ();
 sg13g2_fill_2 FILLER_77_1187 ();
 sg13g2_fill_1 FILLER_77_1189 ();
 sg13g2_fill_1 FILLER_77_1222 ();
 sg13g2_fill_1 FILLER_77_1242 ();
 sg13g2_fill_2 FILLER_77_1249 ();
 sg13g2_fill_1 FILLER_77_1292 ();
 sg13g2_fill_1 FILLER_77_1300 ();
 sg13g2_decap_8 FILLER_77_1339 ();
 sg13g2_decap_4 FILLER_77_1346 ();
 sg13g2_fill_1 FILLER_77_1350 ();
 sg13g2_fill_2 FILLER_77_1381 ();
 sg13g2_fill_1 FILLER_77_1383 ();
 sg13g2_fill_1 FILLER_77_1400 ();
 sg13g2_fill_2 FILLER_77_1432 ();
 sg13g2_fill_1 FILLER_77_1434 ();
 sg13g2_fill_2 FILLER_77_1445 ();
 sg13g2_fill_1 FILLER_77_1469 ();
 sg13g2_decap_4 FILLER_77_1477 ();
 sg13g2_fill_1 FILLER_77_1500 ();
 sg13g2_fill_1 FILLER_77_1504 ();
 sg13g2_decap_8 FILLER_77_1510 ();
 sg13g2_decap_4 FILLER_77_1517 ();
 sg13g2_fill_1 FILLER_77_1521 ();
 sg13g2_fill_2 FILLER_77_1556 ();
 sg13g2_fill_1 FILLER_77_1558 ();
 sg13g2_fill_2 FILLER_77_1564 ();
 sg13g2_fill_1 FILLER_77_1566 ();
 sg13g2_fill_1 FILLER_77_1574 ();
 sg13g2_fill_1 FILLER_77_1609 ();
 sg13g2_decap_8 FILLER_77_1615 ();
 sg13g2_decap_8 FILLER_77_1622 ();
 sg13g2_decap_8 FILLER_77_1629 ();
 sg13g2_decap_8 FILLER_77_1636 ();
 sg13g2_fill_1 FILLER_77_1643 ();
 sg13g2_decap_8 FILLER_77_1653 ();
 sg13g2_decap_8 FILLER_77_1660 ();
 sg13g2_decap_4 FILLER_77_1667 ();
 sg13g2_fill_2 FILLER_77_1671 ();
 sg13g2_decap_8 FILLER_77_1679 ();
 sg13g2_fill_2 FILLER_77_1686 ();
 sg13g2_fill_1 FILLER_77_1688 ();
 sg13g2_decap_8 FILLER_77_1701 ();
 sg13g2_decap_8 FILLER_77_1708 ();
 sg13g2_decap_8 FILLER_77_1715 ();
 sg13g2_decap_4 FILLER_77_1731 ();
 sg13g2_fill_1 FILLER_77_1735 ();
 sg13g2_decap_8 FILLER_77_1748 ();
 sg13g2_decap_8 FILLER_77_1755 ();
 sg13g2_fill_1 FILLER_77_1762 ();
 sg13g2_fill_1 FILLER_77_1773 ();
 sg13g2_decap_4 FILLER_77_1792 ();
 sg13g2_decap_4 FILLER_77_1800 ();
 sg13g2_fill_2 FILLER_77_1804 ();
 sg13g2_decap_8 FILLER_77_1837 ();
 sg13g2_decap_8 FILLER_77_1844 ();
 sg13g2_decap_8 FILLER_77_1851 ();
 sg13g2_decap_8 FILLER_77_1858 ();
 sg13g2_decap_8 FILLER_77_1865 ();
 sg13g2_fill_2 FILLER_77_1872 ();
 sg13g2_decap_4 FILLER_77_1878 ();
 sg13g2_fill_2 FILLER_77_1882 ();
 sg13g2_decap_8 FILLER_77_1892 ();
 sg13g2_decap_8 FILLER_77_1899 ();
 sg13g2_fill_1 FILLER_77_1906 ();
 sg13g2_decap_8 FILLER_77_1910 ();
 sg13g2_decap_8 FILLER_77_1917 ();
 sg13g2_decap_8 FILLER_77_1924 ();
 sg13g2_fill_2 FILLER_77_1931 ();
 sg13g2_fill_1 FILLER_77_1933 ();
 sg13g2_fill_2 FILLER_77_1955 ();
 sg13g2_decap_8 FILLER_77_1961 ();
 sg13g2_decap_8 FILLER_77_1968 ();
 sg13g2_decap_8 FILLER_77_1975 ();
 sg13g2_decap_8 FILLER_77_1982 ();
 sg13g2_decap_4 FILLER_77_1989 ();
 sg13g2_fill_1 FILLER_77_1993 ();
 sg13g2_decap_4 FILLER_77_2000 ();
 sg13g2_fill_1 FILLER_77_2004 ();
 sg13g2_decap_8 FILLER_77_2010 ();
 sg13g2_fill_2 FILLER_77_2017 ();
 sg13g2_fill_1 FILLER_77_2019 ();
 sg13g2_decap_8 FILLER_77_2032 ();
 sg13g2_decap_8 FILLER_77_2039 ();
 sg13g2_decap_8 FILLER_77_2046 ();
 sg13g2_decap_8 FILLER_77_2053 ();
 sg13g2_decap_8 FILLER_77_2060 ();
 sg13g2_decap_8 FILLER_77_2067 ();
 sg13g2_decap_8 FILLER_77_2074 ();
 sg13g2_decap_4 FILLER_77_2081 ();
 sg13g2_fill_2 FILLER_77_2085 ();
 sg13g2_decap_8 FILLER_77_2097 ();
 sg13g2_fill_2 FILLER_77_2104 ();
 sg13g2_decap_4 FILLER_77_2176 ();
 sg13g2_fill_1 FILLER_77_2180 ();
 sg13g2_fill_2 FILLER_77_2223 ();
 sg13g2_fill_1 FILLER_77_2256 ();
 sg13g2_fill_1 FILLER_77_2322 ();
 sg13g2_fill_1 FILLER_77_2389 ();
 sg13g2_fill_2 FILLER_77_2398 ();
 sg13g2_fill_1 FILLER_77_2408 ();
 sg13g2_fill_2 FILLER_77_2442 ();
 sg13g2_fill_2 FILLER_77_2515 ();
 sg13g2_fill_1 FILLER_77_2553 ();
 sg13g2_decap_8 FILLER_77_2595 ();
 sg13g2_decap_8 FILLER_77_2602 ();
 sg13g2_decap_8 FILLER_77_2609 ();
 sg13g2_decap_8 FILLER_77_2616 ();
 sg13g2_decap_8 FILLER_77_2623 ();
 sg13g2_decap_8 FILLER_77_2630 ();
 sg13g2_decap_8 FILLER_77_2637 ();
 sg13g2_decap_8 FILLER_77_2644 ();
 sg13g2_decap_8 FILLER_77_2651 ();
 sg13g2_decap_8 FILLER_77_2658 ();
 sg13g2_decap_4 FILLER_77_2665 ();
 sg13g2_fill_1 FILLER_77_2669 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_4 FILLER_78_18 ();
 sg13g2_fill_1 FILLER_78_53 ();
 sg13g2_fill_2 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_82 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_fill_2 FILLER_78_187 ();
 sg13g2_fill_2 FILLER_78_236 ();
 sg13g2_fill_2 FILLER_78_310 ();
 sg13g2_fill_1 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_decap_4 FILLER_78_356 ();
 sg13g2_fill_1 FILLER_78_360 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_fill_1 FILLER_78_567 ();
 sg13g2_fill_2 FILLER_78_607 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_fill_1 FILLER_78_682 ();
 sg13g2_fill_2 FILLER_78_709 ();
 sg13g2_fill_1 FILLER_78_711 ();
 sg13g2_fill_1 FILLER_78_726 ();
 sg13g2_fill_1 FILLER_78_732 ();
 sg13g2_fill_1 FILLER_78_795 ();
 sg13g2_fill_1 FILLER_78_840 ();
 sg13g2_fill_1 FILLER_78_847 ();
 sg13g2_fill_1 FILLER_78_858 ();
 sg13g2_fill_2 FILLER_78_869 ();
 sg13g2_decap_4 FILLER_78_905 ();
 sg13g2_fill_1 FILLER_78_933 ();
 sg13g2_fill_2 FILLER_78_964 ();
 sg13g2_decap_8 FILLER_78_1018 ();
 sg13g2_fill_1 FILLER_78_1025 ();
 sg13g2_decap_8 FILLER_78_1040 ();
 sg13g2_fill_1 FILLER_78_1047 ();
 sg13g2_fill_1 FILLER_78_1074 ();
 sg13g2_fill_1 FILLER_78_1101 ();
 sg13g2_fill_1 FILLER_78_1112 ();
 sg13g2_fill_1 FILLER_78_1123 ();
 sg13g2_decap_8 FILLER_78_1186 ();
 sg13g2_fill_1 FILLER_78_1193 ();
 sg13g2_fill_2 FILLER_78_1198 ();
 sg13g2_fill_1 FILLER_78_1236 ();
 sg13g2_fill_2 FILLER_78_1318 ();
 sg13g2_fill_2 FILLER_78_1357 ();
 sg13g2_fill_2 FILLER_78_1364 ();
 sg13g2_fill_2 FILLER_78_1371 ();
 sg13g2_fill_1 FILLER_78_1373 ();
 sg13g2_fill_2 FILLER_78_1379 ();
 sg13g2_fill_1 FILLER_78_1393 ();
 sg13g2_fill_2 FILLER_78_1420 ();
 sg13g2_fill_2 FILLER_78_1427 ();
 sg13g2_decap_8 FILLER_78_1488 ();
 sg13g2_fill_1 FILLER_78_1495 ();
 sg13g2_fill_1 FILLER_78_1513 ();
 sg13g2_decap_4 FILLER_78_1549 ();
 sg13g2_fill_1 FILLER_78_1563 ();
 sg13g2_fill_1 FILLER_78_1574 ();
 sg13g2_fill_1 FILLER_78_1592 ();
 sg13g2_decap_8 FILLER_78_1616 ();
 sg13g2_decap_8 FILLER_78_1623 ();
 sg13g2_decap_8 FILLER_78_1630 ();
 sg13g2_decap_8 FILLER_78_1637 ();
 sg13g2_decap_8 FILLER_78_1644 ();
 sg13g2_decap_8 FILLER_78_1651 ();
 sg13g2_decap_8 FILLER_78_1658 ();
 sg13g2_decap_8 FILLER_78_1665 ();
 sg13g2_decap_8 FILLER_78_1672 ();
 sg13g2_decap_8 FILLER_78_1679 ();
 sg13g2_decap_8 FILLER_78_1686 ();
 sg13g2_decap_8 FILLER_78_1693 ();
 sg13g2_decap_8 FILLER_78_1700 ();
 sg13g2_decap_8 FILLER_78_1707 ();
 sg13g2_decap_8 FILLER_78_1714 ();
 sg13g2_fill_1 FILLER_78_1721 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_8 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1754 ();
 sg13g2_decap_8 FILLER_78_1761 ();
 sg13g2_decap_8 FILLER_78_1768 ();
 sg13g2_decap_8 FILLER_78_1775 ();
 sg13g2_decap_8 FILLER_78_1782 ();
 sg13g2_decap_8 FILLER_78_1789 ();
 sg13g2_decap_8 FILLER_78_1796 ();
 sg13g2_decap_8 FILLER_78_1803 ();
 sg13g2_decap_8 FILLER_78_1810 ();
 sg13g2_decap_8 FILLER_78_1817 ();
 sg13g2_decap_8 FILLER_78_1824 ();
 sg13g2_decap_8 FILLER_78_1831 ();
 sg13g2_decap_8 FILLER_78_1838 ();
 sg13g2_decap_8 FILLER_78_1845 ();
 sg13g2_decap_8 FILLER_78_1852 ();
 sg13g2_decap_8 FILLER_78_1859 ();
 sg13g2_fill_2 FILLER_78_1866 ();
 sg13g2_decap_8 FILLER_78_1872 ();
 sg13g2_decap_8 FILLER_78_1879 ();
 sg13g2_decap_8 FILLER_78_1886 ();
 sg13g2_decap_8 FILLER_78_1893 ();
 sg13g2_decap_8 FILLER_78_1900 ();
 sg13g2_decap_8 FILLER_78_1907 ();
 sg13g2_decap_8 FILLER_78_1914 ();
 sg13g2_decap_8 FILLER_78_1921 ();
 sg13g2_decap_8 FILLER_78_1928 ();
 sg13g2_decap_8 FILLER_78_1935 ();
 sg13g2_decap_8 FILLER_78_1942 ();
 sg13g2_decap_8 FILLER_78_1949 ();
 sg13g2_decap_8 FILLER_78_1956 ();
 sg13g2_decap_8 FILLER_78_1963 ();
 sg13g2_decap_8 FILLER_78_1970 ();
 sg13g2_fill_2 FILLER_78_1977 ();
 sg13g2_decap_8 FILLER_78_1984 ();
 sg13g2_decap_8 FILLER_78_1991 ();
 sg13g2_decap_8 FILLER_78_1998 ();
 sg13g2_decap_4 FILLER_78_2005 ();
 sg13g2_fill_1 FILLER_78_2009 ();
 sg13g2_decap_8 FILLER_78_2014 ();
 sg13g2_decap_8 FILLER_78_2021 ();
 sg13g2_decap_8 FILLER_78_2028 ();
 sg13g2_decap_8 FILLER_78_2035 ();
 sg13g2_decap_8 FILLER_78_2042 ();
 sg13g2_decap_8 FILLER_78_2049 ();
 sg13g2_decap_8 FILLER_78_2056 ();
 sg13g2_decap_8 FILLER_78_2063 ();
 sg13g2_decap_8 FILLER_78_2070 ();
 sg13g2_decap_8 FILLER_78_2077 ();
 sg13g2_fill_1 FILLER_78_2084 ();
 sg13g2_fill_2 FILLER_78_2111 ();
 sg13g2_fill_1 FILLER_78_2130 ();
 sg13g2_fill_2 FILLER_78_2161 ();
 sg13g2_fill_1 FILLER_78_2193 ();
 sg13g2_fill_2 FILLER_78_2225 ();
 sg13g2_fill_1 FILLER_78_2227 ();
 sg13g2_fill_2 FILLER_78_2254 ();
 sg13g2_fill_1 FILLER_78_2260 ();
 sg13g2_fill_1 FILLER_78_2374 ();
 sg13g2_fill_2 FILLER_78_2440 ();
 sg13g2_fill_1 FILLER_78_2468 ();
 sg13g2_fill_2 FILLER_78_2495 ();
 sg13g2_fill_1 FILLER_78_2523 ();
 sg13g2_fill_2 FILLER_78_2550 ();
 sg13g2_decap_8 FILLER_78_2581 ();
 sg13g2_decap_8 FILLER_78_2588 ();
 sg13g2_decap_8 FILLER_78_2595 ();
 sg13g2_decap_8 FILLER_78_2602 ();
 sg13g2_decap_8 FILLER_78_2609 ();
 sg13g2_decap_8 FILLER_78_2616 ();
 sg13g2_decap_8 FILLER_78_2623 ();
 sg13g2_decap_8 FILLER_78_2630 ();
 sg13g2_decap_8 FILLER_78_2637 ();
 sg13g2_decap_8 FILLER_78_2644 ();
 sg13g2_decap_8 FILLER_78_2651 ();
 sg13g2_decap_8 FILLER_78_2658 ();
 sg13g2_decap_4 FILLER_78_2665 ();
 sg13g2_fill_1 FILLER_78_2669 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_34 ();
 sg13g2_fill_2 FILLER_79_39 ();
 sg13g2_fill_1 FILLER_79_46 ();
 sg13g2_fill_2 FILLER_79_73 ();
 sg13g2_fill_1 FILLER_79_80 ();
 sg13g2_fill_1 FILLER_79_96 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_118 ();
 sg13g2_fill_1 FILLER_79_132 ();
 sg13g2_fill_1 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_142 ();
 sg13g2_fill_1 FILLER_79_148 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_2 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_2 FILLER_79_258 ();
 sg13g2_decap_8 FILLER_79_268 ();
 sg13g2_decap_4 FILLER_79_275 ();
 sg13g2_fill_2 FILLER_79_279 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_4 FILLER_79_317 ();
 sg13g2_fill_2 FILLER_79_321 ();
 sg13g2_fill_2 FILLER_79_328 ();
 sg13g2_decap_4 FILLER_79_334 ();
 sg13g2_fill_1 FILLER_79_338 ();
 sg13g2_fill_1 FILLER_79_366 ();
 sg13g2_fill_1 FILLER_79_380 ();
 sg13g2_fill_2 FILLER_79_385 ();
 sg13g2_fill_1 FILLER_79_450 ();
 sg13g2_fill_1 FILLER_79_465 ();
 sg13g2_decap_4 FILLER_79_492 ();
 sg13g2_decap_8 FILLER_79_537 ();
 sg13g2_decap_4 FILLER_79_544 ();
 sg13g2_fill_1 FILLER_79_556 ();
 sg13g2_fill_1 FILLER_79_562 ();
 sg13g2_fill_1 FILLER_79_568 ();
 sg13g2_fill_1 FILLER_79_574 ();
 sg13g2_fill_1 FILLER_79_601 ();
 sg13g2_fill_1 FILLER_79_612 ();
 sg13g2_fill_2 FILLER_79_644 ();
 sg13g2_fill_1 FILLER_79_646 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_fill_2 FILLER_79_687 ();
 sg13g2_fill_1 FILLER_79_720 ();
 sg13g2_fill_2 FILLER_79_750 ();
 sg13g2_fill_1 FILLER_79_848 ();
 sg13g2_fill_1 FILLER_79_875 ();
 sg13g2_fill_1 FILLER_79_985 ();
 sg13g2_fill_1 FILLER_79_1067 ();
 sg13g2_decap_4 FILLER_79_1116 ();
 sg13g2_fill_2 FILLER_79_1154 ();
 sg13g2_fill_1 FILLER_79_1156 ();
 sg13g2_decap_8 FILLER_79_1174 ();
 sg13g2_fill_1 FILLER_79_1181 ();
 sg13g2_fill_2 FILLER_79_1258 ();
 sg13g2_fill_2 FILLER_79_1346 ();
 sg13g2_decap_8 FILLER_79_1379 ();
 sg13g2_decap_4 FILLER_79_1386 ();
 sg13g2_fill_2 FILLER_79_1403 ();
 sg13g2_fill_1 FILLER_79_1405 ();
 sg13g2_fill_1 FILLER_79_1411 ();
 sg13g2_fill_2 FILLER_79_1416 ();
 sg13g2_fill_1 FILLER_79_1418 ();
 sg13g2_decap_8 FILLER_79_1424 ();
 sg13g2_decap_4 FILLER_79_1431 ();
 sg13g2_fill_2 FILLER_79_1435 ();
 sg13g2_decap_4 FILLER_79_1447 ();
 sg13g2_decap_4 FILLER_79_1456 ();
 sg13g2_decap_4 FILLER_79_1486 ();
 sg13g2_fill_2 FILLER_79_1490 ();
 sg13g2_fill_2 FILLER_79_1518 ();
 sg13g2_fill_1 FILLER_79_1528 ();
 sg13g2_decap_4 FILLER_79_1557 ();
 sg13g2_fill_1 FILLER_79_1561 ();
 sg13g2_decap_4 FILLER_79_1567 ();
 sg13g2_fill_1 FILLER_79_1571 ();
 sg13g2_fill_1 FILLER_79_1576 ();
 sg13g2_fill_1 FILLER_79_1586 ();
 sg13g2_fill_1 FILLER_79_1592 ();
 sg13g2_decap_8 FILLER_79_1597 ();
 sg13g2_decap_8 FILLER_79_1604 ();
 sg13g2_decap_8 FILLER_79_1611 ();
 sg13g2_decap_8 FILLER_79_1618 ();
 sg13g2_decap_8 FILLER_79_1625 ();
 sg13g2_decap_8 FILLER_79_1632 ();
 sg13g2_decap_8 FILLER_79_1639 ();
 sg13g2_decap_8 FILLER_79_1646 ();
 sg13g2_decap_8 FILLER_79_1653 ();
 sg13g2_decap_8 FILLER_79_1660 ();
 sg13g2_decap_8 FILLER_79_1667 ();
 sg13g2_decap_8 FILLER_79_1674 ();
 sg13g2_decap_8 FILLER_79_1681 ();
 sg13g2_decap_8 FILLER_79_1688 ();
 sg13g2_decap_8 FILLER_79_1695 ();
 sg13g2_decap_8 FILLER_79_1702 ();
 sg13g2_decap_8 FILLER_79_1709 ();
 sg13g2_decap_8 FILLER_79_1716 ();
 sg13g2_decap_8 FILLER_79_1723 ();
 sg13g2_decap_8 FILLER_79_1730 ();
 sg13g2_decap_8 FILLER_79_1737 ();
 sg13g2_decap_8 FILLER_79_1744 ();
 sg13g2_decap_8 FILLER_79_1751 ();
 sg13g2_decap_8 FILLER_79_1758 ();
 sg13g2_decap_8 FILLER_79_1765 ();
 sg13g2_decap_8 FILLER_79_1772 ();
 sg13g2_decap_8 FILLER_79_1779 ();
 sg13g2_decap_8 FILLER_79_1786 ();
 sg13g2_decap_8 FILLER_79_1793 ();
 sg13g2_decap_8 FILLER_79_1800 ();
 sg13g2_decap_8 FILLER_79_1807 ();
 sg13g2_decap_8 FILLER_79_1814 ();
 sg13g2_decap_8 FILLER_79_1821 ();
 sg13g2_decap_8 FILLER_79_1828 ();
 sg13g2_decap_8 FILLER_79_1835 ();
 sg13g2_decap_8 FILLER_79_1842 ();
 sg13g2_decap_8 FILLER_79_1849 ();
 sg13g2_decap_8 FILLER_79_1856 ();
 sg13g2_decap_8 FILLER_79_1863 ();
 sg13g2_decap_8 FILLER_79_1870 ();
 sg13g2_decap_8 FILLER_79_1877 ();
 sg13g2_decap_8 FILLER_79_1884 ();
 sg13g2_decap_8 FILLER_79_1891 ();
 sg13g2_decap_8 FILLER_79_1898 ();
 sg13g2_decap_8 FILLER_79_1905 ();
 sg13g2_decap_8 FILLER_79_1912 ();
 sg13g2_decap_8 FILLER_79_1919 ();
 sg13g2_decap_8 FILLER_79_1926 ();
 sg13g2_decap_8 FILLER_79_1933 ();
 sg13g2_decap_8 FILLER_79_1940 ();
 sg13g2_decap_8 FILLER_79_1947 ();
 sg13g2_decap_8 FILLER_79_1954 ();
 sg13g2_decap_8 FILLER_79_1961 ();
 sg13g2_decap_8 FILLER_79_1968 ();
 sg13g2_decap_8 FILLER_79_1975 ();
 sg13g2_decap_8 FILLER_79_1982 ();
 sg13g2_decap_8 FILLER_79_1989 ();
 sg13g2_decap_8 FILLER_79_1996 ();
 sg13g2_decap_8 FILLER_79_2003 ();
 sg13g2_decap_8 FILLER_79_2010 ();
 sg13g2_decap_8 FILLER_79_2017 ();
 sg13g2_decap_8 FILLER_79_2024 ();
 sg13g2_decap_8 FILLER_79_2031 ();
 sg13g2_decap_8 FILLER_79_2038 ();
 sg13g2_decap_8 FILLER_79_2045 ();
 sg13g2_decap_8 FILLER_79_2052 ();
 sg13g2_decap_8 FILLER_79_2059 ();
 sg13g2_decap_8 FILLER_79_2066 ();
 sg13g2_decap_8 FILLER_79_2073 ();
 sg13g2_fill_2 FILLER_79_2080 ();
 sg13g2_fill_2 FILLER_79_2108 ();
 sg13g2_fill_1 FILLER_79_2110 ();
 sg13g2_fill_2 FILLER_79_2121 ();
 sg13g2_fill_1 FILLER_79_2123 ();
 sg13g2_fill_2 FILLER_79_2150 ();
 sg13g2_fill_1 FILLER_79_2152 ();
 sg13g2_fill_2 FILLER_79_2157 ();
 sg13g2_fill_1 FILLER_79_2159 ();
 sg13g2_fill_2 FILLER_79_2186 ();
 sg13g2_fill_1 FILLER_79_2193 ();
 sg13g2_fill_1 FILLER_79_2225 ();
 sg13g2_fill_2 FILLER_79_2239 ();
 sg13g2_fill_2 FILLER_79_2267 ();
 sg13g2_fill_1 FILLER_79_2295 ();
 sg13g2_fill_2 FILLER_79_2306 ();
 sg13g2_fill_1 FILLER_79_2360 ();
 sg13g2_fill_1 FILLER_79_2437 ();
 sg13g2_fill_1 FILLER_79_2469 ();
 sg13g2_fill_1 FILLER_79_2502 ();
 sg13g2_fill_2 FILLER_79_2507 ();
 sg13g2_fill_2 FILLER_79_2513 ();
 sg13g2_fill_2 FILLER_79_2565 ();
 sg13g2_decap_8 FILLER_79_2583 ();
 sg13g2_decap_8 FILLER_79_2590 ();
 sg13g2_decap_8 FILLER_79_2597 ();
 sg13g2_decap_8 FILLER_79_2604 ();
 sg13g2_decap_8 FILLER_79_2611 ();
 sg13g2_decap_8 FILLER_79_2618 ();
 sg13g2_decap_8 FILLER_79_2625 ();
 sg13g2_decap_8 FILLER_79_2632 ();
 sg13g2_decap_8 FILLER_79_2639 ();
 sg13g2_decap_8 FILLER_79_2646 ();
 sg13g2_decap_8 FILLER_79_2653 ();
 sg13g2_decap_8 FILLER_79_2660 ();
 sg13g2_fill_2 FILLER_79_2667 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_32 ();
 sg13g2_decap_8 FILLER_80_37 ();
 sg13g2_decap_8 FILLER_80_44 ();
 sg13g2_fill_2 FILLER_80_51 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_fill_1 FILLER_80_161 ();
 sg13g2_fill_2 FILLER_80_169 ();
 sg13g2_fill_1 FILLER_80_171 ();
 sg13g2_fill_1 FILLER_80_203 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_2 FILLER_80_244 ();
 sg13g2_decap_4 FILLER_80_250 ();
 sg13g2_fill_1 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_259 ();
 sg13g2_fill_2 FILLER_80_266 ();
 sg13g2_decap_4 FILLER_80_273 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_4 FILLER_80_313 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_344 ();
 sg13g2_fill_1 FILLER_80_352 ();
 sg13g2_fill_2 FILLER_80_364 ();
 sg13g2_fill_2 FILLER_80_400 ();
 sg13g2_fill_1 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_420 ();
 sg13g2_fill_2 FILLER_80_443 ();
 sg13g2_fill_2 FILLER_80_457 ();
 sg13g2_fill_1 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_fill_1 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_decap_8 FILLER_80_545 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_decap_4 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_4 FILLER_80_575 ();
 sg13g2_fill_2 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_4 FILLER_80_613 ();
 sg13g2_fill_1 FILLER_80_621 ();
 sg13g2_fill_2 FILLER_80_626 ();
 sg13g2_fill_1 FILLER_80_633 ();
 sg13g2_fill_2 FILLER_80_647 ();
 sg13g2_fill_1 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_fill_2 FILLER_80_691 ();
 sg13g2_fill_1 FILLER_80_693 ();
 sg13g2_fill_2 FILLER_80_707 ();
 sg13g2_fill_1 FILLER_80_709 ();
 sg13g2_fill_2 FILLER_80_720 ();
 sg13g2_fill_2 FILLER_80_742 ();
 sg13g2_fill_1 FILLER_80_754 ();
 sg13g2_fill_1 FILLER_80_771 ();
 sg13g2_fill_2 FILLER_80_775 ();
 sg13g2_fill_1 FILLER_80_814 ();
 sg13g2_fill_1 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_4 FILLER_80_849 ();
 sg13g2_fill_2 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_862 ();
 sg13g2_fill_1 FILLER_80_864 ();
 sg13g2_fill_1 FILLER_80_874 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_fill_1 FILLER_80_910 ();
 sg13g2_decap_4 FILLER_80_925 ();
 sg13g2_fill_2 FILLER_80_929 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_fill_1 FILLER_80_942 ();
 sg13g2_decap_4 FILLER_80_947 ();
 sg13g2_fill_1 FILLER_80_951 ();
 sg13g2_fill_2 FILLER_80_977 ();
 sg13g2_fill_1 FILLER_80_998 ();
 sg13g2_fill_1 FILLER_80_1006 ();
 sg13g2_decap_8 FILLER_80_1014 ();
 sg13g2_decap_8 FILLER_80_1021 ();
 sg13g2_fill_2 FILLER_80_1028 ();
 sg13g2_fill_1 FILLER_80_1030 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_4 FILLER_80_1082 ();
 sg13g2_decap_8 FILLER_80_1094 ();
 sg13g2_decap_8 FILLER_80_1101 ();
 sg13g2_decap_4 FILLER_80_1108 ();
 sg13g2_fill_1 FILLER_80_1112 ();
 sg13g2_decap_8 FILLER_80_1143 ();
 sg13g2_decap_8 FILLER_80_1150 ();
 sg13g2_decap_8 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1171 ();
 sg13g2_fill_2 FILLER_80_1178 ();
 sg13g2_decap_4 FILLER_80_1206 ();
 sg13g2_fill_2 FILLER_80_1210 ();
 sg13g2_decap_8 FILLER_80_1220 ();
 sg13g2_decap_4 FILLER_80_1227 ();
 sg13g2_fill_1 FILLER_80_1231 ();
 sg13g2_fill_1 FILLER_80_1246 ();
 sg13g2_fill_2 FILLER_80_1295 ();
 sg13g2_fill_2 FILLER_80_1318 ();
 sg13g2_fill_1 FILLER_80_1337 ();
 sg13g2_fill_2 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_decap_8 FILLER_80_1376 ();
 sg13g2_decap_8 FILLER_80_1383 ();
 sg13g2_decap_8 FILLER_80_1390 ();
 sg13g2_decap_4 FILLER_80_1397 ();
 sg13g2_fill_1 FILLER_80_1401 ();
 sg13g2_decap_8 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1413 ();
 sg13g2_decap_8 FILLER_80_1420 ();
 sg13g2_decap_8 FILLER_80_1427 ();
 sg13g2_decap_8 FILLER_80_1434 ();
 sg13g2_decap_8 FILLER_80_1441 ();
 sg13g2_decap_8 FILLER_80_1448 ();
 sg13g2_decap_8 FILLER_80_1455 ();
 sg13g2_decap_4 FILLER_80_1462 ();
 sg13g2_fill_1 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1471 ();
 sg13g2_decap_8 FILLER_80_1478 ();
 sg13g2_decap_8 FILLER_80_1485 ();
 sg13g2_decap_4 FILLER_80_1492 ();
 sg13g2_fill_2 FILLER_80_1496 ();
 sg13g2_decap_8 FILLER_80_1502 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_decap_8 FILLER_80_1516 ();
 sg13g2_decap_8 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1530 ();
 sg13g2_decap_8 FILLER_80_1537 ();
 sg13g2_decap_8 FILLER_80_1544 ();
 sg13g2_decap_8 FILLER_80_1551 ();
 sg13g2_decap_8 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1572 ();
 sg13g2_decap_8 FILLER_80_1579 ();
 sg13g2_decap_8 FILLER_80_1586 ();
 sg13g2_decap_8 FILLER_80_1593 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_8 FILLER_80_1607 ();
 sg13g2_decap_8 FILLER_80_1614 ();
 sg13g2_decap_8 FILLER_80_1621 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_8 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1691 ();
 sg13g2_decap_8 FILLER_80_1698 ();
 sg13g2_decap_8 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1712 ();
 sg13g2_decap_8 FILLER_80_1719 ();
 sg13g2_decap_8 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_80_1768 ();
 sg13g2_decap_8 FILLER_80_1775 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_8 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1803 ();
 sg13g2_decap_8 FILLER_80_1810 ();
 sg13g2_decap_8 FILLER_80_1817 ();
 sg13g2_decap_8 FILLER_80_1824 ();
 sg13g2_decap_8 FILLER_80_1831 ();
 sg13g2_decap_8 FILLER_80_1838 ();
 sg13g2_decap_8 FILLER_80_1845 ();
 sg13g2_decap_8 FILLER_80_1852 ();
 sg13g2_decap_8 FILLER_80_1859 ();
 sg13g2_decap_8 FILLER_80_1866 ();
 sg13g2_decap_8 FILLER_80_1873 ();
 sg13g2_decap_8 FILLER_80_1880 ();
 sg13g2_decap_8 FILLER_80_1887 ();
 sg13g2_decap_8 FILLER_80_1894 ();
 sg13g2_decap_8 FILLER_80_1901 ();
 sg13g2_decap_8 FILLER_80_1908 ();
 sg13g2_decap_8 FILLER_80_1915 ();
 sg13g2_decap_8 FILLER_80_1922 ();
 sg13g2_decap_8 FILLER_80_1929 ();
 sg13g2_decap_8 FILLER_80_1936 ();
 sg13g2_decap_8 FILLER_80_1943 ();
 sg13g2_decap_8 FILLER_80_1950 ();
 sg13g2_decap_8 FILLER_80_1957 ();
 sg13g2_decap_8 FILLER_80_1964 ();
 sg13g2_decap_8 FILLER_80_1971 ();
 sg13g2_decap_8 FILLER_80_1978 ();
 sg13g2_decap_8 FILLER_80_1985 ();
 sg13g2_decap_8 FILLER_80_1992 ();
 sg13g2_decap_8 FILLER_80_1999 ();
 sg13g2_decap_8 FILLER_80_2006 ();
 sg13g2_decap_8 FILLER_80_2013 ();
 sg13g2_decap_8 FILLER_80_2020 ();
 sg13g2_decap_8 FILLER_80_2027 ();
 sg13g2_decap_8 FILLER_80_2034 ();
 sg13g2_decap_8 FILLER_80_2041 ();
 sg13g2_decap_8 FILLER_80_2048 ();
 sg13g2_decap_8 FILLER_80_2055 ();
 sg13g2_decap_8 FILLER_80_2062 ();
 sg13g2_decap_8 FILLER_80_2069 ();
 sg13g2_decap_8 FILLER_80_2076 ();
 sg13g2_decap_4 FILLER_80_2083 ();
 sg13g2_fill_2 FILLER_80_2091 ();
 sg13g2_decap_8 FILLER_80_2097 ();
 sg13g2_decap_4 FILLER_80_2104 ();
 sg13g2_decap_4 FILLER_80_2122 ();
 sg13g2_fill_2 FILLER_80_2126 ();
 sg13g2_fill_2 FILLER_80_2132 ();
 sg13g2_fill_1 FILLER_80_2134 ();
 sg13g2_decap_4 FILLER_80_2161 ();
 sg13g2_fill_2 FILLER_80_2165 ();
 sg13g2_fill_2 FILLER_80_2179 ();
 sg13g2_fill_1 FILLER_80_2181 ();
 sg13g2_decap_4 FILLER_80_2186 ();
 sg13g2_fill_1 FILLER_80_2190 ();
 sg13g2_decap_4 FILLER_80_2195 ();
 sg13g2_decap_8 FILLER_80_2207 ();
 sg13g2_decap_4 FILLER_80_2214 ();
 sg13g2_fill_1 FILLER_80_2218 ();
 sg13g2_fill_1 FILLER_80_2251 ();
 sg13g2_fill_2 FILLER_80_2286 ();
 sg13g2_fill_1 FILLER_80_2294 ();
 sg13g2_fill_1 FILLER_80_2322 ();
 sg13g2_fill_1 FILLER_80_2342 ();
 sg13g2_fill_1 FILLER_80_2351 ();
 sg13g2_fill_1 FILLER_80_2359 ();
 sg13g2_fill_2 FILLER_80_2373 ();
 sg13g2_fill_1 FILLER_80_2402 ();
 sg13g2_fill_2 FILLER_80_2432 ();
 sg13g2_fill_1 FILLER_80_2490 ();
 sg13g2_fill_1 FILLER_80_2507 ();
 sg13g2_fill_2 FILLER_80_2541 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_4 FILLER_80_2665 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
