module tt_um_tommythorn_maxbw (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire net199;
 wire \tokenflow_inst.i1.c.q ;
 wire \tokenflow_inst.i10.cg.b ;
 wire \tokenflow_inst.i10.d0.inv_chain[0] ;
 wire \tokenflow_inst.i10.d0.inv_chain[1] ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[0] ;
 wire \tokenflow_inst.i11.i.d0.inv_chain[1] ;
 wire \tokenflow_inst.i2.cg1.a ;
 wire \tokenflow_inst.i2.cg1.q ;
 wire \tokenflow_inst.i2.cg2.a ;
 wire \tokenflow_inst.i2.cg2.q ;
 wire \tokenflow_inst.i3.cg_elem.a ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i3.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i3.ydata[0] ;
 wire \tokenflow_inst.i3.ydata[10] ;
 wire \tokenflow_inst.i3.ydata[11] ;
 wire \tokenflow_inst.i3.ydata[12] ;
 wire \tokenflow_inst.i3.ydata[13] ;
 wire \tokenflow_inst.i3.ydata[14] ;
 wire \tokenflow_inst.i3.ydata[15] ;
 wire \tokenflow_inst.i3.ydata[16] ;
 wire \tokenflow_inst.i3.ydata[17] ;
 wire \tokenflow_inst.i3.ydata[18] ;
 wire \tokenflow_inst.i3.ydata[19] ;
 wire \tokenflow_inst.i3.ydata[1] ;
 wire \tokenflow_inst.i3.ydata[20] ;
 wire \tokenflow_inst.i3.ydata[21] ;
 wire \tokenflow_inst.i3.ydata[22] ;
 wire \tokenflow_inst.i3.ydata[23] ;
 wire \tokenflow_inst.i3.ydata[24] ;
 wire \tokenflow_inst.i3.ydata[25] ;
 wire \tokenflow_inst.i3.ydata[26] ;
 wire \tokenflow_inst.i3.ydata[27] ;
 wire \tokenflow_inst.i3.ydata[28] ;
 wire \tokenflow_inst.i3.ydata[29] ;
 wire \tokenflow_inst.i3.ydata[2] ;
 wire \tokenflow_inst.i3.ydata[30] ;
 wire \tokenflow_inst.i3.ydata[31] ;
 wire \tokenflow_inst.i3.ydata[32] ;
 wire \tokenflow_inst.i3.ydata[33] ;
 wire \tokenflow_inst.i3.ydata[34] ;
 wire \tokenflow_inst.i3.ydata[35] ;
 wire \tokenflow_inst.i3.ydata[36] ;
 wire \tokenflow_inst.i3.ydata[37] ;
 wire \tokenflow_inst.i3.ydata[38] ;
 wire \tokenflow_inst.i3.ydata[39] ;
 wire \tokenflow_inst.i3.ydata[3] ;
 wire \tokenflow_inst.i3.ydata[40] ;
 wire \tokenflow_inst.i3.ydata[41] ;
 wire \tokenflow_inst.i3.ydata[42] ;
 wire \tokenflow_inst.i3.ydata[43] ;
 wire \tokenflow_inst.i3.ydata[44] ;
 wire \tokenflow_inst.i3.ydata[45] ;
 wire \tokenflow_inst.i3.ydata[46] ;
 wire \tokenflow_inst.i3.ydata[47] ;
 wire \tokenflow_inst.i3.ydata[48] ;
 wire \tokenflow_inst.i3.ydata[49] ;
 wire \tokenflow_inst.i3.ydata[4] ;
 wire \tokenflow_inst.i3.ydata[50] ;
 wire \tokenflow_inst.i3.ydata[51] ;
 wire \tokenflow_inst.i3.ydata[52] ;
 wire \tokenflow_inst.i3.ydata[53] ;
 wire \tokenflow_inst.i3.ydata[54] ;
 wire \tokenflow_inst.i3.ydata[55] ;
 wire \tokenflow_inst.i3.ydata[56] ;
 wire \tokenflow_inst.i3.ydata[57] ;
 wire \tokenflow_inst.i3.ydata[58] ;
 wire \tokenflow_inst.i3.ydata[59] ;
 wire \tokenflow_inst.i3.ydata[5] ;
 wire \tokenflow_inst.i3.ydata[60] ;
 wire \tokenflow_inst.i3.ydata[61] ;
 wire \tokenflow_inst.i3.ydata[62] ;
 wire \tokenflow_inst.i3.ydata[63] ;
 wire \tokenflow_inst.i3.ydata[64] ;
 wire \tokenflow_inst.i3.ydata[65] ;
 wire \tokenflow_inst.i3.ydata[66] ;
 wire \tokenflow_inst.i3.ydata[67] ;
 wire \tokenflow_inst.i3.ydata[68] ;
 wire \tokenflow_inst.i3.ydata[69] ;
 wire \tokenflow_inst.i3.ydata[6] ;
 wire \tokenflow_inst.i3.ydata[70] ;
 wire \tokenflow_inst.i3.ydata[71] ;
 wire \tokenflow_inst.i3.ydata[72] ;
 wire \tokenflow_inst.i3.ydata[73] ;
 wire \tokenflow_inst.i3.ydata[74] ;
 wire \tokenflow_inst.i3.ydata[75] ;
 wire \tokenflow_inst.i3.ydata[76] ;
 wire \tokenflow_inst.i3.ydata[77] ;
 wire \tokenflow_inst.i3.ydata[7] ;
 wire \tokenflow_inst.i3.ydata[8] ;
 wire \tokenflow_inst.i3.ydata[9] ;
 wire \tokenflow_inst.i6.cg_elem.a ;
 wire \tokenflow_inst.i6.cg_elem.q ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i6.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i6.ydata[0] ;
 wire \tokenflow_inst.i6.ydata[10] ;
 wire \tokenflow_inst.i6.ydata[11] ;
 wire \tokenflow_inst.i6.ydata[12] ;
 wire \tokenflow_inst.i6.ydata[13] ;
 wire \tokenflow_inst.i6.ydata[14] ;
 wire \tokenflow_inst.i6.ydata[15] ;
 wire \tokenflow_inst.i6.ydata[16] ;
 wire \tokenflow_inst.i6.ydata[17] ;
 wire \tokenflow_inst.i6.ydata[18] ;
 wire \tokenflow_inst.i6.ydata[19] ;
 wire \tokenflow_inst.i6.ydata[1] ;
 wire \tokenflow_inst.i6.ydata[20] ;
 wire \tokenflow_inst.i6.ydata[21] ;
 wire \tokenflow_inst.i6.ydata[22] ;
 wire \tokenflow_inst.i6.ydata[23] ;
 wire \tokenflow_inst.i6.ydata[24] ;
 wire \tokenflow_inst.i6.ydata[25] ;
 wire \tokenflow_inst.i6.ydata[26] ;
 wire \tokenflow_inst.i6.ydata[27] ;
 wire \tokenflow_inst.i6.ydata[28] ;
 wire \tokenflow_inst.i6.ydata[29] ;
 wire \tokenflow_inst.i6.ydata[2] ;
 wire \tokenflow_inst.i6.ydata[30] ;
 wire \tokenflow_inst.i6.ydata[31] ;
 wire \tokenflow_inst.i6.ydata[32] ;
 wire \tokenflow_inst.i6.ydata[33] ;
 wire \tokenflow_inst.i6.ydata[34] ;
 wire \tokenflow_inst.i6.ydata[35] ;
 wire \tokenflow_inst.i6.ydata[36] ;
 wire \tokenflow_inst.i6.ydata[37] ;
 wire \tokenflow_inst.i6.ydata[38] ;
 wire \tokenflow_inst.i6.ydata[39] ;
 wire \tokenflow_inst.i6.ydata[3] ;
 wire \tokenflow_inst.i6.ydata[40] ;
 wire \tokenflow_inst.i6.ydata[41] ;
 wire \tokenflow_inst.i6.ydata[42] ;
 wire \tokenflow_inst.i6.ydata[43] ;
 wire \tokenflow_inst.i6.ydata[44] ;
 wire \tokenflow_inst.i6.ydata[45] ;
 wire \tokenflow_inst.i6.ydata[46] ;
 wire \tokenflow_inst.i6.ydata[47] ;
 wire \tokenflow_inst.i6.ydata[48] ;
 wire \tokenflow_inst.i6.ydata[49] ;
 wire \tokenflow_inst.i6.ydata[4] ;
 wire \tokenflow_inst.i6.ydata[50] ;
 wire \tokenflow_inst.i6.ydata[51] ;
 wire \tokenflow_inst.i6.ydata[52] ;
 wire \tokenflow_inst.i6.ydata[53] ;
 wire \tokenflow_inst.i6.ydata[54] ;
 wire \tokenflow_inst.i6.ydata[55] ;
 wire \tokenflow_inst.i6.ydata[56] ;
 wire \tokenflow_inst.i6.ydata[57] ;
 wire \tokenflow_inst.i6.ydata[58] ;
 wire \tokenflow_inst.i6.ydata[59] ;
 wire \tokenflow_inst.i6.ydata[5] ;
 wire \tokenflow_inst.i6.ydata[60] ;
 wire \tokenflow_inst.i6.ydata[61] ;
 wire \tokenflow_inst.i6.ydata[62] ;
 wire \tokenflow_inst.i6.ydata[63] ;
 wire \tokenflow_inst.i6.ydata[64] ;
 wire \tokenflow_inst.i6.ydata[65] ;
 wire \tokenflow_inst.i6.ydata[66] ;
 wire \tokenflow_inst.i6.ydata[67] ;
 wire \tokenflow_inst.i6.ydata[68] ;
 wire \tokenflow_inst.i6.ydata[69] ;
 wire \tokenflow_inst.i6.ydata[6] ;
 wire \tokenflow_inst.i6.ydata[70] ;
 wire \tokenflow_inst.i6.ydata[71] ;
 wire \tokenflow_inst.i6.ydata[72] ;
 wire \tokenflow_inst.i6.ydata[73] ;
 wire \tokenflow_inst.i6.ydata[74] ;
 wire \tokenflow_inst.i6.ydata[75] ;
 wire \tokenflow_inst.i6.ydata[76] ;
 wire \tokenflow_inst.i6.ydata[77] ;
 wire \tokenflow_inst.i6.ydata[7] ;
 wire \tokenflow_inst.i6.ydata[8] ;
 wire \tokenflow_inst.i6.ydata[9] ;
 wire \tokenflow_inst.i78.cg_elem.a ;
 wire \tokenflow_inst.i78.cg_elem.q ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i78.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i78.ydata[0] ;
 wire \tokenflow_inst.i78.ydata[10] ;
 wire \tokenflow_inst.i78.ydata[11] ;
 wire \tokenflow_inst.i78.ydata[12] ;
 wire \tokenflow_inst.i78.ydata[13] ;
 wire \tokenflow_inst.i78.ydata[14] ;
 wire \tokenflow_inst.i78.ydata[15] ;
 wire \tokenflow_inst.i78.ydata[16] ;
 wire \tokenflow_inst.i78.ydata[17] ;
 wire \tokenflow_inst.i78.ydata[18] ;
 wire \tokenflow_inst.i78.ydata[19] ;
 wire \tokenflow_inst.i78.ydata[1] ;
 wire \tokenflow_inst.i78.ydata[20] ;
 wire \tokenflow_inst.i78.ydata[21] ;
 wire \tokenflow_inst.i78.ydata[22] ;
 wire \tokenflow_inst.i78.ydata[23] ;
 wire \tokenflow_inst.i78.ydata[24] ;
 wire \tokenflow_inst.i78.ydata[25] ;
 wire \tokenflow_inst.i78.ydata[26] ;
 wire \tokenflow_inst.i78.ydata[27] ;
 wire \tokenflow_inst.i78.ydata[28] ;
 wire \tokenflow_inst.i78.ydata[29] ;
 wire \tokenflow_inst.i78.ydata[2] ;
 wire \tokenflow_inst.i78.ydata[30] ;
 wire \tokenflow_inst.i78.ydata[31] ;
 wire \tokenflow_inst.i78.ydata[32] ;
 wire \tokenflow_inst.i78.ydata[33] ;
 wire \tokenflow_inst.i78.ydata[34] ;
 wire \tokenflow_inst.i78.ydata[35] ;
 wire \tokenflow_inst.i78.ydata[36] ;
 wire \tokenflow_inst.i78.ydata[37] ;
 wire \tokenflow_inst.i78.ydata[38] ;
 wire \tokenflow_inst.i78.ydata[39] ;
 wire \tokenflow_inst.i78.ydata[3] ;
 wire \tokenflow_inst.i78.ydata[40] ;
 wire \tokenflow_inst.i78.ydata[41] ;
 wire \tokenflow_inst.i78.ydata[42] ;
 wire \tokenflow_inst.i78.ydata[43] ;
 wire \tokenflow_inst.i78.ydata[44] ;
 wire \tokenflow_inst.i78.ydata[45] ;
 wire \tokenflow_inst.i78.ydata[46] ;
 wire \tokenflow_inst.i78.ydata[47] ;
 wire \tokenflow_inst.i78.ydata[48] ;
 wire \tokenflow_inst.i78.ydata[49] ;
 wire \tokenflow_inst.i78.ydata[4] ;
 wire \tokenflow_inst.i78.ydata[50] ;
 wire \tokenflow_inst.i78.ydata[51] ;
 wire \tokenflow_inst.i78.ydata[52] ;
 wire \tokenflow_inst.i78.ydata[53] ;
 wire \tokenflow_inst.i78.ydata[54] ;
 wire \tokenflow_inst.i78.ydata[55] ;
 wire \tokenflow_inst.i78.ydata[56] ;
 wire \tokenflow_inst.i78.ydata[57] ;
 wire \tokenflow_inst.i78.ydata[58] ;
 wire \tokenflow_inst.i78.ydata[59] ;
 wire \tokenflow_inst.i78.ydata[5] ;
 wire \tokenflow_inst.i78.ydata[60] ;
 wire \tokenflow_inst.i78.ydata[61] ;
 wire \tokenflow_inst.i78.ydata[62] ;
 wire \tokenflow_inst.i78.ydata[63] ;
 wire \tokenflow_inst.i78.ydata[64] ;
 wire \tokenflow_inst.i78.ydata[65] ;
 wire \tokenflow_inst.i78.ydata[66] ;
 wire \tokenflow_inst.i78.ydata[67] ;
 wire \tokenflow_inst.i78.ydata[68] ;
 wire \tokenflow_inst.i78.ydata[69] ;
 wire \tokenflow_inst.i78.ydata[6] ;
 wire \tokenflow_inst.i78.ydata[70] ;
 wire \tokenflow_inst.i78.ydata[71] ;
 wire \tokenflow_inst.i78.ydata[72] ;
 wire \tokenflow_inst.i78.ydata[73] ;
 wire \tokenflow_inst.i78.ydata[74] ;
 wire \tokenflow_inst.i78.ydata[75] ;
 wire \tokenflow_inst.i78.ydata[76] ;
 wire \tokenflow_inst.i78.ydata[77] ;
 wire \tokenflow_inst.i78.ydata[7] ;
 wire \tokenflow_inst.i78.ydata[8] ;
 wire \tokenflow_inst.i78.ydata[9] ;
 wire \tokenflow_inst.i8.cg_elem.a ;
 wire \tokenflow_inst.i8.cg_elem.q ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[10] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[11] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[12] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[13] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[14] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[15] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[16] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[17] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[18] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[19] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[20] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[21] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[22] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[23] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[24] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[25] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[26] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[27] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[28] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[29] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[30] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[31] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[32] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[33] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[34] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[35] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[36] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[37] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[38] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[39] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[3] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[40] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[41] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[42] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[43] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[44] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[45] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[46] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[47] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[48] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[49] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[4] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[50] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[51] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[52] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[5] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[6] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[7] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[8] ;
 wire \tokenflow_inst.i8.d0_elem.inv_chain[9] ;
 wire \tokenflow_inst.i8.ydata[0] ;
 wire \tokenflow_inst.i8.ydata[10] ;
 wire \tokenflow_inst.i8.ydata[11] ;
 wire \tokenflow_inst.i8.ydata[12] ;
 wire \tokenflow_inst.i8.ydata[13] ;
 wire \tokenflow_inst.i8.ydata[14] ;
 wire \tokenflow_inst.i8.ydata[15] ;
 wire \tokenflow_inst.i8.ydata[16] ;
 wire \tokenflow_inst.i8.ydata[17] ;
 wire \tokenflow_inst.i8.ydata[18] ;
 wire \tokenflow_inst.i8.ydata[19] ;
 wire \tokenflow_inst.i8.ydata[1] ;
 wire \tokenflow_inst.i8.ydata[20] ;
 wire \tokenflow_inst.i8.ydata[21] ;
 wire \tokenflow_inst.i8.ydata[22] ;
 wire \tokenflow_inst.i8.ydata[23] ;
 wire \tokenflow_inst.i8.ydata[24] ;
 wire \tokenflow_inst.i8.ydata[25] ;
 wire \tokenflow_inst.i8.ydata[26] ;
 wire \tokenflow_inst.i8.ydata[27] ;
 wire \tokenflow_inst.i8.ydata[28] ;
 wire \tokenflow_inst.i8.ydata[29] ;
 wire \tokenflow_inst.i8.ydata[2] ;
 wire \tokenflow_inst.i8.ydata[30] ;
 wire \tokenflow_inst.i8.ydata[31] ;
 wire \tokenflow_inst.i8.ydata[32] ;
 wire \tokenflow_inst.i8.ydata[33] ;
 wire \tokenflow_inst.i8.ydata[34] ;
 wire \tokenflow_inst.i8.ydata[35] ;
 wire \tokenflow_inst.i8.ydata[36] ;
 wire \tokenflow_inst.i8.ydata[37] ;
 wire \tokenflow_inst.i8.ydata[38] ;
 wire \tokenflow_inst.i8.ydata[39] ;
 wire \tokenflow_inst.i8.ydata[3] ;
 wire \tokenflow_inst.i8.ydata[40] ;
 wire \tokenflow_inst.i8.ydata[41] ;
 wire \tokenflow_inst.i8.ydata[42] ;
 wire \tokenflow_inst.i8.ydata[43] ;
 wire \tokenflow_inst.i8.ydata[44] ;
 wire \tokenflow_inst.i8.ydata[45] ;
 wire \tokenflow_inst.i8.ydata[46] ;
 wire \tokenflow_inst.i8.ydata[47] ;
 wire \tokenflow_inst.i8.ydata[48] ;
 wire \tokenflow_inst.i8.ydata[49] ;
 wire \tokenflow_inst.i8.ydata[4] ;
 wire \tokenflow_inst.i8.ydata[50] ;
 wire \tokenflow_inst.i8.ydata[51] ;
 wire \tokenflow_inst.i8.ydata[52] ;
 wire \tokenflow_inst.i8.ydata[53] ;
 wire \tokenflow_inst.i8.ydata[54] ;
 wire \tokenflow_inst.i8.ydata[55] ;
 wire \tokenflow_inst.i8.ydata[56] ;
 wire \tokenflow_inst.i8.ydata[57] ;
 wire \tokenflow_inst.i8.ydata[58] ;
 wire \tokenflow_inst.i8.ydata[59] ;
 wire \tokenflow_inst.i8.ydata[5] ;
 wire \tokenflow_inst.i8.ydata[60] ;
 wire \tokenflow_inst.i8.ydata[61] ;
 wire \tokenflow_inst.i8.ydata[62] ;
 wire \tokenflow_inst.i8.ydata[63] ;
 wire \tokenflow_inst.i8.ydata[64] ;
 wire \tokenflow_inst.i8.ydata[65] ;
 wire \tokenflow_inst.i8.ydata[66] ;
 wire \tokenflow_inst.i8.ydata[67] ;
 wire \tokenflow_inst.i8.ydata[68] ;
 wire \tokenflow_inst.i8.ydata[69] ;
 wire \tokenflow_inst.i8.ydata[6] ;
 wire \tokenflow_inst.i8.ydata[70] ;
 wire \tokenflow_inst.i8.ydata[71] ;
 wire \tokenflow_inst.i8.ydata[72] ;
 wire \tokenflow_inst.i8.ydata[73] ;
 wire \tokenflow_inst.i8.ydata[74] ;
 wire \tokenflow_inst.i8.ydata[75] ;
 wire \tokenflow_inst.i8.ydata[76] ;
 wire \tokenflow_inst.i8.ydata[77] ;
 wire \tokenflow_inst.i8.ydata[7] ;
 wire \tokenflow_inst.i8.ydata[8] ;
 wire \tokenflow_inst.i8.ydata[9] ;
 wire \tokenflow_inst.i9.c.q ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii1.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii1.ydata[0] ;
 wire \tokenflow_inst.ii1.ydata[10] ;
 wire \tokenflow_inst.ii1.ydata[11] ;
 wire \tokenflow_inst.ii1.ydata[12] ;
 wire \tokenflow_inst.ii1.ydata[13] ;
 wire \tokenflow_inst.ii1.ydata[14] ;
 wire \tokenflow_inst.ii1.ydata[15] ;
 wire \tokenflow_inst.ii1.ydata[16] ;
 wire \tokenflow_inst.ii1.ydata[17] ;
 wire \tokenflow_inst.ii1.ydata[18] ;
 wire \tokenflow_inst.ii1.ydata[19] ;
 wire \tokenflow_inst.ii1.ydata[1] ;
 wire \tokenflow_inst.ii1.ydata[20] ;
 wire \tokenflow_inst.ii1.ydata[21] ;
 wire \tokenflow_inst.ii1.ydata[22] ;
 wire \tokenflow_inst.ii1.ydata[23] ;
 wire \tokenflow_inst.ii1.ydata[24] ;
 wire \tokenflow_inst.ii1.ydata[25] ;
 wire \tokenflow_inst.ii1.ydata[2] ;
 wire \tokenflow_inst.ii1.ydata[3] ;
 wire \tokenflow_inst.ii1.ydata[4] ;
 wire \tokenflow_inst.ii1.ydata[5] ;
 wire \tokenflow_inst.ii1.ydata[6] ;
 wire \tokenflow_inst.ii1.ydata[7] ;
 wire \tokenflow_inst.ii1.ydata[8] ;
 wire \tokenflow_inst.ii1.ydata[9] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii2.d0_elem.inv_chain[2] ;
 wire \tokenflow_inst.ii2.ydata[0] ;
 wire \tokenflow_inst.ii2.ydata[10] ;
 wire \tokenflow_inst.ii2.ydata[11] ;
 wire \tokenflow_inst.ii2.ydata[12] ;
 wire \tokenflow_inst.ii2.ydata[13] ;
 wire \tokenflow_inst.ii2.ydata[14] ;
 wire \tokenflow_inst.ii2.ydata[15] ;
 wire \tokenflow_inst.ii2.ydata[16] ;
 wire \tokenflow_inst.ii2.ydata[17] ;
 wire \tokenflow_inst.ii2.ydata[18] ;
 wire \tokenflow_inst.ii2.ydata[19] ;
 wire \tokenflow_inst.ii2.ydata[1] ;
 wire \tokenflow_inst.ii2.ydata[20] ;
 wire \tokenflow_inst.ii2.ydata[21] ;
 wire \tokenflow_inst.ii2.ydata[22] ;
 wire \tokenflow_inst.ii2.ydata[23] ;
 wire \tokenflow_inst.ii2.ydata[24] ;
 wire \tokenflow_inst.ii2.ydata[25] ;
 wire \tokenflow_inst.ii2.ydata[2] ;
 wire \tokenflow_inst.ii2.ydata[3] ;
 wire \tokenflow_inst.ii2.ydata[4] ;
 wire \tokenflow_inst.ii2.ydata[5] ;
 wire \tokenflow_inst.ii2.ydata[6] ;
 wire \tokenflow_inst.ii2.ydata[7] ;
 wire \tokenflow_inst.ii2.ydata[8] ;
 wire \tokenflow_inst.ii2.ydata[9] ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ;
 wire \tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ;
 wire \tokenflow_inst.ii3.i.ydata[0] ;
 wire \tokenflow_inst.ii3.i.ydata[10] ;
 wire \tokenflow_inst.ii3.i.ydata[11] ;
 wire \tokenflow_inst.ii3.i.ydata[12] ;
 wire \tokenflow_inst.ii3.i.ydata[13] ;
 wire \tokenflow_inst.ii3.i.ydata[14] ;
 wire \tokenflow_inst.ii3.i.ydata[15] ;
 wire \tokenflow_inst.ii3.i.ydata[16] ;
 wire \tokenflow_inst.ii3.i.ydata[17] ;
 wire \tokenflow_inst.ii3.i.ydata[18] ;
 wire \tokenflow_inst.ii3.i.ydata[19] ;
 wire \tokenflow_inst.ii3.i.ydata[1] ;
 wire \tokenflow_inst.ii3.i.ydata[20] ;
 wire \tokenflow_inst.ii3.i.ydata[21] ;
 wire \tokenflow_inst.ii3.i.ydata[22] ;
 wire \tokenflow_inst.ii3.i.ydata[23] ;
 wire \tokenflow_inst.ii3.i.ydata[24] ;
 wire \tokenflow_inst.ii3.i.ydata[25] ;
 wire \tokenflow_inst.ii3.i.ydata[2] ;
 wire \tokenflow_inst.ii3.i.ydata[3] ;
 wire \tokenflow_inst.ii3.i.ydata[4] ;
 wire \tokenflow_inst.ii3.i.ydata[5] ;
 wire \tokenflow_inst.ii3.i.ydata[6] ;
 wire \tokenflow_inst.ii3.i.ydata[7] ;
 wire \tokenflow_inst.ii3.i.ydata[8] ;
 wire \tokenflow_inst.ii3.i.ydata[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;

 sg13g2_buf_8 _1497_ (.A(net185),
    .X(_1377_));
 sg13g2_buf_1 _1498_ (.A(_1377_),
    .X(_1378_));
 sg13g2_buf_1 _1499_ (.A(net182),
    .X(_1379_));
 sg13g2_buf_1 _1500_ (.A(net181),
    .X(_1380_));
 sg13g2_and2_1 _1501_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[0] ),
    .X(_0086_));
 sg13g2_and2_1 _1502_ (.A(_1380_),
    .B(\tokenflow_inst.i3.ydata[1] ),
    .X(_0097_));
 sg13g2_and2_1 _1503_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[2] ),
    .X(_0108_));
 sg13g2_and2_1 _1504_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[3] ),
    .X(_0119_));
 sg13g2_and2_1 _1505_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[4] ),
    .X(_0130_));
 sg13g2_and2_1 _1506_ (.A(_1380_),
    .B(\tokenflow_inst.i3.ydata[5] ),
    .X(_0141_));
 sg13g2_and2_1 _1507_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[6] ),
    .X(_0152_));
 sg13g2_and2_1 _1508_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[7] ),
    .X(_0161_));
 sg13g2_and2_1 _1509_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[8] ),
    .X(_0162_));
 sg13g2_and2_1 _1510_ (.A(net175),
    .B(\tokenflow_inst.i3.ydata[9] ),
    .X(_0163_));
 sg13g2_buf_1 _1511_ (.A(net181),
    .X(_1381_));
 sg13g2_and2_1 _1512_ (.A(_1381_),
    .B(\tokenflow_inst.i3.ydata[10] ),
    .X(_0087_));
 sg13g2_and2_1 _1513_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[11] ),
    .X(_0088_));
 sg13g2_and2_1 _1514_ (.A(_1381_),
    .B(\tokenflow_inst.i3.ydata[12] ),
    .X(_0089_));
 sg13g2_and2_1 _1515_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[13] ),
    .X(_0090_));
 sg13g2_and2_1 _1516_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[14] ),
    .X(_0091_));
 sg13g2_and2_1 _1517_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[15] ),
    .X(_0092_));
 sg13g2_and2_1 _1518_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[16] ),
    .X(_0093_));
 sg13g2_and2_1 _1519_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[17] ),
    .X(_0094_));
 sg13g2_and2_1 _1520_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[18] ),
    .X(_0095_));
 sg13g2_and2_1 _1521_ (.A(net174),
    .B(\tokenflow_inst.i3.ydata[19] ),
    .X(_0096_));
 sg13g2_buf_1 _1522_ (.A(_1379_),
    .X(_1382_));
 sg13g2_and2_1 _1523_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[20] ),
    .X(_0098_));
 sg13g2_and2_1 _1524_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[21] ),
    .X(_0099_));
 sg13g2_and2_1 _1525_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[22] ),
    .X(_0100_));
 sg13g2_and2_1 _1526_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[23] ),
    .X(_0101_));
 sg13g2_and2_1 _1527_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[24] ),
    .X(_0102_));
 sg13g2_and2_1 _1528_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[25] ),
    .X(_0103_));
 sg13g2_and2_1 _1529_ (.A(_1382_),
    .B(\tokenflow_inst.i3.ydata[26] ),
    .X(_0104_));
 sg13g2_and2_1 _1530_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[27] ),
    .X(_0105_));
 sg13g2_and2_1 _1531_ (.A(net173),
    .B(\tokenflow_inst.i3.ydata[28] ),
    .X(_0106_));
 sg13g2_and2_1 _1532_ (.A(_1382_),
    .B(\tokenflow_inst.i3.ydata[29] ),
    .X(_0107_));
 sg13g2_buf_1 _1533_ (.A(net181),
    .X(_1383_));
 sg13g2_and2_1 _1534_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[30] ),
    .X(_0109_));
 sg13g2_and2_1 _1535_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[31] ),
    .X(_0110_));
 sg13g2_and2_1 _1536_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[32] ),
    .X(_0111_));
 sg13g2_and2_1 _1537_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[33] ),
    .X(_0112_));
 sg13g2_and2_1 _1538_ (.A(_1383_),
    .B(\tokenflow_inst.i3.ydata[34] ),
    .X(_0113_));
 sg13g2_and2_1 _1539_ (.A(_1383_),
    .B(\tokenflow_inst.i3.ydata[35] ),
    .X(_0114_));
 sg13g2_and2_1 _1540_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[36] ),
    .X(_0115_));
 sg13g2_and2_1 _1541_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[37] ),
    .X(_0116_));
 sg13g2_and2_1 _1542_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[38] ),
    .X(_0117_));
 sg13g2_and2_1 _1543_ (.A(net172),
    .B(\tokenflow_inst.i3.ydata[39] ),
    .X(_0118_));
 sg13g2_buf_1 _1544_ (.A(net181),
    .X(_1384_));
 sg13g2_and2_1 _1545_ (.A(_1384_),
    .B(\tokenflow_inst.i3.ydata[40] ),
    .X(_0120_));
 sg13g2_and2_1 _1546_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[41] ),
    .X(_0121_));
 sg13g2_and2_1 _1547_ (.A(_1384_),
    .B(\tokenflow_inst.i3.ydata[42] ),
    .X(_0122_));
 sg13g2_and2_1 _1548_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[43] ),
    .X(_0123_));
 sg13g2_and2_1 _1549_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[44] ),
    .X(_0124_));
 sg13g2_and2_1 _1550_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[45] ),
    .X(_0125_));
 sg13g2_and2_1 _1551_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[46] ),
    .X(_0126_));
 sg13g2_and2_1 _1552_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[47] ),
    .X(_0127_));
 sg13g2_and2_1 _1553_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[48] ),
    .X(_0128_));
 sg13g2_and2_1 _1554_ (.A(net171),
    .B(\tokenflow_inst.i3.ydata[49] ),
    .X(_0129_));
 sg13g2_buf_1 _1555_ (.A(net181),
    .X(_1385_));
 sg13g2_and2_1 _1556_ (.A(_1385_),
    .B(\tokenflow_inst.i3.ydata[50] ),
    .X(_0131_));
 sg13g2_and2_1 _1557_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[51] ),
    .X(_0132_));
 sg13g2_and2_1 _1558_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[52] ),
    .X(_0133_));
 sg13g2_and2_1 _1559_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[53] ),
    .X(_0134_));
 sg13g2_and2_1 _1560_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[54] ),
    .X(_0135_));
 sg13g2_and2_1 _1561_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[55] ),
    .X(_0136_));
 sg13g2_and2_1 _1562_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[56] ),
    .X(_0137_));
 sg13g2_and2_1 _1563_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[57] ),
    .X(_0138_));
 sg13g2_and2_1 _1564_ (.A(_1385_),
    .B(\tokenflow_inst.i3.ydata[58] ),
    .X(_0139_));
 sg13g2_and2_1 _1565_ (.A(net170),
    .B(\tokenflow_inst.i3.ydata[59] ),
    .X(_0140_));
 sg13g2_buf_1 _1566_ (.A(net182),
    .X(_1386_));
 sg13g2_buf_1 _1567_ (.A(_1386_),
    .X(_1387_));
 sg13g2_and2_1 _1568_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[60] ),
    .X(_0142_));
 sg13g2_and2_1 _1569_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[61] ),
    .X(_0143_));
 sg13g2_and2_1 _1570_ (.A(_1387_),
    .B(\tokenflow_inst.i3.ydata[62] ),
    .X(_0144_));
 sg13g2_and2_1 _1571_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[63] ),
    .X(_0145_));
 sg13g2_and2_1 _1572_ (.A(_1387_),
    .B(\tokenflow_inst.i3.ydata[64] ),
    .X(_0146_));
 sg13g2_and2_1 _1573_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[65] ),
    .X(_0147_));
 sg13g2_and2_1 _1574_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[66] ),
    .X(_0148_));
 sg13g2_and2_1 _1575_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[67] ),
    .X(_0149_));
 sg13g2_and2_1 _1576_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[68] ),
    .X(_0150_));
 sg13g2_and2_1 _1577_ (.A(net169),
    .B(\tokenflow_inst.i3.ydata[69] ),
    .X(_0151_));
 sg13g2_buf_1 _1578_ (.A(net180),
    .X(_1388_));
 sg13g2_and2_1 _1579_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[70] ),
    .X(_0153_));
 sg13g2_and2_1 _1580_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[71] ),
    .X(_0154_));
 sg13g2_and2_1 _1581_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[72] ),
    .X(_0155_));
 sg13g2_and2_1 _1582_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[73] ),
    .X(_0156_));
 sg13g2_and2_1 _1583_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[74] ),
    .X(_0157_));
 sg13g2_and2_1 _1584_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[75] ),
    .X(_0158_));
 sg13g2_and2_1 _1585_ (.A(net168),
    .B(\tokenflow_inst.i3.ydata[76] ),
    .X(_0159_));
 sg13g2_and2_1 _1586_ (.A(_1388_),
    .B(\tokenflow_inst.i3.ydata[77] ),
    .X(_0160_));
 sg13g2_buf_8 _1587_ (.A(\tokenflow_inst.ii2.ydata[0] ),
    .X(_1389_));
 sg13g2_and2_1 _1588_ (.A(net168),
    .B(_1389_),
    .X(\tokenflow_inst.ii3.i.ydata[0] ));
 sg13g2_inv_1 _1589_ (.Y(_1390_),
    .A(_1377_));
 sg13g2_buf_1 _1590_ (.A(_1390_),
    .X(_1391_));
 sg13g2_buf_1 _1591_ (.A(net179),
    .X(_1392_));
 sg13g2_buf_1 _1592_ (.A(net167),
    .X(_1393_));
 sg13g2_buf_1 _1593_ (.A(\tokenflow_inst.i2.cg1.q ),
    .X(_1394_));
 sg13g2_buf_1 _1594_ (.A(_1394_),
    .X(_1395_));
 sg13g2_nor2b_1 _1595_ (.A(net29),
    .B_N(_1389_),
    .Y(_1396_));
 sg13g2_a21oi_1 _1596_ (.A1(\tokenflow_inst.i78.ydata[0] ),
    .A2(net29),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_nor2_1 _1597_ (.A(net154),
    .B(_1397_),
    .Y(_0007_));
 sg13g2_buf_8 _1598_ (.A(\tokenflow_inst.ii2.ydata[1] ),
    .X(_1398_));
 sg13g2_and2_1 _1599_ (.A(_1388_),
    .B(_1398_),
    .X(\tokenflow_inst.ii3.i.ydata[1] ));
 sg13g2_buf_1 _1600_ (.A(_1394_),
    .X(_1399_));
 sg13g2_buf_1 _1601_ (.A(net28),
    .X(_1400_));
 sg13g2_nor2b_1 _1602_ (.A(_1395_),
    .B_N(_1398_),
    .Y(_1401_));
 sg13g2_a21oi_1 _1603_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[1] ),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_nor2_1 _1604_ (.A(net154),
    .B(_1402_),
    .Y(_0018_));
 sg13g2_buf_1 _1605_ (.A(net180),
    .X(_1403_));
 sg13g2_buf_8 _1606_ (.A(\tokenflow_inst.ii2.ydata[2] ),
    .X(_1404_));
 sg13g2_and2_1 _1607_ (.A(net166),
    .B(_1404_),
    .X(\tokenflow_inst.ii3.i.ydata[2] ));
 sg13g2_nor2b_1 _1608_ (.A(_1399_),
    .B_N(_1404_),
    .Y(_1405_));
 sg13g2_a21oi_1 _1609_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[2] ),
    .Y(_1406_),
    .B1(_1405_));
 sg13g2_nor2_1 _1610_ (.A(net154),
    .B(_1406_),
    .Y(_0029_));
 sg13g2_and2_1 _1611_ (.A(net166),
    .B(\tokenflow_inst.ii2.ydata[3] ),
    .X(\tokenflow_inst.ii3.i.ydata[3] ));
 sg13g2_buf_1 _1612_ (.A(_1394_),
    .X(_1407_));
 sg13g2_nor2b_1 _1613_ (.A(net27),
    .B_N(\tokenflow_inst.ii2.ydata[3] ),
    .Y(_1408_));
 sg13g2_a21oi_1 _1614_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[3] ),
    .Y(_1409_),
    .B1(_1408_));
 sg13g2_nor2_1 _1615_ (.A(_1393_),
    .B(_1409_),
    .Y(_0040_));
 sg13g2_and2_1 _1616_ (.A(_1377_),
    .B(\tokenflow_inst.ii2.ydata[4] ),
    .X(_1410_));
 sg13g2_buf_1 _1617_ (.A(_1410_),
    .X(\tokenflow_inst.ii3.i.ydata[4] ));
 sg13g2_nor2b_1 _1618_ (.A(net27),
    .B_N(\tokenflow_inst.ii2.ydata[4] ),
    .Y(_1411_));
 sg13g2_a21oi_1 _1619_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[4] ),
    .Y(_1412_),
    .B1(_1411_));
 sg13g2_nor2_1 _1620_ (.A(_1393_),
    .B(_1412_),
    .Y(_0051_));
 sg13g2_buf_2 _1621_ (.A(\tokenflow_inst.ii2.ydata[5] ),
    .X(_1413_));
 sg13g2_and2_1 _1622_ (.A(net166),
    .B(_1413_),
    .X(\tokenflow_inst.ii3.i.ydata[5] ));
 sg13g2_nor2b_1 _1623_ (.A(net27),
    .B_N(_1413_),
    .Y(_1414_));
 sg13g2_a21oi_1 _1624_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[5] ),
    .Y(_1415_),
    .B1(_1414_));
 sg13g2_nor2_1 _1625_ (.A(net154),
    .B(_1415_),
    .Y(_0062_));
 sg13g2_and2_1 _1626_ (.A(_1377_),
    .B(\tokenflow_inst.ii2.ydata[6] ),
    .X(_1416_));
 sg13g2_buf_1 _1627_ (.A(_1416_),
    .X(\tokenflow_inst.ii3.i.ydata[6] ));
 sg13g2_nor2b_1 _1628_ (.A(_1407_),
    .B_N(\tokenflow_inst.ii2.ydata[6] ),
    .Y(_1417_));
 sg13g2_a21oi_1 _1629_ (.A1(_1400_),
    .A2(\tokenflow_inst.i78.ydata[6] ),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_nor2_1 _1630_ (.A(net154),
    .B(_1418_),
    .Y(_0073_));
 sg13g2_buf_1 _1631_ (.A(\tokenflow_inst.ii2.ydata[7] ),
    .X(_1419_));
 sg13g2_and2_1 _1632_ (.A(_1403_),
    .B(_1419_),
    .X(\tokenflow_inst.ii3.i.ydata[7] ));
 sg13g2_nor2b_1 _1633_ (.A(_1407_),
    .B_N(_1419_),
    .Y(_1420_));
 sg13g2_a21oi_1 _1634_ (.A1(_1400_),
    .A2(\tokenflow_inst.i78.ydata[7] ),
    .Y(_1421_),
    .B1(_1420_));
 sg13g2_nor2_1 _1635_ (.A(net154),
    .B(_1421_),
    .Y(_0082_));
 sg13g2_and2_1 _1636_ (.A(_1403_),
    .B(\tokenflow_inst.ii2.ydata[8] ),
    .X(\tokenflow_inst.ii3.i.ydata[8] ));
 sg13g2_nor2b_1 _1637_ (.A(net27),
    .B_N(\tokenflow_inst.ii2.ydata[8] ),
    .Y(_1422_));
 sg13g2_a21oi_1 _1638_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[8] ),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_nor2_1 _1639_ (.A(net154),
    .B(_1423_),
    .Y(_0083_));
 sg13g2_and2_1 _1640_ (.A(_1377_),
    .B(\tokenflow_inst.ii2.ydata[9] ),
    .X(_1424_));
 sg13g2_buf_1 _1641_ (.A(_1424_),
    .X(\tokenflow_inst.ii3.i.ydata[9] ));
 sg13g2_nor2b_1 _1642_ (.A(net27),
    .B_N(\tokenflow_inst.ii2.ydata[9] ),
    .Y(_1425_));
 sg13g2_a21oi_1 _1643_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[9] ),
    .Y(_1426_),
    .B1(_1425_));
 sg13g2_nor2_1 _1644_ (.A(net154),
    .B(_1426_),
    .Y(_0084_));
 sg13g2_buf_1 _1645_ (.A(\tokenflow_inst.ii2.ydata[10] ),
    .X(_1427_));
 sg13g2_and2_1 _1646_ (.A(net166),
    .B(_1427_),
    .X(\tokenflow_inst.ii3.i.ydata[10] ));
 sg13g2_buf_1 _1647_ (.A(net167),
    .X(_1428_));
 sg13g2_nor2b_1 _1648_ (.A(net27),
    .B_N(_1427_),
    .Y(_1429_));
 sg13g2_a21oi_1 _1649_ (.A1(net25),
    .A2(\tokenflow_inst.i78.ydata[10] ),
    .Y(_1430_),
    .B1(_1429_));
 sg13g2_nor2_1 _1650_ (.A(net153),
    .B(_1430_),
    .Y(_0008_));
 sg13g2_inv_1 _1651_ (.Y(_1431_),
    .A(\tokenflow_inst.ii2.ydata[11] ));
 sg13g2_nor2_1 _1652_ (.A(net153),
    .B(_1431_),
    .Y(\tokenflow_inst.ii3.i.ydata[11] ));
 sg13g2_buf_1 _1653_ (.A(net28),
    .X(_1432_));
 sg13g2_nor2_1 _1654_ (.A(net28),
    .B(_1431_),
    .Y(_1433_));
 sg13g2_a21oi_1 _1655_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[11] ),
    .Y(_1434_),
    .B1(_1433_));
 sg13g2_nor2_1 _1656_ (.A(net153),
    .B(_1434_),
    .Y(_0009_));
 sg13g2_buf_1 _1657_ (.A(\tokenflow_inst.ii2.ydata[12] ),
    .X(_1435_));
 sg13g2_and2_1 _1658_ (.A(net166),
    .B(_1435_),
    .X(\tokenflow_inst.ii3.i.ydata[12] ));
 sg13g2_nor2b_1 _1659_ (.A(net27),
    .B_N(_1435_),
    .Y(_1436_));
 sg13g2_a21oi_1 _1660_ (.A1(_1432_),
    .A2(\tokenflow_inst.i78.ydata[12] ),
    .Y(_1437_),
    .B1(_1436_));
 sg13g2_nor2_1 _1661_ (.A(_1428_),
    .B(_1437_),
    .Y(_0010_));
 sg13g2_and2_1 _1662_ (.A(net182),
    .B(\tokenflow_inst.ii2.ydata[13] ),
    .X(\tokenflow_inst.ii3.i.ydata[13] ));
 sg13g2_nor2b_1 _1663_ (.A(net27),
    .B_N(\tokenflow_inst.ii2.ydata[13] ),
    .Y(_1438_));
 sg13g2_a21oi_1 _1664_ (.A1(_1432_),
    .A2(\tokenflow_inst.i78.ydata[13] ),
    .Y(_1439_),
    .B1(_1438_));
 sg13g2_nor2_1 _1665_ (.A(_1428_),
    .B(_1439_),
    .Y(_0011_));
 sg13g2_buf_2 _1666_ (.A(\tokenflow_inst.ii2.ydata[14] ),
    .X(_1440_));
 sg13g2_and2_1 _1667_ (.A(net166),
    .B(_1440_),
    .X(\tokenflow_inst.ii3.i.ydata[14] ));
 sg13g2_buf_1 _1668_ (.A(_1394_),
    .X(_1441_));
 sg13g2_nor2b_1 _1669_ (.A(_1441_),
    .B_N(_1440_),
    .Y(_1442_));
 sg13g2_a21oi_1 _1670_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[14] ),
    .Y(_1443_),
    .B1(_1442_));
 sg13g2_nor2_1 _1671_ (.A(net153),
    .B(_1443_),
    .Y(_0012_));
 sg13g2_and2_1 _1672_ (.A(net166),
    .B(\tokenflow_inst.ii2.ydata[15] ),
    .X(\tokenflow_inst.ii3.i.ydata[15] ));
 sg13g2_nor2b_1 _1673_ (.A(net26),
    .B_N(\tokenflow_inst.ii2.ydata[15] ),
    .Y(_1444_));
 sg13g2_a21oi_1 _1674_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[15] ),
    .Y(_1445_),
    .B1(_1444_));
 sg13g2_nor2_1 _1675_ (.A(net153),
    .B(_1445_),
    .Y(_0013_));
 sg13g2_buf_2 _1676_ (.A(\tokenflow_inst.ii2.ydata[16] ),
    .X(_1446_));
 sg13g2_and2_1 _1677_ (.A(net166),
    .B(_1446_),
    .X(\tokenflow_inst.ii3.i.ydata[16] ));
 sg13g2_nor2b_1 _1678_ (.A(net26),
    .B_N(_1446_),
    .Y(_1447_));
 sg13g2_a21oi_1 _1679_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[16] ),
    .Y(_1448_),
    .B1(_1447_));
 sg13g2_nor2_1 _1680_ (.A(net153),
    .B(_1448_),
    .Y(_0014_));
 sg13g2_buf_1 _1681_ (.A(net180),
    .X(_1449_));
 sg13g2_buf_2 _1682_ (.A(\tokenflow_inst.ii2.ydata[17] ),
    .X(_1450_));
 sg13g2_and2_1 _1683_ (.A(net165),
    .B(_1450_),
    .X(\tokenflow_inst.ii3.i.ydata[17] ));
 sg13g2_nor2b_1 _1684_ (.A(net26),
    .B_N(_1450_),
    .Y(_1451_));
 sg13g2_a21oi_1 _1685_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[17] ),
    .Y(_1452_),
    .B1(_1451_));
 sg13g2_nor2_1 _1686_ (.A(net153),
    .B(_1452_),
    .Y(_0015_));
 sg13g2_and2_1 _1687_ (.A(net165),
    .B(\tokenflow_inst.ii2.ydata[18] ),
    .X(\tokenflow_inst.ii3.i.ydata[18] ));
 sg13g2_nor2b_1 _1688_ (.A(net26),
    .B_N(\tokenflow_inst.ii2.ydata[18] ),
    .Y(_1453_));
 sg13g2_a21oi_1 _1689_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[18] ),
    .Y(_1454_),
    .B1(_1453_));
 sg13g2_nor2_1 _1690_ (.A(net153),
    .B(_1454_),
    .Y(_0016_));
 sg13g2_buf_2 _1691_ (.A(\tokenflow_inst.ii2.ydata[19] ),
    .X(_1455_));
 sg13g2_and2_1 _1692_ (.A(net165),
    .B(_1455_),
    .X(\tokenflow_inst.ii3.i.ydata[19] ));
 sg13g2_buf_1 _1693_ (.A(_1391_),
    .X(_1456_));
 sg13g2_buf_1 _1694_ (.A(net164),
    .X(_1457_));
 sg13g2_nor2b_1 _1695_ (.A(net26),
    .B_N(_1455_),
    .Y(_1458_));
 sg13g2_a21oi_1 _1696_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[19] ),
    .Y(_1459_),
    .B1(_1458_));
 sg13g2_nor2_1 _1697_ (.A(net152),
    .B(_1459_),
    .Y(_0017_));
 sg13g2_buf_2 _1698_ (.A(\tokenflow_inst.ii2.ydata[20] ),
    .X(_1460_));
 sg13g2_and2_1 _1699_ (.A(net165),
    .B(_1460_),
    .X(\tokenflow_inst.ii3.i.ydata[20] ));
 sg13g2_nor2b_1 _1700_ (.A(net26),
    .B_N(_1460_),
    .Y(_1461_));
 sg13g2_a21oi_1 _1701_ (.A1(net24),
    .A2(\tokenflow_inst.i78.ydata[20] ),
    .Y(_1462_),
    .B1(_1461_));
 sg13g2_nor2_1 _1702_ (.A(net152),
    .B(_1462_),
    .Y(_0019_));
 sg13g2_and2_1 _1703_ (.A(_1377_),
    .B(\tokenflow_inst.ii2.ydata[21] ),
    .X(_1463_));
 sg13g2_buf_1 _1704_ (.A(_1463_),
    .X(\tokenflow_inst.ii3.i.ydata[21] ));
 sg13g2_buf_1 _1705_ (.A(net28),
    .X(_1464_));
 sg13g2_nor2b_1 _1706_ (.A(_1441_),
    .B_N(\tokenflow_inst.ii2.ydata[21] ),
    .Y(_1465_));
 sg13g2_a21oi_1 _1707_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[21] ),
    .Y(_1466_),
    .B1(_1465_));
 sg13g2_nor2_1 _1708_ (.A(net152),
    .B(_1466_),
    .Y(_0020_));
 sg13g2_buf_1 _1709_ (.A(\tokenflow_inst.ii2.ydata[22] ),
    .X(_1467_));
 sg13g2_and2_1 _1710_ (.A(net165),
    .B(_1467_),
    .X(\tokenflow_inst.ii3.i.ydata[22] ));
 sg13g2_nor2b_1 _1711_ (.A(net26),
    .B_N(_1467_),
    .Y(_1468_));
 sg13g2_a21oi_1 _1712_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[22] ),
    .Y(_1469_),
    .B1(_1468_));
 sg13g2_nor2_1 _1713_ (.A(net152),
    .B(_1469_),
    .Y(_0021_));
 sg13g2_and2_1 _1714_ (.A(net165),
    .B(\tokenflow_inst.ii2.ydata[23] ),
    .X(\tokenflow_inst.ii3.i.ydata[23] ));
 sg13g2_nor2b_1 _1715_ (.A(net26),
    .B_N(\tokenflow_inst.ii2.ydata[23] ),
    .Y(_1470_));
 sg13g2_a21oi_1 _1716_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[23] ),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_nor2_1 _1717_ (.A(net152),
    .B(_1471_),
    .Y(_0022_));
 sg13g2_buf_2 _1718_ (.A(\tokenflow_inst.ii2.ydata[24] ),
    .X(_1472_));
 sg13g2_and2_1 _1719_ (.A(net165),
    .B(_1472_),
    .X(\tokenflow_inst.ii3.i.ydata[24] ));
 sg13g2_nor2b_1 _1720_ (.A(net29),
    .B_N(_1472_),
    .Y(_1473_));
 sg13g2_a21oi_1 _1721_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[24] ),
    .Y(_1474_),
    .B1(_1473_));
 sg13g2_nor2_1 _1722_ (.A(net152),
    .B(_1474_),
    .Y(_0023_));
 sg13g2_and2_1 _1723_ (.A(net165),
    .B(\tokenflow_inst.ii2.ydata[25] ),
    .X(\tokenflow_inst.ii3.i.ydata[25] ));
 sg13g2_nor2b_1 _1724_ (.A(net29),
    .B_N(\tokenflow_inst.ii2.ydata[25] ),
    .Y(_1475_));
 sg13g2_a21oi_1 _1725_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[25] ),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_nor2_1 _1726_ (.A(_1457_),
    .B(_1476_),
    .Y(_0024_));
 sg13g2_a21oi_1 _1727_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[26] ),
    .Y(_1477_),
    .B1(_1396_));
 sg13g2_nor2_1 _1728_ (.A(net152),
    .B(_1477_),
    .Y(_0025_));
 sg13g2_a21oi_1 _1729_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[27] ),
    .Y(_1478_),
    .B1(_1401_));
 sg13g2_nor2_1 _1730_ (.A(net152),
    .B(_1478_),
    .Y(_0026_));
 sg13g2_a21oi_1 _1731_ (.A1(net23),
    .A2(\tokenflow_inst.i78.ydata[28] ),
    .Y(_1479_),
    .B1(_1405_));
 sg13g2_nor2_1 _1732_ (.A(_1457_),
    .B(_1479_),
    .Y(_0027_));
 sg13g2_buf_1 _1733_ (.A(net164),
    .X(_1480_));
 sg13g2_a21oi_1 _1734_ (.A1(_1464_),
    .A2(\tokenflow_inst.i78.ydata[29] ),
    .Y(_1481_),
    .B1(_1408_));
 sg13g2_nor2_1 _1735_ (.A(net151),
    .B(_1481_),
    .Y(_0028_));
 sg13g2_a21oi_1 _1736_ (.A1(_1464_),
    .A2(\tokenflow_inst.i78.ydata[30] ),
    .Y(_1482_),
    .B1(_1411_));
 sg13g2_nor2_1 _1737_ (.A(net151),
    .B(_1482_),
    .Y(_0030_));
 sg13g2_buf_1 _1738_ (.A(_1399_),
    .X(_1483_));
 sg13g2_a21oi_1 _1739_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[31] ),
    .Y(_1484_),
    .B1(_1414_));
 sg13g2_nor2_1 _1740_ (.A(net151),
    .B(_1484_),
    .Y(_0031_));
 sg13g2_a21oi_1 _1741_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[32] ),
    .Y(_1485_),
    .B1(_1417_));
 sg13g2_nor2_1 _1742_ (.A(net151),
    .B(_1485_),
    .Y(_0032_));
 sg13g2_a21oi_1 _1743_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[33] ),
    .Y(_1486_),
    .B1(_1420_));
 sg13g2_nor2_1 _1744_ (.A(_1480_),
    .B(_1486_),
    .Y(_0033_));
 sg13g2_a21oi_1 _1745_ (.A1(_1483_),
    .A2(\tokenflow_inst.i78.ydata[34] ),
    .Y(_1487_),
    .B1(_1422_));
 sg13g2_nor2_1 _1746_ (.A(_1480_),
    .B(_1487_),
    .Y(_0034_));
 sg13g2_a21oi_1 _1747_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[35] ),
    .Y(_1488_),
    .B1(_1425_));
 sg13g2_nor2_1 _1748_ (.A(net151),
    .B(_1488_),
    .Y(_0035_));
 sg13g2_a21oi_1 _1749_ (.A1(_1483_),
    .A2(\tokenflow_inst.i78.ydata[36] ),
    .Y(_1489_),
    .B1(_1429_));
 sg13g2_nor2_1 _1750_ (.A(net151),
    .B(_1489_),
    .Y(_0036_));
 sg13g2_a21oi_1 _1751_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[37] ),
    .Y(_1490_),
    .B1(_1433_));
 sg13g2_nor2_1 _1752_ (.A(net151),
    .B(_1490_),
    .Y(_0037_));
 sg13g2_a21oi_1 _1753_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[38] ),
    .Y(_1491_),
    .B1(_1436_));
 sg13g2_nor2_1 _1754_ (.A(net151),
    .B(_1491_),
    .Y(_0038_));
 sg13g2_buf_1 _1755_ (.A(net164),
    .X(_1492_));
 sg13g2_a21oi_1 _1756_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[39] ),
    .Y(_1493_),
    .B1(_1438_));
 sg13g2_nor2_1 _1757_ (.A(_1492_),
    .B(_1493_),
    .Y(_0039_));
 sg13g2_a21oi_1 _1758_ (.A1(net22),
    .A2(\tokenflow_inst.i78.ydata[40] ),
    .Y(_1494_),
    .B1(_1442_));
 sg13g2_nor2_1 _1759_ (.A(_1492_),
    .B(_1494_),
    .Y(_0041_));
 sg13g2_buf_1 _1760_ (.A(net28),
    .X(_0317_));
 sg13g2_a21oi_1 _1761_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[41] ),
    .Y(_0318_),
    .B1(_1444_));
 sg13g2_nor2_1 _1762_ (.A(net150),
    .B(_0318_),
    .Y(_0042_));
 sg13g2_a21oi_1 _1763_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[42] ),
    .Y(_0319_),
    .B1(_1447_));
 sg13g2_nor2_1 _1764_ (.A(net150),
    .B(_0319_),
    .Y(_0043_));
 sg13g2_a21oi_1 _1765_ (.A1(_0317_),
    .A2(\tokenflow_inst.i78.ydata[43] ),
    .Y(_0320_),
    .B1(_1451_));
 sg13g2_nor2_1 _1766_ (.A(net150),
    .B(_0320_),
    .Y(_0044_));
 sg13g2_a21oi_1 _1767_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[44] ),
    .Y(_0321_),
    .B1(_1453_));
 sg13g2_nor2_1 _1768_ (.A(net150),
    .B(_0321_),
    .Y(_0045_));
 sg13g2_a21oi_1 _1769_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[45] ),
    .Y(_0322_),
    .B1(_1458_));
 sg13g2_nor2_1 _1770_ (.A(net150),
    .B(_0322_),
    .Y(_0046_));
 sg13g2_a21oi_1 _1771_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[46] ),
    .Y(_0323_),
    .B1(_1461_));
 sg13g2_nor2_1 _1772_ (.A(net150),
    .B(_0323_),
    .Y(_0047_));
 sg13g2_a21oi_1 _1773_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[47] ),
    .Y(_0324_),
    .B1(_1465_));
 sg13g2_nor2_1 _1774_ (.A(net150),
    .B(_0324_),
    .Y(_0048_));
 sg13g2_a21oi_1 _1775_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[48] ),
    .Y(_0325_),
    .B1(_1468_));
 sg13g2_nor2_1 _1776_ (.A(net150),
    .B(_0325_),
    .Y(_0049_));
 sg13g2_buf_1 _1777_ (.A(net164),
    .X(_0326_));
 sg13g2_a21oi_1 _1778_ (.A1(net21),
    .A2(\tokenflow_inst.i78.ydata[49] ),
    .Y(_0327_),
    .B1(_1470_));
 sg13g2_nor2_1 _1779_ (.A(_0326_),
    .B(_0327_),
    .Y(_0050_));
 sg13g2_nor2_1 _1780_ (.A(net179),
    .B(net29),
    .Y(_0328_));
 sg13g2_and2_1 _1781_ (.A(_1472_),
    .B(_0328_),
    .X(_0052_));
 sg13g2_and2_1 _1782_ (.A(\tokenflow_inst.ii2.ydata[25] ),
    .B(_0328_),
    .X(_0053_));
 sg13g2_and2_1 _1783_ (.A(_1389_),
    .B(_0328_),
    .X(_0054_));
 sg13g2_and2_1 _1784_ (.A(_1398_),
    .B(_0328_),
    .X(_0055_));
 sg13g2_a21oi_1 _1785_ (.A1(_0317_),
    .A2(\tokenflow_inst.i78.ydata[54] ),
    .Y(_0329_),
    .B1(_1405_));
 sg13g2_nor2_1 _1786_ (.A(net149),
    .B(_0329_),
    .Y(_0056_));
 sg13g2_buf_1 _1787_ (.A(net28),
    .X(_0330_));
 sg13g2_a21oi_1 _1788_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[55] ),
    .Y(_0331_),
    .B1(_1408_));
 sg13g2_nor2_1 _1789_ (.A(net149),
    .B(_0331_),
    .Y(_0057_));
 sg13g2_a21oi_1 _1790_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[56] ),
    .Y(_0332_),
    .B1(_1411_));
 sg13g2_nor2_1 _1791_ (.A(net149),
    .B(_0332_),
    .Y(_0058_));
 sg13g2_a21oi_1 _1792_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[57] ),
    .Y(_0333_),
    .B1(_1414_));
 sg13g2_nor2_1 _1793_ (.A(net149),
    .B(_0333_),
    .Y(_0059_));
 sg13g2_a21oi_1 _1794_ (.A1(_0330_),
    .A2(\tokenflow_inst.i78.ydata[58] ),
    .Y(_0334_),
    .B1(_1417_));
 sg13g2_nor2_1 _1795_ (.A(net149),
    .B(_0334_),
    .Y(_0060_));
 sg13g2_a21oi_1 _1796_ (.A1(_0330_),
    .A2(\tokenflow_inst.i78.ydata[59] ),
    .Y(_0335_),
    .B1(_1420_));
 sg13g2_nor2_1 _1797_ (.A(_0326_),
    .B(_0335_),
    .Y(_0061_));
 sg13g2_a21oi_1 _1798_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[60] ),
    .Y(_0336_),
    .B1(_1422_));
 sg13g2_nor2_1 _1799_ (.A(net149),
    .B(_0336_),
    .Y(_0063_));
 sg13g2_a21oi_1 _1800_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[61] ),
    .Y(_0337_),
    .B1(_1425_));
 sg13g2_nor2_1 _1801_ (.A(net149),
    .B(_0337_),
    .Y(_0064_));
 sg13g2_a21oi_1 _1802_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[62] ),
    .Y(_0338_),
    .B1(_1429_));
 sg13g2_nor2_1 _1803_ (.A(net149),
    .B(_0338_),
    .Y(_0065_));
 sg13g2_buf_1 _1804_ (.A(_1456_),
    .X(_0339_));
 sg13g2_a21oi_1 _1805_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[63] ),
    .Y(_0340_),
    .B1(_1433_));
 sg13g2_nor2_1 _1806_ (.A(net148),
    .B(_0340_),
    .Y(_0066_));
 sg13g2_a21oi_1 _1807_ (.A1(net20),
    .A2(\tokenflow_inst.i78.ydata[64] ),
    .Y(_0341_),
    .B1(_1436_));
 sg13g2_nor2_1 _1808_ (.A(_0339_),
    .B(_0341_),
    .Y(_0067_));
 sg13g2_buf_1 _1809_ (.A(net28),
    .X(_0342_));
 sg13g2_a21oi_1 _1810_ (.A1(_0342_),
    .A2(\tokenflow_inst.i78.ydata[65] ),
    .Y(_0343_),
    .B1(_1438_));
 sg13g2_nor2_1 _1811_ (.A(_0339_),
    .B(_0343_),
    .Y(_0068_));
 sg13g2_a21oi_1 _1812_ (.A1(_0342_),
    .A2(\tokenflow_inst.i78.ydata[66] ),
    .Y(_0344_),
    .B1(_1442_));
 sg13g2_nor2_1 _1813_ (.A(net148),
    .B(_0344_),
    .Y(_0069_));
 sg13g2_a21oi_1 _1814_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[67] ),
    .Y(_0345_),
    .B1(_1444_));
 sg13g2_nor2_1 _1815_ (.A(net148),
    .B(_0345_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1816_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[68] ),
    .Y(_0346_),
    .B1(_1447_));
 sg13g2_nor2_1 _1817_ (.A(net148),
    .B(_0346_),
    .Y(_0071_));
 sg13g2_a21oi_1 _1818_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[69] ),
    .Y(_0347_),
    .B1(_1451_));
 sg13g2_nor2_1 _1819_ (.A(net148),
    .B(_0347_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1820_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[70] ),
    .Y(_0348_),
    .B1(_1453_));
 sg13g2_nor2_1 _1821_ (.A(net148),
    .B(_0348_),
    .Y(_0074_));
 sg13g2_a21oi_1 _1822_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[71] ),
    .Y(_0349_),
    .B1(_1458_));
 sg13g2_nor2_1 _1823_ (.A(net148),
    .B(_0349_),
    .Y(_0075_));
 sg13g2_a21oi_1 _1824_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[72] ),
    .Y(_0350_),
    .B1(_1461_));
 sg13g2_nor2_1 _1825_ (.A(net148),
    .B(_0350_),
    .Y(_0076_));
 sg13g2_buf_1 _1826_ (.A(net164),
    .X(_0351_));
 sg13g2_a21oi_1 _1827_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[73] ),
    .Y(_0352_),
    .B1(_1465_));
 sg13g2_nor2_1 _1828_ (.A(net147),
    .B(_0352_),
    .Y(_0077_));
 sg13g2_a21oi_1 _1829_ (.A1(net19),
    .A2(\tokenflow_inst.i78.ydata[74] ),
    .Y(_0353_),
    .B1(_1468_));
 sg13g2_nor2_1 _1830_ (.A(net147),
    .B(_0353_),
    .Y(_0078_));
 sg13g2_a21oi_1 _1831_ (.A1(net29),
    .A2(\tokenflow_inst.i78.ydata[75] ),
    .Y(_0354_),
    .B1(_1470_));
 sg13g2_nor2_1 _1832_ (.A(net147),
    .B(_0354_),
    .Y(_0079_));
 sg13g2_a21oi_1 _1833_ (.A1(net29),
    .A2(\tokenflow_inst.i78.ydata[76] ),
    .Y(_0355_),
    .B1(_1473_));
 sg13g2_nor2_1 _1834_ (.A(net147),
    .B(_0355_),
    .Y(_0080_));
 sg13g2_a21oi_1 _1835_ (.A1(net29),
    .A2(\tokenflow_inst.i78.ydata[77] ),
    .Y(_0356_),
    .B1(_1475_));
 sg13g2_nor2_1 _1836_ (.A(net147),
    .B(_0356_),
    .Y(_0081_));
 sg13g2_buf_1 _1837_ (.A(\tokenflow_inst.i6.ydata[26] ),
    .X(_0357_));
 sg13g2_buf_1 _1838_ (.A(_0357_),
    .X(_0358_));
 sg13g2_buf_1 _1839_ (.A(_0358_),
    .X(_0359_));
 sg13g2_buf_1 _1840_ (.A(net90),
    .X(_0360_));
 sg13g2_buf_1 _1841_ (.A(_0360_),
    .X(_0361_));
 sg13g2_buf_1 _1842_ (.A(_0361_),
    .X(_0362_));
 sg13g2_nand2_1 _1843_ (.Y(_0363_),
    .A(net84),
    .B(\tokenflow_inst.i6.ydata[52] ));
 sg13g2_xor2_1 _1844_ (.B(_0363_),
    .A(\tokenflow_inst.i6.ydata[0] ),
    .X(_0364_));
 sg13g2_nor2_1 _1845_ (.A(net147),
    .B(_0364_),
    .Y(_0240_));
 sg13g2_buf_2 _1846_ (.A(\tokenflow_inst.i6.ydata[53] ),
    .X(_0365_));
 sg13g2_nand2_1 _1847_ (.Y(_0366_),
    .A(\tokenflow_inst.i6.ydata[52] ),
    .B(\tokenflow_inst.i6.ydata[0] ));
 sg13g2_xnor2_1 _1848_ (.Y(_0367_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_nand2_1 _1849_ (.Y(_0368_),
    .A(net84),
    .B(_0367_));
 sg13g2_xor2_1 _1850_ (.B(_0368_),
    .A(\tokenflow_inst.i6.ydata[1] ),
    .X(_0369_));
 sg13g2_nor2_1 _1851_ (.A(net147),
    .B(_0369_),
    .Y(_0251_));
 sg13g2_nor2_1 _1852_ (.A(_0365_),
    .B(\tokenflow_inst.i6.ydata[1] ),
    .Y(_0370_));
 sg13g2_a22oi_1 _1853_ (.Y(_0371_),
    .B1(_0365_),
    .B2(\tokenflow_inst.i6.ydata[1] ),
    .A2(\tokenflow_inst.i6.ydata[0] ),
    .A1(\tokenflow_inst.i6.ydata[52] ));
 sg13g2_nor2_1 _1854_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_xor2_1 _1855_ (.B(_0372_),
    .A(\tokenflow_inst.i6.ydata[54] ),
    .X(_0373_));
 sg13g2_nand2_1 _1856_ (.Y(_0374_),
    .A(_0362_),
    .B(_0373_));
 sg13g2_xor2_1 _1857_ (.B(_0374_),
    .A(\tokenflow_inst.i6.ydata[2] ),
    .X(_0375_));
 sg13g2_nor2_1 _1858_ (.A(net147),
    .B(_0375_),
    .Y(_0262_));
 sg13g2_buf_1 _1859_ (.A(\tokenflow_inst.i6.ydata[3] ),
    .X(_0376_));
 sg13g2_inv_1 _1860_ (.Y(_0377_),
    .A(net92));
 sg13g2_buf_1 _1861_ (.A(_0377_),
    .X(_0378_));
 sg13g2_buf_1 _1862_ (.A(net87),
    .X(_0379_));
 sg13g2_buf_1 _1863_ (.A(net85),
    .X(_0380_));
 sg13g2_buf_1 _1864_ (.A(\tokenflow_inst.i6.ydata[55] ),
    .X(_0381_));
 sg13g2_nand2_1 _1865_ (.Y(_0382_),
    .A(\tokenflow_inst.i6.ydata[54] ),
    .B(\tokenflow_inst.i6.ydata[2] ));
 sg13g2_o21ai_1 _1866_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0370_),
    .A2(_0371_));
 sg13g2_or2_1 _1867_ (.X(_0384_),
    .B(\tokenflow_inst.i6.ydata[2] ),
    .A(\tokenflow_inst.i6.ydata[54] ));
 sg13g2_buf_1 _1868_ (.A(_0384_),
    .X(_0385_));
 sg13g2_nand2_1 _1869_ (.Y(_0386_),
    .A(_0383_),
    .B(_0385_));
 sg13g2_xor2_1 _1870_ (.B(_0386_),
    .A(_0381_),
    .X(_0387_));
 sg13g2_nor2_1 _1871_ (.A(net83),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_xnor2_1 _1872_ (.Y(_0389_),
    .A(_0376_),
    .B(_0388_));
 sg13g2_nor2_1 _1873_ (.A(_0351_),
    .B(_0389_),
    .Y(_0273_));
 sg13g2_buf_1 _1874_ (.A(\tokenflow_inst.i6.ydata[4] ),
    .X(_0390_));
 sg13g2_buf_2 _1875_ (.A(\tokenflow_inst.i6.ydata[56] ),
    .X(_0391_));
 sg13g2_or2_1 _1876_ (.X(_0392_),
    .B(_0376_),
    .A(_0381_));
 sg13g2_nand3_1 _1877_ (.B(_0385_),
    .C(_0392_),
    .A(_0383_),
    .Y(_0393_));
 sg13g2_nand2_1 _1878_ (.Y(_0394_),
    .A(_0381_),
    .B(_0376_));
 sg13g2_and2_1 _1879_ (.A(_0393_),
    .B(_0394_),
    .X(_0395_));
 sg13g2_buf_1 _1880_ (.A(_0395_),
    .X(_0396_));
 sg13g2_xor2_1 _1881_ (.B(_0396_),
    .A(_0391_),
    .X(_0397_));
 sg13g2_nor2_1 _1882_ (.A(_0380_),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_xnor2_1 _1883_ (.Y(_0399_),
    .A(_0390_),
    .B(_0398_));
 sg13g2_nor2_1 _1884_ (.A(_0351_),
    .B(_0399_),
    .Y(_0284_));
 sg13g2_buf_1 _1885_ (.A(net164),
    .X(_0400_));
 sg13g2_or2_1 _1886_ (.X(_0401_),
    .B(_0390_),
    .A(_0391_));
 sg13g2_nand3_1 _1887_ (.B(_0392_),
    .C(_0401_),
    .A(net92),
    .Y(_0402_));
 sg13g2_nand3b_1 _1888_ (.B(_0385_),
    .C(_0383_),
    .Y(_0403_),
    .A_N(_0402_));
 sg13g2_inv_1 _1889_ (.Y(_0404_),
    .A(_0390_));
 sg13g2_a21oi_1 _1890_ (.A1(_0381_),
    .A2(_0376_),
    .Y(_0405_),
    .B1(_0391_));
 sg13g2_nand3_1 _1891_ (.B(_0376_),
    .C(_0391_),
    .A(_0381_),
    .Y(_0406_));
 sg13g2_o21ai_1 _1892_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_0404_),
    .A2(_0405_));
 sg13g2_nand2_1 _1893_ (.Y(_0408_),
    .A(net92),
    .B(_0407_));
 sg13g2_nand2_1 _1894_ (.Y(_0409_),
    .A(_0403_),
    .B(_0408_));
 sg13g2_buf_2 _1895_ (.A(\tokenflow_inst.i6.ydata[5] ),
    .X(_0410_));
 sg13g2_buf_1 _1896_ (.A(net86),
    .X(_0411_));
 sg13g2_buf_2 _1897_ (.A(\tokenflow_inst.i6.ydata[57] ),
    .X(_0412_));
 sg13g2_nand2_1 _1898_ (.Y(_0413_),
    .A(net82),
    .B(_0412_));
 sg13g2_xnor2_1 _1899_ (.Y(_0414_),
    .A(_0410_),
    .B(_0413_));
 sg13g2_xnor2_1 _1900_ (.Y(_0415_),
    .A(_0409_),
    .B(_0414_));
 sg13g2_nor2_1 _1901_ (.A(net146),
    .B(_0415_),
    .Y(_0293_));
 sg13g2_buf_1 _1902_ (.A(\tokenflow_inst.i6.ydata[6] ),
    .X(_0416_));
 sg13g2_inv_1 _1903_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_buf_1 _1904_ (.A(\tokenflow_inst.i6.ydata[58] ),
    .X(_0418_));
 sg13g2_inv_1 _1905_ (.Y(_0419_),
    .A(_0418_));
 sg13g2_or2_1 _1906_ (.X(_0420_),
    .B(_0410_),
    .A(_0412_));
 sg13g2_and2_1 _1907_ (.A(_0357_),
    .B(_0391_),
    .X(_0421_));
 sg13g2_and2_1 _1908_ (.A(_0412_),
    .B(_0410_),
    .X(_0422_));
 sg13g2_buf_1 _1909_ (.A(_0422_),
    .X(_0423_));
 sg13g2_a221oi_1 _1910_ (.B2(_0421_),
    .C1(_0423_),
    .B1(_0420_),
    .A1(_0390_),
    .Y(_0424_),
    .A2(_0410_));
 sg13g2_buf_1 _1911_ (.A(_0424_),
    .X(_0425_));
 sg13g2_and2_1 _1912_ (.A(_0391_),
    .B(_0390_),
    .X(_0426_));
 sg13g2_and2_1 _1913_ (.A(_0357_),
    .B(_0390_),
    .X(_0427_));
 sg13g2_o21ai_1 _1914_ (.B1(_0412_),
    .Y(_0428_),
    .A1(_0426_),
    .A2(_0427_));
 sg13g2_buf_1 _1915_ (.A(_0428_),
    .X(_0429_));
 sg13g2_a21oi_1 _1916_ (.A1(_0426_),
    .A2(_0420_),
    .Y(_0430_),
    .B1(_0423_));
 sg13g2_a22oi_1 _1917_ (.Y(_0431_),
    .B1(_0430_),
    .B2(_0396_),
    .A2(_0429_),
    .A1(_0425_));
 sg13g2_xnor2_1 _1918_ (.Y(_0432_),
    .A(_0419_),
    .B(_0431_));
 sg13g2_nand2_1 _1919_ (.Y(_0433_),
    .A(_0362_),
    .B(_0432_));
 sg13g2_xnor2_1 _1920_ (.Y(_0434_),
    .A(_0417_),
    .B(_0433_));
 sg13g2_nor2_1 _1921_ (.A(net146),
    .B(_0434_),
    .Y(_0304_));
 sg13g2_buf_1 _1922_ (.A(net92),
    .X(_0435_));
 sg13g2_nor2b_1 _1923_ (.A(_0410_),
    .B_N(_0412_),
    .Y(_0436_));
 sg13g2_nor2b_1 _1924_ (.A(_0412_),
    .B_N(_0410_),
    .Y(_0437_));
 sg13g2_a21oi_1 _1925_ (.A1(net89),
    .A2(_0436_),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_nor2_1 _1926_ (.A(_0419_),
    .B(_0416_),
    .Y(_0439_));
 sg13g2_nor2_1 _1927_ (.A(_0418_),
    .B(_0417_),
    .Y(_0440_));
 sg13g2_a21oi_1 _1928_ (.A1(net89),
    .A2(_0439_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nor2_1 _1929_ (.A(_0438_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_o21ai_1 _1930_ (.B1(_0416_),
    .Y(_0443_),
    .A1(_0418_),
    .A2(_0423_));
 sg13g2_nand2_1 _1931_ (.Y(_0444_),
    .A(_0418_),
    .B(_0423_));
 sg13g2_a21oi_1 _1932_ (.A1(_0443_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(_0378_));
 sg13g2_a21oi_1 _1933_ (.A1(_0409_),
    .A2(_0442_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_buf_2 _1934_ (.A(\tokenflow_inst.i6.ydata[7] ),
    .X(_0447_));
 sg13g2_buf_2 _1935_ (.A(\tokenflow_inst.i6.ydata[59] ),
    .X(_0448_));
 sg13g2_nand2_1 _1936_ (.Y(_0449_),
    .A(_0361_),
    .B(_0448_));
 sg13g2_xor2_1 _1937_ (.B(_0449_),
    .A(_0447_),
    .X(_0450_));
 sg13g2_xnor2_1 _1938_ (.Y(_0451_),
    .A(_0446_),
    .B(_0450_));
 sg13g2_nor2_1 _1939_ (.A(_0400_),
    .B(_0451_),
    .Y(_0313_));
 sg13g2_buf_2 _1940_ (.A(\tokenflow_inst.i6.ydata[8] ),
    .X(_0452_));
 sg13g2_buf_2 _1941_ (.A(\tokenflow_inst.i6.ydata[60] ),
    .X(_0453_));
 sg13g2_nand2_1 _1942_ (.Y(_0454_),
    .A(_0425_),
    .B(_0429_));
 sg13g2_or2_1 _1943_ (.X(_0455_),
    .B(_0447_),
    .A(_0448_));
 sg13g2_buf_1 _1944_ (.A(_0455_),
    .X(_0456_));
 sg13g2_nand3_1 _1945_ (.B(_0454_),
    .C(_0456_),
    .A(_0416_),
    .Y(_0457_));
 sg13g2_nand3_1 _1946_ (.B(_0454_),
    .C(_0456_),
    .A(_0418_),
    .Y(_0458_));
 sg13g2_a22oi_1 _1947_ (.Y(_0459_),
    .B1(_0457_),
    .B2(_0458_),
    .A2(_0430_),
    .A1(_0396_));
 sg13g2_and2_1 _1948_ (.A(_0448_),
    .B(_0447_),
    .X(_0460_));
 sg13g2_nor2_1 _1949_ (.A(_0419_),
    .B(_0417_),
    .Y(_0461_));
 sg13g2_o21ai_1 _1950_ (.B1(_0456_),
    .Y(_0462_),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_nand2b_1 _1951_ (.Y(_0463_),
    .B(_0462_),
    .A_N(_0459_));
 sg13g2_xnor2_1 _1952_ (.Y(_0464_),
    .A(_0453_),
    .B(_0463_));
 sg13g2_nor2_1 _1953_ (.A(_0380_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_xnor2_1 _1954_ (.Y(_0466_),
    .A(_0452_),
    .B(_0465_));
 sg13g2_nor2_1 _1955_ (.A(_0400_),
    .B(_0466_),
    .Y(_0314_));
 sg13g2_nor2b_1 _1956_ (.A(_0452_),
    .B_N(_0453_),
    .Y(_0467_));
 sg13g2_nor2b_1 _1957_ (.A(_0448_),
    .B_N(_0447_),
    .Y(_0468_));
 sg13g2_xor2_1 _1958_ (.B(_0452_),
    .A(_0453_),
    .X(_0469_));
 sg13g2_nor2b_1 _1959_ (.A(_0447_),
    .B_N(_0448_),
    .Y(_0470_));
 sg13g2_a22oi_1 _1960_ (.Y(_0471_),
    .B1(_0469_),
    .B2(_0470_),
    .A2(_0468_),
    .A1(_0467_));
 sg13g2_nand2b_1 _1961_ (.Y(_0472_),
    .B(_0435_),
    .A_N(_0471_));
 sg13g2_o21ai_1 _1962_ (.B1(_0357_),
    .Y(_0473_),
    .A1(_0448_),
    .A2(_0453_));
 sg13g2_nand3_1 _1963_ (.B(_0452_),
    .C(_0473_),
    .A(_0447_),
    .Y(_0474_));
 sg13g2_a22oi_1 _1964_ (.Y(_0475_),
    .B1(_0472_),
    .B2(_0474_),
    .A2(_0408_),
    .A1(_0403_));
 sg13g2_o21ai_1 _1965_ (.B1(_0474_),
    .Y(_0476_),
    .A1(_0377_),
    .A2(_0471_));
 sg13g2_nand2_1 _1966_ (.Y(_0477_),
    .A(_0448_),
    .B(_0447_));
 sg13g2_nor2_1 _1967_ (.A(_0453_),
    .B(_0452_),
    .Y(_0478_));
 sg13g2_nand2_1 _1968_ (.Y(_0479_),
    .A(_0453_),
    .B(_0452_));
 sg13g2_o21ai_1 _1969_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0477_),
    .A2(_0478_));
 sg13g2_and2_1 _1970_ (.A(net92),
    .B(_0480_),
    .X(_0481_));
 sg13g2_a21o_1 _1971_ (.A2(_0476_),
    .A1(_0445_),
    .B1(_0481_),
    .X(_0482_));
 sg13g2_a21o_1 _1972_ (.A2(_0475_),
    .A1(_0442_),
    .B1(_0482_),
    .X(_0483_));
 sg13g2_buf_1 _1973_ (.A(_0483_),
    .X(_0484_));
 sg13g2_buf_1 _1974_ (.A(\tokenflow_inst.i6.ydata[9] ),
    .X(_0485_));
 sg13g2_buf_1 _1975_ (.A(\tokenflow_inst.i6.ydata[61] ),
    .X(_0486_));
 sg13g2_nand2_1 _1976_ (.Y(_0487_),
    .A(_0411_),
    .B(net116));
 sg13g2_xnor2_1 _1977_ (.Y(_0488_),
    .A(net117),
    .B(_0487_));
 sg13g2_xnor2_1 _1978_ (.Y(_0489_),
    .A(_0484_),
    .B(_0488_));
 sg13g2_nor2_1 _1979_ (.A(net146),
    .B(_0489_),
    .Y(_0315_));
 sg13g2_buf_1 _1980_ (.A(\tokenflow_inst.i6.ydata[10] ),
    .X(_0490_));
 sg13g2_buf_1 _1981_ (.A(\tokenflow_inst.i6.ydata[62] ),
    .X(_0491_));
 sg13g2_nor2_1 _1982_ (.A(net116),
    .B(net117),
    .Y(_0492_));
 sg13g2_a22oi_1 _1983_ (.Y(_0493_),
    .B1(_0486_),
    .B2(net117),
    .A2(_0452_),
    .A1(_0453_));
 sg13g2_or2_1 _1984_ (.X(_0494_),
    .B(_0493_),
    .A(_0492_));
 sg13g2_buf_1 _1985_ (.A(_0494_),
    .X(_0495_));
 sg13g2_and4_1 _1986_ (.A(_0393_),
    .B(_0394_),
    .C(_0430_),
    .D(_0462_),
    .X(_0496_));
 sg13g2_buf_1 _1987_ (.A(_0496_),
    .X(_0497_));
 sg13g2_nand4_1 _1988_ (.B(_0425_),
    .C(_0429_),
    .A(_0417_),
    .Y(_0498_),
    .D(_0477_));
 sg13g2_nand4_1 _1989_ (.B(_0425_),
    .C(_0429_),
    .A(_0419_),
    .Y(_0499_),
    .D(_0477_));
 sg13g2_xor2_1 _1990_ (.B(net117),
    .A(net116),
    .X(_0500_));
 sg13g2_nand4_1 _1991_ (.B(_0456_),
    .C(_0469_),
    .A(_0435_),
    .Y(_0501_),
    .D(_0500_));
 sg13g2_nor3_1 _1992_ (.A(_0418_),
    .B(_0416_),
    .C(_0460_),
    .Y(_0502_));
 sg13g2_nor2_1 _1993_ (.A(_0501_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_nand3_1 _1994_ (.B(_0499_),
    .C(_0503_),
    .A(_0498_),
    .Y(_0504_));
 sg13g2_nor2_1 _1995_ (.A(_0497_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_nand3b_1 _1996_ (.B(_0495_),
    .C(net114),
    .Y(_0506_),
    .A_N(_0505_));
 sg13g2_o21ai_1 _1997_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net114),
    .A2(_0495_));
 sg13g2_nand2_1 _1998_ (.Y(_0508_),
    .A(net84),
    .B(net114));
 sg13g2_a22oi_1 _1999_ (.Y(_0509_),
    .B1(_0508_),
    .B2(_0505_),
    .A2(_0507_),
    .A1(net84));
 sg13g2_xor2_1 _2000_ (.B(_0509_),
    .A(net115),
    .X(_0510_));
 sg13g2_nor2_1 _2001_ (.A(net146),
    .B(_0510_),
    .Y(_0241_));
 sg13g2_buf_1 _2002_ (.A(\tokenflow_inst.i6.ydata[11] ),
    .X(_0511_));
 sg13g2_nor2b_1 _2003_ (.A(net116),
    .B_N(net117),
    .Y(_0512_));
 sg13g2_nor2b_1 _2004_ (.A(\tokenflow_inst.i6.ydata[10] ),
    .B_N(\tokenflow_inst.i6.ydata[62] ),
    .Y(_0513_));
 sg13g2_nor2b_1 _2005_ (.A(net114),
    .B_N(net115),
    .Y(_0514_));
 sg13g2_or2_1 _2006_ (.X(_0515_),
    .B(_0514_),
    .A(_0513_));
 sg13g2_nor2b_1 _2007_ (.A(net117),
    .B_N(net116),
    .Y(_0516_));
 sg13g2_a22oi_1 _2008_ (.Y(_0517_),
    .B1(_0515_),
    .B2(_0516_),
    .A2(_0513_),
    .A1(_0512_));
 sg13g2_o21ai_1 _2009_ (.B1(_0358_),
    .Y(_0518_),
    .A1(net116),
    .A2(net114));
 sg13g2_nand3_1 _2010_ (.B(_0490_),
    .C(_0518_),
    .A(net117),
    .Y(_0519_));
 sg13g2_o21ai_1 _2011_ (.B1(_0519_),
    .Y(_0520_),
    .A1(_0378_),
    .A2(_0517_));
 sg13g2_nand2_1 _2012_ (.Y(_0521_),
    .A(_0476_),
    .B(_0520_));
 sg13g2_nand3_1 _2013_ (.B(_0490_),
    .C(_0481_),
    .A(_0485_),
    .Y(_0522_));
 sg13g2_o21ai_1 _2014_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0446_),
    .A2(_0521_));
 sg13g2_a21o_1 _2015_ (.A2(_0481_),
    .A1(_0485_),
    .B1(_0486_),
    .X(_0524_));
 sg13g2_inv_1 _2016_ (.Y(_0525_),
    .A(_0491_));
 sg13g2_a21oi_1 _2017_ (.A1(_0359_),
    .A2(_0480_),
    .Y(_0526_),
    .B1(net117));
 sg13g2_nor2_1 _2018_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_a21oi_1 _2019_ (.A1(_0524_),
    .A2(_0527_),
    .Y(_0528_),
    .B1(net115));
 sg13g2_nand2b_1 _2020_ (.Y(_0529_),
    .B(net116),
    .A_N(_0526_));
 sg13g2_and2_1 _2021_ (.A(_0525_),
    .B(_0529_),
    .X(_0530_));
 sg13g2_buf_1 _2022_ (.A(\tokenflow_inst.i6.ydata[63] ),
    .X(_0531_));
 sg13g2_buf_1 _2023_ (.A(_0531_),
    .X(_0532_));
 sg13g2_o21ai_1 _2024_ (.B1(net91),
    .Y(_0533_),
    .A1(_0528_),
    .A2(_0530_));
 sg13g2_or3_1 _2025_ (.A(_0532_),
    .B(_0528_),
    .C(_0530_),
    .X(_0534_));
 sg13g2_o21ai_1 _2026_ (.B1(_0534_),
    .Y(_0535_),
    .A1(_0523_),
    .A2(_0533_));
 sg13g2_nand2_1 _2027_ (.Y(_0536_),
    .A(_0411_),
    .B(_0532_));
 sg13g2_a22oi_1 _2028_ (.Y(_0537_),
    .B1(_0536_),
    .B2(_0523_),
    .A2(_0535_),
    .A1(net84));
 sg13g2_xor2_1 _2029_ (.B(_0537_),
    .A(_0511_),
    .X(_0538_));
 sg13g2_nor2_1 _2030_ (.A(net146),
    .B(_0538_),
    .Y(_0242_));
 sg13g2_nor2b_1 _2031_ (.A(net113),
    .B_N(_0531_),
    .Y(_0539_));
 sg13g2_xor2_1 _2032_ (.B(_0511_),
    .A(net91),
    .X(_0540_));
 sg13g2_a22oi_1 _2033_ (.Y(_0541_),
    .B1(_0540_),
    .B2(_0513_),
    .A2(_0539_),
    .A1(_0514_));
 sg13g2_o21ai_1 _2034_ (.B1(net92),
    .Y(_0542_),
    .A1(net114),
    .A2(net91));
 sg13g2_nand3_1 _2035_ (.B(net113),
    .C(_0542_),
    .A(net115),
    .Y(_0543_));
 sg13g2_o21ai_1 _2036_ (.B1(_0543_),
    .Y(_0544_),
    .A1(net87),
    .A2(_0541_));
 sg13g2_or2_1 _2037_ (.X(_0545_),
    .B(net113),
    .A(net91));
 sg13g2_nor2_1 _2038_ (.A(\tokenflow_inst.i6.ydata[62] ),
    .B(net115),
    .Y(_0546_));
 sg13g2_nand2_1 _2039_ (.Y(_0547_),
    .A(net114),
    .B(net115));
 sg13g2_o21ai_1 _2040_ (.B1(_0547_),
    .Y(_0548_),
    .A1(_0495_),
    .A2(_0546_));
 sg13g2_and2_1 _2041_ (.A(net91),
    .B(net113),
    .X(_0549_));
 sg13g2_a21oi_1 _2042_ (.A1(_0545_),
    .A2(_0548_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_nor2_1 _2043_ (.A(net85),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_a21o_1 _2044_ (.A2(_0544_),
    .A1(_0505_),
    .B1(_0551_),
    .X(_0552_));
 sg13g2_buf_2 _2045_ (.A(\tokenflow_inst.i6.ydata[12] ),
    .X(_0553_));
 sg13g2_buf_1 _2046_ (.A(\tokenflow_inst.i6.ydata[64] ),
    .X(_0554_));
 sg13g2_nand2_1 _2047_ (.Y(_0555_),
    .A(net82),
    .B(net112));
 sg13g2_xnor2_1 _2048_ (.Y(_0556_),
    .A(_0553_),
    .B(_0555_));
 sg13g2_xnor2_1 _2049_ (.Y(_0557_),
    .A(_0552_),
    .B(_0556_));
 sg13g2_nor2_1 _2050_ (.A(net146),
    .B(_0557_),
    .Y(_0243_));
 sg13g2_nor2b_1 _2051_ (.A(net91),
    .B_N(net113),
    .Y(_0558_));
 sg13g2_nor2b_1 _2052_ (.A(_0553_),
    .B_N(net112),
    .Y(_0559_));
 sg13g2_nor2b_1 _2053_ (.A(net112),
    .B_N(_0553_),
    .Y(_0560_));
 sg13g2_or2_1 _2054_ (.X(_0561_),
    .B(_0560_),
    .A(_0559_));
 sg13g2_a22oi_1 _2055_ (.Y(_0562_),
    .B1(_0561_),
    .B2(_0539_),
    .A2(_0559_),
    .A1(_0558_));
 sg13g2_o21ai_1 _2056_ (.B1(net89),
    .Y(_0563_),
    .A1(net91),
    .A2(net112));
 sg13g2_nand3_1 _2057_ (.B(_0553_),
    .C(_0563_),
    .A(net113),
    .Y(_0564_));
 sg13g2_o21ai_1 _2058_ (.B1(_0564_),
    .Y(_0565_),
    .A1(net85),
    .A2(_0562_));
 sg13g2_nand3_1 _2059_ (.B(_0520_),
    .C(_0565_),
    .A(_0484_),
    .Y(_0566_));
 sg13g2_a22oi_1 _2060_ (.Y(_0567_),
    .B1(_0491_),
    .B2(net115),
    .A2(\tokenflow_inst.i6.ydata[9] ),
    .A1(\tokenflow_inst.i6.ydata[61] ));
 sg13g2_a22oi_1 _2061_ (.Y(_0568_),
    .B1(net112),
    .B2(_0553_),
    .A2(net113),
    .A1(_0531_));
 sg13g2_o21ai_1 _2062_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_0546_),
    .A2(_0567_));
 sg13g2_nor2_1 _2063_ (.A(_0531_),
    .B(net113),
    .Y(_0570_));
 sg13g2_nor2_1 _2064_ (.A(net112),
    .B(_0553_),
    .Y(_0571_));
 sg13g2_nand2_1 _2065_ (.Y(_0572_),
    .A(net112),
    .B(_0553_));
 sg13g2_o21ai_1 _2066_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_nand3_1 _2067_ (.B(_0569_),
    .C(_0573_),
    .A(net84),
    .Y(_0574_));
 sg13g2_nand2_1 _2068_ (.Y(_0575_),
    .A(_0566_),
    .B(_0574_));
 sg13g2_buf_1 _2069_ (.A(\tokenflow_inst.i6.ydata[13] ),
    .X(_0576_));
 sg13g2_buf_1 _2070_ (.A(\tokenflow_inst.i6.ydata[65] ),
    .X(_0577_));
 sg13g2_nand2_1 _2071_ (.Y(_0578_),
    .A(net82),
    .B(_0577_));
 sg13g2_xnor2_1 _2072_ (.Y(_0579_),
    .A(net111),
    .B(_0578_));
 sg13g2_xnor2_1 _2073_ (.Y(_0580_),
    .A(_0575_),
    .B(_0579_));
 sg13g2_nor2_1 _2074_ (.A(net146),
    .B(_0580_),
    .Y(_0244_));
 sg13g2_buf_1 _2075_ (.A(\tokenflow_inst.i6.ydata[14] ),
    .X(_0581_));
 sg13g2_inv_1 _2076_ (.Y(_0582_),
    .A(net109));
 sg13g2_buf_1 _2077_ (.A(\tokenflow_inst.i6.ydata[66] ),
    .X(_0583_));
 sg13g2_nand2_1 _2078_ (.Y(_0584_),
    .A(net90),
    .B(net108));
 sg13g2_xnor2_1 _2079_ (.Y(_0585_),
    .A(_0582_),
    .B(_0584_));
 sg13g2_nor2_1 _2080_ (.A(net110),
    .B(net111),
    .Y(_0586_));
 sg13g2_nand2_1 _2081_ (.Y(_0587_),
    .A(net110),
    .B(net111));
 sg13g2_o21ai_1 _2082_ (.B1(_0587_),
    .Y(_0588_),
    .A1(_0572_),
    .A2(_0586_));
 sg13g2_nor3_1 _2083_ (.A(net87),
    .B(_0495_),
    .C(_0541_),
    .Y(_0589_));
 sg13g2_and2_1 _2084_ (.A(net114),
    .B(net115),
    .X(_0590_));
 sg13g2_a21oi_1 _2085_ (.A1(_0545_),
    .A2(_0590_),
    .Y(_0591_),
    .B1(_0549_));
 sg13g2_o21ai_1 _2086_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0495_),
    .A2(_0543_));
 sg13g2_nor2b_1 _2087_ (.A(\tokenflow_inst.i6.ydata[13] ),
    .B_N(net110),
    .Y(_0593_));
 sg13g2_xor2_1 _2088_ (.B(_0576_),
    .A(net110),
    .X(_0594_));
 sg13g2_a22oi_1 _2089_ (.Y(_0595_),
    .B1(_0594_),
    .B2(_0559_),
    .A2(_0593_),
    .A1(_0560_));
 sg13g2_o21ai_1 _2090_ (.B1(net92),
    .Y(_0596_),
    .A1(_0554_),
    .A2(net110));
 sg13g2_nand3_1 _2091_ (.B(net111),
    .C(_0596_),
    .A(_0553_),
    .Y(_0597_));
 sg13g2_o21ai_1 _2092_ (.B1(_0597_),
    .Y(_0598_),
    .A1(net87),
    .A2(_0595_));
 sg13g2_o21ai_1 _2093_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0589_),
    .A2(_0592_));
 sg13g2_nand2b_1 _2094_ (.Y(_0600_),
    .B(_0599_),
    .A_N(_0588_));
 sg13g2_nand2_1 _2095_ (.Y(_0601_),
    .A(_0544_),
    .B(_0598_));
 sg13g2_nor3_1 _2096_ (.A(_0497_),
    .B(_0504_),
    .C(_0601_),
    .Y(_0602_));
 sg13g2_a21oi_1 _2097_ (.A1(net84),
    .A2(_0600_),
    .Y(_0603_),
    .B1(_0602_));
 sg13g2_xnor2_1 _2098_ (.Y(_0604_),
    .A(_0585_),
    .B(_0603_));
 sg13g2_nor2_1 _2099_ (.A(net146),
    .B(_0604_),
    .Y(_0245_));
 sg13g2_buf_1 _2100_ (.A(net164),
    .X(_0605_));
 sg13g2_nor2b_1 _2101_ (.A(net110),
    .B_N(net111),
    .Y(_0606_));
 sg13g2_nor2b_1 _2102_ (.A(net109),
    .B_N(net108),
    .Y(_0607_));
 sg13g2_nor2b_1 _2103_ (.A(net108),
    .B_N(net109),
    .Y(_0608_));
 sg13g2_or2_1 _2104_ (.X(_0609_),
    .B(_0608_),
    .A(_0607_));
 sg13g2_a22oi_1 _2105_ (.Y(_0610_),
    .B1(_0609_),
    .B2(_0593_),
    .A2(_0607_),
    .A1(_0606_));
 sg13g2_o21ai_1 _2106_ (.B1(net89),
    .Y(_0611_),
    .A1(net110),
    .A2(net108));
 sg13g2_nand3_1 _2107_ (.B(net109),
    .C(_0611_),
    .A(net111),
    .Y(_0612_));
 sg13g2_o21ai_1 _2108_ (.B1(_0612_),
    .Y(_0613_),
    .A1(net85),
    .A2(_0610_));
 sg13g2_nor2b_1 _2109_ (.A(_0566_),
    .B_N(_0613_),
    .Y(_0614_));
 sg13g2_and3_1 _2110_ (.X(_0615_),
    .A(net89),
    .B(_0569_),
    .C(_0573_));
 sg13g2_nand3_1 _2111_ (.B(_0581_),
    .C(_0615_),
    .A(net111),
    .Y(_0616_));
 sg13g2_nand4_1 _2112_ (.B(_0576_),
    .C(_0569_),
    .A(net90),
    .Y(_0617_),
    .D(_0573_));
 sg13g2_a21o_1 _2113_ (.A2(_0617_),
    .A1(_0582_),
    .B1(_0584_),
    .X(_0618_));
 sg13g2_o21ai_1 _2114_ (.B1(net110),
    .Y(_0619_),
    .A1(net108),
    .A2(_0581_));
 sg13g2_nor2_1 _2115_ (.A(net87),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _2116_ (.B1(_0620_),
    .Y(_0621_),
    .A1(net111),
    .A2(_0615_));
 sg13g2_nand3_1 _2117_ (.B(_0618_),
    .C(_0621_),
    .A(_0616_),
    .Y(_0622_));
 sg13g2_nor2_1 _2118_ (.A(_0614_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_buf_1 _2119_ (.A(\tokenflow_inst.i6.ydata[15] ),
    .X(_0624_));
 sg13g2_buf_1 _2120_ (.A(\tokenflow_inst.i6.ydata[67] ),
    .X(_0625_));
 sg13g2_nand2_1 _2121_ (.Y(_0626_),
    .A(net86),
    .B(net106));
 sg13g2_xor2_1 _2122_ (.B(_0626_),
    .A(net107),
    .X(_0627_));
 sg13g2_xnor2_1 _2123_ (.Y(_0628_),
    .A(_0623_),
    .B(_0627_));
 sg13g2_nor2_1 _2124_ (.A(net145),
    .B(_0628_),
    .Y(_0246_));
 sg13g2_buf_2 _2125_ (.A(\tokenflow_inst.i6.ydata[16] ),
    .X(_0629_));
 sg13g2_nor2b_1 _2126_ (.A(net107),
    .B_N(net106),
    .Y(_0630_));
 sg13g2_xor2_1 _2127_ (.B(net107),
    .A(net106),
    .X(_0631_));
 sg13g2_a22oi_1 _2128_ (.Y(_0632_),
    .B1(_0631_),
    .B2(_0607_),
    .A2(_0630_),
    .A1(_0608_));
 sg13g2_o21ai_1 _2129_ (.B1(net89),
    .Y(_0633_),
    .A1(_0583_),
    .A2(net106));
 sg13g2_nand3_1 _2130_ (.B(net107),
    .C(_0633_),
    .A(net109),
    .Y(_0634_));
 sg13g2_o21ai_1 _2131_ (.B1(_0634_),
    .Y(_0635_),
    .A1(net87),
    .A2(_0632_));
 sg13g2_and2_1 _2132_ (.A(_0598_),
    .B(_0635_),
    .X(_0636_));
 sg13g2_buf_1 _2133_ (.A(\tokenflow_inst.i6.ydata[68] ),
    .X(_0637_));
 sg13g2_inv_1 _2134_ (.Y(_0638_),
    .A(net105));
 sg13g2_a21oi_1 _2135_ (.A1(_0552_),
    .A2(_0636_),
    .Y(_0639_),
    .B1(_0638_));
 sg13g2_nor2_1 _2136_ (.A(net106),
    .B(net107),
    .Y(_0640_));
 sg13g2_a21o_1 _2137_ (.A2(_0588_),
    .A1(net109),
    .B1(net108),
    .X(_0641_));
 sg13g2_o21ai_1 _2138_ (.B1(_0641_),
    .Y(_0642_),
    .A1(net109),
    .A2(_0588_));
 sg13g2_nand2_1 _2139_ (.Y(_0643_),
    .A(net106),
    .B(net107));
 sg13g2_o21ai_1 _2140_ (.B1(_0643_),
    .Y(_0644_),
    .A1(_0640_),
    .A2(_0642_));
 sg13g2_nor2_1 _2141_ (.A(net83),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_nor2_1 _2142_ (.A(net83),
    .B(net105),
    .Y(_0646_));
 sg13g2_nand2_1 _2143_ (.Y(_0647_),
    .A(net86),
    .B(net105));
 sg13g2_and3_1 _2144_ (.X(_0648_),
    .A(_0552_),
    .B(_0636_),
    .C(_0647_));
 sg13g2_a221oi_1 _2145_ (.B2(_0644_),
    .C1(_0648_),
    .B1(_0646_),
    .A1(_0639_),
    .Y(_0649_),
    .A2(_0645_));
 sg13g2_xor2_1 _2146_ (.B(_0649_),
    .A(_0629_),
    .X(_0650_));
 sg13g2_nor2_1 _2147_ (.A(net145),
    .B(_0650_),
    .Y(_0247_));
 sg13g2_buf_2 _2148_ (.A(\tokenflow_inst.i6.ydata[17] ),
    .X(_0651_));
 sg13g2_nor2b_1 _2149_ (.A(net106),
    .B_N(_0624_),
    .Y(_0652_));
 sg13g2_nor2b_1 _2150_ (.A(_0629_),
    .B_N(_0637_),
    .Y(_0653_));
 sg13g2_nor2b_1 _2151_ (.A(_0637_),
    .B_N(_0629_),
    .Y(_0654_));
 sg13g2_or2_1 _2152_ (.X(_0655_),
    .B(_0654_),
    .A(_0653_));
 sg13g2_a22oi_1 _2153_ (.Y(_0656_),
    .B1(_0655_),
    .B2(_0630_),
    .A2(_0653_),
    .A1(_0652_));
 sg13g2_o21ai_1 _2154_ (.B1(net92),
    .Y(_0657_),
    .A1(_0625_),
    .A2(net105));
 sg13g2_nand3_1 _2155_ (.B(_0629_),
    .C(_0657_),
    .A(net107),
    .Y(_0658_));
 sg13g2_o21ai_1 _2156_ (.B1(_0658_),
    .Y(_0659_),
    .A1(net87),
    .A2(_0656_));
 sg13g2_and4_1 _2157_ (.A(_0520_),
    .B(_0565_),
    .C(_0613_),
    .D(_0659_),
    .X(_0660_));
 sg13g2_a22oi_1 _2158_ (.Y(_0661_),
    .B1(_0660_),
    .B2(_0484_),
    .A2(_0659_),
    .A1(_0622_));
 sg13g2_buf_1 _2159_ (.A(_0661_),
    .X(_0662_));
 sg13g2_nor2_1 _2160_ (.A(net105),
    .B(_0629_),
    .Y(_0663_));
 sg13g2_nand2_1 _2161_ (.Y(_0664_),
    .A(net105),
    .B(_0629_));
 sg13g2_o21ai_1 _2162_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_0643_),
    .A2(_0663_));
 sg13g2_buf_1 _2163_ (.A(_0665_),
    .X(_0666_));
 sg13g2_buf_1 _2164_ (.A(\tokenflow_inst.i6.ydata[69] ),
    .X(_0667_));
 sg13g2_nor2b_1 _2165_ (.A(_0666_),
    .B_N(net104),
    .Y(_0668_));
 sg13g2_nor2b_1 _2166_ (.A(net104),
    .B_N(_0666_),
    .Y(_0669_));
 sg13g2_a21o_1 _2167_ (.A2(_0668_),
    .A1(_0662_),
    .B1(_0669_),
    .X(_0670_));
 sg13g2_a21oi_1 _2168_ (.A1(net82),
    .A2(net104),
    .Y(_0671_),
    .B1(_0662_));
 sg13g2_a21oi_1 _2169_ (.A1(net84),
    .A2(_0670_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_xor2_1 _2170_ (.B(_0672_),
    .A(_0651_),
    .X(_0673_));
 sg13g2_nor2_1 _2171_ (.A(net145),
    .B(_0673_),
    .Y(_0248_));
 sg13g2_nor2_1 _2172_ (.A(\tokenflow_inst.i6.ydata[69] ),
    .B(_0651_),
    .Y(_0674_));
 sg13g2_a22oi_1 _2173_ (.Y(_0675_),
    .B1(_0625_),
    .B2(net107),
    .A2(net109),
    .A1(net108));
 sg13g2_nor3_1 _2174_ (.A(_0640_),
    .B(_0663_),
    .C(_0675_),
    .Y(_0676_));
 sg13g2_a21oi_1 _2175_ (.A1(net105),
    .A2(_0629_),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_nand2_1 _2176_ (.Y(_0678_),
    .A(net104),
    .B(_0651_));
 sg13g2_o21ai_1 _2177_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0674_),
    .A2(_0677_));
 sg13g2_nor2b_1 _2178_ (.A(_0651_),
    .B_N(net104),
    .Y(_0680_));
 sg13g2_xor2_1 _2179_ (.B(_0651_),
    .A(net104),
    .X(_0681_));
 sg13g2_a22oi_1 _2180_ (.Y(_0682_),
    .B1(_0681_),
    .B2(_0653_),
    .A2(_0680_),
    .A1(_0654_));
 sg13g2_o21ai_1 _2181_ (.B1(net89),
    .Y(_0683_),
    .A1(net105),
    .A2(net104));
 sg13g2_nand3_1 _2182_ (.B(_0651_),
    .C(_0683_),
    .A(_0629_),
    .Y(_0684_));
 sg13g2_o21ai_1 _2183_ (.B1(_0684_),
    .Y(_0685_),
    .A1(net85),
    .A2(_0682_));
 sg13g2_nand2_1 _2184_ (.Y(_0686_),
    .A(_0635_),
    .B(_0685_));
 sg13g2_nor2_1 _2185_ (.A(_0379_),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_nor4_1 _2186_ (.A(_0497_),
    .B(_0504_),
    .C(_0601_),
    .D(_0686_),
    .Y(_0688_));
 sg13g2_a221oi_1 _2187_ (.B2(_0600_),
    .C1(_0688_),
    .B1(_0687_),
    .A1(_0360_),
    .Y(_0689_),
    .A2(_0679_));
 sg13g2_buf_1 _2188_ (.A(_0689_),
    .X(_0690_));
 sg13g2_buf_1 _2189_ (.A(\tokenflow_inst.i6.ydata[70] ),
    .X(_0691_));
 sg13g2_buf_1 _2190_ (.A(\tokenflow_inst.i6.ydata[18] ),
    .X(_0692_));
 sg13g2_a21oi_1 _2191_ (.A1(net82),
    .A2(net103),
    .Y(_0693_),
    .B1(net102));
 sg13g2_and3_1 _2192_ (.X(_0694_),
    .A(net89),
    .B(net103),
    .C(net102));
 sg13g2_nor2_1 _2193_ (.A(_0693_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_xor2_1 _2194_ (.B(_0695_),
    .A(_0690_),
    .X(_0696_));
 sg13g2_nor2_1 _2195_ (.A(net145),
    .B(_0696_),
    .Y(_0249_));
 sg13g2_nor2_1 _2196_ (.A(_0691_),
    .B(\tokenflow_inst.i6.ydata[18] ),
    .Y(_0697_));
 sg13g2_nor3_1 _2197_ (.A(net87),
    .B(_0674_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_nand2_1 _2198_ (.Y(_0699_),
    .A(_0666_),
    .B(_0698_));
 sg13g2_nor2_1 _2199_ (.A(_0678_),
    .B(_0697_),
    .Y(_0700_));
 sg13g2_nand2_1 _2200_ (.Y(_0701_),
    .A(net90),
    .B(_0700_));
 sg13g2_nand3b_1 _2201_ (.B(_0699_),
    .C(_0701_),
    .Y(_0702_),
    .A_N(_0694_));
 sg13g2_nor2b_1 _2202_ (.A(_0667_),
    .B_N(_0651_),
    .Y(_0703_));
 sg13g2_nor2b_1 _2203_ (.A(net102),
    .B_N(net103),
    .Y(_0704_));
 sg13g2_xor2_1 _2204_ (.B(_0692_),
    .A(net103),
    .X(_0705_));
 sg13g2_a22oi_1 _2205_ (.Y(_0706_),
    .B1(_0705_),
    .B2(_0680_),
    .A2(_0704_),
    .A1(_0703_));
 sg13g2_o21ai_1 _2206_ (.B1(net90),
    .Y(_0707_),
    .A1(_0667_),
    .A2(net103));
 sg13g2_nand3_1 _2207_ (.B(_0692_),
    .C(_0707_),
    .A(_0651_),
    .Y(_0708_));
 sg13g2_o21ai_1 _2208_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_0379_),
    .A2(_0706_));
 sg13g2_nor2b_1 _2209_ (.A(_0662_),
    .B_N(_0709_),
    .Y(_0710_));
 sg13g2_nor2_1 _2210_ (.A(_0702_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_buf_1 _2211_ (.A(\tokenflow_inst.i6.ydata[19] ),
    .X(_0712_));
 sg13g2_inv_1 _2212_ (.Y(_0713_),
    .A(net101));
 sg13g2_buf_1 _2213_ (.A(\tokenflow_inst.i6.ydata[71] ),
    .X(_0714_));
 sg13g2_nand2_1 _2214_ (.Y(_0715_),
    .A(net82),
    .B(net100));
 sg13g2_xnor2_1 _2215_ (.Y(_0716_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_xnor2_1 _2216_ (.Y(_0717_),
    .A(_0711_),
    .B(_0716_));
 sg13g2_nor2_1 _2217_ (.A(net145),
    .B(_0717_),
    .Y(_0250_));
 sg13g2_o21ai_1 _2218_ (.B1(net103),
    .Y(_0718_),
    .A1(net100),
    .A2(net101));
 sg13g2_or2_1 _2219_ (.X(_0719_),
    .B(_0718_),
    .A(net83));
 sg13g2_nand3_1 _2220_ (.B(net102),
    .C(net100),
    .A(net88),
    .Y(_0720_));
 sg13g2_a21oi_1 _2221_ (.A1(_0719_),
    .A2(_0720_),
    .Y(_0721_),
    .B1(_0690_));
 sg13g2_inv_1 _2222_ (.Y(_0722_),
    .A(net102));
 sg13g2_nor3_1 _2223_ (.A(_0722_),
    .B(_0713_),
    .C(_0690_),
    .Y(_0723_));
 sg13g2_nand2_1 _2224_ (.Y(_0724_),
    .A(net88),
    .B(net102));
 sg13g2_nand3_1 _2225_ (.B(net100),
    .C(net101),
    .A(net88),
    .Y(_0725_));
 sg13g2_o21ai_1 _2226_ (.B1(_0725_),
    .Y(_0726_),
    .A1(_0718_),
    .A2(_0724_));
 sg13g2_nor3_2 _2227_ (.A(_0721_),
    .B(_0723_),
    .C(_0726_),
    .Y(_0727_));
 sg13g2_buf_1 _2228_ (.A(\tokenflow_inst.i6.ydata[20] ),
    .X(_0728_));
 sg13g2_buf_1 _2229_ (.A(\tokenflow_inst.i6.ydata[72] ),
    .X(_0729_));
 sg13g2_nand2_1 _2230_ (.Y(_0730_),
    .A(net86),
    .B(_0729_));
 sg13g2_xor2_1 _2231_ (.B(_0730_),
    .A(net99),
    .X(_0731_));
 sg13g2_xnor2_1 _2232_ (.Y(_0732_),
    .A(_0727_),
    .B(_0731_));
 sg13g2_nor2_1 _2233_ (.A(net145),
    .B(_0732_),
    .Y(_0252_));
 sg13g2_nor2b_1 _2234_ (.A(_0728_),
    .B_N(\tokenflow_inst.i6.ydata[72] ),
    .Y(_0733_));
 sg13g2_nor2_1 _2235_ (.A(\tokenflow_inst.i6.ydata[71] ),
    .B(_0713_),
    .Y(_0734_));
 sg13g2_nor2b_1 _2236_ (.A(net98),
    .B_N(net99),
    .Y(_0735_));
 sg13g2_or2_1 _2237_ (.X(_0736_),
    .B(_0735_),
    .A(_0733_));
 sg13g2_nor2b_1 _2238_ (.A(net101),
    .B_N(\tokenflow_inst.i6.ydata[71] ),
    .Y(_0737_));
 sg13g2_a22oi_1 _2239_ (.Y(_0738_),
    .B1(_0736_),
    .B2(_0737_),
    .A2(_0734_),
    .A1(_0733_));
 sg13g2_o21ai_1 _2240_ (.B1(net90),
    .Y(_0739_),
    .A1(net100),
    .A2(net98));
 sg13g2_nand3_1 _2241_ (.B(net99),
    .C(_0739_),
    .A(net101),
    .Y(_0740_));
 sg13g2_o21ai_1 _2242_ (.B1(_0740_),
    .Y(_0741_),
    .A1(net85),
    .A2(_0738_));
 sg13g2_nand2_1 _2243_ (.Y(_0742_),
    .A(_0709_),
    .B(_0741_));
 sg13g2_a221oi_1 _2244_ (.B2(_0359_),
    .C1(_0694_),
    .B1(_0700_),
    .A1(_0666_),
    .Y(_0743_),
    .A2(_0698_));
 sg13g2_nand2_1 _2245_ (.Y(_0744_),
    .A(net101),
    .B(net98));
 sg13g2_nand2_1 _2246_ (.Y(_0745_),
    .A(net98),
    .B(net99));
 sg13g2_o21ai_1 _2247_ (.B1(_0745_),
    .Y(_0746_),
    .A1(_0743_),
    .A2(_0744_));
 sg13g2_o21ai_1 _2248_ (.B1(_0714_),
    .Y(_0747_),
    .A1(_0729_),
    .A2(_0728_));
 sg13g2_a21oi_1 _2249_ (.A1(_0713_),
    .A2(_0743_),
    .Y(_0748_),
    .B1(_0747_));
 sg13g2_o21ai_1 _2250_ (.B1(net88),
    .Y(_0749_),
    .A1(_0746_),
    .A2(_0748_));
 sg13g2_nand3_1 _2251_ (.B(net99),
    .C(_0702_),
    .A(net101),
    .Y(_0750_));
 sg13g2_and2_1 _2252_ (.A(_0749_),
    .B(_0750_),
    .X(_0751_));
 sg13g2_o21ai_1 _2253_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0662_),
    .A2(_0742_));
 sg13g2_buf_2 _2254_ (.A(\tokenflow_inst.i6.ydata[21] ),
    .X(_0753_));
 sg13g2_buf_1 _2255_ (.A(\tokenflow_inst.i6.ydata[73] ),
    .X(_0754_));
 sg13g2_nand2_1 _2256_ (.Y(_0755_),
    .A(net82),
    .B(net97));
 sg13g2_xnor2_1 _2257_ (.Y(_0756_),
    .A(_0753_),
    .B(_0755_));
 sg13g2_xnor2_1 _2258_ (.Y(_0757_),
    .A(_0752_),
    .B(_0756_));
 sg13g2_nor2_1 _2259_ (.A(net145),
    .B(_0757_),
    .Y(_0253_));
 sg13g2_and2_1 _2260_ (.A(net99),
    .B(_0753_),
    .X(_0758_));
 sg13g2_o21ai_1 _2261_ (.B1(net88),
    .Y(_0759_),
    .A1(net98),
    .A2(net97));
 sg13g2_nor2b_1 _2262_ (.A(_0753_),
    .B_N(net97),
    .Y(_0760_));
 sg13g2_xor2_1 _2263_ (.B(_0753_),
    .A(net97),
    .X(_0761_));
 sg13g2_a22oi_1 _2264_ (.Y(_0762_),
    .B1(_0761_),
    .B2(_0733_),
    .A2(_0760_),
    .A1(_0735_));
 sg13g2_nor2_1 _2265_ (.A(net85),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_a21oi_1 _2266_ (.A1(_0758_),
    .A2(_0759_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_buf_1 _2267_ (.A(\tokenflow_inst.i6.ydata[22] ),
    .X(_0765_));
 sg13g2_buf_1 _2268_ (.A(\tokenflow_inst.i6.ydata[74] ),
    .X(_0766_));
 sg13g2_nand2_1 _2269_ (.Y(_0767_),
    .A(net88),
    .B(net95));
 sg13g2_xor2_1 _2270_ (.B(_0767_),
    .A(_0765_),
    .X(_0768_));
 sg13g2_and2_1 _2271_ (.A(net182),
    .B(_0768_),
    .X(_0769_));
 sg13g2_nor2b_1 _2272_ (.A(_0764_),
    .B_N(_0769_),
    .Y(_0770_));
 sg13g2_inv_1 _2273_ (.Y(_0771_),
    .A(_0753_));
 sg13g2_a21oi_1 _2274_ (.A1(net98),
    .A2(net99),
    .Y(_0772_),
    .B1(net97));
 sg13g2_nand3_1 _2275_ (.B(net99),
    .C(net97),
    .A(net98),
    .Y(_0773_));
 sg13g2_o21ai_1 _2276_ (.B1(_0773_),
    .Y(_0774_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_and2_1 _2277_ (.A(net90),
    .B(_0774_),
    .X(_0775_));
 sg13g2_buf_1 _2278_ (.A(_0775_),
    .X(_0776_));
 sg13g2_nor3_1 _2279_ (.A(net179),
    .B(_0768_),
    .C(_0776_),
    .Y(_0777_));
 sg13g2_mux2_1 _2280_ (.A0(_0770_),
    .A1(_0777_),
    .S(_0727_),
    .X(_0778_));
 sg13g2_a22oi_1 _2281_ (.Y(_0779_),
    .B1(_0769_),
    .B2(_0776_),
    .A2(_0777_),
    .A1(_0764_));
 sg13g2_nand2b_1 _2282_ (.Y(_0254_),
    .B(_0779_),
    .A_N(_0778_));
 sg13g2_buf_1 _2283_ (.A(\tokenflow_inst.i6.ydata[23] ),
    .X(_0780_));
 sg13g2_nor2_1 _2284_ (.A(net167),
    .B(net94),
    .Y(_0781_));
 sg13g2_and2_1 _2285_ (.A(net182),
    .B(net94),
    .X(_0782_));
 sg13g2_buf_1 _2286_ (.A(\tokenflow_inst.i6.ydata[75] ),
    .X(_0783_));
 sg13g2_inv_1 _2287_ (.Y(_0784_),
    .A(net93));
 sg13g2_nor2_1 _2288_ (.A(_0754_),
    .B(_0771_),
    .Y(_0785_));
 sg13g2_nor2b_1 _2289_ (.A(net96),
    .B_N(net95),
    .Y(_0786_));
 sg13g2_nor2b_1 _2290_ (.A(net95),
    .B_N(net96),
    .Y(_0787_));
 sg13g2_or2_1 _2291_ (.X(_0788_),
    .B(_0787_),
    .A(_0786_));
 sg13g2_a22oi_1 _2292_ (.Y(_0789_),
    .B1(_0788_),
    .B2(_0760_),
    .A2(_0786_),
    .A1(_0785_));
 sg13g2_o21ai_1 _2293_ (.B1(net88),
    .Y(_0790_),
    .A1(net97),
    .A2(net95));
 sg13g2_nand3_1 _2294_ (.B(net96),
    .C(_0790_),
    .A(_0753_),
    .Y(_0791_));
 sg13g2_o21ai_1 _2295_ (.B1(_0791_),
    .Y(_0792_),
    .A1(net83),
    .A2(_0789_));
 sg13g2_and2_1 _2296_ (.A(_0752_),
    .B(_0792_),
    .X(_0793_));
 sg13g2_nor2_1 _2297_ (.A(net95),
    .B(net96),
    .Y(_0794_));
 sg13g2_a22oi_1 _2298_ (.Y(_0795_),
    .B1(net95),
    .B2(net96),
    .A2(_0753_),
    .A1(net97));
 sg13g2_nor2_1 _2299_ (.A(_0794_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_nor2_1 _2300_ (.A(net83),
    .B(net93),
    .Y(_0797_));
 sg13g2_nand3b_1 _2301_ (.B(net93),
    .C(net86),
    .Y(_0798_),
    .A_N(_0796_));
 sg13g2_a21oi_1 _2302_ (.A1(_0752_),
    .A2(_0792_),
    .Y(_0799_),
    .B1(_0798_));
 sg13g2_a221oi_1 _2303_ (.B2(_0797_),
    .C1(_0799_),
    .B1(_0796_),
    .A1(_0784_),
    .Y(_0800_),
    .A2(_0793_));
 sg13g2_mux2_1 _2304_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0800_),
    .X(_0255_));
 sg13g2_nor2b_1 _2305_ (.A(net94),
    .B_N(\tokenflow_inst.i6.ydata[75] ),
    .Y(_0801_));
 sg13g2_nor2b_1 _2306_ (.A(net93),
    .B_N(net94),
    .Y(_0802_));
 sg13g2_or2_1 _2307_ (.X(_0803_),
    .B(_0802_),
    .A(_0801_));
 sg13g2_a22oi_1 _2308_ (.Y(_0804_),
    .B1(_0803_),
    .B2(_0786_),
    .A2(_0801_),
    .A1(_0787_));
 sg13g2_and2_1 _2309_ (.A(net96),
    .B(_0780_),
    .X(_0805_));
 sg13g2_o21ai_1 _2310_ (.B1(net90),
    .Y(_0806_),
    .A1(net95),
    .A2(_0783_));
 sg13g2_nand2_1 _2311_ (.Y(_0807_),
    .A(_0805_),
    .B(_0806_));
 sg13g2_o21ai_1 _2312_ (.B1(_0807_),
    .Y(_0808_),
    .A1(net85),
    .A2(_0804_));
 sg13g2_nor2b_1 _2313_ (.A(_0764_),
    .B_N(_0808_),
    .Y(_0809_));
 sg13g2_nand2_1 _2314_ (.Y(_0810_),
    .A(_0723_),
    .B(_0809_));
 sg13g2_nor2_1 _2315_ (.A(net96),
    .B(_0776_),
    .Y(_0811_));
 sg13g2_o21ai_1 _2316_ (.B1(_0766_),
    .Y(_0812_),
    .A1(net93),
    .A2(_0780_));
 sg13g2_a21oi_1 _2317_ (.A1(net96),
    .A2(_0776_),
    .Y(_0813_),
    .B1(net94));
 sg13g2_nand2b_1 _2318_ (.Y(_0814_),
    .B(_0783_),
    .A_N(_0813_));
 sg13g2_o21ai_1 _2319_ (.B1(_0814_),
    .Y(_0815_),
    .A1(_0811_),
    .A2(_0812_));
 sg13g2_nand2_1 _2320_ (.Y(_0816_),
    .A(_0713_),
    .B(_0718_));
 sg13g2_a22oi_1 _2321_ (.Y(_0817_),
    .B1(_0816_),
    .B2(net102),
    .A2(_0712_),
    .A1(net100));
 sg13g2_o21ai_1 _2322_ (.B1(net88),
    .Y(_0818_),
    .A1(net103),
    .A2(net100));
 sg13g2_or2_1 _2323_ (.X(_0819_),
    .B(net102),
    .A(net103));
 sg13g2_a21oi_1 _2324_ (.A1(_0714_),
    .A2(_0819_),
    .Y(_0820_),
    .B1(net101));
 sg13g2_nor2_1 _2325_ (.A(_0818_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_nand2_1 _2326_ (.Y(_0822_),
    .A(_0809_),
    .B(_0821_));
 sg13g2_a21oi_1 _2327_ (.A1(_0690_),
    .A2(_0817_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_a221oi_1 _2328_ (.B2(net82),
    .C1(_0823_),
    .B1(_0815_),
    .A1(_0776_),
    .Y(_0824_),
    .A2(_0805_));
 sg13g2_buf_2 _2329_ (.A(\tokenflow_inst.i6.ydata[24] ),
    .X(_0825_));
 sg13g2_buf_2 _2330_ (.A(\tokenflow_inst.i6.ydata[76] ),
    .X(_0826_));
 sg13g2_nand2_1 _2331_ (.Y(_0827_),
    .A(net86),
    .B(_0826_));
 sg13g2_xnor2_1 _2332_ (.Y(_0828_),
    .A(_0825_),
    .B(_0827_));
 sg13g2_a21o_1 _2333_ (.A2(_0824_),
    .A1(_0810_),
    .B1(_0828_),
    .X(_0829_));
 sg13g2_nand3_1 _2334_ (.B(_0824_),
    .C(_0828_),
    .A(_0810_),
    .Y(_0830_));
 sg13g2_a21oi_1 _2335_ (.A1(_0829_),
    .A2(_0830_),
    .Y(_0256_),
    .B1(net167));
 sg13g2_nand2_1 _2336_ (.Y(_0831_),
    .A(net86),
    .B(\tokenflow_inst.i6.ydata[77] ));
 sg13g2_xor2_1 _2337_ (.B(_0831_),
    .A(\tokenflow_inst.i6.ydata[25] ),
    .X(_0832_));
 sg13g2_and2_1 _2338_ (.A(net182),
    .B(_0832_),
    .X(_0833_));
 sg13g2_nor2_1 _2339_ (.A(net179),
    .B(_0832_),
    .Y(_0834_));
 sg13g2_nor2b_1 _2340_ (.A(_0825_),
    .B_N(_0826_),
    .Y(_0835_));
 sg13g2_xor2_1 _2341_ (.B(_0825_),
    .A(_0826_),
    .X(_0836_));
 sg13g2_a22oi_1 _2342_ (.Y(_0837_),
    .B1(_0836_),
    .B2(_0801_),
    .A2(_0835_),
    .A1(_0802_));
 sg13g2_o21ai_1 _2343_ (.B1(net86),
    .Y(_0838_),
    .A1(net93),
    .A2(_0826_));
 sg13g2_nand3_1 _2344_ (.B(_0825_),
    .C(_0838_),
    .A(net94),
    .Y(_0839_));
 sg13g2_o21ai_1 _2345_ (.B1(_0839_),
    .Y(_0840_),
    .A1(net83),
    .A2(_0837_));
 sg13g2_nor2_1 _2346_ (.A(_0826_),
    .B(_0825_),
    .Y(_0841_));
 sg13g2_o21ai_1 _2347_ (.B1(_0796_),
    .Y(_0842_),
    .A1(net93),
    .A2(net94));
 sg13g2_inv_1 _2348_ (.Y(_0843_),
    .A(_0842_));
 sg13g2_a221oi_1 _2349_ (.B2(_0825_),
    .C1(_0843_),
    .B1(_0826_),
    .A1(net93),
    .Y(_0844_),
    .A2(net94));
 sg13g2_nor3_1 _2350_ (.A(net83),
    .B(_0841_),
    .C(_0844_),
    .Y(_0845_));
 sg13g2_a21oi_1 _2351_ (.A1(_0793_),
    .A2(_0840_),
    .Y(_0846_),
    .B1(_0845_));
 sg13g2_mux2_1 _2352_ (.A0(_0833_),
    .A1(_0834_),
    .S(_0846_),
    .X(_0257_));
 sg13g2_and2_1 _2353_ (.A(_1449_),
    .B(\tokenflow_inst.i6.ydata[27] ),
    .X(_0258_));
 sg13g2_and2_1 _2354_ (.A(_1449_),
    .B(\tokenflow_inst.i6.ydata[28] ),
    .X(_0259_));
 sg13g2_buf_1 _2355_ (.A(net180),
    .X(_0847_));
 sg13g2_and2_1 _2356_ (.A(_0847_),
    .B(\tokenflow_inst.i6.ydata[29] ),
    .X(_0260_));
 sg13g2_and2_1 _2357_ (.A(_0847_),
    .B(\tokenflow_inst.i6.ydata[30] ),
    .X(_0261_));
 sg13g2_and2_1 _2358_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[31] ),
    .X(_0263_));
 sg13g2_and2_1 _2359_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[32] ),
    .X(_0264_));
 sg13g2_and2_1 _2360_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[33] ),
    .X(_0265_));
 sg13g2_and2_1 _2361_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[34] ),
    .X(_0266_));
 sg13g2_and2_1 _2362_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[35] ),
    .X(_0267_));
 sg13g2_and2_1 _2363_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[36] ),
    .X(_0268_));
 sg13g2_and2_1 _2364_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[37] ),
    .X(_0269_));
 sg13g2_and2_1 _2365_ (.A(net163),
    .B(\tokenflow_inst.i6.ydata[38] ),
    .X(_0270_));
 sg13g2_buf_1 _2366_ (.A(net180),
    .X(_0848_));
 sg13g2_and2_1 _2367_ (.A(_0848_),
    .B(\tokenflow_inst.i6.ydata[39] ),
    .X(_0271_));
 sg13g2_and2_1 _2368_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[40] ),
    .X(_0272_));
 sg13g2_and2_1 _2369_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[41] ),
    .X(_0274_));
 sg13g2_and2_1 _2370_ (.A(_0848_),
    .B(\tokenflow_inst.i6.ydata[42] ),
    .X(_0275_));
 sg13g2_and2_1 _2371_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[43] ),
    .X(_0276_));
 sg13g2_and2_1 _2372_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[44] ),
    .X(_0277_));
 sg13g2_and2_1 _2373_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[45] ),
    .X(_0278_));
 sg13g2_and2_1 _2374_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[46] ),
    .X(_0279_));
 sg13g2_and2_1 _2375_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[47] ),
    .X(_0280_));
 sg13g2_and2_1 _2376_ (.A(net162),
    .B(\tokenflow_inst.i6.ydata[48] ),
    .X(_0281_));
 sg13g2_buf_1 _2377_ (.A(net180),
    .X(_0849_));
 sg13g2_and2_1 _2378_ (.A(net161),
    .B(\tokenflow_inst.i6.ydata[49] ),
    .X(_0282_));
 sg13g2_and2_1 _2379_ (.A(net161),
    .B(\tokenflow_inst.i6.ydata[50] ),
    .X(_0283_));
 sg13g2_and2_1 _2380_ (.A(_0849_),
    .B(\tokenflow_inst.i6.ydata[51] ),
    .X(_0285_));
 sg13g2_and2_1 _2381_ (.A(net161),
    .B(\tokenflow_inst.i6.ydata[52] ),
    .X(_0286_));
 sg13g2_and2_1 _2382_ (.A(net161),
    .B(_0365_),
    .X(_0287_));
 sg13g2_and2_1 _2383_ (.A(net161),
    .B(\tokenflow_inst.i6.ydata[54] ),
    .X(_0288_));
 sg13g2_and2_1 _2384_ (.A(net161),
    .B(_0381_),
    .X(_0289_));
 sg13g2_and2_1 _2385_ (.A(net161),
    .B(_0391_),
    .X(_0290_));
 sg13g2_and2_1 _2386_ (.A(net161),
    .B(_0412_),
    .X(_0291_));
 sg13g2_nor2_1 _2387_ (.A(_0605_),
    .B(_0419_),
    .Y(_0292_));
 sg13g2_and2_1 _2388_ (.A(_0849_),
    .B(_0448_),
    .X(_0294_));
 sg13g2_buf_1 _2389_ (.A(_1386_),
    .X(_0850_));
 sg13g2_and2_1 _2390_ (.A(_0850_),
    .B(_0453_),
    .X(_0295_));
 sg13g2_and2_1 _2391_ (.A(net160),
    .B(net116),
    .X(_0296_));
 sg13g2_nor2_1 _2392_ (.A(_0605_),
    .B(_0525_),
    .Y(_0297_));
 sg13g2_and2_1 _2393_ (.A(net160),
    .B(net91),
    .X(_0298_));
 sg13g2_and2_1 _2394_ (.A(_0850_),
    .B(net112),
    .X(_0299_));
 sg13g2_and2_1 _2395_ (.A(net160),
    .B(_0577_),
    .X(_0300_));
 sg13g2_and2_1 _2396_ (.A(net160),
    .B(net108),
    .X(_0301_));
 sg13g2_and2_1 _2397_ (.A(net160),
    .B(net106),
    .X(_0302_));
 sg13g2_nor2_1 _2398_ (.A(net145),
    .B(_0638_),
    .Y(_0303_));
 sg13g2_and2_1 _2399_ (.A(net160),
    .B(net104),
    .X(_0305_));
 sg13g2_and2_1 _2400_ (.A(net160),
    .B(_0691_),
    .X(_0306_));
 sg13g2_and2_1 _2401_ (.A(net160),
    .B(net100),
    .X(_0307_));
 sg13g2_buf_1 _2402_ (.A(net180),
    .X(_0851_));
 sg13g2_and2_1 _2403_ (.A(net159),
    .B(net98),
    .X(_0308_));
 sg13g2_and2_1 _2404_ (.A(net159),
    .B(_0754_),
    .X(_0309_));
 sg13g2_and2_1 _2405_ (.A(net159),
    .B(net95),
    .X(_0310_));
 sg13g2_buf_1 _2406_ (.A(net164),
    .X(_0852_));
 sg13g2_nor2_1 _2407_ (.A(net144),
    .B(_0784_),
    .Y(_0311_));
 sg13g2_and2_1 _2408_ (.A(net159),
    .B(_0826_),
    .X(_0312_));
 sg13g2_and2_1 _2409_ (.A(net159),
    .B(\tokenflow_inst.i8.ydata[0] ),
    .X(_0165_));
 sg13g2_buf_1 _2410_ (.A(\tokenflow_inst.i8.ydata[26] ),
    .X(_0853_));
 sg13g2_buf_1 _2411_ (.A(net68),
    .X(_0854_));
 sg13g2_buf_1 _2412_ (.A(net50),
    .X(_0855_));
 sg13g2_buf_1 _2413_ (.A(net48),
    .X(_0856_));
 sg13g2_buf_1 _2414_ (.A(_0856_),
    .X(_0857_));
 sg13g2_nand2_1 _2415_ (.Y(_0858_),
    .A(net44),
    .B(\tokenflow_inst.i8.ydata[53] ));
 sg13g2_xor2_1 _2416_ (.B(_0858_),
    .A(\tokenflow_inst.i8.ydata[1] ),
    .X(_0859_));
 sg13g2_nor2_1 _2417_ (.A(net144),
    .B(_0859_),
    .Y(_0176_));
 sg13g2_buf_2 _2418_ (.A(\tokenflow_inst.i8.ydata[54] ),
    .X(_0860_));
 sg13g2_nand2_1 _2419_ (.Y(_0861_),
    .A(\tokenflow_inst.i8.ydata[53] ),
    .B(\tokenflow_inst.i8.ydata[1] ));
 sg13g2_xnor2_1 _2420_ (.Y(_0862_),
    .A(_0860_),
    .B(_0861_));
 sg13g2_nand2_1 _2421_ (.Y(_0863_),
    .A(net44),
    .B(_0862_));
 sg13g2_xor2_1 _2422_ (.B(_0863_),
    .A(\tokenflow_inst.i8.ydata[2] ),
    .X(_0864_));
 sg13g2_nor2_1 _2423_ (.A(net144),
    .B(_0864_),
    .Y(_0187_));
 sg13g2_inv_2 _2424_ (.Y(_0865_),
    .A(net68));
 sg13g2_buf_1 _2425_ (.A(_0865_),
    .X(_0866_));
 sg13g2_buf_1 _2426_ (.A(net47),
    .X(_0867_));
 sg13g2_nor2_1 _2427_ (.A(_0860_),
    .B(\tokenflow_inst.i8.ydata[2] ),
    .Y(_0868_));
 sg13g2_a22oi_1 _2428_ (.Y(_0869_),
    .B1(_0860_),
    .B2(\tokenflow_inst.i8.ydata[2] ),
    .A2(\tokenflow_inst.i8.ydata[1] ),
    .A1(\tokenflow_inst.i8.ydata[53] ));
 sg13g2_nor2_1 _2429_ (.A(_0868_),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_xnor2_1 _2430_ (.Y(_0871_),
    .A(\tokenflow_inst.i8.ydata[55] ),
    .B(_0870_));
 sg13g2_nor2_1 _2431_ (.A(net45),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_xnor2_1 _2432_ (.Y(_0873_),
    .A(\tokenflow_inst.i8.ydata[3] ),
    .B(_0872_));
 sg13g2_nor2_1 _2433_ (.A(net144),
    .B(_0873_),
    .Y(_0198_));
 sg13g2_inv_1 _2434_ (.Y(_0874_),
    .A(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_and2_1 _2435_ (.A(\tokenflow_inst.i8.ydata[55] ),
    .B(\tokenflow_inst.i8.ydata[3] ),
    .X(_0875_));
 sg13g2_buf_1 _2436_ (.A(_0875_),
    .X(_0876_));
 sg13g2_nor2_1 _2437_ (.A(\tokenflow_inst.i8.ydata[55] ),
    .B(\tokenflow_inst.i8.ydata[3] ),
    .Y(_0877_));
 sg13g2_nor3_2 _2438_ (.A(_0868_),
    .B(_0869_),
    .C(_0877_),
    .Y(_0878_));
 sg13g2_o21ai_1 _2439_ (.B1(\tokenflow_inst.i8.ydata[56] ),
    .Y(_0879_),
    .A1(_0876_),
    .A2(_0878_));
 sg13g2_or3_1 _2440_ (.A(\tokenflow_inst.i8.ydata[56] ),
    .B(_0876_),
    .C(_0878_),
    .X(_0880_));
 sg13g2_nand3_1 _2441_ (.B(_0879_),
    .C(_0880_),
    .A(_0857_),
    .Y(_0881_));
 sg13g2_xnor2_1 _2442_ (.Y(_0882_),
    .A(_0874_),
    .B(_0881_));
 sg13g2_nor2_1 _2443_ (.A(_0852_),
    .B(_0882_),
    .Y(_0209_));
 sg13g2_buf_1 _2444_ (.A(\tokenflow_inst.i8.ydata[5] ),
    .X(_0883_));
 sg13g2_buf_1 _2445_ (.A(\tokenflow_inst.i8.ydata[57] ),
    .X(_0884_));
 sg13g2_inv_1 _2446_ (.Y(_0885_),
    .A(\tokenflow_inst.i8.ydata[56] ));
 sg13g2_o21ai_1 _2447_ (.B1(\tokenflow_inst.i8.ydata[4] ),
    .Y(_0886_),
    .A1(_0876_),
    .A2(_0878_));
 sg13g2_nor3_1 _2448_ (.A(\tokenflow_inst.i8.ydata[4] ),
    .B(_0876_),
    .C(_0878_),
    .Y(_0887_));
 sg13g2_a21o_1 _2449_ (.A2(_0886_),
    .A1(_0885_),
    .B1(_0887_),
    .X(_0888_));
 sg13g2_xnor2_1 _2450_ (.Y(_0889_),
    .A(_0884_),
    .B(_0888_));
 sg13g2_nand2_1 _2451_ (.Y(_0890_),
    .A(_0857_),
    .B(_0889_));
 sg13g2_xor2_1 _2452_ (.B(_0890_),
    .A(_0883_),
    .X(_0891_));
 sg13g2_nor2_1 _2453_ (.A(_0852_),
    .B(_0891_),
    .Y(_0216_));
 sg13g2_nor2_1 _2454_ (.A(_0884_),
    .B(_0883_),
    .Y(_0892_));
 sg13g2_o21ai_1 _2455_ (.B1(net68),
    .Y(_0893_),
    .A1(\tokenflow_inst.i8.ydata[56] ),
    .A2(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_nor2_1 _2456_ (.A(_0892_),
    .B(_0893_),
    .Y(_0894_));
 sg13g2_o21ai_1 _2457_ (.B1(_0894_),
    .Y(_0895_),
    .A1(_0876_),
    .A2(_0878_));
 sg13g2_and2_1 _2458_ (.A(_0884_),
    .B(_0883_),
    .X(_0896_));
 sg13g2_nor3_1 _2459_ (.A(_0885_),
    .B(_0874_),
    .C(_0892_),
    .Y(_0897_));
 sg13g2_o21ai_1 _2460_ (.B1(net68),
    .Y(_0898_),
    .A1(_0896_),
    .A2(_0897_));
 sg13g2_nand2_1 _2461_ (.Y(_0899_),
    .A(_0895_),
    .B(_0898_));
 sg13g2_buf_2 _2462_ (.A(\tokenflow_inst.i8.ydata[6] ),
    .X(_0900_));
 sg13g2_buf_1 _2463_ (.A(net46),
    .X(_0901_));
 sg13g2_buf_2 _2464_ (.A(\tokenflow_inst.i8.ydata[58] ),
    .X(_0902_));
 sg13g2_nand2_1 _2465_ (.Y(_0903_),
    .A(net43),
    .B(_0902_));
 sg13g2_xnor2_1 _2466_ (.Y(_0904_),
    .A(_0900_),
    .B(_0903_));
 sg13g2_xnor2_1 _2467_ (.Y(_0905_),
    .A(_0899_),
    .B(_0904_));
 sg13g2_nor2_1 _2468_ (.A(net144),
    .B(_0905_),
    .Y(_0227_));
 sg13g2_buf_1 _2469_ (.A(\tokenflow_inst.i8.ydata[7] ),
    .X(_0906_));
 sg13g2_buf_2 _2470_ (.A(\tokenflow_inst.i8.ydata[59] ),
    .X(_0907_));
 sg13g2_nor2_1 _2471_ (.A(_0902_),
    .B(_0900_),
    .Y(_0908_));
 sg13g2_and2_1 _2472_ (.A(_0902_),
    .B(_0900_),
    .X(_0909_));
 sg13g2_buf_1 _2473_ (.A(_0909_),
    .X(_0910_));
 sg13g2_nor2_1 _2474_ (.A(_0896_),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_or2_1 _2475_ (.X(_0912_),
    .B(_0911_),
    .A(_0908_));
 sg13g2_nand2_1 _2476_ (.Y(_0913_),
    .A(_0883_),
    .B(_0902_));
 sg13g2_o21ai_1 _2477_ (.B1(_0884_),
    .Y(_0914_),
    .A1(_0902_),
    .A2(_0900_));
 sg13g2_a21oi_1 _2478_ (.A1(_0913_),
    .A2(_0914_),
    .Y(_0915_),
    .B1(_0865_));
 sg13g2_a21o_1 _2479_ (.A2(_0902_),
    .A1(_0884_),
    .B1(_0900_),
    .X(_0916_));
 sg13g2_a21o_1 _2480_ (.A2(_0916_),
    .A1(_0883_),
    .B1(_0910_),
    .X(_0917_));
 sg13g2_nor2_1 _2481_ (.A(_0915_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_a21oi_1 _2482_ (.A1(_0888_),
    .A2(_0912_),
    .Y(_0919_),
    .B1(_0918_));
 sg13g2_xnor2_1 _2483_ (.Y(_0920_),
    .A(_0907_),
    .B(_0919_));
 sg13g2_nor2_1 _2484_ (.A(net45),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_xnor2_1 _2485_ (.Y(_0922_),
    .A(net67),
    .B(_0921_));
 sg13g2_nor2_1 _2486_ (.A(net144),
    .B(_0922_),
    .Y(_0236_));
 sg13g2_and2_1 _2487_ (.A(_0900_),
    .B(_0907_),
    .X(_0923_));
 sg13g2_nand3b_1 _2488_ (.B(_0895_),
    .C(_0898_),
    .Y(_0924_),
    .A_N(_0900_));
 sg13g2_nor2_1 _2489_ (.A(_0907_),
    .B(net67),
    .Y(_0925_));
 sg13g2_nor2b_1 _2490_ (.A(_0925_),
    .B_N(_0902_),
    .Y(_0926_));
 sg13g2_and2_1 _2491_ (.A(_0907_),
    .B(net67),
    .X(_0927_));
 sg13g2_a221oi_1 _2492_ (.B2(_0926_),
    .C1(_0927_),
    .B1(_0924_),
    .A1(_0899_),
    .Y(_0928_),
    .A2(_0923_));
 sg13g2_and2_1 _2493_ (.A(_0900_),
    .B(net67),
    .X(_0929_));
 sg13g2_nand2_1 _2494_ (.Y(_0930_),
    .A(_0899_),
    .B(_0929_));
 sg13g2_o21ai_1 _2495_ (.B1(_0930_),
    .Y(_0931_),
    .A1(_0867_),
    .A2(_0928_));
 sg13g2_buf_2 _2496_ (.A(\tokenflow_inst.i8.ydata[8] ),
    .X(_0932_));
 sg13g2_buf_2 _2497_ (.A(\tokenflow_inst.i8.ydata[60] ),
    .X(_0933_));
 sg13g2_nand2_1 _2498_ (.Y(_0934_),
    .A(net43),
    .B(_0933_));
 sg13g2_xnor2_1 _2499_ (.Y(_0935_),
    .A(_0932_),
    .B(_0934_));
 sg13g2_xnor2_1 _2500_ (.Y(_0936_),
    .A(_0931_),
    .B(_0935_));
 sg13g2_nor2_1 _2501_ (.A(net144),
    .B(_0936_),
    .Y(_0237_));
 sg13g2_nor2_1 _2502_ (.A(net67),
    .B(_0919_),
    .Y(_0937_));
 sg13g2_a21oi_1 _2503_ (.A1(net67),
    .A2(_0919_),
    .Y(_0938_),
    .B1(_0907_));
 sg13g2_nand2_2 _2504_ (.Y(_0939_),
    .A(_0933_),
    .B(_0932_));
 sg13g2_o21ai_1 _2505_ (.B1(_0939_),
    .Y(_0940_),
    .A1(_0937_),
    .A2(_0938_));
 sg13g2_or2_1 _2506_ (.X(_0941_),
    .B(_0932_),
    .A(_0933_));
 sg13g2_buf_1 _2507_ (.A(_0941_),
    .X(_0942_));
 sg13g2_nand2_1 _2508_ (.Y(_0943_),
    .A(_1377_),
    .B(_0856_));
 sg13g2_buf_2 _2509_ (.A(\tokenflow_inst.i8.ydata[61] ),
    .X(_0944_));
 sg13g2_buf_1 _2510_ (.A(\tokenflow_inst.i8.ydata[9] ),
    .X(_0945_));
 sg13g2_nor2_1 _2511_ (.A(_0944_),
    .B(net66),
    .Y(_0946_));
 sg13g2_nor2b_1 _2512_ (.A(_0943_),
    .B_N(_0946_),
    .Y(_0947_));
 sg13g2_nand3_1 _2513_ (.B(_0942_),
    .C(_0947_),
    .A(_0940_),
    .Y(_0948_));
 sg13g2_and2_1 _2514_ (.A(_1378_),
    .B(_0944_),
    .X(_0219_));
 sg13g2_nand4_1 _2515_ (.B(_0940_),
    .C(_0942_),
    .A(net66),
    .Y(_0949_),
    .D(_0219_));
 sg13g2_nor2b_1 _2516_ (.A(net66),
    .B_N(_0944_),
    .Y(_0950_));
 sg13g2_nand2b_1 _2517_ (.Y(_0951_),
    .B(_0950_),
    .A_N(_0943_));
 sg13g2_nor2_1 _2518_ (.A(net179),
    .B(_0944_),
    .Y(_0952_));
 sg13g2_nand2_1 _2519_ (.Y(_0953_),
    .A(net66),
    .B(_0952_));
 sg13g2_a21o_1 _2520_ (.A2(_0953_),
    .A1(_0951_),
    .B1(_0940_),
    .X(_0954_));
 sg13g2_nor2_1 _2521_ (.A(net179),
    .B(net44),
    .Y(_0955_));
 sg13g2_nor2_1 _2522_ (.A(_0933_),
    .B(_0932_),
    .Y(_0956_));
 sg13g2_nand3_1 _2523_ (.B(_0956_),
    .C(_0952_),
    .A(net66),
    .Y(_0957_));
 sg13g2_o21ai_1 _2524_ (.B1(_0957_),
    .Y(_0958_),
    .A1(_0942_),
    .A2(_0951_));
 sg13g2_a21oi_1 _2525_ (.A1(net66),
    .A2(_0955_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nand4_1 _2526_ (.B(_0949_),
    .C(_0954_),
    .A(_0948_),
    .Y(_0238_),
    .D(_0959_));
 sg13g2_nand2_1 _2527_ (.Y(_0960_),
    .A(_0944_),
    .B(net66));
 sg13g2_o21ai_1 _2528_ (.B1(_0960_),
    .Y(_0961_),
    .A1(_0939_),
    .A2(_0946_));
 sg13g2_nor2b_1 _2529_ (.A(_0933_),
    .B_N(_0932_),
    .Y(_0962_));
 sg13g2_xor2_1 _2530_ (.B(_0945_),
    .A(_0944_),
    .X(_0963_));
 sg13g2_nor2b_1 _2531_ (.A(_0932_),
    .B_N(_0933_),
    .Y(_0964_));
 sg13g2_a22oi_1 _2532_ (.Y(_0965_),
    .B1(_0963_),
    .B2(_0964_),
    .A2(_0962_),
    .A1(_0950_));
 sg13g2_o21ai_1 _2533_ (.B1(\tokenflow_inst.i8.ydata[26] ),
    .Y(_0966_),
    .A1(_0933_),
    .A2(_0944_));
 sg13g2_nand3_1 _2534_ (.B(net66),
    .C(_0966_),
    .A(_0932_),
    .Y(_0967_));
 sg13g2_o21ai_1 _2535_ (.B1(_0906_),
    .Y(_0968_),
    .A1(_0907_),
    .A2(_0910_));
 sg13g2_nand2_1 _2536_ (.Y(_0969_),
    .A(_0907_),
    .B(_0910_));
 sg13g2_a221oi_1 _2537_ (.B2(_0969_),
    .C1(net47),
    .B1(_0968_),
    .A1(_0965_),
    .Y(_0970_),
    .A2(_0967_));
 sg13g2_a21o_1 _2538_ (.A2(_0961_),
    .A1(_0854_),
    .B1(_0970_),
    .X(_0971_));
 sg13g2_nand2b_1 _2539_ (.Y(_0972_),
    .B(net68),
    .A_N(_0965_));
 sg13g2_nor4_1 _2540_ (.A(_0908_),
    .B(_0910_),
    .C(_0927_),
    .D(_0925_),
    .Y(_0973_));
 sg13g2_a21oi_1 _2541_ (.A1(net47),
    .A2(_0929_),
    .Y(_0974_),
    .B1(_0973_));
 sg13g2_a221oi_1 _2542_ (.B2(_0967_),
    .C1(_0974_),
    .B1(_0972_),
    .A1(_0895_),
    .Y(_0975_),
    .A2(_0898_));
 sg13g2_nor2_1 _2543_ (.A(_0971_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_buf_1 _2544_ (.A(\tokenflow_inst.i8.ydata[10] ),
    .X(_0977_));
 sg13g2_buf_1 _2545_ (.A(\tokenflow_inst.i8.ydata[62] ),
    .X(_0978_));
 sg13g2_nand2_1 _2546_ (.Y(_0979_),
    .A(_0901_),
    .B(_0978_));
 sg13g2_xor2_1 _2547_ (.B(_0979_),
    .A(_0977_),
    .X(_0980_));
 sg13g2_xnor2_1 _2548_ (.Y(_0981_),
    .A(_0976_),
    .B(_0980_));
 sg13g2_nor2_1 _2549_ (.A(net144),
    .B(_0981_),
    .Y(_0166_));
 sg13g2_buf_1 _2550_ (.A(_1456_),
    .X(_0982_));
 sg13g2_buf_2 _2551_ (.A(\tokenflow_inst.i8.ydata[11] ),
    .X(_0983_));
 sg13g2_nand2b_1 _2552_ (.Y(_0984_),
    .B(_0939_),
    .A_N(_0927_));
 sg13g2_nor2_1 _2553_ (.A(_0908_),
    .B(_0911_),
    .Y(_0985_));
 sg13g2_a21oi_1 _2554_ (.A1(_0942_),
    .A2(_0984_),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_nor2b_1 _2555_ (.A(_0978_),
    .B_N(_0977_),
    .Y(_0987_));
 sg13g2_nor2b_1 _2556_ (.A(_0977_),
    .B_N(_0978_),
    .Y(_0988_));
 sg13g2_or2_1 _2557_ (.X(_0989_),
    .B(_0988_),
    .A(_0987_));
 sg13g2_nand3_1 _2558_ (.B(_0963_),
    .C(_0989_),
    .A(net50),
    .Y(_0990_));
 sg13g2_a21oi_1 _2559_ (.A1(_0888_),
    .A2(_0986_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_inv_1 _2560_ (.Y(_0992_),
    .A(_0907_));
 sg13g2_o21ai_1 _2561_ (.B1(net67),
    .Y(_0993_),
    .A1(_0915_),
    .A2(_0917_));
 sg13g2_nor3_1 _2562_ (.A(net67),
    .B(_0915_),
    .C(_0917_),
    .Y(_0994_));
 sg13g2_a21o_1 _2563_ (.A2(_0993_),
    .A1(_0992_),
    .B1(_0994_),
    .X(_0995_));
 sg13g2_a21oi_1 _2564_ (.A1(_0939_),
    .A2(_0995_),
    .Y(_0996_),
    .B1(_0956_));
 sg13g2_nand2_1 _2565_ (.Y(_0997_),
    .A(_0991_),
    .B(_0996_));
 sg13g2_nor2_1 _2566_ (.A(_0978_),
    .B(_0977_),
    .Y(_0998_));
 sg13g2_nand2_1 _2567_ (.Y(_0999_),
    .A(_0978_),
    .B(_0977_));
 sg13g2_o21ai_1 _2568_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_0960_),
    .A2(_0998_));
 sg13g2_buf_1 _2569_ (.A(_1000_),
    .X(_1001_));
 sg13g2_buf_1 _2570_ (.A(\tokenflow_inst.i8.ydata[63] ),
    .X(_1002_));
 sg13g2_nor2b_1 _2571_ (.A(_1001_),
    .B_N(net65),
    .Y(_1003_));
 sg13g2_nor2b_1 _2572_ (.A(net65),
    .B_N(_1001_),
    .Y(_1004_));
 sg13g2_a21o_1 _2573_ (.A2(_1003_),
    .A1(_0997_),
    .B1(_1004_),
    .X(_1005_));
 sg13g2_a21oi_1 _2574_ (.A1(net43),
    .A2(net65),
    .Y(_1006_),
    .B1(_0997_));
 sg13g2_a21oi_1 _2575_ (.A1(net44),
    .A2(_1005_),
    .Y(_1007_),
    .B1(_1006_));
 sg13g2_xor2_1 _2576_ (.B(_1007_),
    .A(_0983_),
    .X(_1008_));
 sg13g2_nor2_1 _2577_ (.A(net143),
    .B(_1008_),
    .Y(_0167_));
 sg13g2_nand2_1 _2578_ (.Y(_1009_),
    .A(_0972_),
    .B(_0967_));
 sg13g2_nor2b_1 _2579_ (.A(_0983_),
    .B_N(\tokenflow_inst.i8.ydata[63] ),
    .Y(_1010_));
 sg13g2_xor2_1 _2580_ (.B(_0983_),
    .A(net65),
    .X(_1011_));
 sg13g2_a22oi_1 _2581_ (.Y(_1012_),
    .B1(_1011_),
    .B2(_0988_),
    .A2(_1010_),
    .A1(_0987_));
 sg13g2_o21ai_1 _2582_ (.B1(_0853_),
    .Y(_1013_),
    .A1(_0978_),
    .A2(net65));
 sg13g2_nand3_1 _2583_ (.B(_0983_),
    .C(_1013_),
    .A(_0977_),
    .Y(_1014_));
 sg13g2_o21ai_1 _2584_ (.B1(_1014_),
    .Y(_1015_),
    .A1(_0865_),
    .A2(_1012_));
 sg13g2_buf_1 _2585_ (.A(_1015_),
    .X(_1016_));
 sg13g2_and2_1 _2586_ (.A(_1009_),
    .B(_1016_),
    .X(_1017_));
 sg13g2_nor2_1 _2587_ (.A(net65),
    .B(_0983_),
    .Y(_1018_));
 sg13g2_nand2_1 _2588_ (.Y(_1019_),
    .A(net65),
    .B(_0983_));
 sg13g2_o21ai_1 _2589_ (.B1(_1019_),
    .Y(_1020_),
    .A1(_0999_),
    .A2(_1018_));
 sg13g2_a21oi_1 _2590_ (.A1(_0961_),
    .A2(_1016_),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_nor2_1 _2591_ (.A(_0867_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_a21o_1 _2592_ (.A2(_1017_),
    .A1(_0931_),
    .B1(_1022_),
    .X(_1023_));
 sg13g2_buf_1 _2593_ (.A(\tokenflow_inst.i8.ydata[64] ),
    .X(_1024_));
 sg13g2_buf_1 _2594_ (.A(\tokenflow_inst.i8.ydata[12] ),
    .X(_1025_));
 sg13g2_and2_1 _2595_ (.A(net64),
    .B(net63),
    .X(_1026_));
 sg13g2_buf_1 _2596_ (.A(_1026_),
    .X(_1027_));
 sg13g2_a21oi_1 _2597_ (.A1(net44),
    .A2(net64),
    .Y(_1028_),
    .B1(net63));
 sg13g2_a21oi_1 _2598_ (.A1(net44),
    .A2(_1027_),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_xnor2_1 _2599_ (.Y(_1030_),
    .A(_1023_),
    .B(_1029_));
 sg13g2_nor2_1 _2600_ (.A(net143),
    .B(_1030_),
    .Y(_0168_));
 sg13g2_nor2_1 _2601_ (.A(net64),
    .B(net63),
    .Y(_1031_));
 sg13g2_nor3_1 _2602_ (.A(_0865_),
    .B(_1018_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_nand2_1 _2603_ (.Y(_1033_),
    .A(_1001_),
    .B(_1032_));
 sg13g2_nor3_1 _2604_ (.A(net47),
    .B(_1019_),
    .C(_1031_),
    .Y(_1034_));
 sg13g2_a21oi_1 _2605_ (.A1(net50),
    .A2(_1027_),
    .Y(_1035_),
    .B1(_1034_));
 sg13g2_nand2_1 _2606_ (.Y(_1036_),
    .A(_1033_),
    .B(_1035_));
 sg13g2_nor2b_1 _2607_ (.A(_1002_),
    .B_N(_0983_),
    .Y(_1037_));
 sg13g2_nor2b_1 _2608_ (.A(_1025_),
    .B_N(net64),
    .Y(_1038_));
 sg13g2_xor2_1 _2609_ (.B(net63),
    .A(net64),
    .X(_1039_));
 sg13g2_a22oi_1 _2610_ (.Y(_1040_),
    .B1(_1039_),
    .B2(_1010_),
    .A2(_1038_),
    .A1(_1037_));
 sg13g2_o21ai_1 _2611_ (.B1(_0853_),
    .Y(_1041_),
    .A1(_1002_),
    .A2(_1024_));
 sg13g2_nand3_1 _2612_ (.B(net63),
    .C(_1041_),
    .A(_0983_),
    .Y(_1042_));
 sg13g2_o21ai_1 _2613_ (.B1(_1042_),
    .Y(_1043_),
    .A1(net47),
    .A2(_1040_));
 sg13g2_nor2b_1 _2614_ (.A(_0997_),
    .B_N(_1043_),
    .Y(_1044_));
 sg13g2_nor2_1 _2615_ (.A(_1036_),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_buf_1 _2616_ (.A(\tokenflow_inst.i8.ydata[13] ),
    .X(_1046_));
 sg13g2_buf_1 _2617_ (.A(\tokenflow_inst.i8.ydata[65] ),
    .X(_1047_));
 sg13g2_nand2_1 _2618_ (.Y(_1048_),
    .A(_0901_),
    .B(net61));
 sg13g2_xor2_1 _2619_ (.B(_1048_),
    .A(net62),
    .X(_1049_));
 sg13g2_xnor2_1 _2620_ (.Y(_1050_),
    .A(_1045_),
    .B(_1049_));
 sg13g2_nor2_1 _2621_ (.A(_0982_),
    .B(_1050_),
    .Y(_0169_));
 sg13g2_nor2b_1 _2622_ (.A(net64),
    .B_N(net63),
    .Y(_1051_));
 sg13g2_nor2b_1 _2623_ (.A(net62),
    .B_N(\tokenflow_inst.i8.ydata[65] ),
    .Y(_1052_));
 sg13g2_xor2_1 _2624_ (.B(net62),
    .A(net61),
    .X(_1053_));
 sg13g2_a22oi_1 _2625_ (.Y(_1054_),
    .B1(_1053_),
    .B2(_1038_),
    .A2(_1052_),
    .A1(_1051_));
 sg13g2_o21ai_1 _2626_ (.B1(net68),
    .Y(_1055_),
    .A1(net64),
    .A2(_1047_));
 sg13g2_nand3_1 _2627_ (.B(_1046_),
    .C(_1055_),
    .A(net63),
    .Y(_1056_));
 sg13g2_o21ai_1 _2628_ (.B1(_1056_),
    .Y(_1057_),
    .A1(_0865_),
    .A2(_1054_));
 sg13g2_nand2_1 _2629_ (.Y(_1058_),
    .A(_1016_),
    .B(_1057_));
 sg13g2_nor2_1 _2630_ (.A(net61),
    .B(net62),
    .Y(_1059_));
 sg13g2_or2_1 _2631_ (.X(_1060_),
    .B(net63),
    .A(net64));
 sg13g2_a21oi_1 _2632_ (.A1(_1020_),
    .A2(_1060_),
    .Y(_1061_),
    .B1(_1027_));
 sg13g2_nand2_1 _2633_ (.Y(_1062_),
    .A(net61),
    .B(net62));
 sg13g2_o21ai_1 _2634_ (.B1(_1062_),
    .Y(_1063_),
    .A1(_1059_),
    .A2(_1061_));
 sg13g2_nand2_1 _2635_ (.Y(_1064_),
    .A(net44),
    .B(_1063_));
 sg13g2_o21ai_1 _2636_ (.B1(_1064_),
    .Y(_1065_),
    .A1(_0976_),
    .A2(_1058_));
 sg13g2_buf_1 _2637_ (.A(\tokenflow_inst.i8.ydata[14] ),
    .X(_1066_));
 sg13g2_buf_1 _2638_ (.A(\tokenflow_inst.i8.ydata[66] ),
    .X(_1067_));
 sg13g2_buf_1 _2639_ (.A(_1067_),
    .X(_1068_));
 sg13g2_nand2_1 _2640_ (.Y(_1069_),
    .A(net43),
    .B(net49));
 sg13g2_xnor2_1 _2641_ (.Y(_1070_),
    .A(net60),
    .B(_1069_));
 sg13g2_xnor2_1 _2642_ (.Y(_1071_),
    .A(_1065_),
    .B(_1070_));
 sg13g2_nor2_1 _2643_ (.A(_0982_),
    .B(_1071_),
    .Y(_0170_));
 sg13g2_and2_1 _2644_ (.A(net62),
    .B(net60),
    .X(_1072_));
 sg13g2_nor2b_1 _2645_ (.A(net61),
    .B_N(_1046_),
    .Y(_1073_));
 sg13g2_nor2b_1 _2646_ (.A(net60),
    .B_N(_1067_),
    .Y(_1074_));
 sg13g2_xor2_1 _2647_ (.B(net60),
    .A(net49),
    .X(_1075_));
 sg13g2_a22oi_1 _2648_ (.Y(_1076_),
    .B1(_1075_),
    .B2(_1052_),
    .A2(_1074_),
    .A1(_1073_));
 sg13g2_o21ai_1 _2649_ (.B1(_0854_),
    .Y(_1077_),
    .A1(net61),
    .A2(net49));
 sg13g2_nand2_1 _2650_ (.Y(_1078_),
    .A(_1072_),
    .B(_1077_));
 sg13g2_o21ai_1 _2651_ (.B1(_1078_),
    .Y(_1079_),
    .A1(_0866_),
    .A2(_1076_));
 sg13g2_nand3_1 _2652_ (.B(_1043_),
    .C(_1079_),
    .A(_0942_),
    .Y(_1080_));
 sg13g2_a21oi_1 _2653_ (.A1(_0939_),
    .A2(_0995_),
    .Y(_1081_),
    .B1(_1080_));
 sg13g2_nand2_1 _2654_ (.Y(_1082_),
    .A(net62),
    .B(net49));
 sg13g2_o21ai_1 _2655_ (.B1(net61),
    .Y(_1083_),
    .A1(net49),
    .A2(net60));
 sg13g2_a221oi_1 _2656_ (.B2(_1001_),
    .C1(_1034_),
    .B1(_1032_),
    .A1(net50),
    .Y(_1084_),
    .A2(_1027_));
 sg13g2_a21o_1 _2657_ (.A2(_1083_),
    .A1(_1082_),
    .B1(_1084_),
    .X(_1085_));
 sg13g2_nor2_1 _2658_ (.A(_1068_),
    .B(_1066_),
    .Y(_1086_));
 sg13g2_nor2b_1 _2659_ (.A(_1086_),
    .B_N(_1047_),
    .Y(_1087_));
 sg13g2_a22oi_1 _2660_ (.Y(_1088_),
    .B1(_1087_),
    .B2(net62),
    .A2(_1066_),
    .A1(_1068_));
 sg13g2_a21oi_1 _2661_ (.A1(_1085_),
    .A2(_1088_),
    .Y(_1089_),
    .B1(_0866_));
 sg13g2_a221oi_1 _2662_ (.B2(_0991_),
    .C1(_1089_),
    .B1(_1081_),
    .A1(_1036_),
    .Y(_1090_),
    .A2(_1072_));
 sg13g2_buf_1 _2663_ (.A(_1090_),
    .X(_1091_));
 sg13g2_buf_1 _2664_ (.A(\tokenflow_inst.i8.ydata[15] ),
    .X(_1092_));
 sg13g2_buf_2 _2665_ (.A(\tokenflow_inst.i8.ydata[67] ),
    .X(_1093_));
 sg13g2_nand2_1 _2666_ (.Y(_1094_),
    .A(net48),
    .B(_1093_));
 sg13g2_xor2_1 _2667_ (.B(_1094_),
    .A(net59),
    .X(_1095_));
 sg13g2_xnor2_1 _2668_ (.Y(_1096_),
    .A(_1091_),
    .B(_1095_));
 sg13g2_nor2_1 _2669_ (.A(net143),
    .B(_1096_),
    .Y(_0171_));
 sg13g2_nor2_1 _2670_ (.A(_1093_),
    .B(net59),
    .Y(_1097_));
 sg13g2_nor2b_1 _2671_ (.A(_1027_),
    .B_N(_1062_),
    .Y(_1098_));
 sg13g2_nor3_1 _2672_ (.A(_1059_),
    .B(_1086_),
    .C(_1098_),
    .Y(_1099_));
 sg13g2_a21oi_1 _2673_ (.A1(net49),
    .A2(net60),
    .Y(_1100_),
    .B1(_1099_));
 sg13g2_nand2_1 _2674_ (.Y(_1101_),
    .A(_1093_),
    .B(net59));
 sg13g2_o21ai_1 _2675_ (.B1(_1101_),
    .Y(_1102_),
    .A1(_1097_),
    .A2(_1100_));
 sg13g2_nor2b_1 _2676_ (.A(_1067_),
    .B_N(\tokenflow_inst.i8.ydata[14] ),
    .Y(_1103_));
 sg13g2_nor2b_1 _2677_ (.A(net59),
    .B_N(_1093_),
    .Y(_1104_));
 sg13g2_xor2_1 _2678_ (.B(net59),
    .A(_1093_),
    .X(_1105_));
 sg13g2_a22oi_1 _2679_ (.Y(_1106_),
    .B1(_1105_),
    .B2(_1074_),
    .A2(_1104_),
    .A1(_1103_));
 sg13g2_o21ai_1 _2680_ (.B1(net68),
    .Y(_1107_),
    .A1(_1067_),
    .A2(_1093_));
 sg13g2_nand3_1 _2681_ (.B(net59),
    .C(_1107_),
    .A(net60),
    .Y(_1108_));
 sg13g2_o21ai_1 _2682_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_0865_),
    .A2(_1106_));
 sg13g2_and2_1 _2683_ (.A(_1057_),
    .B(_1109_),
    .X(_1110_));
 sg13g2_a22oi_1 _2684_ (.Y(_1111_),
    .B1(_1110_),
    .B2(_1023_),
    .A2(_1102_),
    .A1(net44));
 sg13g2_buf_2 _2685_ (.A(\tokenflow_inst.i8.ydata[16] ),
    .X(_1112_));
 sg13g2_buf_1 _2686_ (.A(\tokenflow_inst.i8.ydata[68] ),
    .X(_1113_));
 sg13g2_and2_1 _2687_ (.A(net48),
    .B(_1113_),
    .X(_1114_));
 sg13g2_xnor2_1 _2688_ (.Y(_1115_),
    .A(_1112_),
    .B(_1114_));
 sg13g2_xnor2_1 _2689_ (.Y(_1116_),
    .A(_1111_),
    .B(_1115_));
 sg13g2_nor2_1 _2690_ (.A(net143),
    .B(_1116_),
    .Y(_0172_));
 sg13g2_nor2_1 _2691_ (.A(_1113_),
    .B(_1112_),
    .Y(_1117_));
 sg13g2_nor2_1 _2692_ (.A(_1094_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_a22oi_1 _2693_ (.Y(_1119_),
    .B1(_1118_),
    .B2(net59),
    .A2(_1114_),
    .A1(_1112_));
 sg13g2_nand2_1 _2694_ (.Y(_1120_),
    .A(net59),
    .B(_1112_));
 sg13g2_nand2_1 _2695_ (.Y(_1121_),
    .A(_1113_),
    .B(_1112_));
 sg13g2_a22oi_1 _2696_ (.Y(_1122_),
    .B1(_1121_),
    .B2(_1097_),
    .A2(_1120_),
    .A1(net47));
 sg13g2_nand2b_1 _2697_ (.Y(_1123_),
    .B(_1122_),
    .A_N(_1117_));
 sg13g2_a21oi_1 _2698_ (.A1(_1091_),
    .A2(_1119_),
    .Y(_1124_),
    .B1(_1123_));
 sg13g2_buf_1 _2699_ (.A(\tokenflow_inst.i8.ydata[17] ),
    .X(_1125_));
 sg13g2_buf_1 _2700_ (.A(\tokenflow_inst.i8.ydata[69] ),
    .X(_1126_));
 sg13g2_nand2_1 _2701_ (.Y(_1127_),
    .A(net43),
    .B(net57));
 sg13g2_xnor2_1 _2702_ (.Y(_1128_),
    .A(net58),
    .B(_1127_));
 sg13g2_xnor2_1 _2703_ (.Y(_1129_),
    .A(_1124_),
    .B(_1128_));
 sg13g2_nor2_1 _2704_ (.A(net143),
    .B(_1129_),
    .Y(_0173_));
 sg13g2_a22oi_1 _2705_ (.Y(_1130_),
    .B1(_1093_),
    .B2(_1092_),
    .A2(net60),
    .A1(net49));
 sg13g2_o21ai_1 _2706_ (.B1(_1121_),
    .Y(_1131_),
    .A1(_1097_),
    .A2(_1130_));
 sg13g2_nor2_1 _2707_ (.A(net57),
    .B(_1125_),
    .Y(_1132_));
 sg13g2_nor2_1 _2708_ (.A(_1117_),
    .B(_1132_),
    .Y(_1133_));
 sg13g2_a22oi_1 _2709_ (.Y(_1134_),
    .B1(_1131_),
    .B2(_1133_),
    .A2(_1125_),
    .A1(net57));
 sg13g2_nor2_1 _2710_ (.A(net47),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_nor2b_1 _2711_ (.A(net58),
    .B_N(\tokenflow_inst.i8.ydata[69] ),
    .Y(_1136_));
 sg13g2_nor2b_1 _2712_ (.A(_1113_),
    .B_N(_1112_),
    .Y(_1137_));
 sg13g2_xor2_1 _2713_ (.B(net58),
    .A(net57),
    .X(_1138_));
 sg13g2_nor2b_1 _2714_ (.A(_1112_),
    .B_N(_1113_),
    .Y(_1139_));
 sg13g2_a22oi_1 _2715_ (.Y(_1140_),
    .B1(_1138_),
    .B2(_1139_),
    .A2(_1137_),
    .A1(_1136_));
 sg13g2_o21ai_1 _2716_ (.B1(net68),
    .Y(_1141_),
    .A1(_1113_),
    .A2(_1126_));
 sg13g2_nand3_1 _2717_ (.B(net58),
    .C(_1141_),
    .A(_1112_),
    .Y(_1142_));
 sg13g2_o21ai_1 _2718_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_0865_),
    .A2(_1140_));
 sg13g2_and4_1 _2719_ (.A(_1016_),
    .B(_1057_),
    .C(_1109_),
    .D(_1143_),
    .X(_1144_));
 sg13g2_o21ai_1 _2720_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_0971_),
    .A2(_0975_));
 sg13g2_nand4_1 _2721_ (.B(_1063_),
    .C(_1109_),
    .A(net50),
    .Y(_1146_),
    .D(_1143_));
 sg13g2_nand3b_1 _2722_ (.B(_1145_),
    .C(_1146_),
    .Y(_1147_),
    .A_N(_1135_));
 sg13g2_buf_1 _2723_ (.A(_1147_),
    .X(_1148_));
 sg13g2_buf_2 _2724_ (.A(\tokenflow_inst.i8.ydata[18] ),
    .X(_1149_));
 sg13g2_buf_2 _2725_ (.A(\tokenflow_inst.i8.ydata[70] ),
    .X(_1150_));
 sg13g2_nand2_1 _2726_ (.Y(_1151_),
    .A(net48),
    .B(_1150_));
 sg13g2_xnor2_1 _2727_ (.Y(_1152_),
    .A(_1149_),
    .B(_1151_));
 sg13g2_xnor2_1 _2728_ (.Y(_1153_),
    .A(_1148_),
    .B(_1152_));
 sg13g2_nor2_1 _2729_ (.A(net143),
    .B(_1153_),
    .Y(_0174_));
 sg13g2_inv_1 _2730_ (.Y(_1154_),
    .A(_1149_));
 sg13g2_a21oi_1 _2731_ (.A1(net57),
    .A2(net58),
    .Y(_1155_),
    .B1(_1150_));
 sg13g2_nand3_1 _2732_ (.B(net58),
    .C(_1150_),
    .A(net57),
    .Y(_1156_));
 sg13g2_o21ai_1 _2733_ (.B1(_1156_),
    .Y(_1157_),
    .A1(_1154_),
    .A2(_1155_));
 sg13g2_nand2_1 _2734_ (.Y(_1158_),
    .A(_0855_),
    .B(_1157_));
 sg13g2_nor2b_1 _2735_ (.A(net57),
    .B_N(net58),
    .Y(_1159_));
 sg13g2_nor2b_1 _2736_ (.A(_1149_),
    .B_N(_1150_),
    .Y(_1160_));
 sg13g2_xor2_1 _2737_ (.B(_1149_),
    .A(_1150_),
    .X(_1161_));
 sg13g2_a22oi_1 _2738_ (.Y(_1162_),
    .B1(_1161_),
    .B2(_1136_),
    .A2(_1160_),
    .A1(_1159_));
 sg13g2_o21ai_1 _2739_ (.B1(_0855_),
    .Y(_1163_),
    .A1(net57),
    .A2(_1150_));
 sg13g2_nand3_1 _2740_ (.B(_1149_),
    .C(_1163_),
    .A(net58),
    .Y(_1164_));
 sg13g2_o21ai_1 _2741_ (.B1(_1164_),
    .Y(_1165_),
    .A1(net45),
    .A2(_1162_));
 sg13g2_nand2b_1 _2742_ (.Y(_1166_),
    .B(_1165_),
    .A_N(_1123_));
 sg13g2_a21o_1 _2743_ (.A2(_1119_),
    .A1(_1091_),
    .B1(_1166_),
    .X(_1167_));
 sg13g2_nand2_1 _2744_ (.Y(_1168_),
    .A(_1158_),
    .B(_1167_));
 sg13g2_buf_1 _2745_ (.A(\tokenflow_inst.i8.ydata[19] ),
    .X(_1169_));
 sg13g2_inv_1 _2746_ (.Y(_1170_),
    .A(_1169_));
 sg13g2_buf_1 _2747_ (.A(\tokenflow_inst.i8.ydata[71] ),
    .X(_1171_));
 sg13g2_and2_1 _2748_ (.A(net50),
    .B(_1171_),
    .X(_1172_));
 sg13g2_buf_1 _2749_ (.A(_1172_),
    .X(_1173_));
 sg13g2_xnor2_1 _2750_ (.Y(_1174_),
    .A(_1170_),
    .B(_1173_));
 sg13g2_xnor2_1 _2751_ (.Y(_1175_),
    .A(_1168_),
    .B(_1174_));
 sg13g2_nor2_1 _2752_ (.A(net143),
    .B(_1175_),
    .Y(_0175_));
 sg13g2_nor2_1 _2753_ (.A(_1171_),
    .B(_1169_),
    .Y(_1176_));
 sg13g2_nor2_1 _2754_ (.A(_1151_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_and2_1 _2755_ (.A(_1149_),
    .B(_1173_),
    .X(_1178_));
 sg13g2_o21ai_1 _2756_ (.B1(_1148_),
    .Y(_1179_),
    .A1(_1177_),
    .A2(_1178_));
 sg13g2_nor2_1 _2757_ (.A(_1154_),
    .B(_1170_),
    .Y(_1180_));
 sg13g2_nor3_1 _2758_ (.A(_1154_),
    .B(_1151_),
    .C(_1176_),
    .Y(_1181_));
 sg13g2_a221oi_1 _2759_ (.B2(_1148_),
    .C1(_1181_),
    .B1(_1180_),
    .A1(_1169_),
    .Y(_1182_),
    .A2(_1173_));
 sg13g2_nand2_1 _2760_ (.Y(_1183_),
    .A(_1179_),
    .B(_1182_));
 sg13g2_buf_1 _2761_ (.A(\tokenflow_inst.i8.ydata[20] ),
    .X(_1184_));
 sg13g2_buf_1 _2762_ (.A(\tokenflow_inst.i8.ydata[72] ),
    .X(_1185_));
 sg13g2_nand2_1 _2763_ (.Y(_1186_),
    .A(net43),
    .B(net55));
 sg13g2_xnor2_1 _2764_ (.Y(_1187_),
    .A(_1184_),
    .B(_1186_));
 sg13g2_xnor2_1 _2765_ (.Y(_1188_),
    .A(_1183_),
    .B(_1187_));
 sg13g2_nor2_1 _2766_ (.A(net143),
    .B(_1188_),
    .Y(_0177_));
 sg13g2_buf_1 _2767_ (.A(net179),
    .X(_1189_));
 sg13g2_a21oi_1 _2768_ (.A1(_1091_),
    .A2(_1119_),
    .Y(_1190_),
    .B1(_1166_));
 sg13g2_nor2b_1 _2769_ (.A(net56),
    .B_N(net55),
    .Y(_1191_));
 sg13g2_nor2_1 _2770_ (.A(_1171_),
    .B(_1170_),
    .Y(_1192_));
 sg13g2_nor2b_1 _2771_ (.A(net55),
    .B_N(net56),
    .Y(_1193_));
 sg13g2_or2_1 _2772_ (.X(_1194_),
    .B(_1193_),
    .A(_1191_));
 sg13g2_nor2b_1 _2773_ (.A(_1169_),
    .B_N(_1171_),
    .Y(_1195_));
 sg13g2_a22oi_1 _2774_ (.Y(_1196_),
    .B1(_1194_),
    .B2(_1195_),
    .A2(_1192_),
    .A1(_1191_));
 sg13g2_o21ai_1 _2775_ (.B1(net48),
    .Y(_1197_),
    .A1(_1171_),
    .A2(net55));
 sg13g2_nand3_1 _2776_ (.B(net56),
    .C(_1197_),
    .A(_1169_),
    .Y(_1198_));
 sg13g2_o21ai_1 _2777_ (.B1(_1198_),
    .Y(_1199_),
    .A1(net45),
    .A2(_1196_));
 sg13g2_and2_1 _2778_ (.A(net50),
    .B(_1157_),
    .X(_1200_));
 sg13g2_a21o_1 _2779_ (.A2(_1200_),
    .A1(_1169_),
    .B1(net56),
    .X(_1201_));
 sg13g2_o21ai_1 _2780_ (.B1(_1171_),
    .Y(_1202_),
    .A1(net55),
    .A2(_1184_));
 sg13g2_a21oi_1 _2781_ (.A1(_1170_),
    .A2(_1158_),
    .Y(_1203_),
    .B1(_1202_));
 sg13g2_a21oi_1 _2782_ (.A1(_1185_),
    .A2(_1201_),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_nand3_1 _2783_ (.B(net56),
    .C(_1200_),
    .A(_1169_),
    .Y(_1205_));
 sg13g2_o21ai_1 _2784_ (.B1(_1205_),
    .Y(_1206_),
    .A1(net45),
    .A2(_1204_));
 sg13g2_a21oi_1 _2785_ (.A1(_1190_),
    .A2(_1199_),
    .Y(_1207_),
    .B1(_1206_));
 sg13g2_buf_1 _2786_ (.A(\tokenflow_inst.i8.ydata[21] ),
    .X(_1208_));
 sg13g2_inv_1 _2787_ (.Y(_1209_),
    .A(_1208_));
 sg13g2_buf_1 _2788_ (.A(\tokenflow_inst.i8.ydata[73] ),
    .X(_1210_));
 sg13g2_nand2_1 _2789_ (.Y(_1211_),
    .A(net43),
    .B(net54));
 sg13g2_xnor2_1 _2790_ (.Y(_1212_),
    .A(_1209_),
    .B(_1211_));
 sg13g2_xnor2_1 _2791_ (.Y(_1213_),
    .A(_1207_),
    .B(_1212_));
 sg13g2_nor2_1 _2792_ (.A(net158),
    .B(_1213_),
    .Y(_0178_));
 sg13g2_a21oi_1 _2793_ (.A1(net55),
    .A2(net56),
    .Y(_1214_),
    .B1(net54));
 sg13g2_nand3_1 _2794_ (.B(net56),
    .C(net54),
    .A(net55),
    .Y(_1215_));
 sg13g2_o21ai_1 _2795_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1209_),
    .A2(_1214_));
 sg13g2_nand2_1 _2796_ (.Y(_1217_),
    .A(net48),
    .B(_1216_));
 sg13g2_inv_1 _2797_ (.Y(_1218_),
    .A(_1217_));
 sg13g2_nor2b_1 _2798_ (.A(_1208_),
    .B_N(net54),
    .Y(_1219_));
 sg13g2_nor2_1 _2799_ (.A(net54),
    .B(_1209_),
    .Y(_1220_));
 sg13g2_or2_1 _2800_ (.X(_1221_),
    .B(_1220_),
    .A(_1219_));
 sg13g2_a22oi_1 _2801_ (.Y(_1222_),
    .B1(_1221_),
    .B2(_1191_),
    .A2(_1219_),
    .A1(_1193_));
 sg13g2_o21ai_1 _2802_ (.B1(net46),
    .Y(_1223_),
    .A1(net55),
    .A2(net54));
 sg13g2_nand3_1 _2803_ (.B(_1208_),
    .C(_1223_),
    .A(net56),
    .Y(_1224_));
 sg13g2_o21ai_1 _2804_ (.B1(_1224_),
    .Y(_1225_),
    .A1(net45),
    .A2(_1222_));
 sg13g2_inv_1 _2805_ (.Y(_1226_),
    .A(_1225_));
 sg13g2_a21oi_1 _2806_ (.A1(_1179_),
    .A2(_1182_),
    .Y(_1227_),
    .B1(_1226_));
 sg13g2_buf_1 _2807_ (.A(\tokenflow_inst.i8.ydata[22] ),
    .X(_1228_));
 sg13g2_inv_1 _2808_ (.Y(_1229_),
    .A(_1228_));
 sg13g2_buf_1 _2809_ (.A(\tokenflow_inst.i8.ydata[74] ),
    .X(_1230_));
 sg13g2_nand2_1 _2810_ (.Y(_1231_),
    .A(net46),
    .B(net53));
 sg13g2_xnor2_1 _2811_ (.Y(_1232_),
    .A(_1229_),
    .B(_1231_));
 sg13g2_o21ai_1 _2812_ (.B1(_1232_),
    .Y(_1233_),
    .A1(_1218_),
    .A2(_1227_));
 sg13g2_or3_1 _2813_ (.A(_1218_),
    .B(_1227_),
    .C(_1232_),
    .X(_1234_));
 sg13g2_a21oi_1 _2814_ (.A1(_1233_),
    .A2(_1234_),
    .Y(_0179_),
    .B1(net167));
 sg13g2_nor2b_1 _2815_ (.A(_1228_),
    .B_N(net53),
    .Y(_1235_));
 sg13g2_nor2_1 _2816_ (.A(net53),
    .B(_1229_),
    .Y(_1236_));
 sg13g2_or2_1 _2817_ (.X(_1237_),
    .B(_1236_),
    .A(_1235_));
 sg13g2_a22oi_1 _2818_ (.Y(_1238_),
    .B1(_1237_),
    .B2(_1219_),
    .A2(_1235_),
    .A1(_1220_));
 sg13g2_o21ai_1 _2819_ (.B1(net48),
    .Y(_1239_),
    .A1(_1210_),
    .A2(_1230_));
 sg13g2_nand3_1 _2820_ (.B(_1228_),
    .C(_1239_),
    .A(_1208_),
    .Y(_1240_));
 sg13g2_o21ai_1 _2821_ (.B1(_1240_),
    .Y(_1241_),
    .A1(net47),
    .A2(_1238_));
 sg13g2_buf_1 _2822_ (.A(_1241_),
    .X(_1242_));
 sg13g2_nand2_1 _2823_ (.Y(_1243_),
    .A(_1199_),
    .B(_1242_));
 sg13g2_a21oi_1 _2824_ (.A1(net54),
    .A2(_1208_),
    .Y(_1244_),
    .B1(net53));
 sg13g2_nand3_1 _2825_ (.B(_1208_),
    .C(net53),
    .A(net54),
    .Y(_1245_));
 sg13g2_o21ai_1 _2826_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_1229_),
    .A2(_1244_));
 sg13g2_and2_1 _2827_ (.A(net50),
    .B(_1246_),
    .X(_1247_));
 sg13g2_buf_1 _2828_ (.A(_1247_),
    .X(_1248_));
 sg13g2_a21oi_1 _2829_ (.A1(_1206_),
    .A2(_1242_),
    .Y(_1249_),
    .B1(_1248_));
 sg13g2_o21ai_1 _2830_ (.B1(_1249_),
    .Y(_1250_),
    .A1(_1167_),
    .A2(_1243_));
 sg13g2_buf_1 _2831_ (.A(\tokenflow_inst.i8.ydata[23] ),
    .X(_1251_));
 sg13g2_buf_1 _2832_ (.A(\tokenflow_inst.i8.ydata[75] ),
    .X(_1252_));
 sg13g2_nand2_1 _2833_ (.Y(_1253_),
    .A(net46),
    .B(net51));
 sg13g2_xor2_1 _2834_ (.B(_1253_),
    .A(_1251_),
    .X(_1254_));
 sg13g2_xnor2_1 _2835_ (.Y(_1255_),
    .A(_1250_),
    .B(_1254_));
 sg13g2_and2_1 _2836_ (.A(net159),
    .B(_1255_),
    .X(_0180_));
 sg13g2_a21o_1 _2837_ (.A2(_1218_),
    .A1(_1228_),
    .B1(net52),
    .X(_1256_));
 sg13g2_o21ai_1 _2838_ (.B1(net53),
    .Y(_1257_),
    .A1(net51),
    .A2(net52));
 sg13g2_a21oi_1 _2839_ (.A1(_1229_),
    .A2(_1217_),
    .Y(_1258_),
    .B1(_1257_));
 sg13g2_a21oi_1 _2840_ (.A1(net51),
    .A2(_1256_),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_nand2_1 _2841_ (.Y(_1260_),
    .A(_1228_),
    .B(net52));
 sg13g2_or2_1 _2842_ (.X(_1261_),
    .B(_1260_),
    .A(_1217_));
 sg13g2_o21ai_1 _2843_ (.B1(_1261_),
    .Y(_1262_),
    .A1(net45),
    .A2(_1259_));
 sg13g2_nor2b_1 _2844_ (.A(net52),
    .B_N(net51),
    .Y(_1263_));
 sg13g2_nor2b_1 _2845_ (.A(net51),
    .B_N(net52),
    .Y(_1264_));
 sg13g2_or2_1 _2846_ (.X(_1265_),
    .B(_1264_),
    .A(_1263_));
 sg13g2_a22oi_1 _2847_ (.Y(_1266_),
    .B1(_1265_),
    .B2(_1235_),
    .A2(_1263_),
    .A1(_1236_));
 sg13g2_nand2b_1 _2848_ (.Y(_1267_),
    .B(net46),
    .A_N(_1266_));
 sg13g2_o21ai_1 _2849_ (.B1(net46),
    .Y(_1268_),
    .A1(net53),
    .A2(net51));
 sg13g2_nand2b_1 _2850_ (.Y(_1269_),
    .B(_1268_),
    .A_N(_1260_));
 sg13g2_a221oi_1 _2851_ (.B2(_1269_),
    .C1(_1226_),
    .B1(_1267_),
    .A1(_1179_),
    .Y(_1270_),
    .A2(_1182_));
 sg13g2_buf_2 _2852_ (.A(\tokenflow_inst.i8.ydata[24] ),
    .X(_1271_));
 sg13g2_buf_2 _2853_ (.A(\tokenflow_inst.i8.ydata[76] ),
    .X(_1272_));
 sg13g2_nand2_1 _2854_ (.Y(_1273_),
    .A(net46),
    .B(_1272_));
 sg13g2_xor2_1 _2855_ (.B(_1273_),
    .A(_1271_),
    .X(_1274_));
 sg13g2_o21ai_1 _2856_ (.B1(_1274_),
    .Y(_1275_),
    .A1(_1262_),
    .A2(_1270_));
 sg13g2_or3_1 _2857_ (.A(_1274_),
    .B(_1262_),
    .C(_1270_),
    .X(_1276_));
 sg13g2_a21oi_1 _2858_ (.A1(_1275_),
    .A2(_1276_),
    .Y(_0181_),
    .B1(net167));
 sg13g2_nor2b_1 _2859_ (.A(_1271_),
    .B_N(_1272_),
    .Y(_1277_));
 sg13g2_xor2_1 _2860_ (.B(_1271_),
    .A(_1272_),
    .X(_1278_));
 sg13g2_a22oi_1 _2861_ (.Y(_1279_),
    .B1(_1278_),
    .B2(_1263_),
    .A2(_1277_),
    .A1(_1264_));
 sg13g2_o21ai_1 _2862_ (.B1(net48),
    .Y(_1280_),
    .A1(_1252_),
    .A2(_1272_));
 sg13g2_nand3_1 _2863_ (.B(_1271_),
    .C(_1280_),
    .A(net52),
    .Y(_1281_));
 sg13g2_o21ai_1 _2864_ (.B1(_1281_),
    .Y(_1282_),
    .A1(net45),
    .A2(_1279_));
 sg13g2_nand3_1 _2865_ (.B(_1242_),
    .C(_1282_),
    .A(_1199_),
    .Y(_1283_));
 sg13g2_nor2_1 _2866_ (.A(net52),
    .B(_1248_),
    .Y(_1284_));
 sg13g2_o21ai_1 _2867_ (.B1(net51),
    .Y(_1285_),
    .A1(_1272_),
    .A2(_1271_));
 sg13g2_a21oi_1 _2868_ (.A1(net52),
    .A2(_1248_),
    .Y(_1286_),
    .B1(_1271_));
 sg13g2_nand2b_1 _2869_ (.Y(_1287_),
    .B(_1272_),
    .A_N(_1286_));
 sg13g2_o21ai_1 _2870_ (.B1(_1287_),
    .Y(_1288_),
    .A1(_1284_),
    .A2(_1285_));
 sg13g2_and2_1 _2871_ (.A(_1242_),
    .B(_1282_),
    .X(_1289_));
 sg13g2_and3_1 _2872_ (.X(_1290_),
    .A(_1251_),
    .B(_1271_),
    .C(_1248_));
 sg13g2_a221oi_1 _2873_ (.B2(_1206_),
    .C1(_1290_),
    .B1(_1289_),
    .A1(net46),
    .Y(_1291_),
    .A2(_1288_));
 sg13g2_o21ai_1 _2874_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_1167_),
    .A2(_1283_));
 sg13g2_nand2_1 _2875_ (.Y(_1293_),
    .A(net43),
    .B(\tokenflow_inst.i8.ydata[77] ));
 sg13g2_xnor2_1 _2876_ (.Y(_1294_),
    .A(\tokenflow_inst.i8.ydata[25] ),
    .B(_1293_));
 sg13g2_xnor2_1 _2877_ (.Y(_1295_),
    .A(_1292_),
    .B(_1294_));
 sg13g2_nor2_1 _2878_ (.A(net158),
    .B(_1295_),
    .Y(_0182_));
 sg13g2_and2_1 _2879_ (.A(net159),
    .B(\tokenflow_inst.i8.ydata[27] ),
    .X(_0183_));
 sg13g2_and2_1 _2880_ (.A(net159),
    .B(\tokenflow_inst.i8.ydata[28] ),
    .X(_0184_));
 sg13g2_and2_1 _2881_ (.A(_0851_),
    .B(\tokenflow_inst.i8.ydata[29] ),
    .X(_0185_));
 sg13g2_and2_1 _2882_ (.A(_0851_),
    .B(\tokenflow_inst.i8.ydata[30] ),
    .X(_0186_));
 sg13g2_buf_1 _2883_ (.A(net180),
    .X(_1296_));
 sg13g2_and2_1 _2884_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[31] ),
    .X(_0188_));
 sg13g2_and2_1 _2885_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[32] ),
    .X(_0189_));
 sg13g2_and2_1 _2886_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[33] ),
    .X(_0190_));
 sg13g2_and2_1 _2887_ (.A(_1296_),
    .B(\tokenflow_inst.i8.ydata[34] ),
    .X(_0191_));
 sg13g2_and2_1 _2888_ (.A(_1296_),
    .B(\tokenflow_inst.i8.ydata[35] ),
    .X(_0192_));
 sg13g2_and2_1 _2889_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[36] ),
    .X(_0193_));
 sg13g2_and2_1 _2890_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[37] ),
    .X(_0194_));
 sg13g2_and2_1 _2891_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[38] ),
    .X(_0195_));
 sg13g2_and2_1 _2892_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[39] ),
    .X(_0196_));
 sg13g2_and2_1 _2893_ (.A(net157),
    .B(\tokenflow_inst.i8.ydata[40] ),
    .X(_0197_));
 sg13g2_buf_1 _2894_ (.A(net182),
    .X(_1297_));
 sg13g2_and2_1 _2895_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[41] ),
    .X(_0199_));
 sg13g2_and2_1 _2896_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[42] ),
    .X(_0200_));
 sg13g2_and2_1 _2897_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[43] ),
    .X(_0201_));
 sg13g2_and2_1 _2898_ (.A(_1297_),
    .B(\tokenflow_inst.i8.ydata[44] ),
    .X(_0202_));
 sg13g2_and2_1 _2899_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[45] ),
    .X(_0203_));
 sg13g2_and2_1 _2900_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[46] ),
    .X(_0204_));
 sg13g2_and2_1 _2901_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[47] ),
    .X(_0205_));
 sg13g2_and2_1 _2902_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[48] ),
    .X(_0206_));
 sg13g2_and2_1 _2903_ (.A(net178),
    .B(\tokenflow_inst.i8.ydata[49] ),
    .X(_0207_));
 sg13g2_and2_1 _2904_ (.A(_1297_),
    .B(\tokenflow_inst.i8.ydata[50] ),
    .X(_0208_));
 sg13g2_buf_1 _2905_ (.A(_1378_),
    .X(_1298_));
 sg13g2_and2_1 _2906_ (.A(net177),
    .B(\tokenflow_inst.i8.ydata[53] ),
    .X(_0210_));
 sg13g2_and2_1 _2907_ (.A(net177),
    .B(_0860_),
    .X(_0211_));
 sg13g2_and2_1 _2908_ (.A(net177),
    .B(\tokenflow_inst.i8.ydata[55] ),
    .X(_0212_));
 sg13g2_nor2_1 _2909_ (.A(net158),
    .B(_0885_),
    .Y(_0213_));
 sg13g2_and2_1 _2910_ (.A(net177),
    .B(_0884_),
    .X(_0214_));
 sg13g2_and2_1 _2911_ (.A(_1298_),
    .B(_0902_),
    .X(_0215_));
 sg13g2_nor2_1 _2912_ (.A(net158),
    .B(_0992_),
    .Y(_0217_));
 sg13g2_and2_1 _2913_ (.A(_1298_),
    .B(_0933_),
    .X(_0218_));
 sg13g2_and2_1 _2914_ (.A(net177),
    .B(_0978_),
    .X(_0220_));
 sg13g2_and2_1 _2915_ (.A(net177),
    .B(net65),
    .X(_0221_));
 sg13g2_and2_1 _2916_ (.A(net177),
    .B(_1024_),
    .X(_0222_));
 sg13g2_and2_1 _2917_ (.A(net177),
    .B(net61),
    .X(_0223_));
 sg13g2_buf_1 _2918_ (.A(net182),
    .X(_1299_));
 sg13g2_and2_1 _2919_ (.A(net176),
    .B(net49),
    .X(_0224_));
 sg13g2_and2_1 _2920_ (.A(net176),
    .B(_1093_),
    .X(_0225_));
 sg13g2_and2_1 _2921_ (.A(net176),
    .B(_1113_),
    .X(_0226_));
 sg13g2_and2_1 _2922_ (.A(net176),
    .B(_1126_),
    .X(_0228_));
 sg13g2_and2_1 _2923_ (.A(_1299_),
    .B(_1150_),
    .X(_0229_));
 sg13g2_and2_1 _2924_ (.A(_1299_),
    .B(_1171_),
    .X(_0230_));
 sg13g2_and2_1 _2925_ (.A(net176),
    .B(_1185_),
    .X(_0231_));
 sg13g2_and2_1 _2926_ (.A(net176),
    .B(_1210_),
    .X(_0232_));
 sg13g2_and2_1 _2927_ (.A(net176),
    .B(net53),
    .X(_0233_));
 sg13g2_and2_1 _2928_ (.A(net176),
    .B(net51),
    .X(_0234_));
 sg13g2_and2_1 _2929_ (.A(net181),
    .B(_1272_),
    .X(_0235_));
 sg13g2_nor2_1 _2930_ (.A(net158),
    .B(\tokenflow_inst.i6.cg_elem.q ),
    .Y(_0164_));
 sg13g2_and2_1 _2931_ (.A(\tokenflow_inst.i78.cg_elem.q ),
    .B(\tokenflow_inst.i78.d0_elem.inv_chain[3] ),
    .X(_1300_));
 sg13g2_buf_1 _2932_ (.A(_1300_),
    .X(\tokenflow_inst.i2.cg1.a ));
 sg13g2_nor2_1 _2933_ (.A(\tokenflow_inst.i6.cg_elem.q ),
    .B(\tokenflow_inst.i9.c.q ),
    .Y(\tokenflow_inst.i3.cg_elem.a ));
 sg13g2_nor2b_1 _2934_ (.A(net28),
    .B_N(\tokenflow_inst.i1.c.q ),
    .Y(_1301_));
 sg13g2_a21oi_1 _2935_ (.A1(_1395_),
    .A2(\tokenflow_inst.i2.cg1.a ),
    .Y(_1302_),
    .B1(_1301_));
 sg13g2_xnor2_1 _2936_ (.Y(_0000_),
    .A(\tokenflow_inst.i3.cg_elem.a ),
    .B(_1302_));
 sg13g2_buf_1 _2937_ (.A(\tokenflow_inst.i2.cg2.a ),
    .X(_1303_));
 sg13g2_nor2_1 _2938_ (.A(net158),
    .B(_1303_),
    .Y(_0085_));
 sg13g2_xnor2_1 _2939_ (.Y(_0001_),
    .A(\tokenflow_inst.i1.c.q ),
    .B(\tokenflow_inst.i2.cg1.a ));
 sg13g2_xor2_1 _2940_ (.B(\tokenflow_inst.i2.cg1.a ),
    .A(_1303_),
    .X(_0002_));
 sg13g2_xor2_1 _2941_ (.B(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ),
    .A(\tokenflow_inst.i11.i.d0.inv_chain[1] ),
    .X(_0003_));
 sg13g2_inv_1 _2942_ (.Y(\tokenflow_inst.i8.cg_elem.a ),
    .A(\tokenflow_inst.i78.cg_elem.q ));
 sg13g2_nand2_1 _2943_ (.Y(_1304_),
    .A(\tokenflow_inst.i6.cg_elem.q ),
    .B(\tokenflow_inst.i6.d0_elem.inv_chain[52] ));
 sg13g2_xnor2_1 _2944_ (.Y(_0004_),
    .A(\tokenflow_inst.i8.cg_elem.a ),
    .B(_1304_));
 sg13g2_nor2_1 _2945_ (.A(net158),
    .B(\tokenflow_inst.i8.cg_elem.q ),
    .Y(_0316_));
 sg13g2_inv_1 _2946_ (.Y(\tokenflow_inst.i78.cg_elem.a ),
    .A(\tokenflow_inst.i2.cg2.q ));
 sg13g2_nand2_1 _2947_ (.Y(_1305_),
    .A(\tokenflow_inst.i8.cg_elem.q ),
    .B(\tokenflow_inst.i8.d0_elem.inv_chain[52] ));
 sg13g2_xnor2_1 _2948_ (.Y(_0005_),
    .A(\tokenflow_inst.i78.cg_elem.a ),
    .B(_1305_));
 sg13g2_nor2_1 _2949_ (.A(net158),
    .B(\tokenflow_inst.i78.cg_elem.q ),
    .Y(_0239_));
 sg13g2_inv_1 _2950_ (.Y(\tokenflow_inst.i6.cg_elem.a ),
    .A(\tokenflow_inst.i8.cg_elem.q ));
 sg13g2_nor2_1 _2951_ (.A(\tokenflow_inst.i3.ydata[36] ),
    .B(\tokenflow_inst.i3.ydata[37] ),
    .Y(_1306_));
 sg13g2_nor4_1 _2952_ (.A(\tokenflow_inst.i3.ydata[32] ),
    .B(\tokenflow_inst.i3.ydata[33] ),
    .C(\tokenflow_inst.i3.ydata[34] ),
    .D(\tokenflow_inst.i3.ydata[35] ),
    .Y(_1307_));
 sg13g2_nor4_1 _2953_ (.A(\tokenflow_inst.i3.ydata[29] ),
    .B(\tokenflow_inst.i3.ydata[30] ),
    .C(\tokenflow_inst.i3.ydata[31] ),
    .D(\tokenflow_inst.i3.ydata[38] ),
    .Y(_1308_));
 sg13g2_nor4_1 _2954_ (.A(\tokenflow_inst.i3.ydata[26] ),
    .B(\tokenflow_inst.i3.ydata[27] ),
    .C(\tokenflow_inst.i3.ydata[28] ),
    .D(\tokenflow_inst.i3.ydata[51] ),
    .Y(_1309_));
 sg13g2_nand4_1 _2955_ (.B(_1307_),
    .C(_1308_),
    .A(_1306_),
    .Y(_1310_),
    .D(_1309_));
 sg13g2_nor4_1 _2956_ (.A(\tokenflow_inst.i3.ydata[45] ),
    .B(\tokenflow_inst.i3.ydata[48] ),
    .C(\tokenflow_inst.i3.ydata[49] ),
    .D(\tokenflow_inst.i3.ydata[50] ),
    .Y(_1311_));
 sg13g2_nor4_1 _2957_ (.A(\tokenflow_inst.i3.ydata[39] ),
    .B(\tokenflow_inst.i3.ydata[44] ),
    .C(\tokenflow_inst.i3.ydata[46] ),
    .D(\tokenflow_inst.i3.ydata[47] ),
    .Y(_1312_));
 sg13g2_nor4_1 _2958_ (.A(\tokenflow_inst.i3.ydata[40] ),
    .B(\tokenflow_inst.i3.ydata[41] ),
    .C(\tokenflow_inst.i3.ydata[42] ),
    .D(\tokenflow_inst.i3.ydata[43] ),
    .Y(_1313_));
 sg13g2_nand3_1 _2959_ (.B(_1312_),
    .C(_1313_),
    .A(_1311_),
    .Y(_1314_));
 sg13g2_nor2_1 _2960_ (.A(_1310_),
    .B(_1314_),
    .Y(_1315_));
 sg13g2_nand3b_1 _2961_ (.B(\tokenflow_inst.i3.d0_elem.inv_chain[3] ),
    .C(_1303_),
    .Y(_1316_),
    .A_N(_1315_));
 sg13g2_xnor2_1 _2962_ (.Y(_0006_),
    .A(\tokenflow_inst.i6.cg_elem.a ),
    .B(_1316_));
 sg13g2_and3_1 _2963_ (.X(\tokenflow_inst.i10.cg.b ),
    .A(_1303_),
    .B(\tokenflow_inst.i3.d0_elem.inv_chain[3] ),
    .C(_1315_));
 sg13g2_and2_1 _2964_ (.A(_1379_),
    .B(_1303_),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[0] ));
 sg13g2_and2_1 _2965_ (.A(net181),
    .B(\tokenflow_inst.i6.cg_elem.q ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[0] ));
 sg13g2_nor2_1 _2966_ (.A(_1189_),
    .B(\tokenflow_inst.i8.cg_elem.a ),
    .Y(\tokenflow_inst.i78.d0_elem.inv_chain[0] ));
 sg13g2_nor2_1 _2967_ (.A(_1189_),
    .B(\tokenflow_inst.i6.cg_elem.a ),
    .Y(\tokenflow_inst.i8.d0_elem.inv_chain[0] ));
 sg13g2_buf_1 _2968_ (.A(_1391_),
    .X(_1317_));
 sg13g2_nor2_1 _2969_ (.A(_1317_),
    .B(_1389_),
    .Y(\tokenflow_inst.ii1.ydata[0] ));
 sg13g2_and4_1 _2970_ (.A(_1389_),
    .B(_1398_),
    .C(_1404_),
    .D(\tokenflow_inst.ii2.ydata[3] ),
    .X(_1318_));
 sg13g2_buf_8 _2971_ (.A(_1318_),
    .X(_1319_));
 sg13g2_nand3_1 _2972_ (.B(\tokenflow_inst.ii3.i.ydata[4] ),
    .C(_1319_),
    .A(_1413_),
    .Y(_1320_));
 sg13g2_nand3_1 _2973_ (.B(_1419_),
    .C(\tokenflow_inst.ii2.ydata[8] ),
    .A(\tokenflow_inst.ii2.ydata[6] ),
    .Y(_1321_));
 sg13g2_nor2_1 _2974_ (.A(_1320_),
    .B(_1321_),
    .Y(_1322_));
 sg13g2_nand2_1 _2975_ (.Y(_1323_),
    .A(\tokenflow_inst.ii2.ydata[9] ),
    .B(_1322_));
 sg13g2_xor2_1 _2976_ (.B(_1323_),
    .A(_1427_),
    .X(_1324_));
 sg13g2_nor2_1 _2977_ (.A(net156),
    .B(_1324_),
    .Y(\tokenflow_inst.ii1.ydata[10] ));
 sg13g2_nand3_1 _2978_ (.B(\tokenflow_inst.ii3.i.ydata[9] ),
    .C(_1322_),
    .A(_1427_),
    .Y(_1325_));
 sg13g2_xnor2_1 _2979_ (.Y(_1326_),
    .A(_1431_),
    .B(_1325_));
 sg13g2_nor2_1 _2980_ (.A(_1317_),
    .B(_1326_),
    .Y(\tokenflow_inst.ii1.ydata[11] ));
 sg13g2_nand2_1 _2981_ (.Y(_1327_),
    .A(_1427_),
    .B(\tokenflow_inst.ii3.i.ydata[9] ));
 sg13g2_nor4_2 _2982_ (.A(_1431_),
    .B(_1320_),
    .C(_1321_),
    .Y(_1328_),
    .D(_1327_));
 sg13g2_xnor2_1 _2983_ (.Y(_1329_),
    .A(_1435_),
    .B(_1328_));
 sg13g2_nor2_1 _2984_ (.A(net156),
    .B(_1329_),
    .Y(\tokenflow_inst.ii1.ydata[12] ));
 sg13g2_nand2_1 _2985_ (.Y(_1330_),
    .A(_1435_),
    .B(_1328_));
 sg13g2_nand2_1 _2986_ (.Y(_1331_),
    .A(\tokenflow_inst.ii3.i.ydata[13] ),
    .B(_1330_));
 sg13g2_o21ai_1 _2987_ (.B1(_1331_),
    .Y(\tokenflow_inst.ii1.ydata[13] ),
    .A1(\tokenflow_inst.ii2.ydata[13] ),
    .A2(_1330_));
 sg13g2_and3_1 _2988_ (.X(_1332_),
    .A(_1435_),
    .B(\tokenflow_inst.ii2.ydata[13] ),
    .C(_1328_));
 sg13g2_buf_1 _2989_ (.A(_1332_),
    .X(_1333_));
 sg13g2_xnor2_1 _2990_ (.Y(_1334_),
    .A(_1440_),
    .B(_1333_));
 sg13g2_nor2_1 _2991_ (.A(net156),
    .B(_1334_),
    .Y(\tokenflow_inst.ii1.ydata[14] ));
 sg13g2_nand2_1 _2992_ (.Y(_1335_),
    .A(_1440_),
    .B(_1333_));
 sg13g2_xor2_1 _2993_ (.B(_1335_),
    .A(\tokenflow_inst.ii2.ydata[15] ),
    .X(_1336_));
 sg13g2_nor2_1 _2994_ (.A(net156),
    .B(_1336_),
    .Y(\tokenflow_inst.ii1.ydata[15] ));
 sg13g2_and3_1 _2995_ (.X(_1337_),
    .A(_1440_),
    .B(\tokenflow_inst.ii2.ydata[15] ),
    .C(_1333_));
 sg13g2_buf_8 _2996_ (.A(_1337_),
    .X(_1338_));
 sg13g2_xnor2_1 _2997_ (.Y(_1339_),
    .A(_1446_),
    .B(_1338_));
 sg13g2_nor2_1 _2998_ (.A(net156),
    .B(_1339_),
    .Y(\tokenflow_inst.ii1.ydata[16] ));
 sg13g2_nand2_1 _2999_ (.Y(_1340_),
    .A(_1446_),
    .B(_1338_));
 sg13g2_xor2_1 _3000_ (.B(_1340_),
    .A(_1450_),
    .X(_1341_));
 sg13g2_nor2_1 _3001_ (.A(net156),
    .B(_1341_),
    .Y(\tokenflow_inst.ii1.ydata[17] ));
 sg13g2_nand3_1 _3002_ (.B(_1450_),
    .C(_1338_),
    .A(_1446_),
    .Y(_1342_));
 sg13g2_xor2_1 _3003_ (.B(_1342_),
    .A(\tokenflow_inst.ii2.ydata[18] ),
    .X(_1343_));
 sg13g2_nor2_1 _3004_ (.A(net156),
    .B(_1343_),
    .Y(\tokenflow_inst.ii1.ydata[18] ));
 sg13g2_and4_1 _3005_ (.A(_1446_),
    .B(_1450_),
    .C(\tokenflow_inst.ii2.ydata[18] ),
    .D(_1338_),
    .X(_1344_));
 sg13g2_buf_8 _3006_ (.A(_1344_),
    .X(_1345_));
 sg13g2_xnor2_1 _3007_ (.Y(_1346_),
    .A(_1455_),
    .B(_1345_));
 sg13g2_nor2_1 _3008_ (.A(net156),
    .B(_1346_),
    .Y(\tokenflow_inst.ii1.ydata[19] ));
 sg13g2_buf_1 _3009_ (.A(net179),
    .X(_1347_));
 sg13g2_xnor2_1 _3010_ (.Y(_1348_),
    .A(_1389_),
    .B(_1398_));
 sg13g2_nor2_1 _3011_ (.A(net155),
    .B(_1348_),
    .Y(\tokenflow_inst.ii1.ydata[1] ));
 sg13g2_nand2_1 _3012_ (.Y(_1349_),
    .A(_1455_),
    .B(_1345_));
 sg13g2_xor2_1 _3013_ (.B(_1349_),
    .A(_1460_),
    .X(_1350_));
 sg13g2_nor2_1 _3014_ (.A(net155),
    .B(_1350_),
    .Y(\tokenflow_inst.ii1.ydata[20] ));
 sg13g2_nand3_1 _3015_ (.B(_1460_),
    .C(_1345_),
    .A(_1455_),
    .Y(_1351_));
 sg13g2_xnor2_1 _3016_ (.Y(_1352_),
    .A(\tokenflow_inst.ii2.ydata[21] ),
    .B(_1351_));
 sg13g2_and2_1 _3017_ (.A(net181),
    .B(_1352_),
    .X(\tokenflow_inst.ii1.ydata[21] ));
 sg13g2_nand4_1 _3018_ (.B(_1460_),
    .C(\tokenflow_inst.ii2.ydata[21] ),
    .A(_1455_),
    .Y(_1353_),
    .D(_1345_));
 sg13g2_xor2_1 _3019_ (.B(_1353_),
    .A(_1467_),
    .X(_1354_));
 sg13g2_nor2_1 _3020_ (.A(net155),
    .B(_1354_),
    .Y(\tokenflow_inst.ii1.ydata[22] ));
 sg13g2_nand2_1 _3021_ (.Y(_1355_),
    .A(_1467_),
    .B(\tokenflow_inst.ii3.i.ydata[21] ));
 sg13g2_nor2_1 _3022_ (.A(_1351_),
    .B(_1355_),
    .Y(_1356_));
 sg13g2_xnor2_1 _3023_ (.Y(_1357_),
    .A(\tokenflow_inst.ii2.ydata[23] ),
    .B(_1356_));
 sg13g2_nor2_1 _3024_ (.A(net155),
    .B(_1357_),
    .Y(\tokenflow_inst.ii1.ydata[23] ));
 sg13g2_and3_1 _3025_ (.X(_1358_),
    .A(_1467_),
    .B(\tokenflow_inst.ii2.ydata[23] ),
    .C(\tokenflow_inst.ii3.i.ydata[21] ));
 sg13g2_and4_1 _3026_ (.A(_1455_),
    .B(_1460_),
    .C(_1345_),
    .D(_1358_),
    .X(_1359_));
 sg13g2_xnor2_1 _3027_ (.Y(_1360_),
    .A(_1472_),
    .B(_1359_));
 sg13g2_nor2_1 _3028_ (.A(net155),
    .B(_1360_),
    .Y(\tokenflow_inst.ii1.ydata[24] ));
 sg13g2_nand2_1 _3029_ (.Y(_1361_),
    .A(_1472_),
    .B(_1359_));
 sg13g2_xor2_1 _3030_ (.B(_1361_),
    .A(\tokenflow_inst.ii2.ydata[25] ),
    .X(_1362_));
 sg13g2_nor2_1 _3031_ (.A(net155),
    .B(_1362_),
    .Y(\tokenflow_inst.ii1.ydata[25] ));
 sg13g2_nand2_1 _3032_ (.Y(_1363_),
    .A(_1389_),
    .B(_1398_));
 sg13g2_xor2_1 _3033_ (.B(_1363_),
    .A(_1404_),
    .X(_1364_));
 sg13g2_nor2_1 _3034_ (.A(net155),
    .B(_1364_),
    .Y(\tokenflow_inst.ii1.ydata[2] ));
 sg13g2_nand3_1 _3035_ (.B(_1398_),
    .C(_1404_),
    .A(_1389_),
    .Y(_1365_));
 sg13g2_xor2_1 _3036_ (.B(_1365_),
    .A(\tokenflow_inst.ii2.ydata[3] ),
    .X(_1366_));
 sg13g2_nor2_1 _3037_ (.A(net155),
    .B(_1366_),
    .Y(\tokenflow_inst.ii1.ydata[3] ));
 sg13g2_xnor2_1 _3038_ (.Y(_1367_),
    .A(\tokenflow_inst.ii2.ydata[4] ),
    .B(_1319_));
 sg13g2_nor2_1 _3039_ (.A(_1347_),
    .B(_1367_),
    .Y(\tokenflow_inst.ii1.ydata[4] ));
 sg13g2_and2_1 _3040_ (.A(\tokenflow_inst.ii3.i.ydata[4] ),
    .B(_1319_),
    .X(_1368_));
 sg13g2_xnor2_1 _3041_ (.Y(_1369_),
    .A(_1413_),
    .B(_1368_));
 sg13g2_nor2_1 _3042_ (.A(_1347_),
    .B(_1369_),
    .Y(\tokenflow_inst.ii1.ydata[5] ));
 sg13g2_xor2_1 _3043_ (.B(_1320_),
    .A(\tokenflow_inst.ii2.ydata[6] ),
    .X(_1370_));
 sg13g2_nor2_1 _3044_ (.A(net167),
    .B(_1370_),
    .Y(\tokenflow_inst.ii1.ydata[6] ));
 sg13g2_and2_1 _3045_ (.A(_1413_),
    .B(_1368_),
    .X(_1371_));
 sg13g2_nand2_1 _3046_ (.Y(_1372_),
    .A(\tokenflow_inst.ii3.i.ydata[6] ),
    .B(_1371_));
 sg13g2_xor2_1 _3047_ (.B(_1372_),
    .A(_1419_),
    .X(_1373_));
 sg13g2_nor2_1 _3048_ (.A(net167),
    .B(_1373_),
    .Y(\tokenflow_inst.ii1.ydata[7] ));
 sg13g2_nand3_1 _3049_ (.B(\tokenflow_inst.ii3.i.ydata[6] ),
    .C(_1371_),
    .A(_1419_),
    .Y(_1374_));
 sg13g2_xor2_1 _3050_ (.B(_1374_),
    .A(\tokenflow_inst.ii2.ydata[8] ),
    .X(_1375_));
 sg13g2_nor2_1 _3051_ (.A(_1392_),
    .B(_1375_),
    .Y(\tokenflow_inst.ii1.ydata[8] ));
 sg13g2_xnor2_1 _3052_ (.Y(_1376_),
    .A(\tokenflow_inst.ii2.ydata[9] ),
    .B(_1322_));
 sg13g2_nor2_1 _3053_ (.A(_1392_),
    .B(_1376_),
    .Y(\tokenflow_inst.ii1.ydata[9] ));
 sg13g2_xor2_1 _3054_ (.B(\tokenflow_inst.i3.ydata[22] ),
    .A(\tokenflow_inst.i3.ydata[7] ),
    .X(net3));
 sg13g2_xor2_1 _3055_ (.B(\tokenflow_inst.i3.ydata[23] ),
    .A(\tokenflow_inst.i3.ydata[8] ),
    .X(net4));
 sg13g2_xor2_1 _3056_ (.B(\tokenflow_inst.i3.ydata[24] ),
    .A(\tokenflow_inst.i3.ydata[9] ),
    .X(net5));
 sg13g2_xor2_1 _3057_ (.B(\tokenflow_inst.i3.ydata[25] ),
    .A(\tokenflow_inst.i3.ydata[10] ),
    .X(net6));
 sg13g2_xor2_1 _3058_ (.B(\tokenflow_inst.i3.ydata[15] ),
    .A(\tokenflow_inst.i3.ydata[0] ),
    .X(net12));
 sg13g2_xor2_1 _3059_ (.B(\tokenflow_inst.i3.ydata[16] ),
    .A(\tokenflow_inst.i3.ydata[1] ),
    .X(net13));
 sg13g2_xor2_1 _3060_ (.B(\tokenflow_inst.i3.ydata[17] ),
    .A(\tokenflow_inst.i3.ydata[2] ),
    .X(net14));
 sg13g2_xor2_1 _3061_ (.B(\tokenflow_inst.i3.ydata[18] ),
    .A(\tokenflow_inst.i3.ydata[3] ),
    .X(net15));
 sg13g2_xor2_1 _3062_ (.B(\tokenflow_inst.i3.ydata[19] ),
    .A(\tokenflow_inst.i3.ydata[4] ),
    .X(net16));
 sg13g2_xor2_1 _3063_ (.B(\tokenflow_inst.i3.ydata[20] ),
    .A(\tokenflow_inst.i3.ydata[5] ),
    .X(net17));
 sg13g2_xor2_1 _3064_ (.B(\tokenflow_inst.i3.ydata[21] ),
    .A(\tokenflow_inst.i3.ydata[6] ),
    .X(net18));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tiehi _3078__199 (.L_HI(net199));
 sg13g2_buf_1 _3067_ (.A(net187),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[0] ));
 sg13g2_buf_1 _3068_ (.A(net189),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[0] ));
 sg13g2_buf_1 _3069_ (.A(net187),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[0] ));
 sg13g2_buf_1 _3070_ (.A(net190),
    .X(\tokenflow_inst.i8.ydata[51] ));
 sg13g2_buf_1 _3071_ (.A(net191),
    .X(\tokenflow_inst.i8.ydata[52] ));
 sg13g2_buf_1 _3072_ (.A(net192),
    .X(\tokenflow_inst.i10.d0.inv_chain[0] ));
 sg13g2_buf_1 _3073_ (.A(net187),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[0] ));
 sg13g2_buf_1 _3074_ (.A(net193),
    .X(\tokenflow_inst.i78.ydata[50] ));
 sg13g2_buf_1 _3075_ (.A(net194),
    .X(\tokenflow_inst.i78.ydata[51] ));
 sg13g2_buf_1 _3076_ (.A(net195),
    .X(\tokenflow_inst.i78.ydata[52] ));
 sg13g2_buf_1 _3077_ (.A(net196),
    .X(\tokenflow_inst.i78.ydata[53] ));
 sg13g2_buf_1 _3078_ (.A(net199),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3079_ (.A(net200),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3080_ (.A(net201),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3081_ (.A(net202),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3082_ (.A(net203),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3083_ (.A(net204),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3084_ (.A(net205),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3085_ (.A(net206),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3086_ (.A(\tokenflow_inst.i3.ydata[11] ),
    .X(net7));
 sg13g2_buf_1 _3087_ (.A(\tokenflow_inst.i3.ydata[12] ),
    .X(net8));
 sg13g2_buf_1 _3088_ (.A(\tokenflow_inst.i3.ydata[13] ),
    .X(net9));
 sg13g2_buf_1 _3089_ (.A(\tokenflow_inst.i3.ydata[14] ),
    .X(net10));
 sg13g2_buf_1 _3090_ (.A(\tokenflow_inst.i10.cg.b ),
    .X(net11));
 sg13g2_dllrq_1 \tokenflow_inst.i1.c.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ),
    .GATE_N(_0003_),
    .RESET_B(net207),
    .Q(\tokenflow_inst.i1.c.q ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i10.d0.genblk1[0].min_delay_inst.d0  (.A(net197),
    .X(\tokenflow_inst.i10.d0.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i11.i.d0.genblk1[0].min_delay_inst.d0  (.A(net186),
    .X(\tokenflow_inst.i11.i.d0.inv_chain[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.i2.cg1.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i2.cg1.a ),
    .GATE_N(_0001_),
    .RESET_B(net208),
    .Q(\tokenflow_inst.i2.cg1.q ));
 sg13g2_dllrq_1 \tokenflow_inst.i2.cg2.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i2.cg2.a ),
    .GATE_N(_0002_),
    .RESET_B(net209),
    .Q(\tokenflow_inst.i2.cg2.q ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i3.cg_elem.a ),
    .GATE_N(_0000_),
    .RESET_B(net210),
    .Q(\tokenflow_inst.i2.cg2.a ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i3.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i3.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[2] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i3.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i3.d0_elem.inv_chain[2] ),
    .X(\tokenflow_inst.i3.d0_elem.inv_chain[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(net139),
    .RESET_B(net211),
    .Q(\tokenflow_inst.i3.ydata[0] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(net140),
    .RESET_B(net212),
    .Q(\tokenflow_inst.i3.ydata[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0009_),
    .GATE_N(net135),
    .RESET_B(net213),
    .Q(\tokenflow_inst.i3.ydata[11] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(net135),
    .RESET_B(net214),
    .Q(\tokenflow_inst.i3.ydata[12] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0011_),
    .GATE_N(net135),
    .RESET_B(net215),
    .Q(\tokenflow_inst.i3.ydata[13] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0012_),
    .GATE_N(net135),
    .RESET_B(net216),
    .Q(\tokenflow_inst.i3.ydata[14] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(net134),
    .RESET_B(net217),
    .Q(\tokenflow_inst.i3.ydata[15] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0014_),
    .GATE_N(net134),
    .RESET_B(net218),
    .Q(\tokenflow_inst.i3.ydata[16] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0015_),
    .GATE_N(net133),
    .RESET_B(net219),
    .Q(\tokenflow_inst.i3.ydata[17] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0016_),
    .GATE_N(net133),
    .RESET_B(net220),
    .Q(\tokenflow_inst.i3.ydata[18] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0017_),
    .GATE_N(net135),
    .RESET_B(net221),
    .Q(\tokenflow_inst.i3.ydata[19] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0018_),
    .GATE_N(net141),
    .RESET_B(net222),
    .Q(\tokenflow_inst.i3.ydata[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0019_),
    .GATE_N(net135),
    .RESET_B(net223),
    .Q(\tokenflow_inst.i3.ydata[20] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0020_),
    .GATE_N(net135),
    .RESET_B(net224),
    .Q(\tokenflow_inst.i3.ydata[21] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0021_),
    .GATE_N(net132),
    .RESET_B(net225),
    .Q(\tokenflow_inst.i3.ydata[22] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0022_),
    .GATE_N(net132),
    .RESET_B(net226),
    .Q(\tokenflow_inst.i3.ydata[23] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0023_),
    .GATE_N(net132),
    .RESET_B(net227),
    .Q(\tokenflow_inst.i3.ydata[24] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0024_),
    .GATE_N(net137),
    .RESET_B(net228),
    .Q(\tokenflow_inst.i3.ydata[25] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0025_),
    .GATE_N(net138),
    .RESET_B(net229),
    .Q(\tokenflow_inst.i3.ydata[26] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0026_),
    .GATE_N(net138),
    .RESET_B(net230),
    .Q(\tokenflow_inst.i3.ydata[27] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0027_),
    .GATE_N(net138),
    .RESET_B(net231),
    .Q(\tokenflow_inst.i3.ydata[28] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0028_),
    .GATE_N(net139),
    .RESET_B(net232),
    .Q(\tokenflow_inst.i3.ydata[29] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0029_),
    .GATE_N(net141),
    .RESET_B(net233),
    .Q(\tokenflow_inst.i3.ydata[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0030_),
    .GATE_N(net139),
    .RESET_B(net234),
    .Q(\tokenflow_inst.i3.ydata[30] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0031_),
    .GATE_N(net137),
    .RESET_B(net235),
    .Q(\tokenflow_inst.i3.ydata[31] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0032_),
    .GATE_N(net137),
    .RESET_B(net236),
    .Q(\tokenflow_inst.i3.ydata[32] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0033_),
    .GATE_N(net137),
    .RESET_B(net237),
    .Q(\tokenflow_inst.i3.ydata[33] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0034_),
    .GATE_N(net137),
    .RESET_B(net238),
    .Q(\tokenflow_inst.i3.ydata[34] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0035_),
    .GATE_N(net137),
    .RESET_B(net239),
    .Q(\tokenflow_inst.i3.ydata[35] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0036_),
    .GATE_N(net137),
    .RESET_B(net240),
    .Q(\tokenflow_inst.i3.ydata[36] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0037_),
    .GATE_N(net137),
    .RESET_B(net241),
    .Q(\tokenflow_inst.i3.ydata[37] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0038_),
    .GATE_N(net132),
    .RESET_B(net242),
    .Q(\tokenflow_inst.i3.ydata[38] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0039_),
    .GATE_N(net132),
    .RESET_B(net243),
    .Q(\tokenflow_inst.i3.ydata[39] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0040_),
    .GATE_N(net141),
    .RESET_B(net244),
    .Q(\tokenflow_inst.i3.ydata[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0041_),
    .GATE_N(net132),
    .RESET_B(net245),
    .Q(\tokenflow_inst.i3.ydata[40] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0042_),
    .GATE_N(net131),
    .RESET_B(net246),
    .Q(\tokenflow_inst.i3.ydata[41] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0043_),
    .GATE_N(net130),
    .RESET_B(net247),
    .Q(\tokenflow_inst.i3.ydata[42] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0044_),
    .GATE_N(net131),
    .RESET_B(net248),
    .Q(\tokenflow_inst.i3.ydata[43] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0045_),
    .GATE_N(net130),
    .RESET_B(net249),
    .Q(\tokenflow_inst.i3.ydata[44] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0046_),
    .GATE_N(net130),
    .RESET_B(net250),
    .Q(\tokenflow_inst.i3.ydata[45] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0047_),
    .GATE_N(net130),
    .RESET_B(net251),
    .Q(\tokenflow_inst.i3.ydata[46] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0048_),
    .GATE_N(net130),
    .RESET_B(net252),
    .Q(\tokenflow_inst.i3.ydata[47] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0049_),
    .GATE_N(net130),
    .RESET_B(net253),
    .Q(\tokenflow_inst.i3.ydata[48] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0050_),
    .GATE_N(net130),
    .RESET_B(net254),
    .Q(\tokenflow_inst.i3.ydata[49] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0051_),
    .GATE_N(net141),
    .RESET_B(net255),
    .Q(\tokenflow_inst.i3.ydata[4] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0052_),
    .GATE_N(net130),
    .RESET_B(net256),
    .Q(\tokenflow_inst.i3.ydata[50] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[51]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0053_),
    .GATE_N(net138),
    .RESET_B(net257),
    .Q(\tokenflow_inst.i3.ydata[51] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[52]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0054_),
    .GATE_N(net139),
    .RESET_B(net258),
    .Q(\tokenflow_inst.i3.ydata[52] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0055_),
    .GATE_N(net139),
    .RESET_B(net259),
    .Q(\tokenflow_inst.i3.ydata[53] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0056_),
    .GATE_N(net139),
    .RESET_B(net260),
    .Q(\tokenflow_inst.i3.ydata[54] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0057_),
    .GATE_N(net141),
    .RESET_B(net261),
    .Q(\tokenflow_inst.i3.ydata[55] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0058_),
    .GATE_N(net142),
    .RESET_B(net262),
    .Q(\tokenflow_inst.i3.ydata[56] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0059_),
    .GATE_N(net141),
    .RESET_B(net263),
    .Q(\tokenflow_inst.i3.ydata[57] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0060_),
    .GATE_N(net141),
    .RESET_B(net264),
    .Q(\tokenflow_inst.i3.ydata[58] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0061_),
    .GATE_N(net142),
    .RESET_B(net265),
    .Q(\tokenflow_inst.i3.ydata[59] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0062_),
    .GATE_N(net141),
    .RESET_B(net266),
    .Q(\tokenflow_inst.i3.ydata[5] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0063_),
    .GATE_N(net140),
    .RESET_B(net267),
    .Q(\tokenflow_inst.i3.ydata[60] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0064_),
    .GATE_N(net140),
    .RESET_B(net268),
    .Q(\tokenflow_inst.i3.ydata[61] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0065_),
    .GATE_N(net140),
    .RESET_B(net269),
    .Q(\tokenflow_inst.i3.ydata[62] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0066_),
    .GATE_N(net136),
    .RESET_B(net270),
    .Q(\tokenflow_inst.i3.ydata[63] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0067_),
    .GATE_N(net135),
    .RESET_B(net271),
    .Q(\tokenflow_inst.i3.ydata[64] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0068_),
    .GATE_N(net133),
    .RESET_B(net272),
    .Q(\tokenflow_inst.i3.ydata[65] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0069_),
    .GATE_N(net133),
    .RESET_B(net273),
    .Q(\tokenflow_inst.i3.ydata[66] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0070_),
    .GATE_N(net133),
    .RESET_B(net274),
    .Q(\tokenflow_inst.i3.ydata[67] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0071_),
    .GATE_N(net133),
    .RESET_B(net275),
    .Q(\tokenflow_inst.i3.ydata[68] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0072_),
    .GATE_N(net133),
    .RESET_B(net276),
    .Q(\tokenflow_inst.i3.ydata[69] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0073_),
    .GATE_N(net140),
    .RESET_B(net277),
    .Q(\tokenflow_inst.i3.ydata[6] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0074_),
    .GATE_N(net133),
    .RESET_B(net278),
    .Q(\tokenflow_inst.i3.ydata[70] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0075_),
    .GATE_N(net134),
    .RESET_B(net279),
    .Q(\tokenflow_inst.i3.ydata[71] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0076_),
    .GATE_N(net134),
    .RESET_B(net280),
    .Q(\tokenflow_inst.i3.ydata[72] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0077_),
    .GATE_N(net131),
    .RESET_B(net281),
    .Q(\tokenflow_inst.i3.ydata[73] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0078_),
    .GATE_N(net131),
    .RESET_B(net282),
    .Q(\tokenflow_inst.i3.ydata[74] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0079_),
    .GATE_N(net131),
    .RESET_B(net283),
    .Q(\tokenflow_inst.i3.ydata[75] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0080_),
    .GATE_N(net131),
    .RESET_B(net284),
    .Q(\tokenflow_inst.i3.ydata[76] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0081_),
    .GATE_N(net132),
    .RESET_B(net285),
    .Q(\tokenflow_inst.i3.ydata[77] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0082_),
    .GATE_N(net140),
    .RESET_B(net286),
    .Q(\tokenflow_inst.i3.ydata[7] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0083_),
    .GATE_N(net140),
    .RESET_B(net287),
    .Q(\tokenflow_inst.i3.ydata[8] ));
 sg13g2_dllrq_1 \tokenflow_inst.i3.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0084_),
    .GATE_N(net140),
    .RESET_B(net288),
    .Q(\tokenflow_inst.i3.ydata[9] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i6.cg_elem.a ),
    .GATE_N(_0006_),
    .RESET_B(net289),
    .Q(\tokenflow_inst.i6.cg_elem.q ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[10].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[10] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[11] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[11].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[11] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[12] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[12].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[12] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[13] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[13].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[13] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[14] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[14].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[14] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[15] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[15].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[15] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[16] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[16].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[16] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[17] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[17].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[17] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[18] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[18].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[18] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[19] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[19].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[19] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[20] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[2] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[20].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[20] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[21] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[21].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[21] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[22] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[22].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[22] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[23] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[23].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[23] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[24] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[24].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[24] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[25] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[25].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[25] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[26] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[26].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[26] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[27] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[27].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[27] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[28] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[28].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[28] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[29] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[29].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[29] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[30] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[2] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[3] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[30].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[30] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[31] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[31].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[31] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[32] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[32].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[32] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[33] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[33].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[33] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[34] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[34].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[34] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[35] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[35].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[35] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[36] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[36].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[36] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[37] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[37].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[37] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[38] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[38].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[38] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[39] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[39].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[39] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[40] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[3].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[3] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[4] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[40].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[40] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[41] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[41].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[41] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[42] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[42].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[42] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[43] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[43].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[43] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[44] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[44].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[44] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[45] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[45].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[45] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[46] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[46].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[46] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[47] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[47].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[47] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[48] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[48].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[48] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[49] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[49].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[49] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[50] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[4].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[4] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[5] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[50].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[50] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[51] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[51].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[51] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[52] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[5].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[5] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[6] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[6].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[6] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[7] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[7].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[7] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[8] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[8].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[8] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[9] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i6.d0_elem.genblk1[9].min_delay_inst.d0  (.A(\tokenflow_inst.i6.d0_elem.inv_chain[9] ),
    .X(\tokenflow_inst.i6.d0_elem.inv_chain[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0086_),
    .GATE_N(net125),
    .RESET_B(net290),
    .Q(\tokenflow_inst.i6.ydata[0] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0087_),
    .GATE_N(net128),
    .RESET_B(net291),
    .Q(\tokenflow_inst.i6.ydata[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0088_),
    .GATE_N(net122),
    .RESET_B(net292),
    .Q(\tokenflow_inst.i6.ydata[11] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0089_),
    .GATE_N(net122),
    .RESET_B(net293),
    .Q(\tokenflow_inst.i6.ydata[12] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0090_),
    .GATE_N(net123),
    .RESET_B(net294),
    .Q(\tokenflow_inst.i6.ydata[13] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0091_),
    .GATE_N(net122),
    .RESET_B(net295),
    .Q(\tokenflow_inst.i6.ydata[14] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0092_),
    .GATE_N(net121),
    .RESET_B(net296),
    .Q(\tokenflow_inst.i6.ydata[15] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0093_),
    .GATE_N(net121),
    .RESET_B(net297),
    .Q(\tokenflow_inst.i6.ydata[16] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0094_),
    .GATE_N(net121),
    .RESET_B(net298),
    .Q(\tokenflow_inst.i6.ydata[17] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0095_),
    .GATE_N(net121),
    .RESET_B(net299),
    .Q(\tokenflow_inst.i6.ydata[18] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0096_),
    .GATE_N(net122),
    .RESET_B(net300),
    .Q(\tokenflow_inst.i6.ydata[19] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0097_),
    .GATE_N(net126),
    .RESET_B(net301),
    .Q(\tokenflow_inst.i6.ydata[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0098_),
    .GATE_N(net122),
    .RESET_B(net302),
    .Q(\tokenflow_inst.i6.ydata[20] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0099_),
    .GATE_N(net122),
    .RESET_B(net303),
    .Q(\tokenflow_inst.i6.ydata[21] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0100_),
    .GATE_N(net120),
    .RESET_B(net304),
    .Q(\tokenflow_inst.i6.ydata[22] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0101_),
    .GATE_N(net120),
    .RESET_B(net305),
    .Q(\tokenflow_inst.i6.ydata[23] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0102_),
    .GATE_N(net120),
    .RESET_B(net306),
    .Q(\tokenflow_inst.i6.ydata[24] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0103_),
    .GATE_N(net126),
    .RESET_B(net307),
    .Q(\tokenflow_inst.i6.ydata[25] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0104_),
    .GATE_N(net129),
    .RESET_B(net308),
    .Q(\tokenflow_inst.i6.ydata[26] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0105_),
    .GATE_N(net124),
    .RESET_B(net309),
    .Q(\tokenflow_inst.i6.ydata[27] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0106_),
    .GATE_N(net124),
    .RESET_B(net310),
    .Q(\tokenflow_inst.i6.ydata[28] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0107_),
    .GATE_N(net125),
    .RESET_B(net311),
    .Q(\tokenflow_inst.i6.ydata[29] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0108_),
    .GATE_N(net127),
    .RESET_B(net312),
    .Q(\tokenflow_inst.i6.ydata[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0109_),
    .GATE_N(net125),
    .RESET_B(net313),
    .Q(\tokenflow_inst.i6.ydata[30] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0110_),
    .GATE_N(net125),
    .RESET_B(net314),
    .Q(\tokenflow_inst.i6.ydata[31] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0111_),
    .GATE_N(net125),
    .RESET_B(net315),
    .Q(\tokenflow_inst.i6.ydata[32] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0112_),
    .GATE_N(net125),
    .RESET_B(net316),
    .Q(\tokenflow_inst.i6.ydata[33] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0113_),
    .GATE_N(net124),
    .RESET_B(net317),
    .Q(\tokenflow_inst.i6.ydata[34] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0114_),
    .GATE_N(net124),
    .RESET_B(net318),
    .Q(\tokenflow_inst.i6.ydata[35] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0115_),
    .GATE_N(net124),
    .RESET_B(net319),
    .Q(\tokenflow_inst.i6.ydata[36] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0116_),
    .GATE_N(net124),
    .RESET_B(net320),
    .Q(\tokenflow_inst.i6.ydata[37] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0117_),
    .GATE_N(net124),
    .RESET_B(net321),
    .Q(\tokenflow_inst.i6.ydata[38] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0118_),
    .GATE_N(net120),
    .RESET_B(net322),
    .Q(\tokenflow_inst.i6.ydata[39] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0119_),
    .GATE_N(net127),
    .RESET_B(net323),
    .Q(\tokenflow_inst.i6.ydata[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0120_),
    .GATE_N(net120),
    .RESET_B(net324),
    .Q(\tokenflow_inst.i6.ydata[40] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0121_),
    .GATE_N(net120),
    .RESET_B(net325),
    .Q(\tokenflow_inst.i6.ydata[41] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0122_),
    .GATE_N(net118),
    .RESET_B(net326),
    .Q(\tokenflow_inst.i6.ydata[42] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0123_),
    .GATE_N(net118),
    .RESET_B(net327),
    .Q(\tokenflow_inst.i6.ydata[43] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0124_),
    .GATE_N(net118),
    .RESET_B(net328),
    .Q(\tokenflow_inst.i6.ydata[44] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0125_),
    .GATE_N(net118),
    .RESET_B(net329),
    .Q(\tokenflow_inst.i6.ydata[45] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0126_),
    .GATE_N(net118),
    .RESET_B(net330),
    .Q(\tokenflow_inst.i6.ydata[46] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0127_),
    .GATE_N(net118),
    .RESET_B(net331),
    .Q(\tokenflow_inst.i6.ydata[47] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0128_),
    .GATE_N(net118),
    .RESET_B(net332),
    .Q(\tokenflow_inst.i6.ydata[48] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0129_),
    .GATE_N(net119),
    .RESET_B(net333),
    .Q(\tokenflow_inst.i6.ydata[49] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0130_),
    .GATE_N(net127),
    .RESET_B(net334),
    .Q(\tokenflow_inst.i6.ydata[4] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0131_),
    .GATE_N(net118),
    .RESET_B(net335),
    .Q(\tokenflow_inst.i6.ydata[50] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[51]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0132_),
    .GATE_N(net124),
    .RESET_B(net336),
    .Q(\tokenflow_inst.i6.ydata[51] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[52]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0133_),
    .GATE_N(net126),
    .RESET_B(net337),
    .Q(\tokenflow_inst.i6.ydata[52] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0134_),
    .GATE_N(net125),
    .RESET_B(net338),
    .Q(\tokenflow_inst.i6.ydata[53] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0135_),
    .GATE_N(net125),
    .RESET_B(net339),
    .Q(\tokenflow_inst.i6.ydata[54] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0136_),
    .GATE_N(net127),
    .RESET_B(net340),
    .Q(\tokenflow_inst.i6.ydata[55] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0137_),
    .GATE_N(net127),
    .RESET_B(net341),
    .Q(\tokenflow_inst.i6.ydata[56] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0138_),
    .GATE_N(net129),
    .RESET_B(net342),
    .Q(\tokenflow_inst.i6.ydata[57] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0139_),
    .GATE_N(net129),
    .RESET_B(net343),
    .Q(\tokenflow_inst.i6.ydata[58] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0140_),
    .GATE_N(net127),
    .RESET_B(net344),
    .Q(\tokenflow_inst.i6.ydata[59] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0141_),
    .GATE_N(net127),
    .RESET_B(net345),
    .Q(\tokenflow_inst.i6.ydata[5] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0142_),
    .GATE_N(net128),
    .RESET_B(net346),
    .Q(\tokenflow_inst.i6.ydata[60] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0143_),
    .GATE_N(net128),
    .RESET_B(net347),
    .Q(\tokenflow_inst.i6.ydata[61] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0144_),
    .GATE_N(net128),
    .RESET_B(net348),
    .Q(\tokenflow_inst.i6.ydata[62] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0145_),
    .GATE_N(net122),
    .RESET_B(net349),
    .Q(\tokenflow_inst.i6.ydata[63] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0146_),
    .GATE_N(net122),
    .RESET_B(net350),
    .Q(\tokenflow_inst.i6.ydata[64] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0147_),
    .GATE_N(net123),
    .RESET_B(net351),
    .Q(\tokenflow_inst.i6.ydata[65] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0148_),
    .GATE_N(net121),
    .RESET_B(net352),
    .Q(\tokenflow_inst.i6.ydata[66] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0149_),
    .GATE_N(net123),
    .RESET_B(net353),
    .Q(\tokenflow_inst.i6.ydata[67] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0150_),
    .GATE_N(net123),
    .RESET_B(net354),
    .Q(\tokenflow_inst.i6.ydata[68] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0151_),
    .GATE_N(net123),
    .RESET_B(net355),
    .Q(\tokenflow_inst.i6.ydata[69] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0152_),
    .GATE_N(net127),
    .RESET_B(net356),
    .Q(\tokenflow_inst.i6.ydata[6] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0153_),
    .GATE_N(net121),
    .RESET_B(net357),
    .Q(\tokenflow_inst.i6.ydata[70] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0154_),
    .GATE_N(net121),
    .RESET_B(net358),
    .Q(\tokenflow_inst.i6.ydata[71] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0155_),
    .GATE_N(net121),
    .RESET_B(net359),
    .Q(\tokenflow_inst.i6.ydata[72] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0156_),
    .GATE_N(net119),
    .RESET_B(net360),
    .Q(\tokenflow_inst.i6.ydata[73] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0157_),
    .GATE_N(net119),
    .RESET_B(net361),
    .Q(\tokenflow_inst.i6.ydata[74] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0158_),
    .GATE_N(net119),
    .RESET_B(net362),
    .Q(\tokenflow_inst.i6.ydata[75] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0159_),
    .GATE_N(net119),
    .RESET_B(net363),
    .Q(\tokenflow_inst.i6.ydata[76] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0160_),
    .GATE_N(net126),
    .RESET_B(net364),
    .Q(\tokenflow_inst.i6.ydata[77] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0161_),
    .GATE_N(net128),
    .RESET_B(net365),
    .Q(\tokenflow_inst.i6.ydata[7] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0162_),
    .GATE_N(net128),
    .RESET_B(net366),
    .Q(\tokenflow_inst.i6.ydata[8] ));
 sg13g2_dllrq_1 \tokenflow_inst.i6.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0163_),
    .GATE_N(net128),
    .RESET_B(net367),
    .Q(\tokenflow_inst.i6.ydata[9] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i78.cg_elem.a ),
    .GATE_N(_0005_),
    .RESET_B(net368),
    .Q(\tokenflow_inst.i78.cg_elem.q ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i78.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i78.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[2] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i78.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i78.d0_elem.inv_chain[2] ),
    .X(\tokenflow_inst.i78.d0_elem.inv_chain[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0165_),
    .GATE_N(net38),
    .RESET_B(net369),
    .Q(\tokenflow_inst.i78.ydata[0] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0166_),
    .GATE_N(net36),
    .RESET_B(net370),
    .Q(\tokenflow_inst.i78.ydata[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0167_),
    .GATE_N(net36),
    .RESET_B(net371),
    .Q(\tokenflow_inst.i78.ydata[11] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0168_),
    .GATE_N(net36),
    .RESET_B(net372),
    .Q(\tokenflow_inst.i78.ydata[12] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0169_),
    .GATE_N(net34),
    .RESET_B(net373),
    .Q(\tokenflow_inst.i78.ydata[13] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0170_),
    .GATE_N(net35),
    .RESET_B(net374),
    .Q(\tokenflow_inst.i78.ydata[14] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0171_),
    .GATE_N(net32),
    .RESET_B(net375),
    .Q(\tokenflow_inst.i78.ydata[15] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0172_),
    .GATE_N(net34),
    .RESET_B(net376),
    .Q(\tokenflow_inst.i78.ydata[16] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0173_),
    .GATE_N(net32),
    .RESET_B(net377),
    .Q(\tokenflow_inst.i78.ydata[17] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0174_),
    .GATE_N(net32),
    .RESET_B(net378),
    .Q(\tokenflow_inst.i78.ydata[18] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0175_),
    .GATE_N(net33),
    .RESET_B(net379),
    .Q(\tokenflow_inst.i78.ydata[19] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0176_),
    .GATE_N(net40),
    .RESET_B(net380),
    .Q(\tokenflow_inst.i78.ydata[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0177_),
    .GATE_N(net32),
    .RESET_B(net381),
    .Q(\tokenflow_inst.i78.ydata[20] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0178_),
    .GATE_N(net34),
    .RESET_B(net382),
    .Q(\tokenflow_inst.i78.ydata[21] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0179_),
    .GATE_N(net30),
    .RESET_B(net383),
    .Q(\tokenflow_inst.i78.ydata[22] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0180_),
    .GATE_N(net31),
    .RESET_B(net384),
    .Q(\tokenflow_inst.i78.ydata[23] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0181_),
    .GATE_N(net30),
    .RESET_B(net385),
    .Q(\tokenflow_inst.i78.ydata[24] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0182_),
    .GATE_N(net37),
    .RESET_B(net386),
    .Q(\tokenflow_inst.i78.ydata[25] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0183_),
    .GATE_N(net38),
    .RESET_B(net387),
    .Q(\tokenflow_inst.i78.ydata[26] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0184_),
    .GATE_N(net41),
    .RESET_B(net388),
    .Q(\tokenflow_inst.i78.ydata[27] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0185_),
    .GATE_N(net38),
    .RESET_B(net389),
    .Q(\tokenflow_inst.i78.ydata[28] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0186_),
    .GATE_N(net41),
    .RESET_B(net390),
    .Q(\tokenflow_inst.i78.ydata[29] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0187_),
    .GATE_N(net40),
    .RESET_B(net391),
    .Q(\tokenflow_inst.i78.ydata[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0188_),
    .GATE_N(net38),
    .RESET_B(net392),
    .Q(\tokenflow_inst.i78.ydata[30] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0189_),
    .GATE_N(net38),
    .RESET_B(net393),
    .Q(\tokenflow_inst.i78.ydata[31] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0190_),
    .GATE_N(net38),
    .RESET_B(net394),
    .Q(\tokenflow_inst.i78.ydata[32] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0191_),
    .GATE_N(net38),
    .RESET_B(net395),
    .Q(\tokenflow_inst.i78.ydata[33] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0192_),
    .GATE_N(net37),
    .RESET_B(net396),
    .Q(\tokenflow_inst.i78.ydata[34] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0193_),
    .GATE_N(net37),
    .RESET_B(net397),
    .Q(\tokenflow_inst.i78.ydata[35] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0194_),
    .GATE_N(net37),
    .RESET_B(net398),
    .Q(\tokenflow_inst.i78.ydata[36] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0195_),
    .GATE_N(net37),
    .RESET_B(net399),
    .Q(\tokenflow_inst.i78.ydata[37] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0196_),
    .GATE_N(net37),
    .RESET_B(net400),
    .Q(\tokenflow_inst.i78.ydata[38] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0197_),
    .GATE_N(net34),
    .RESET_B(net401),
    .Q(\tokenflow_inst.i78.ydata[39] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0198_),
    .GATE_N(net40),
    .RESET_B(net402),
    .Q(\tokenflow_inst.i78.ydata[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0199_),
    .GATE_N(net34),
    .RESET_B(net403),
    .Q(\tokenflow_inst.i78.ydata[40] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0200_),
    .GATE_N(net34),
    .RESET_B(net404),
    .Q(\tokenflow_inst.i78.ydata[41] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0201_),
    .GATE_N(net31),
    .RESET_B(net405),
    .Q(\tokenflow_inst.i78.ydata[42] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0202_),
    .GATE_N(net31),
    .RESET_B(net406),
    .Q(\tokenflow_inst.i78.ydata[43] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0203_),
    .GATE_N(net30),
    .RESET_B(net407),
    .Q(\tokenflow_inst.i78.ydata[44] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0204_),
    .GATE_N(net30),
    .RESET_B(net408),
    .Q(\tokenflow_inst.i78.ydata[45] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0205_),
    .GATE_N(net30),
    .RESET_B(net409),
    .Q(\tokenflow_inst.i78.ydata[46] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0206_),
    .GATE_N(net31),
    .RESET_B(net410),
    .Q(\tokenflow_inst.i78.ydata[47] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0207_),
    .GATE_N(net31),
    .RESET_B(net411),
    .Q(\tokenflow_inst.i78.ydata[48] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0208_),
    .GATE_N(net34),
    .RESET_B(net412),
    .Q(\tokenflow_inst.i78.ydata[49] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0209_),
    .GATE_N(net40),
    .RESET_B(net413),
    .Q(\tokenflow_inst.i78.ydata[4] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0210_),
    .GATE_N(net38),
    .RESET_B(net414),
    .Q(\tokenflow_inst.i78.ydata[54] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0211_),
    .GATE_N(net40),
    .RESET_B(net415),
    .Q(\tokenflow_inst.i78.ydata[55] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0212_),
    .GATE_N(net39),
    .RESET_B(net416),
    .Q(\tokenflow_inst.i78.ydata[56] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0213_),
    .GATE_N(net39),
    .RESET_B(net417),
    .Q(\tokenflow_inst.i78.ydata[57] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0214_),
    .GATE_N(net39),
    .RESET_B(net418),
    .Q(\tokenflow_inst.i78.ydata[58] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0215_),
    .GATE_N(net39),
    .RESET_B(net419),
    .Q(\tokenflow_inst.i78.ydata[59] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0216_),
    .GATE_N(net39),
    .RESET_B(net420),
    .Q(\tokenflow_inst.i78.ydata[5] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0217_),
    .GATE_N(net39),
    .RESET_B(net421),
    .Q(\tokenflow_inst.i78.ydata[60] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0218_),
    .GATE_N(net36),
    .RESET_B(net422),
    .Q(\tokenflow_inst.i78.ydata[61] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0219_),
    .GATE_N(net36),
    .RESET_B(net423),
    .Q(\tokenflow_inst.i78.ydata[62] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0220_),
    .GATE_N(net36),
    .RESET_B(net424),
    .Q(\tokenflow_inst.i78.ydata[63] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0221_),
    .GATE_N(net36),
    .RESET_B(net425),
    .Q(\tokenflow_inst.i78.ydata[64] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0222_),
    .GATE_N(net34),
    .RESET_B(net426),
    .Q(\tokenflow_inst.i78.ydata[65] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0223_),
    .GATE_N(net35),
    .RESET_B(net427),
    .Q(\tokenflow_inst.i78.ydata[66] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0224_),
    .GATE_N(net33),
    .RESET_B(net428),
    .Q(\tokenflow_inst.i78.ydata[67] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0225_),
    .GATE_N(net33),
    .RESET_B(net429),
    .Q(\tokenflow_inst.i78.ydata[68] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0226_),
    .GATE_N(net32),
    .RESET_B(net430),
    .Q(\tokenflow_inst.i78.ydata[69] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0227_),
    .GATE_N(net39),
    .RESET_B(net431),
    .Q(\tokenflow_inst.i78.ydata[6] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0228_),
    .GATE_N(net32),
    .RESET_B(net432),
    .Q(\tokenflow_inst.i78.ydata[70] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0229_),
    .GATE_N(net32),
    .RESET_B(net433),
    .Q(\tokenflow_inst.i78.ydata[71] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0230_),
    .GATE_N(net32),
    .RESET_B(net434),
    .Q(\tokenflow_inst.i78.ydata[72] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0231_),
    .GATE_N(net30),
    .RESET_B(net435),
    .Q(\tokenflow_inst.i78.ydata[73] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0232_),
    .GATE_N(net31),
    .RESET_B(net436),
    .Q(\tokenflow_inst.i78.ydata[74] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0233_),
    .GATE_N(net30),
    .RESET_B(net437),
    .Q(\tokenflow_inst.i78.ydata[75] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0234_),
    .GATE_N(net30),
    .RESET_B(net438),
    .Q(\tokenflow_inst.i78.ydata[76] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0235_),
    .GATE_N(net37),
    .RESET_B(net439),
    .Q(\tokenflow_inst.i78.ydata[77] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0236_),
    .GATE_N(net39),
    .RESET_B(net440),
    .Q(\tokenflow_inst.i78.ydata[7] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0237_),
    .GATE_N(net42),
    .RESET_B(net441),
    .Q(\tokenflow_inst.i78.ydata[8] ));
 sg13g2_dllrq_1 \tokenflow_inst.i78.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0238_),
    .GATE_N(net36),
    .RESET_B(net442),
    .Q(\tokenflow_inst.i78.ydata[9] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.i8.cg_elem.a ),
    .GATE_N(_0004_),
    .RESET_B(net443),
    .Q(\tokenflow_inst.i8.cg_elem.q ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[0].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[0] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[10].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[10] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[11] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[11].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[11] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[12] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[12].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[12] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[13] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[13].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[13] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[14] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[14].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[14] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[15] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[15].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[15] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[16] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[16].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[16] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[17] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[17].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[17] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[18] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[18].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[18] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[19] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[19].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[19] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[20] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[2] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[20].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[20] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[21] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[21].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[21] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[22] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[22].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[22] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[23] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[23].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[23] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[24] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[24].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[24] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[25] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[25].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[25] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[26] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[26].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[26] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[27] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[27].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[27] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[28] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[28].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[28] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[29] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[29].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[29] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[30] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[2].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[2] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[3] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[30].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[30] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[31] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[31].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[31] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[32] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[32].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[32] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[33] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[33].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[33] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[34] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[34].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[34] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[35] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[35].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[35] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[36] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[36].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[36] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[37] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[37].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[37] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[38] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[38].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[38] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[39] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[39].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[39] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[40] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[3].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[3] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[4] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[40].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[40] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[41] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[41].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[41] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[42] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[42].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[42] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[43] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[43].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[43] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[44] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[44].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[44] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[45] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[45].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[45] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[46] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[46].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[46] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[47] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[47].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[47] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[48] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[48].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[48] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[49] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[49].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[49] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[50] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[4].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[4] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[5] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[50].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[50] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[51] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[51].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[51] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[52] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[5].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[5] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[6] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[6].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[6] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[7] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[7].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[7] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[8] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[8].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[8] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[9] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.i8.d0_elem.genblk1[9].min_delay_inst.d0  (.A(\tokenflow_inst.i8.d0_elem.inv_chain[9] ),
    .X(\tokenflow_inst.i8.d0_elem.inv_chain[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0240_),
    .GATE_N(net77),
    .RESET_B(net444),
    .Q(\tokenflow_inst.i8.ydata[0] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0241_),
    .GATE_N(net80),
    .RESET_B(net445),
    .Q(\tokenflow_inst.i8.ydata[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0242_),
    .GATE_N(net80),
    .RESET_B(net446),
    .Q(\tokenflow_inst.i8.ydata[11] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0243_),
    .GATE_N(net74),
    .RESET_B(net447),
    .Q(\tokenflow_inst.i8.ydata[12] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0244_),
    .GATE_N(net74),
    .RESET_B(net448),
    .Q(\tokenflow_inst.i8.ydata[13] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0245_),
    .GATE_N(net72),
    .RESET_B(net449),
    .Q(\tokenflow_inst.i8.ydata[14] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0246_),
    .GATE_N(net72),
    .RESET_B(net450),
    .Q(\tokenflow_inst.i8.ydata[15] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0247_),
    .GATE_N(net72),
    .RESET_B(net451),
    .Q(\tokenflow_inst.i8.ydata[16] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0248_),
    .GATE_N(net72),
    .RESET_B(net452),
    .Q(\tokenflow_inst.i8.ydata[17] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0249_),
    .GATE_N(net72),
    .RESET_B(net453),
    .Q(\tokenflow_inst.i8.ydata[18] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0250_),
    .GATE_N(net73),
    .RESET_B(net454),
    .Q(\tokenflow_inst.i8.ydata[19] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0251_),
    .GATE_N(net76),
    .RESET_B(net455),
    .Q(\tokenflow_inst.i8.ydata[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0252_),
    .GATE_N(net73),
    .RESET_B(net456),
    .Q(\tokenflow_inst.i8.ydata[20] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0253_),
    .GATE_N(net70),
    .RESET_B(net457),
    .Q(\tokenflow_inst.i8.ydata[21] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0254_),
    .GATE_N(net73),
    .RESET_B(net458),
    .Q(\tokenflow_inst.i8.ydata[22] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0255_),
    .GATE_N(net70),
    .RESET_B(net459),
    .Q(\tokenflow_inst.i8.ydata[23] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0256_),
    .GATE_N(net70),
    .RESET_B(net460),
    .Q(\tokenflow_inst.i8.ydata[24] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0257_),
    .GATE_N(net75),
    .RESET_B(net461),
    .Q(\tokenflow_inst.i8.ydata[25] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0258_),
    .GATE_N(net75),
    .RESET_B(net462),
    .Q(\tokenflow_inst.i8.ydata[26] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0259_),
    .GATE_N(net77),
    .RESET_B(net463),
    .Q(\tokenflow_inst.i8.ydata[27] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0260_),
    .GATE_N(net76),
    .RESET_B(net464),
    .Q(\tokenflow_inst.i8.ydata[28] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0261_),
    .GATE_N(net76),
    .RESET_B(net465),
    .Q(\tokenflow_inst.i8.ydata[29] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0262_),
    .GATE_N(net78),
    .RESET_B(net466),
    .Q(\tokenflow_inst.i8.ydata[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0263_),
    .GATE_N(net76),
    .RESET_B(net467),
    .Q(\tokenflow_inst.i8.ydata[30] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0264_),
    .GATE_N(net76),
    .RESET_B(net468),
    .Q(\tokenflow_inst.i8.ydata[31] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0265_),
    .GATE_N(net76),
    .RESET_B(net469),
    .Q(\tokenflow_inst.i8.ydata[32] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0266_),
    .GATE_N(net76),
    .RESET_B(net470),
    .Q(\tokenflow_inst.i8.ydata[33] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0267_),
    .GATE_N(net75),
    .RESET_B(net471),
    .Q(\tokenflow_inst.i8.ydata[34] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0268_),
    .GATE_N(net75),
    .RESET_B(net472),
    .Q(\tokenflow_inst.i8.ydata[35] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0269_),
    .GATE_N(net75),
    .RESET_B(net473),
    .Q(\tokenflow_inst.i8.ydata[36] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0270_),
    .GATE_N(net75),
    .RESET_B(net474),
    .Q(\tokenflow_inst.i8.ydata[37] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0271_),
    .GATE_N(net75),
    .RESET_B(net475),
    .Q(\tokenflow_inst.i8.ydata[38] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0272_),
    .GATE_N(net71),
    .RESET_B(net476),
    .Q(\tokenflow_inst.i8.ydata[39] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0273_),
    .GATE_N(net78),
    .RESET_B(net477),
    .Q(\tokenflow_inst.i8.ydata[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0274_),
    .GATE_N(net71),
    .RESET_B(net478),
    .Q(\tokenflow_inst.i8.ydata[40] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0275_),
    .GATE_N(net71),
    .RESET_B(net479),
    .Q(\tokenflow_inst.i8.ydata[41] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0276_),
    .GATE_N(net69),
    .RESET_B(net480),
    .Q(\tokenflow_inst.i8.ydata[42] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0277_),
    .GATE_N(net69),
    .RESET_B(net481),
    .Q(\tokenflow_inst.i8.ydata[43] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0278_),
    .GATE_N(net69),
    .RESET_B(net482),
    .Q(\tokenflow_inst.i8.ydata[44] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0279_),
    .GATE_N(net69),
    .RESET_B(net483),
    .Q(\tokenflow_inst.i8.ydata[45] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0280_),
    .GATE_N(net69),
    .RESET_B(net484),
    .Q(\tokenflow_inst.i8.ydata[46] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0281_),
    .GATE_N(net69),
    .RESET_B(net485),
    .Q(\tokenflow_inst.i8.ydata[47] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0282_),
    .GATE_N(net69),
    .RESET_B(net486),
    .Q(\tokenflow_inst.i8.ydata[48] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0283_),
    .GATE_N(net69),
    .RESET_B(net487),
    .Q(\tokenflow_inst.i8.ydata[49] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0284_),
    .GATE_N(net78),
    .RESET_B(net488),
    .Q(\tokenflow_inst.i8.ydata[4] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0285_),
    .GATE_N(net75),
    .RESET_B(net489),
    .Q(\tokenflow_inst.i8.ydata[50] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0286_),
    .GATE_N(net77),
    .RESET_B(net490),
    .Q(\tokenflow_inst.i8.ydata[53] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0287_),
    .GATE_N(net76),
    .RESET_B(net491),
    .Q(\tokenflow_inst.i8.ydata[54] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0288_),
    .GATE_N(net78),
    .RESET_B(net492),
    .Q(\tokenflow_inst.i8.ydata[55] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0289_),
    .GATE_N(net78),
    .RESET_B(net493),
    .Q(\tokenflow_inst.i8.ydata[56] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0290_),
    .GATE_N(net78),
    .RESET_B(net494),
    .Q(\tokenflow_inst.i8.ydata[57] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0291_),
    .GATE_N(net78),
    .RESET_B(net495),
    .Q(\tokenflow_inst.i8.ydata[58] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0292_),
    .GATE_N(net80),
    .RESET_B(net496),
    .Q(\tokenflow_inst.i8.ydata[59] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0293_),
    .GATE_N(net78),
    .RESET_B(net497),
    .Q(\tokenflow_inst.i8.ydata[5] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0294_),
    .GATE_N(net79),
    .RESET_B(net498),
    .Q(\tokenflow_inst.i8.ydata[60] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0295_),
    .GATE_N(net80),
    .RESET_B(net499),
    .Q(\tokenflow_inst.i8.ydata[61] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0296_),
    .GATE_N(net80),
    .RESET_B(net500),
    .Q(\tokenflow_inst.i8.ydata[62] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0297_),
    .GATE_N(net80),
    .RESET_B(net501),
    .Q(\tokenflow_inst.i8.ydata[63] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0298_),
    .GATE_N(net80),
    .RESET_B(net502),
    .Q(\tokenflow_inst.i8.ydata[64] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0299_),
    .GATE_N(net74),
    .RESET_B(net503),
    .Q(\tokenflow_inst.i8.ydata[65] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0300_),
    .GATE_N(net72),
    .RESET_B(net504),
    .Q(\tokenflow_inst.i8.ydata[66] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0301_),
    .GATE_N(net73),
    .RESET_B(net505),
    .Q(\tokenflow_inst.i8.ydata[67] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0302_),
    .GATE_N(net73),
    .RESET_B(net506),
    .Q(\tokenflow_inst.i8.ydata[68] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0303_),
    .GATE_N(net72),
    .RESET_B(net507),
    .Q(\tokenflow_inst.i8.ydata[69] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0304_),
    .GATE_N(net79),
    .RESET_B(net508),
    .Q(\tokenflow_inst.i8.ydata[6] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0305_),
    .GATE_N(net72),
    .RESET_B(net509),
    .Q(\tokenflow_inst.i8.ydata[70] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0306_),
    .GATE_N(net73),
    .RESET_B(net510),
    .Q(\tokenflow_inst.i8.ydata[71] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0307_),
    .GATE_N(net73),
    .RESET_B(net511),
    .Q(\tokenflow_inst.i8.ydata[72] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0308_),
    .GATE_N(net70),
    .RESET_B(net512),
    .Q(\tokenflow_inst.i8.ydata[73] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0309_),
    .GATE_N(net70),
    .RESET_B(net513),
    .Q(\tokenflow_inst.i8.ydata[74] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0310_),
    .GATE_N(net70),
    .RESET_B(net514),
    .Q(\tokenflow_inst.i8.ydata[75] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0311_),
    .GATE_N(net77),
    .RESET_B(net515),
    .Q(\tokenflow_inst.i8.ydata[76] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0312_),
    .GATE_N(net71),
    .RESET_B(net516),
    .Q(\tokenflow_inst.i8.ydata[77] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0313_),
    .GATE_N(net79),
    .RESET_B(net517),
    .Q(\tokenflow_inst.i8.ydata[7] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0314_),
    .GATE_N(net79),
    .RESET_B(net518),
    .Q(\tokenflow_inst.i8.ydata[8] ));
 sg13g2_dllrq_1 \tokenflow_inst.i8.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0315_),
    .GATE_N(net80),
    .RESET_B(net519),
    .Q(\tokenflow_inst.i8.ydata[9] ));
 sg13g2_dllrq_1 \tokenflow_inst.i9.c.q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net2),
    .GATE_N(net2),
    .RESET_B(net520),
    .Q(\tokenflow_inst.i9.c.q ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.ii1.d0_elem.genblk1[0].min_delay_inst.d0  (.A(net186),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.ii1.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.ii1.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.ii1.d0_elem.inv_chain[2] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.ii2.d0_elem.genblk1[0].min_delay_inst.d0  (.A(net198),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[1] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.ii2.d0_elem.genblk1[1].min_delay_inst.d0  (.A(\tokenflow_inst.ii2.d0_elem.inv_chain[1] ),
    .X(\tokenflow_inst.ii2.d0_elem.inv_chain[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[0] ),
    .GATE_N(net186),
    .RESET_B(net521),
    .Q(\tokenflow_inst.ii2.ydata[0] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[10] ),
    .GATE_N(net185),
    .RESET_B(net522),
    .Q(\tokenflow_inst.ii2.ydata[10] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[11] ),
    .GATE_N(net185),
    .RESET_B(net523),
    .Q(\tokenflow_inst.ii2.ydata[11] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[12] ),
    .GATE_N(net185),
    .RESET_B(net524),
    .Q(\tokenflow_inst.ii2.ydata[12] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[13] ),
    .GATE_N(net185),
    .RESET_B(net525),
    .Q(\tokenflow_inst.ii2.ydata[13] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[14] ),
    .GATE_N(net183),
    .RESET_B(net526),
    .Q(\tokenflow_inst.ii2.ydata[14] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[15] ),
    .GATE_N(net184),
    .RESET_B(net527),
    .Q(\tokenflow_inst.ii2.ydata[15] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[16] ),
    .GATE_N(net183),
    .RESET_B(net528),
    .Q(\tokenflow_inst.ii2.ydata[16] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[17] ),
    .GATE_N(net183),
    .RESET_B(net529),
    .Q(\tokenflow_inst.ii2.ydata[17] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[18] ),
    .GATE_N(net183),
    .RESET_B(net530),
    .Q(\tokenflow_inst.ii2.ydata[18] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[19] ),
    .GATE_N(net183),
    .RESET_B(net531),
    .Q(\tokenflow_inst.ii2.ydata[19] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[1] ),
    .GATE_N(net186),
    .RESET_B(net532),
    .Q(\tokenflow_inst.ii2.ydata[1] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[20] ),
    .GATE_N(net183),
    .RESET_B(net533),
    .Q(\tokenflow_inst.ii2.ydata[20] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[21] ),
    .GATE_N(net184),
    .RESET_B(net534),
    .Q(\tokenflow_inst.ii2.ydata[21] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[22] ),
    .GATE_N(net183),
    .RESET_B(net535),
    .Q(\tokenflow_inst.ii2.ydata[22] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[23] ),
    .GATE_N(net183),
    .RESET_B(net536),
    .Q(\tokenflow_inst.ii2.ydata[23] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[24] ),
    .GATE_N(net184),
    .RESET_B(net537),
    .Q(\tokenflow_inst.ii2.ydata[24] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[25] ),
    .GATE_N(net185),
    .RESET_B(net538),
    .Q(\tokenflow_inst.ii2.ydata[25] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[2] ),
    .GATE_N(net187),
    .RESET_B(net539),
    .Q(\tokenflow_inst.ii2.ydata[2] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[3] ),
    .GATE_N(net186),
    .RESET_B(net540),
    .Q(\tokenflow_inst.ii2.ydata[3] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[4] ),
    .GATE_N(net186),
    .RESET_B(net541),
    .Q(\tokenflow_inst.ii2.ydata[4] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[5] ),
    .GATE_N(net186),
    .RESET_B(net542),
    .Q(\tokenflow_inst.ii2.ydata[5] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[6] ),
    .GATE_N(net185),
    .RESET_B(net543),
    .Q(\tokenflow_inst.ii2.ydata[6] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[7] ),
    .GATE_N(net186),
    .RESET_B(net544),
    .Q(\tokenflow_inst.ii2.ydata[7] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[8] ),
    .GATE_N(net185),
    .RESET_B(net545),
    .Q(\tokenflow_inst.ii2.ydata[8] ));
 sg13g2_dllrq_1 \tokenflow_inst.ii2.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\tokenflow_inst.ii1.ydata[9] ),
    .GATE_N(net188),
    .RESET_B(net546),
    .Q(\tokenflow_inst.ii2.ydata[9] ));
 sg13g2_dlygate4sd3_1 \tokenflow_inst.ii3.i.d0_elem.genblk1[0].min_delay_inst.d0  (.A(net187),
    .X(\tokenflow_inst.ii3.i.d0_elem.inv_chain[1] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_0342_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0330_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0317_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1483_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1464_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1432_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1400_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1441_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1407_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1399_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1395_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(net31),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net35),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net35),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(net35),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net42),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(net37),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(net42),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(net41),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(net41),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net42),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(_0239_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0901_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0857_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0867_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0856_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0866_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0855_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1068_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0854_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1252_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1251_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1230_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1210_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1185_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1184_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1126_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1125_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1092_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1066_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1047_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1046_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1025_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1024_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1002_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0945_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0906_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0853_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net71),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net71),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(_0316_),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(_0316_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net77),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net81),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net81),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net81),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(_0316_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0411_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0380_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0362_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0379_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0361_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0378_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0360_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0435_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0359_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0532_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0358_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0783_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0780_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0766_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0765_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0754_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0729_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0728_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0714_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0712_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0692_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0691_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0667_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0637_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0625_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0624_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0583_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0581_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0577_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0576_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0554_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0511_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0491_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0490_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0486_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0485_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(_0164_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net123),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(_0164_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net126),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(net129),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(_0164_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net136),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(_0085_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net139),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0085_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net142),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(_0085_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0982_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0852_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0605_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0400_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0351_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0339_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0326_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1492_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_1480_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_1457_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_1428_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_1393_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_1347_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_1317_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_1296_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_1189_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0851_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0850_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0849_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0848_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0847_),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(_1456_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_1449_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_1403_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1392_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_1388_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_1387_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_1385_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_1384_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_1383_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_1382_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_1381_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_1380_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_1299_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_1298_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_1297_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_1391_),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(_1386_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_1379_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_1378_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net188),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net188),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net1),
    .X(net188));
 sg13g2_tielo _3068__189 (.L_LO(net189));
 sg13g2_tielo _3070__190 (.L_LO(net190));
 sg13g2_tielo _3071__191 (.L_LO(net191));
 sg13g2_tielo _3072__192 (.L_LO(net192));
 sg13g2_tielo _3074__193 (.L_LO(net193));
 sg13g2_tielo _3075__194 (.L_LO(net194));
 sg13g2_tielo _3076__195 (.L_LO(net195));
 sg13g2_tielo _3077__196 (.L_LO(net196));
 sg13g2_tielo \tokenflow_inst.i10.d0.genblk1[0].min_delay_inst.d0_197  (.L_LO(net197));
 sg13g2_tielo \tokenflow_inst.ii2.d0_elem.genblk1[0].min_delay_inst.d0_198  (.L_LO(net198));
 sg13g2_tiehi _3079__200 (.L_HI(net200));
 sg13g2_tiehi _3080__201 (.L_HI(net201));
 sg13g2_tiehi _3081__202 (.L_HI(net202));
 sg13g2_tiehi _3082__203 (.L_HI(net203));
 sg13g2_tiehi _3083__204 (.L_HI(net204));
 sg13g2_tiehi _3084__205 (.L_HI(net205));
 sg13g2_tiehi _3085__206 (.L_HI(net206));
 sg13g2_tiehi \tokenflow_inst.i1.c.q$_DLATCH_N_._TECHMAP_DLATCH_N_207  (.L_HI(net207));
 sg13g2_tiehi \tokenflow_inst.i2.cg1.q$_DLATCH_N_._TECHMAP_DLATCH_N_208  (.L_HI(net208));
 sg13g2_tiehi \tokenflow_inst.i2.cg2.q$_DLATCH_N_._TECHMAP_DLATCH_N_209  (.L_HI(net209));
 sg13g2_tiehi \tokenflow_inst.i3.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N_210  (.L_HI(net210));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N_211  (.L_HI(net211));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N_212  (.L_HI(net212));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N_213  (.L_HI(net213));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N_214  (.L_HI(net214));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N_215  (.L_HI(net215));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N_216  (.L_HI(net216));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N_217  (.L_HI(net217));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N_218  (.L_HI(net218));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N_219  (.L_HI(net219));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N_220  (.L_HI(net220));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N_221  (.L_HI(net221));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N_222  (.L_HI(net222));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N_223  (.L_HI(net223));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N_224  (.L_HI(net224));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N_225  (.L_HI(net225));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N_226  (.L_HI(net226));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N_227  (.L_HI(net227));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N_228  (.L_HI(net228));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N_229  (.L_HI(net229));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N_230  (.L_HI(net230));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N_231  (.L_HI(net231));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N_232  (.L_HI(net232));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N_233  (.L_HI(net233));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N_234  (.L_HI(net234));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N_235  (.L_HI(net235));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N_236  (.L_HI(net236));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N_237  (.L_HI(net237));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N_238  (.L_HI(net238));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N_239  (.L_HI(net239));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N_240  (.L_HI(net240));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N_241  (.L_HI(net241));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N_242  (.L_HI(net242));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N_243  (.L_HI(net243));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N_244  (.L_HI(net244));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N_245  (.L_HI(net245));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N_246  (.L_HI(net246));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N_247  (.L_HI(net247));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N_248  (.L_HI(net248));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N_249  (.L_HI(net249));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N_250  (.L_HI(net250));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N_251  (.L_HI(net251));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N_252  (.L_HI(net252));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N_253  (.L_HI(net253));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N_254  (.L_HI(net254));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N_255  (.L_HI(net255));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N_256  (.L_HI(net256));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[51]$_DLATCH_N_._TECHMAP_DLATCH_N_257  (.L_HI(net257));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[52]$_DLATCH_N_._TECHMAP_DLATCH_N_258  (.L_HI(net258));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N_259  (.L_HI(net259));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N_260  (.L_HI(net260));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N_261  (.L_HI(net261));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N_262  (.L_HI(net262));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N_263  (.L_HI(net263));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N_264  (.L_HI(net264));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N_265  (.L_HI(net265));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N_266  (.L_HI(net266));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N_267  (.L_HI(net267));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N_268  (.L_HI(net268));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N_269  (.L_HI(net269));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N_270  (.L_HI(net270));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N_271  (.L_HI(net271));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N_272  (.L_HI(net272));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N_273  (.L_HI(net273));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N_274  (.L_HI(net274));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N_275  (.L_HI(net275));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N_276  (.L_HI(net276));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N_277  (.L_HI(net277));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N_278  (.L_HI(net278));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N_279  (.L_HI(net279));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N_280  (.L_HI(net280));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N_281  (.L_HI(net281));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N_282  (.L_HI(net282));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N_283  (.L_HI(net283));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N_284  (.L_HI(net284));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N_285  (.L_HI(net285));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N_286  (.L_HI(net286));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N_287  (.L_HI(net287));
 sg13g2_tiehi \tokenflow_inst.i3.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N_288  (.L_HI(net288));
 sg13g2_tiehi \tokenflow_inst.i6.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N_289  (.L_HI(net289));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N_290  (.L_HI(net290));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N_291  (.L_HI(net291));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N_292  (.L_HI(net292));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N_293  (.L_HI(net293));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N_294  (.L_HI(net294));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N_295  (.L_HI(net295));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N_296  (.L_HI(net296));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N_297  (.L_HI(net297));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N_298  (.L_HI(net298));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N_299  (.L_HI(net299));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N_300  (.L_HI(net300));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N_301  (.L_HI(net301));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N_302  (.L_HI(net302));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N_303  (.L_HI(net303));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N_304  (.L_HI(net304));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N_305  (.L_HI(net305));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N_306  (.L_HI(net306));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N_307  (.L_HI(net307));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N_308  (.L_HI(net308));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N_309  (.L_HI(net309));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N_310  (.L_HI(net310));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N_311  (.L_HI(net311));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N_312  (.L_HI(net312));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N_313  (.L_HI(net313));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N_314  (.L_HI(net314));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N_315  (.L_HI(net315));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N_316  (.L_HI(net316));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N_317  (.L_HI(net317));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N_318  (.L_HI(net318));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N_319  (.L_HI(net319));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N_320  (.L_HI(net320));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N_321  (.L_HI(net321));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N_322  (.L_HI(net322));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N_323  (.L_HI(net323));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N_324  (.L_HI(net324));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N_325  (.L_HI(net325));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N_326  (.L_HI(net326));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N_327  (.L_HI(net327));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N_328  (.L_HI(net328));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N_329  (.L_HI(net329));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N_330  (.L_HI(net330));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N_331  (.L_HI(net331));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N_332  (.L_HI(net332));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N_333  (.L_HI(net333));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N_334  (.L_HI(net334));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N_335  (.L_HI(net335));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[51]$_DLATCH_N_._TECHMAP_DLATCH_N_336  (.L_HI(net336));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[52]$_DLATCH_N_._TECHMAP_DLATCH_N_337  (.L_HI(net337));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N_338  (.L_HI(net338));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N_339  (.L_HI(net339));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N_340  (.L_HI(net340));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N_341  (.L_HI(net341));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N_342  (.L_HI(net342));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N_343  (.L_HI(net343));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N_344  (.L_HI(net344));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N_345  (.L_HI(net345));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N_346  (.L_HI(net346));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N_347  (.L_HI(net347));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N_348  (.L_HI(net348));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N_349  (.L_HI(net349));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N_350  (.L_HI(net350));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N_351  (.L_HI(net351));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N_352  (.L_HI(net352));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N_353  (.L_HI(net353));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N_354  (.L_HI(net354));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N_355  (.L_HI(net355));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N_356  (.L_HI(net356));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N_357  (.L_HI(net357));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N_358  (.L_HI(net358));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N_359  (.L_HI(net359));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N_360  (.L_HI(net360));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N_361  (.L_HI(net361));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N_362  (.L_HI(net362));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N_363  (.L_HI(net363));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N_364  (.L_HI(net364));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N_365  (.L_HI(net365));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N_366  (.L_HI(net366));
 sg13g2_tiehi \tokenflow_inst.i6.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N_367  (.L_HI(net367));
 sg13g2_tiehi \tokenflow_inst.i78.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N_368  (.L_HI(net368));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N_369  (.L_HI(net369));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N_370  (.L_HI(net370));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N_371  (.L_HI(net371));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N_372  (.L_HI(net372));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N_373  (.L_HI(net373));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N_374  (.L_HI(net374));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N_375  (.L_HI(net375));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N_376  (.L_HI(net376));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N_377  (.L_HI(net377));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N_378  (.L_HI(net378));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N_379  (.L_HI(net379));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N_380  (.L_HI(net380));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N_381  (.L_HI(net381));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N_382  (.L_HI(net382));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N_383  (.L_HI(net383));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N_384  (.L_HI(net384));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N_385  (.L_HI(net385));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N_386  (.L_HI(net386));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N_387  (.L_HI(net387));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N_388  (.L_HI(net388));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N_389  (.L_HI(net389));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N_390  (.L_HI(net390));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N_391  (.L_HI(net391));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N_392  (.L_HI(net392));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N_393  (.L_HI(net393));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N_394  (.L_HI(net394));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N_395  (.L_HI(net395));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N_396  (.L_HI(net396));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N_397  (.L_HI(net397));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N_398  (.L_HI(net398));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N_399  (.L_HI(net399));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N_400  (.L_HI(net400));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N_401  (.L_HI(net401));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N_402  (.L_HI(net402));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N_403  (.L_HI(net403));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N_404  (.L_HI(net404));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N_405  (.L_HI(net405));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N_406  (.L_HI(net406));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N_407  (.L_HI(net407));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N_408  (.L_HI(net408));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N_409  (.L_HI(net409));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N_410  (.L_HI(net410));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N_411  (.L_HI(net411));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N_412  (.L_HI(net412));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N_413  (.L_HI(net413));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N_414  (.L_HI(net414));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N_415  (.L_HI(net415));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N_416  (.L_HI(net416));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N_417  (.L_HI(net417));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N_418  (.L_HI(net418));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N_419  (.L_HI(net419));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N_420  (.L_HI(net420));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N_421  (.L_HI(net421));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N_422  (.L_HI(net422));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N_423  (.L_HI(net423));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N_424  (.L_HI(net424));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N_425  (.L_HI(net425));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N_426  (.L_HI(net426));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N_427  (.L_HI(net427));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N_428  (.L_HI(net428));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N_429  (.L_HI(net429));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N_430  (.L_HI(net430));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N_431  (.L_HI(net431));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N_432  (.L_HI(net432));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N_433  (.L_HI(net433));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N_434  (.L_HI(net434));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N_435  (.L_HI(net435));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N_436  (.L_HI(net436));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N_437  (.L_HI(net437));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N_438  (.L_HI(net438));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N_439  (.L_HI(net439));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N_440  (.L_HI(net440));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N_441  (.L_HI(net441));
 sg13g2_tiehi \tokenflow_inst.i78.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N_442  (.L_HI(net442));
 sg13g2_tiehi \tokenflow_inst.i8.cg_elem.q$_DLATCH_N_._TECHMAP_DLATCH_N_443  (.L_HI(net443));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N_444  (.L_HI(net444));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N_445  (.L_HI(net445));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N_446  (.L_HI(net446));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N_447  (.L_HI(net447));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N_448  (.L_HI(net448));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N_449  (.L_HI(net449));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N_450  (.L_HI(net450));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N_451  (.L_HI(net451));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N_452  (.L_HI(net452));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N_453  (.L_HI(net453));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N_454  (.L_HI(net454));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N_455  (.L_HI(net455));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N_456  (.L_HI(net456));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N_457  (.L_HI(net457));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N_458  (.L_HI(net458));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N_459  (.L_HI(net459));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N_460  (.L_HI(net460));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N_461  (.L_HI(net461));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[26]$_DLATCH_N_._TECHMAP_DLATCH_N_462  (.L_HI(net462));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[27]$_DLATCH_N_._TECHMAP_DLATCH_N_463  (.L_HI(net463));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[28]$_DLATCH_N_._TECHMAP_DLATCH_N_464  (.L_HI(net464));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[29]$_DLATCH_N_._TECHMAP_DLATCH_N_465  (.L_HI(net465));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N_466  (.L_HI(net466));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[30]$_DLATCH_N_._TECHMAP_DLATCH_N_467  (.L_HI(net467));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[31]$_DLATCH_N_._TECHMAP_DLATCH_N_468  (.L_HI(net468));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[32]$_DLATCH_N_._TECHMAP_DLATCH_N_469  (.L_HI(net469));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[33]$_DLATCH_N_._TECHMAP_DLATCH_N_470  (.L_HI(net470));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[34]$_DLATCH_N_._TECHMAP_DLATCH_N_471  (.L_HI(net471));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[35]$_DLATCH_N_._TECHMAP_DLATCH_N_472  (.L_HI(net472));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[36]$_DLATCH_N_._TECHMAP_DLATCH_N_473  (.L_HI(net473));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[37]$_DLATCH_N_._TECHMAP_DLATCH_N_474  (.L_HI(net474));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[38]$_DLATCH_N_._TECHMAP_DLATCH_N_475  (.L_HI(net475));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[39]$_DLATCH_N_._TECHMAP_DLATCH_N_476  (.L_HI(net476));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N_477  (.L_HI(net477));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[40]$_DLATCH_N_._TECHMAP_DLATCH_N_478  (.L_HI(net478));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[41]$_DLATCH_N_._TECHMAP_DLATCH_N_479  (.L_HI(net479));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[42]$_DLATCH_N_._TECHMAP_DLATCH_N_480  (.L_HI(net480));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[43]$_DLATCH_N_._TECHMAP_DLATCH_N_481  (.L_HI(net481));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[44]$_DLATCH_N_._TECHMAP_DLATCH_N_482  (.L_HI(net482));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[45]$_DLATCH_N_._TECHMAP_DLATCH_N_483  (.L_HI(net483));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[46]$_DLATCH_N_._TECHMAP_DLATCH_N_484  (.L_HI(net484));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[47]$_DLATCH_N_._TECHMAP_DLATCH_N_485  (.L_HI(net485));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[48]$_DLATCH_N_._TECHMAP_DLATCH_N_486  (.L_HI(net486));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[49]$_DLATCH_N_._TECHMAP_DLATCH_N_487  (.L_HI(net487));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N_488  (.L_HI(net488));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[50]$_DLATCH_N_._TECHMAP_DLATCH_N_489  (.L_HI(net489));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[53]$_DLATCH_N_._TECHMAP_DLATCH_N_490  (.L_HI(net490));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[54]$_DLATCH_N_._TECHMAP_DLATCH_N_491  (.L_HI(net491));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[55]$_DLATCH_N_._TECHMAP_DLATCH_N_492  (.L_HI(net492));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[56]$_DLATCH_N_._TECHMAP_DLATCH_N_493  (.L_HI(net493));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[57]$_DLATCH_N_._TECHMAP_DLATCH_N_494  (.L_HI(net494));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[58]$_DLATCH_N_._TECHMAP_DLATCH_N_495  (.L_HI(net495));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[59]$_DLATCH_N_._TECHMAP_DLATCH_N_496  (.L_HI(net496));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N_497  (.L_HI(net497));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[60]$_DLATCH_N_._TECHMAP_DLATCH_N_498  (.L_HI(net498));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[61]$_DLATCH_N_._TECHMAP_DLATCH_N_499  (.L_HI(net499));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[62]$_DLATCH_N_._TECHMAP_DLATCH_N_500  (.L_HI(net500));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[63]$_DLATCH_N_._TECHMAP_DLATCH_N_501  (.L_HI(net501));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[64]$_DLATCH_N_._TECHMAP_DLATCH_N_502  (.L_HI(net502));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[65]$_DLATCH_N_._TECHMAP_DLATCH_N_503  (.L_HI(net503));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[66]$_DLATCH_N_._TECHMAP_DLATCH_N_504  (.L_HI(net504));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[67]$_DLATCH_N_._TECHMAP_DLATCH_N_505  (.L_HI(net505));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[68]$_DLATCH_N_._TECHMAP_DLATCH_N_506  (.L_HI(net506));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[69]$_DLATCH_N_._TECHMAP_DLATCH_N_507  (.L_HI(net507));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N_508  (.L_HI(net508));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[70]$_DLATCH_N_._TECHMAP_DLATCH_N_509  (.L_HI(net509));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[71]$_DLATCH_N_._TECHMAP_DLATCH_N_510  (.L_HI(net510));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[72]$_DLATCH_N_._TECHMAP_DLATCH_N_511  (.L_HI(net511));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[73]$_DLATCH_N_._TECHMAP_DLATCH_N_512  (.L_HI(net512));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[74]$_DLATCH_N_._TECHMAP_DLATCH_N_513  (.L_HI(net513));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[75]$_DLATCH_N_._TECHMAP_DLATCH_N_514  (.L_HI(net514));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[76]$_DLATCH_N_._TECHMAP_DLATCH_N_515  (.L_HI(net515));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[77]$_DLATCH_N_._TECHMAP_DLATCH_N_516  (.L_HI(net516));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N_517  (.L_HI(net517));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N_518  (.L_HI(net518));
 sg13g2_tiehi \tokenflow_inst.i8.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N_519  (.L_HI(net519));
 sg13g2_tiehi \tokenflow_inst.i9.c.q$_DLATCH_N_._TECHMAP_DLATCH_N_520  (.L_HI(net520));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[0]$_DLATCH_N_._TECHMAP_DLATCH_N_521  (.L_HI(net521));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[10]$_DLATCH_N_._TECHMAP_DLATCH_N_522  (.L_HI(net522));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[11]$_DLATCH_N_._TECHMAP_DLATCH_N_523  (.L_HI(net523));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[12]$_DLATCH_N_._TECHMAP_DLATCH_N_524  (.L_HI(net524));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[13]$_DLATCH_N_._TECHMAP_DLATCH_N_525  (.L_HI(net525));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[14]$_DLATCH_N_._TECHMAP_DLATCH_N_526  (.L_HI(net526));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[15]$_DLATCH_N_._TECHMAP_DLATCH_N_527  (.L_HI(net527));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[16]$_DLATCH_N_._TECHMAP_DLATCH_N_528  (.L_HI(net528));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[17]$_DLATCH_N_._TECHMAP_DLATCH_N_529  (.L_HI(net529));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[18]$_DLATCH_N_._TECHMAP_DLATCH_N_530  (.L_HI(net530));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[19]$_DLATCH_N_._TECHMAP_DLATCH_N_531  (.L_HI(net531));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[1]$_DLATCH_N_._TECHMAP_DLATCH_N_532  (.L_HI(net532));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[20]$_DLATCH_N_._TECHMAP_DLATCH_N_533  (.L_HI(net533));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[21]$_DLATCH_N_._TECHMAP_DLATCH_N_534  (.L_HI(net534));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[22]$_DLATCH_N_._TECHMAP_DLATCH_N_535  (.L_HI(net535));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[23]$_DLATCH_N_._TECHMAP_DLATCH_N_536  (.L_HI(net536));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[24]$_DLATCH_N_._TECHMAP_DLATCH_N_537  (.L_HI(net537));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[25]$_DLATCH_N_._TECHMAP_DLATCH_N_538  (.L_HI(net538));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[2]$_DLATCH_N_._TECHMAP_DLATCH_N_539  (.L_HI(net539));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[3]$_DLATCH_N_._TECHMAP_DLATCH_N_540  (.L_HI(net540));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[4]$_DLATCH_N_._TECHMAP_DLATCH_N_541  (.L_HI(net541));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[5]$_DLATCH_N_._TECHMAP_DLATCH_N_542  (.L_HI(net542));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[6]$_DLATCH_N_._TECHMAP_DLATCH_N_543  (.L_HI(net543));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[7]$_DLATCH_N_._TECHMAP_DLATCH_N_544  (.L_HI(net544));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[8]$_DLATCH_N_._TECHMAP_DLATCH_N_545  (.L_HI(net545));
 sg13g2_tiehi \tokenflow_inst.ii2.ydata[9]$_DLATCH_N_._TECHMAP_DLATCH_N_546  (.L_HI(net546));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_fill_2 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_fill_2 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_4 FILLER_1_159 ();
 sg13g2_fill_2 FILLER_1_172 ();
 sg13g2_fill_1 FILLER_1_174 ();
 sg13g2_fill_2 FILLER_1_179 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_decap_4 FILLER_1_198 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_fill_2 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_fill_2 FILLER_1_233 ();
 sg13g2_fill_1 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_4 FILLER_1_319 ();
 sg13g2_fill_1 FILLER_1_323 ();
 sg13g2_fill_2 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_4 FILLER_2_150 ();
 sg13g2_fill_2 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_fill_1 FILLER_2_197 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_232 ();
 sg13g2_fill_2 FILLER_2_237 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_278 ();
 sg13g2_decap_8 FILLER_2_285 ();
 sg13g2_fill_2 FILLER_2_292 ();
 sg13g2_decap_4 FILLER_2_302 ();
 sg13g2_decap_4 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_4 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_123 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_144 ();
 sg13g2_fill_1 FILLER_3_153 ();
 sg13g2_fill_1 FILLER_3_181 ();
 sg13g2_decap_4 FILLER_3_188 ();
 sg13g2_fill_2 FILLER_3_197 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_fill_2 FILLER_3_262 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_274 ();
 sg13g2_decap_4 FILLER_3_290 ();
 sg13g2_fill_1 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_fill_2 FILLER_3_318 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_decap_4 FILLER_3_329 ();
 sg13g2_fill_2 FILLER_3_333 ();
 sg13g2_fill_1 FILLER_3_343 ();
 sg13g2_fill_1 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_decap_8 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_157 ();
 sg13g2_decap_4 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_fill_2 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_226 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_fill_1 FILLER_4_255 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_4 FILLER_4_306 ();
 sg13g2_fill_1 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_4 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_136 ();
 sg13g2_fill_2 FILLER_5_143 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_fill_2 FILLER_5_154 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_167 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_fill_2 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_4 FILLER_5_242 ();
 sg13g2_fill_2 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_4 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_fill_2 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_151 ();
 sg13g2_fill_2 FILLER_6_182 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_201 ();
 sg13g2_decap_4 FILLER_6_208 ();
 sg13g2_decap_4 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_225 ();
 sg13g2_decap_4 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_234 ();
 sg13g2_decap_4 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_260 ();
 sg13g2_decap_4 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_4 FILLER_6_424 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_143 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_fill_1 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_decap_4 FILLER_7_309 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_decap_4 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_decap_4 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_299 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_313 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_8 FILLER_8_404 ();
 sg13g2_decap_8 FILLER_8_411 ();
 sg13g2_decap_8 FILLER_8_418 ();
 sg13g2_decap_4 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_76 ();
 sg13g2_fill_2 FILLER_9_80 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_4 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_decap_4 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_decap_4 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_fill_2 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_decap_4 FILLER_10_152 ();
 sg13g2_decap_4 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_decap_4 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_275 ();
 sg13g2_fill_2 FILLER_10_280 ();
 sg13g2_fill_1 FILLER_10_282 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_291 ();
 sg13g2_decap_4 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_302 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_fill_1 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_118 ();
 sg13g2_decap_4 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_4 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_4 FILLER_11_308 ();
 sg13g2_fill_2 FILLER_11_312 ();
 sg13g2_decap_4 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_68 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_82 ();
 sg13g2_decap_4 FILLER_12_113 ();
 sg13g2_fill_1 FILLER_12_117 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_decap_8 FILLER_12_141 ();
 sg13g2_fill_2 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_78 ();
 sg13g2_fill_2 FILLER_13_83 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_decap_8 FILLER_13_106 ();
 sg13g2_decap_8 FILLER_13_113 ();
 sg13g2_decap_4 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_271 ();
 sg13g2_decap_4 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_decap_8 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_13_414 ();
 sg13g2_decap_8 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_4 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_74 ();
 sg13g2_fill_1 FILLER_14_95 ();
 sg13g2_fill_2 FILLER_14_100 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_107 ();
 sg13g2_decap_4 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_decap_4 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_decap_4 FILLER_14_172 ();
 sg13g2_decap_4 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_64 ();
 sg13g2_decap_8 FILLER_15_72 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_decap_4 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_decap_4 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_decap_4 FILLER_15_154 ();
 sg13g2_decap_4 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_208 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_278 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_411 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_fill_2 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_4 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_decap_4 FILLER_17_108 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_4 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_58 ();
 sg13g2_decap_4 FILLER_18_67 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_1 FILLER_18_148 ();
 sg13g2_fill_2 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_227 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_decap_4 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_decap_4 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_decap_8 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_68 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_decap_4 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_215 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_318 ();
 sg13g2_decap_4 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_8 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_62 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_decap_8 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_4 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_decap_4 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_decap_4 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_decap_8 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_decap_8 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_decap_8 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_decap_4 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_25_409 ();
 sg13g2_decap_8 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_4 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_4 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_4 FILLER_27_287 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_decap_4 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_51 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_decap_8 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_4 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_decap_4 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_decap_4 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_197 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_4 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_decap_8 FILLER_30_411 ();
 sg13g2_decap_8 FILLER_30_418 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_8 FILLER_31_404 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_decap_4 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_83 ();
 sg13g2_decap_4 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_decap_8 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_8 FILLER_33_404 ();
 sg13g2_decap_8 FILLER_33_411 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_86 ();
 sg13g2_fill_1 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_4 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_decap_4 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_decap_4 FILLER_35_255 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_4 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_decap_8 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_4 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_239 ();
 sg13g2_decap_4 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_274 ();
 sg13g2_decap_4 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_decap_4 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_decap_4 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_decap_4 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_229 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_4 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_decap_8 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_414 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_64 ();
 sg13g2_fill_1 FILLER_38_66 ();
 sg13g2_decap_8 FILLER_38_83 ();
 sg13g2_decap_8 FILLER_38_90 ();
 sg13g2_decap_8 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_decap_4 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_171 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_336 ();
 sg13g2_decap_4 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_416 ();
 sg13g2_decap_8 FILLER_38_423 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_76 ();
 sg13g2_decap_8 FILLER_39_82 ();
 sg13g2_fill_2 FILLER_39_89 ();
 sg13g2_fill_1 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_104 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_decap_4 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_127 ();
 sg13g2_decap_4 FILLER_39_141 ();
 sg13g2_fill_2 FILLER_39_174 ();
 sg13g2_fill_2 FILLER_39_219 ();
 sg13g2_decap_4 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_251 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_2 FILLER_39_280 ();
 sg13g2_decap_4 FILLER_39_292 ();
 sg13g2_decap_8 FILLER_39_304 ();
 sg13g2_decap_4 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_decap_4 FILLER_39_327 ();
 sg13g2_fill_2 FILLER_39_331 ();
 sg13g2_decap_4 FILLER_39_338 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_fill_2 FILLER_39_427 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_fill_2 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_62 ();
 sg13g2_decap_4 FILLER_40_85 ();
 sg13g2_decap_8 FILLER_40_93 ();
 sg13g2_fill_2 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_134 ();
 sg13g2_decap_4 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_158 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_fill_1 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_191 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_2 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_decap_4 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_decap_4 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_fill_2 FILLER_40_290 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_decap_4 FILLER_40_317 ();
 sg13g2_decap_4 FILLER_40_337 ();
 sg13g2_fill_2 FILLER_40_341 ();
 sg13g2_fill_1 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_377 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_419 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_4 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_53 ();
 sg13g2_decap_4 FILLER_41_59 ();
 sg13g2_fill_2 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_96 ();
 sg13g2_fill_2 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_119 ();
 sg13g2_fill_2 FILLER_41_125 ();
 sg13g2_decap_4 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_fill_2 FILLER_41_171 ();
 sg13g2_fill_1 FILLER_41_173 ();
 sg13g2_decap_4 FILLER_41_178 ();
 sg13g2_fill_2 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_205 ();
 sg13g2_fill_1 FILLER_41_207 ();
 sg13g2_decap_4 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_262 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_fill_2 FILLER_41_273 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_4 FILLER_41_308 ();
 sg13g2_fill_2 FILLER_41_316 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_8 FILLER_41_403 ();
 sg13g2_decap_8 FILLER_41_410 ();
 sg13g2_decap_8 FILLER_41_417 ();
 sg13g2_decap_4 FILLER_41_424 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_60 ();
 sg13g2_fill_2 FILLER_42_67 ();
 sg13g2_decap_4 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_fill_1 FILLER_42_129 ();
 sg13g2_decap_4 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_146 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_42_154 ();
 sg13g2_fill_2 FILLER_42_181 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_decap_8 FILLER_42_218 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_decap_4 FILLER_42_231 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_2 FILLER_42_249 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_decap_4 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_decap_8 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_decap_4 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_46 ();
 sg13g2_fill_1 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_decap_4 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_102 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_decap_8 FILLER_43_120 ();
 sg13g2_decap_4 FILLER_43_127 ();
 sg13g2_fill_1 FILLER_43_131 ();
 sg13g2_decap_8 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_150 ();
 sg13g2_decap_4 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_234 ();
 sg13g2_decap_8 FILLER_43_241 ();
 sg13g2_decap_8 FILLER_43_248 ();
 sg13g2_decap_8 FILLER_43_255 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_fill_1 FILLER_43_292 ();
 sg13g2_decap_4 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_fill_2 FILLER_43_324 ();
 sg13g2_fill_2 FILLER_43_330 ();
 sg13g2_fill_2 FILLER_43_336 ();
 sg13g2_fill_1 FILLER_43_338 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_354 ();
 sg13g2_fill_1 FILLER_43_356 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_fill_2 FILLER_43_427 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_89 ();
 sg13g2_decap_4 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_104 ();
 sg13g2_decap_4 FILLER_44_111 ();
 sg13g2_fill_2 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_137 ();
 sg13g2_fill_2 FILLER_44_153 ();
 sg13g2_fill_1 FILLER_44_155 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_188 ();
 sg13g2_fill_2 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_decap_8 FILLER_44_240 ();
 sg13g2_decap_4 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_4 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_309 ();
 sg13g2_fill_2 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_334 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_decap_4 FILLER_44_352 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_4 FILLER_44_424 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_55 ();
 sg13g2_decap_8 FILLER_45_62 ();
 sg13g2_decap_8 FILLER_45_69 ();
 sg13g2_decap_4 FILLER_45_80 ();
 sg13g2_decap_8 FILLER_45_89 ();
 sg13g2_fill_1 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_101 ();
 sg13g2_fill_1 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_128 ();
 sg13g2_fill_2 FILLER_45_133 ();
 sg13g2_fill_2 FILLER_45_139 ();
 sg13g2_decap_8 FILLER_45_145 ();
 sg13g2_decap_4 FILLER_45_152 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_decap_4 FILLER_45_223 ();
 sg13g2_fill_1 FILLER_45_236 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_258 ();
 sg13g2_decap_8 FILLER_45_265 ();
 sg13g2_fill_1 FILLER_45_272 ();
 sg13g2_decap_4 FILLER_45_282 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_decap_4 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_decap_8 FILLER_45_317 ();
 sg13g2_decap_4 FILLER_45_344 ();
 sg13g2_fill_1 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_369 ();
 sg13g2_decap_8 FILLER_45_376 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_8 FILLER_45_404 ();
 sg13g2_decap_8 FILLER_45_411 ();
 sg13g2_decap_8 FILLER_45_418 ();
 sg13g2_decap_4 FILLER_45_425 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_58 ();
 sg13g2_fill_1 FILLER_46_60 ();
 sg13g2_fill_1 FILLER_46_90 ();
 sg13g2_fill_2 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_129 ();
 sg13g2_decap_4 FILLER_46_149 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_decap_8 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_170 ();
 sg13g2_decap_4 FILLER_46_183 ();
 sg13g2_fill_2 FILLER_46_192 ();
 sg13g2_fill_1 FILLER_46_202 ();
 sg13g2_fill_1 FILLER_46_208 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_fill_2 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_decap_4 FILLER_46_258 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_decap_4 FILLER_46_278 ();
 sg13g2_fill_1 FILLER_46_282 ();
 sg13g2_decap_4 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_321 ();
 sg13g2_fill_1 FILLER_46_347 ();
 sg13g2_decap_4 FILLER_46_358 ();
 sg13g2_fill_2 FILLER_46_362 ();
 sg13g2_decap_8 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_418 ();
 sg13g2_decap_4 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_68 ();
 sg13g2_decap_8 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_82 ();
 sg13g2_decap_8 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_decap_4 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_decap_8 FILLER_47_202 ();
 sg13g2_decap_8 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_216 ();
 sg13g2_fill_1 FILLER_47_218 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_4 FILLER_47_287 ();
 sg13g2_fill_2 FILLER_47_291 ();
 sg13g2_decap_4 FILLER_47_313 ();
 sg13g2_fill_1 FILLER_47_317 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_fill_1 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_369 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_8 FILLER_47_404 ();
 sg13g2_decap_8 FILLER_47_411 ();
 sg13g2_decap_8 FILLER_47_418 ();
 sg13g2_decap_4 FILLER_47_425 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_39 ();
 sg13g2_fill_1 FILLER_48_57 ();
 sg13g2_decap_4 FILLER_48_62 ();
 sg13g2_fill_1 FILLER_48_66 ();
 sg13g2_decap_4 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_125 ();
 sg13g2_decap_4 FILLER_48_131 ();
 sg13g2_decap_4 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_143 ();
 sg13g2_fill_2 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_197 ();
 sg13g2_decap_8 FILLER_48_204 ();
 sg13g2_decap_4 FILLER_48_211 ();
 sg13g2_decap_8 FILLER_48_220 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_decap_8 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_246 ();
 sg13g2_decap_4 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_303 ();
 sg13g2_decap_8 FILLER_48_310 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_decap_8 FILLER_48_338 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_8 FILLER_48_403 ();
 sg13g2_decap_8 FILLER_48_410 ();
 sg13g2_decap_8 FILLER_48_417 ();
 sg13g2_decap_4 FILLER_48_424 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_70 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_96 ();
 sg13g2_decap_8 FILLER_49_103 ();
 sg13g2_decap_8 FILLER_49_110 ();
 sg13g2_decap_8 FILLER_49_117 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_fill_1 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_fill_2 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_225 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_246 ();
 sg13g2_decap_4 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_257 ();
 sg13g2_decap_8 FILLER_49_278 ();
 sg13g2_decap_8 FILLER_49_285 ();
 sg13g2_decap_4 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_296 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_4 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_decap_8 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_330 ();
 sg13g2_decap_4 FILLER_49_337 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_359 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_decap_8 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_421 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_48 ();
 sg13g2_decap_4 FILLER_50_55 ();
 sg13g2_fill_2 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_decap_8 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_99 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_decap_8 FILLER_50_127 ();
 sg13g2_decap_8 FILLER_50_134 ();
 sg13g2_decap_8 FILLER_50_145 ();
 sg13g2_fill_2 FILLER_50_152 ();
 sg13g2_fill_1 FILLER_50_154 ();
 sg13g2_fill_1 FILLER_50_175 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_decap_4 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_212 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_223 ();
 sg13g2_fill_2 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_247 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_fill_2 FILLER_50_264 ();
 sg13g2_fill_1 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_344 ();
 sg13g2_fill_2 FILLER_50_350 ();
 sg13g2_fill_1 FILLER_50_352 ();
 sg13g2_decap_8 FILLER_50_365 ();
 sg13g2_decap_8 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_decap_8 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_decap_8 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_50_414 ();
 sg13g2_decap_8 FILLER_50_421 ();
 sg13g2_fill_2 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_32 ();
 sg13g2_decap_8 FILLER_51_71 ();
 sg13g2_decap_4 FILLER_51_78 ();
 sg13g2_fill_2 FILLER_51_82 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_129 ();
 sg13g2_decap_8 FILLER_51_146 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_fill_2 FILLER_51_172 ();
 sg13g2_fill_1 FILLER_51_174 ();
 sg13g2_fill_2 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_197 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_decap_4 FILLER_51_248 ();
 sg13g2_fill_2 FILLER_51_252 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_decap_4 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_290 ();
 sg13g2_fill_2 FILLER_51_296 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_fill_1 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_367 ();
 sg13g2_decap_8 FILLER_51_374 ();
 sg13g2_decap_8 FILLER_51_381 ();
 sg13g2_decap_8 FILLER_51_388 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_decap_8 FILLER_51_416 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_4 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_51 ();
 sg13g2_fill_2 FILLER_52_58 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_85 ();
 sg13g2_decap_8 FILLER_52_92 ();
 sg13g2_decap_4 FILLER_52_99 ();
 sg13g2_fill_2 FILLER_52_103 ();
 sg13g2_decap_4 FILLER_52_110 ();
 sg13g2_fill_1 FILLER_52_114 ();
 sg13g2_decap_4 FILLER_52_129 ();
 sg13g2_fill_2 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_189 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_236 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_281 ();
 sg13g2_fill_2 FILLER_52_287 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_decap_4 FILLER_52_318 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_332 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_8 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_52_412 ();
 sg13g2_decap_8 FILLER_52_419 ();
 sg13g2_decap_4 FILLER_52_426 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_104 ();
 sg13g2_fill_1 FILLER_53_106 ();
 sg13g2_decap_8 FILLER_53_134 ();
 sg13g2_decap_4 FILLER_53_141 ();
 sg13g2_decap_8 FILLER_53_169 ();
 sg13g2_decap_8 FILLER_53_176 ();
 sg13g2_fill_1 FILLER_53_183 ();
 sg13g2_decap_4 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_fill_2 FILLER_53_258 ();
 sg13g2_decap_4 FILLER_53_268 ();
 sg13g2_fill_2 FILLER_53_272 ();
 sg13g2_decap_8 FILLER_53_279 ();
 sg13g2_decap_8 FILLER_53_286 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_304 ();
 sg13g2_decap_4 FILLER_53_349 ();
 sg13g2_decap_8 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_366 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_decap_8 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_53_415 ();
 sg13g2_decap_8 FILLER_53_422 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_75 ();
 sg13g2_decap_4 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_2 FILLER_54_122 ();
 sg13g2_fill_1 FILLER_54_124 ();
 sg13g2_fill_2 FILLER_54_130 ();
 sg13g2_fill_1 FILLER_54_132 ();
 sg13g2_fill_2 FILLER_54_138 ();
 sg13g2_fill_2 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_169 ();
 sg13g2_decap_8 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_181 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_decap_8 FILLER_54_236 ();
 sg13g2_decap_8 FILLER_54_243 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_255 ();
 sg13g2_fill_1 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_273 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_284 ();
 sg13g2_fill_1 FILLER_54_302 ();
 sg13g2_decap_4 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_2 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_decap_8 FILLER_54_353 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_374 ();
 sg13g2_decap_8 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_54_409 ();
 sg13g2_decap_8 FILLER_54_416 ();
 sg13g2_decap_8 FILLER_54_423 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_67 ();
 sg13g2_decap_8 FILLER_55_94 ();
 sg13g2_decap_4 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_117 ();
 sg13g2_fill_1 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_fill_1 FILLER_55_177 ();
 sg13g2_decap_4 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_239 ();
 sg13g2_fill_1 FILLER_55_241 ();
 sg13g2_decap_8 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_fill_1 FILLER_55_256 ();
 sg13g2_fill_1 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_274 ();
 sg13g2_decap_4 FILLER_55_281 ();
 sg13g2_decap_8 FILLER_55_289 ();
 sg13g2_decap_4 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_300 ();
 sg13g2_decap_4 FILLER_55_306 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_323 ();
 sg13g2_fill_2 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_338 ();
 sg13g2_decap_8 FILLER_55_344 ();
 sg13g2_decap_8 FILLER_55_351 ();
 sg13g2_decap_8 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_decap_8 FILLER_55_372 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_55_414 ();
 sg13g2_decap_8 FILLER_55_421 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_4 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_46 ();
 sg13g2_fill_2 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_78 ();
 sg13g2_fill_1 FILLER_56_87 ();
 sg13g2_decap_8 FILLER_56_93 ();
 sg13g2_decap_8 FILLER_56_100 ();
 sg13g2_decap_4 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_111 ();
 sg13g2_fill_2 FILLER_56_120 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_132 ();
 sg13g2_decap_4 FILLER_56_137 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_decap_4 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_178 ();
 sg13g2_fill_1 FILLER_56_183 ();
 sg13g2_fill_2 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_198 ();
 sg13g2_decap_4 FILLER_56_216 ();
 sg13g2_decap_4 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_268 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_fill_2 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_309 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_fill_1 FILLER_56_317 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_345 ();
 sg13g2_fill_1 FILLER_56_347 ();
 sg13g2_decap_8 FILLER_56_353 ();
 sg13g2_decap_8 FILLER_56_360 ();
 sg13g2_decap_8 FILLER_56_367 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_56_409 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_4 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_46 ();
 sg13g2_fill_2 FILLER_57_68 ();
 sg13g2_fill_1 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_92 ();
 sg13g2_decap_8 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_fill_1 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_decap_8 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_143 ();
 sg13g2_fill_1 FILLER_57_145 ();
 sg13g2_decap_4 FILLER_57_150 ();
 sg13g2_fill_2 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_177 ();
 sg13g2_decap_8 FILLER_57_184 ();
 sg13g2_decap_8 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_decap_4 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_221 ();
 sg13g2_decap_4 FILLER_57_232 ();
 sg13g2_fill_1 FILLER_57_236 ();
 sg13g2_decap_4 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_249 ();
 sg13g2_decap_8 FILLER_57_261 ();
 sg13g2_decap_4 FILLER_57_268 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_299 ();
 sg13g2_decap_8 FILLER_57_324 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_1 FILLER_57_345 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_fill_2 FILLER_57_427 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_50 ();
 sg13g2_fill_1 FILLER_58_57 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_132 ();
 sg13g2_decap_8 FILLER_58_171 ();
 sg13g2_decap_8 FILLER_58_178 ();
 sg13g2_decap_8 FILLER_58_185 ();
 sg13g2_decap_4 FILLER_58_192 ();
 sg13g2_fill_2 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_fill_2 FILLER_58_224 ();
 sg13g2_decap_4 FILLER_58_246 ();
 sg13g2_fill_2 FILLER_58_250 ();
 sg13g2_decap_8 FILLER_58_268 ();
 sg13g2_decap_4 FILLER_58_280 ();
 sg13g2_fill_1 FILLER_58_284 ();
 sg13g2_fill_1 FILLER_58_289 ();
 sg13g2_decap_8 FILLER_58_310 ();
 sg13g2_decap_4 FILLER_58_321 ();
 sg13g2_fill_2 FILLER_58_325 ();
 sg13g2_fill_2 FILLER_58_331 ();
 sg13g2_decap_8 FILLER_58_340 ();
 sg13g2_decap_8 FILLER_58_347 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_361 ();
 sg13g2_decap_8 FILLER_58_368 ();
 sg13g2_decap_8 FILLER_58_375 ();
 sg13g2_decap_8 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_389 ();
 sg13g2_decap_8 FILLER_58_396 ();
 sg13g2_decap_8 FILLER_58_403 ();
 sg13g2_decap_8 FILLER_58_410 ();
 sg13g2_decap_8 FILLER_58_417 ();
 sg13g2_decap_4 FILLER_58_424 ();
 sg13g2_fill_2 FILLER_58_428 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_decap_4 FILLER_59_157 ();
 sg13g2_fill_2 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_fill_1 FILLER_59_173 ();
 sg13g2_fill_2 FILLER_59_179 ();
 sg13g2_decap_8 FILLER_59_185 ();
 sg13g2_decap_4 FILLER_59_192 ();
 sg13g2_fill_2 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_202 ();
 sg13g2_decap_8 FILLER_59_214 ();
 sg13g2_decap_8 FILLER_59_221 ();
 sg13g2_decap_8 FILLER_59_228 ();
 sg13g2_fill_2 FILLER_59_235 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_decap_8 FILLER_59_247 ();
 sg13g2_fill_2 FILLER_59_254 ();
 sg13g2_fill_1 FILLER_59_281 ();
 sg13g2_fill_1 FILLER_59_298 ();
 sg13g2_fill_1 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_333 ();
 sg13g2_fill_1 FILLER_59_344 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_8 FILLER_59_388 ();
 sg13g2_decap_8 FILLER_59_395 ();
 sg13g2_decap_8 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_409 ();
 sg13g2_decap_8 FILLER_59_416 ();
 sg13g2_decap_8 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_59 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_fill_2 FILLER_60_123 ();
 sg13g2_fill_1 FILLER_60_125 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_4 FILLER_60_159 ();
 sg13g2_fill_1 FILLER_60_163 ();
 sg13g2_fill_1 FILLER_60_180 ();
 sg13g2_fill_1 FILLER_60_197 ();
 sg13g2_decap_4 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_fill_2 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_328 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_375 ();
 sg13g2_decap_8 FILLER_60_382 ();
 sg13g2_decap_8 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_396 ();
 sg13g2_decap_8 FILLER_60_403 ();
 sg13g2_decap_8 FILLER_60_410 ();
 sg13g2_decap_8 FILLER_60_417 ();
 sg13g2_decap_4 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_4 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_46 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_4 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_85 ();
 sg13g2_decap_8 FILLER_61_107 ();
 sg13g2_decap_4 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_decap_8 FILLER_61_131 ();
 sg13g2_fill_2 FILLER_61_138 ();
 sg13g2_fill_1 FILLER_61_140 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_decap_4 FILLER_61_159 ();
 sg13g2_fill_2 FILLER_61_163 ();
 sg13g2_decap_8 FILLER_61_233 ();
 sg13g2_decap_8 FILLER_61_240 ();
 sg13g2_fill_1 FILLER_61_247 ();
 sg13g2_fill_2 FILLER_61_268 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_fill_2 FILLER_61_351 ();
 sg13g2_fill_1 FILLER_61_353 ();
 sg13g2_decap_8 FILLER_61_358 ();
 sg13g2_decap_8 FILLER_61_365 ();
 sg13g2_decap_8 FILLER_61_372 ();
 sg13g2_decap_8 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_393 ();
 sg13g2_decap_8 FILLER_61_400 ();
 sg13g2_decap_8 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_61_414 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_4 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_53 ();
 sg13g2_decap_4 FILLER_62_63 ();
 sg13g2_fill_2 FILLER_62_67 ();
 sg13g2_fill_2 FILLER_62_73 ();
 sg13g2_decap_4 FILLER_62_80 ();
 sg13g2_fill_2 FILLER_62_100 ();
 sg13g2_decap_4 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_116 ();
 sg13g2_fill_1 FILLER_62_118 ();
 sg13g2_fill_2 FILLER_62_142 ();
 sg13g2_fill_2 FILLER_62_164 ();
 sg13g2_fill_1 FILLER_62_179 ();
 sg13g2_fill_1 FILLER_62_185 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_2 FILLER_62_198 ();
 sg13g2_fill_2 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_206 ();
 sg13g2_fill_1 FILLER_62_217 ();
 sg13g2_fill_1 FILLER_62_227 ();
 sg13g2_decap_4 FILLER_62_241 ();
 sg13g2_fill_2 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_251 ();
 sg13g2_decap_8 FILLER_62_265 ();
 sg13g2_decap_8 FILLER_62_272 ();
 sg13g2_decap_8 FILLER_62_279 ();
 sg13g2_decap_8 FILLER_62_286 ();
 sg13g2_decap_8 FILLER_62_293 ();
 sg13g2_decap_8 FILLER_62_300 ();
 sg13g2_decap_8 FILLER_62_307 ();
 sg13g2_fill_2 FILLER_62_323 ();
 sg13g2_decap_8 FILLER_62_348 ();
 sg13g2_decap_8 FILLER_62_355 ();
 sg13g2_decap_8 FILLER_62_362 ();
 sg13g2_decap_8 FILLER_62_369 ();
 sg13g2_decap_8 FILLER_62_376 ();
 sg13g2_decap_8 FILLER_62_383 ();
 sg13g2_decap_8 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_decap_8 FILLER_62_404 ();
 sg13g2_decap_8 FILLER_62_411 ();
 sg13g2_decap_8 FILLER_62_418 ();
 sg13g2_decap_4 FILLER_62_425 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_4 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_decap_4 FILLER_63_90 ();
 sg13g2_fill_1 FILLER_63_94 ();
 sg13g2_decap_8 FILLER_63_99 ();
 sg13g2_decap_8 FILLER_63_106 ();
 sg13g2_fill_2 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_139 ();
 sg13g2_decap_8 FILLER_63_146 ();
 sg13g2_decap_8 FILLER_63_157 ();
 sg13g2_decap_8 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_185 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_1 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_222 ();
 sg13g2_fill_2 FILLER_63_232 ();
 sg13g2_fill_1 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_240 ();
 sg13g2_decap_4 FILLER_63_246 ();
 sg13g2_fill_2 FILLER_63_250 ();
 sg13g2_decap_8 FILLER_63_256 ();
 sg13g2_decap_8 FILLER_63_263 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_decap_4 FILLER_63_275 ();
 sg13g2_fill_1 FILLER_63_304 ();
 sg13g2_fill_2 FILLER_63_309 ();
 sg13g2_decap_4 FILLER_63_315 ();
 sg13g2_decap_4 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_341 ();
 sg13g2_decap_8 FILLER_63_348 ();
 sg13g2_decap_8 FILLER_63_355 ();
 sg13g2_decap_8 FILLER_63_362 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_383 ();
 sg13g2_decap_8 FILLER_63_390 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_decap_8 FILLER_63_404 ();
 sg13g2_decap_8 FILLER_63_411 ();
 sg13g2_decap_8 FILLER_63_418 ();
 sg13g2_decap_4 FILLER_63_425 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_fill_2 FILLER_64_70 ();
 sg13g2_fill_1 FILLER_64_72 ();
 sg13g2_decap_4 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_decap_4 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_123 ();
 sg13g2_fill_1 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_207 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_fill_2 FILLER_64_240 ();
 sg13g2_fill_1 FILLER_64_242 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_fill_2 FILLER_64_266 ();
 sg13g2_fill_1 FILLER_64_268 ();
 sg13g2_decap_4 FILLER_64_294 ();
 sg13g2_fill_2 FILLER_64_298 ();
 sg13g2_fill_1 FILLER_64_315 ();
 sg13g2_fill_2 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_347 ();
 sg13g2_decap_8 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_decap_8 FILLER_64_375 ();
 sg13g2_decap_8 FILLER_64_382 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_8 FILLER_64_403 ();
 sg13g2_decap_8 FILLER_64_410 ();
 sg13g2_decap_8 FILLER_64_417 ();
 sg13g2_decap_4 FILLER_64_424 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_1 FILLER_65_60 ();
 sg13g2_decap_4 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_102 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_147 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_decap_8 FILLER_65_190 ();
 sg13g2_decap_4 FILLER_65_201 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_215 ();
 sg13g2_decap_4 FILLER_65_222 ();
 sg13g2_fill_2 FILLER_65_226 ();
 sg13g2_fill_1 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_237 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_fill_2 FILLER_65_251 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_2 FILLER_65_270 ();
 sg13g2_fill_1 FILLER_65_272 ();
 sg13g2_decap_4 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_fill_2 FILLER_65_427 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_116 ();
 sg13g2_fill_1 FILLER_66_118 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_decap_4 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_147 ();
 sg13g2_decap_4 FILLER_66_195 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_fill_2 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_206 ();
 sg13g2_fill_1 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_276 ();
 sg13g2_decap_8 FILLER_66_282 ();
 sg13g2_decap_8 FILLER_66_289 ();
 sg13g2_fill_2 FILLER_66_296 ();
 sg13g2_decap_4 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_307 ();
 sg13g2_fill_2 FILLER_66_312 ();
 sg13g2_fill_1 FILLER_66_314 ();
 sg13g2_decap_4 FILLER_66_340 ();
 sg13g2_fill_1 FILLER_66_344 ();
 sg13g2_decap_8 FILLER_66_354 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_66_368 ();
 sg13g2_decap_8 FILLER_66_375 ();
 sg13g2_decap_8 FILLER_66_382 ();
 sg13g2_decap_8 FILLER_66_389 ();
 sg13g2_decap_8 FILLER_66_396 ();
 sg13g2_decap_8 FILLER_66_403 ();
 sg13g2_decap_8 FILLER_66_410 ();
 sg13g2_decap_8 FILLER_66_417 ();
 sg13g2_decap_4 FILLER_66_424 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_117 ();
 sg13g2_fill_1 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_fill_1 FILLER_67_140 ();
 sg13g2_fill_1 FILLER_67_161 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_decap_8 FILLER_67_213 ();
 sg13g2_decap_4 FILLER_67_220 ();
 sg13g2_fill_1 FILLER_67_224 ();
 sg13g2_fill_2 FILLER_67_257 ();
 sg13g2_fill_1 FILLER_67_271 ();
 sg13g2_decap_8 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_decap_8 FILLER_67_292 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_decap_4 FILLER_67_367 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_decap_8 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_422 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_107 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_fill_2 FILLER_68_119 ();
 sg13g2_decap_4 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_137 ();
 sg13g2_decap_4 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_148 ();
 sg13g2_decap_4 FILLER_68_154 ();
 sg13g2_fill_2 FILLER_68_158 ();
 sg13g2_decap_8 FILLER_68_172 ();
 sg13g2_fill_1 FILLER_68_183 ();
 sg13g2_fill_1 FILLER_68_192 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_199 ();
 sg13g2_decap_8 FILLER_68_208 ();
 sg13g2_decap_4 FILLER_68_215 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_decap_8 FILLER_68_244 ();
 sg13g2_decap_4 FILLER_68_251 ();
 sg13g2_decap_4 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_fill_2 FILLER_68_285 ();
 sg13g2_decap_4 FILLER_68_292 ();
 sg13g2_fill_2 FILLER_68_308 ();
 sg13g2_fill_2 FILLER_68_315 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_decap_8 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_8 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_68_412 ();
 sg13g2_decap_8 FILLER_68_419 ();
 sg13g2_decap_4 FILLER_68_426 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_161 ();
 sg13g2_fill_1 FILLER_69_174 ();
 sg13g2_decap_4 FILLER_69_189 ();
 sg13g2_fill_2 FILLER_69_193 ();
 sg13g2_fill_2 FILLER_69_199 ();
 sg13g2_fill_2 FILLER_69_206 ();
 sg13g2_decap_4 FILLER_69_213 ();
 sg13g2_fill_2 FILLER_69_217 ();
 sg13g2_fill_2 FILLER_69_223 ();
 sg13g2_decap_4 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_238 ();
 sg13g2_decap_4 FILLER_69_260 ();
 sg13g2_decap_4 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_312 ();
 sg13g2_decap_8 FILLER_69_319 ();
 sg13g2_decap_8 FILLER_69_326 ();
 sg13g2_decap_8 FILLER_69_333 ();
 sg13g2_decap_8 FILLER_69_340 ();
 sg13g2_decap_4 FILLER_69_347 ();
 sg13g2_decap_4 FILLER_69_360 ();
 sg13g2_fill_1 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_69_409 ();
 sg13g2_decap_8 FILLER_69_416 ();
 sg13g2_decap_8 FILLER_69_423 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_4 FILLER_70_105 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_2 FILLER_70_134 ();
 sg13g2_decap_8 FILLER_70_172 ();
 sg13g2_fill_1 FILLER_70_179 ();
 sg13g2_decap_4 FILLER_70_188 ();
 sg13g2_decap_8 FILLER_70_208 ();
 sg13g2_fill_2 FILLER_70_231 ();
 sg13g2_decap_4 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_257 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_decap_4 FILLER_70_276 ();
 sg13g2_fill_2 FILLER_70_280 ();
 sg13g2_decap_4 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_313 ();
 sg13g2_decap_8 FILLER_70_320 ();
 sg13g2_fill_2 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_338 ();
 sg13g2_decap_8 FILLER_70_354 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_70_412 ();
 sg13g2_decap_8 FILLER_70_419 ();
 sg13g2_decap_4 FILLER_70_426 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_fill_2 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_decap_8 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_142 ();
 sg13g2_fill_2 FILLER_71_148 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_1 FILLER_71_172 ();
 sg13g2_decap_8 FILLER_71_193 ();
 sg13g2_decap_4 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_204 ();
 sg13g2_fill_2 FILLER_71_225 ();
 sg13g2_fill_1 FILLER_71_227 ();
 sg13g2_decap_4 FILLER_71_237 ();
 sg13g2_fill_1 FILLER_71_277 ();
 sg13g2_fill_2 FILLER_71_282 ();
 sg13g2_decap_8 FILLER_71_289 ();
 sg13g2_decap_8 FILLER_71_296 ();
 sg13g2_decap_8 FILLER_71_307 ();
 sg13g2_decap_8 FILLER_71_314 ();
 sg13g2_decap_4 FILLER_71_321 ();
 sg13g2_fill_1 FILLER_71_325 ();
 sg13g2_decap_8 FILLER_71_335 ();
 sg13g2_decap_8 FILLER_71_342 ();
 sg13g2_decap_8 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_decap_8 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_71_414 ();
 sg13g2_decap_8 FILLER_71_421 ();
 sg13g2_fill_2 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_fill_2 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_179 ();
 sg13g2_decap_4 FILLER_72_211 ();
 sg13g2_fill_2 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_243 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_275 ();
 sg13g2_decap_8 FILLER_72_296 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_fill_2 FILLER_72_310 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_decap_8 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_365 ();
 sg13g2_fill_1 FILLER_72_367 ();
 sg13g2_decap_4 FILLER_72_377 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_decap_8 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_72_414 ();
 sg13g2_decap_8 FILLER_72_421 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_4 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_204 ();
 sg13g2_fill_1 FILLER_73_206 ();
 sg13g2_decap_8 FILLER_73_236 ();
 sg13g2_decap_8 FILLER_73_243 ();
 sg13g2_fill_2 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_260 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_322 ();
 sg13g2_fill_1 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_8 FILLER_73_404 ();
 sg13g2_decap_8 FILLER_73_411 ();
 sg13g2_decap_8 FILLER_73_418 ();
 sg13g2_decap_4 FILLER_73_425 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_4 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_165 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_decap_4 FILLER_74_235 ();
 sg13g2_fill_2 FILLER_74_248 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_decap_4 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_decap_4 FILLER_74_316 ();
 sg13g2_fill_2 FILLER_74_320 ();
 sg13g2_decap_8 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_4 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_74_410 ();
 sg13g2_decap_8 FILLER_74_417 ();
 sg13g2_decap_4 FILLER_74_424 ();
 sg13g2_fill_2 FILLER_74_428 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_4 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_148 ();
 sg13g2_decap_4 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_163 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_4 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_198 ();
 sg13g2_fill_2 FILLER_75_203 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_decap_8 FILLER_75_215 ();
 sg13g2_decap_8 FILLER_75_222 ();
 sg13g2_decap_8 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_1 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_282 ();
 sg13g2_decap_4 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_293 ();
 sg13g2_decap_8 FILLER_75_304 ();
 sg13g2_decap_8 FILLER_75_311 ();
 sg13g2_decap_8 FILLER_75_318 ();
 sg13g2_decap_8 FILLER_75_325 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_decap_8 FILLER_75_363 ();
 sg13g2_decap_8 FILLER_75_370 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_decap_4 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_8 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_75_412 ();
 sg13g2_decap_8 FILLER_75_419 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_fill_2 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_135 ();
 sg13g2_decap_4 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_164 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_189 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_decap_4 FILLER_76_208 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_4 FILLER_76_329 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_decap_8 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_351 ();
 sg13g2_decap_8 FILLER_76_358 ();
 sg13g2_decap_8 FILLER_76_365 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_decap_8 FILLER_76_416 ();
 sg13g2_decap_8 FILLER_76_423 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_4 FILLER_77_119 ();
 sg13g2_fill_2 FILLER_77_123 ();
 sg13g2_decap_4 FILLER_77_129 ();
 sg13g2_fill_2 FILLER_77_150 ();
 sg13g2_fill_1 FILLER_77_152 ();
 sg13g2_fill_1 FILLER_77_157 ();
 sg13g2_fill_2 FILLER_77_178 ();
 sg13g2_fill_1 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_198 ();
 sg13g2_fill_1 FILLER_77_202 ();
 sg13g2_fill_1 FILLER_77_219 ();
 sg13g2_fill_2 FILLER_77_224 ();
 sg13g2_fill_2 FILLER_77_233 ();
 sg13g2_fill_1 FILLER_77_235 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_259 ();
 sg13g2_fill_1 FILLER_77_261 ();
 sg13g2_decap_4 FILLER_77_280 ();
 sg13g2_fill_1 FILLER_77_284 ();
 sg13g2_decap_4 FILLER_77_294 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_327 ();
 sg13g2_fill_1 FILLER_77_329 ();
 sg13g2_fill_2 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_368 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_414 ();
 sg13g2_decap_8 FILLER_77_421 ();
 sg13g2_fill_2 FILLER_77_428 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_112 ();
 sg13g2_fill_1 FILLER_78_116 ();
 sg13g2_decap_8 FILLER_78_121 ();
 sg13g2_decap_8 FILLER_78_128 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_fill_1 FILLER_78_142 ();
 sg13g2_fill_2 FILLER_78_159 ();
 sg13g2_fill_1 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_207 ();
 sg13g2_fill_1 FILLER_78_225 ();
 sg13g2_fill_2 FILLER_78_242 ();
 sg13g2_fill_2 FILLER_78_253 ();
 sg13g2_fill_1 FILLER_78_255 ();
 sg13g2_fill_1 FILLER_78_265 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_fill_2 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_decap_8 FILLER_79_128 ();
 sg13g2_decap_8 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_142 ();
 sg13g2_fill_1 FILLER_79_144 ();
 sg13g2_decap_8 FILLER_79_149 ();
 sg13g2_fill_2 FILLER_79_156 ();
 sg13g2_decap_4 FILLER_79_162 ();
 sg13g2_fill_1 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_1 FILLER_79_226 ();
 sg13g2_fill_1 FILLER_79_242 ();
 sg13g2_fill_2 FILLER_79_247 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_2 FILLER_79_270 ();
 sg13g2_fill_1 FILLER_79_272 ();
 sg13g2_fill_1 FILLER_79_309 ();
 sg13g2_fill_1 FILLER_79_319 ();
 sg13g2_fill_1 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_339 ();
 sg13g2_decap_4 FILLER_79_346 ();
 sg13g2_fill_1 FILLER_79_350 ();
 sg13g2_fill_1 FILLER_79_360 ();
 sg13g2_fill_1 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_380 ();
 sg13g2_decap_4 FILLER_79_390 ();
 sg13g2_fill_2 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_414 ();
 sg13g2_decap_8 FILLER_79_421 ();
 sg13g2_fill_2 FILLER_79_428 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_74 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_1 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_89 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_fill_2 FILLER_80_103 ();
 sg13g2_fill_1 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_110 ();
 sg13g2_fill_1 FILLER_80_117 ();
 sg13g2_decap_4 FILLER_80_139 ();
 sg13g2_fill_2 FILLER_80_143 ();
 sg13g2_decap_8 FILLER_80_149 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_2 FILLER_80_173 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_4 FILLER_80_184 ();
 sg13g2_decap_4 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_4 FILLER_80_211 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_222 ();
 sg13g2_fill_2 FILLER_80_230 ();
 sg13g2_decap_4 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_244 ();
 sg13g2_fill_2 FILLER_80_249 ();
 sg13g2_fill_2 FILLER_80_255 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_275 ();
 sg13g2_decap_8 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_8 FILLER_80_324 ();
 sg13g2_decap_8 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_338 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_4 FILLER_80_352 ();
 sg13g2_fill_1 FILLER_80_368 ();
 sg13g2_decap_4 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_fill_2 FILLER_80_394 ();
 sg13g2_fill_1 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
