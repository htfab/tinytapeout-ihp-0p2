module tt_um_snow (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire clknet_0_clk;
 wire net56;
 wire \main._w_demo_video_hs ;
 wire \main._w_demo_video_vs ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[0] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[1] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[2] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[3] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[4] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[5] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[6] ;
 wire \main.demo._d___pip_24_1_1___stage___block_3_y[7] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[0] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[1] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[2] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[3] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[4] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[5] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[6] ;
 wire \main.demo._d___pip_24_1_2___stage___block_3_y[7] ;
 wire \main.demo._q___pip_24_1_2___stage___block_3_s[0] ;
 wire \main.demo._q___pip_24_1_2___stage___block_3_s[1] ;
 wire \main.demo._q_frame[0] ;
 wire \main.demo._q_frame[10] ;
 wire \main.demo._q_frame[11] ;
 wire \main.demo._q_frame[12] ;
 wire \main.demo._q_frame[13] ;
 wire \main.demo._q_frame[14] ;
 wire \main.demo._q_frame[15] ;
 wire \main.demo._q_frame[1] ;
 wire \main.demo._q_frame[2] ;
 wire \main.demo._q_frame[3] ;
 wire \main.demo._q_frame[4] ;
 wire \main.demo._q_frame[5] ;
 wire \main.demo._q_frame[6] ;
 wire \main.demo._q_frame[7] ;
 wire \main.demo._q_frame[8] ;
 wire \main.demo._q_frame[9] ;
 wire \main.demo._q_modulo_0[0] ;
 wire \main.demo._q_modulo_0[10] ;
 wire \main.demo._q_modulo_0[11] ;
 wire \main.demo._q_modulo_0[12] ;
 wire \main.demo._q_modulo_0[13] ;
 wire \main.demo._q_modulo_0[14] ;
 wire \main.demo._q_modulo_0[15] ;
 wire \main.demo._q_modulo_0[1] ;
 wire \main.demo._q_modulo_0[2] ;
 wire \main.demo._q_modulo_0[3] ;
 wire \main.demo._q_modulo_0[4] ;
 wire \main.demo._q_modulo_0[5] ;
 wire \main.demo._q_modulo_0[6] ;
 wire \main.demo._q_modulo_0[7] ;
 wire \main.demo._q_modulo_0[8] ;
 wire \main.demo._q_modulo_0[9] ;
 wire \main.demo._q_modulo_1[0] ;
 wire \main.demo._q_modulo_1[10] ;
 wire \main.demo._q_modulo_1[11] ;
 wire \main.demo._q_modulo_1[12] ;
 wire \main.demo._q_modulo_1[13] ;
 wire \main.demo._q_modulo_1[14] ;
 wire \main.demo._q_modulo_1[15] ;
 wire \main.demo._q_modulo_1[1] ;
 wire \main.demo._q_modulo_1[2] ;
 wire \main.demo._q_modulo_1[3] ;
 wire \main.demo._q_modulo_1[4] ;
 wire \main.demo._q_modulo_1[5] ;
 wire \main.demo._q_modulo_1[6] ;
 wire \main.demo._q_modulo_1[7] ;
 wire \main.demo._q_modulo_1[8] ;
 wire \main.demo._q_modulo_1[9] ;
 wire \main.demo._q_pix_x[0] ;
 wire \main.demo._q_pix_x[1] ;
 wire \main.demo._q_pix_x[2] ;
 wire \main.demo._q_pix_x[3] ;
 wire \main.demo._q_pix_x[4] ;
 wire \main.demo._q_pix_x[5] ;
 wire \main.demo._q_pix_x[6] ;
 wire \main.demo._q_pix_x[7] ;
 wire \main.demo._q_pix_x[8] ;
 wire \main.demo._q_pix_x[9] ;
 wire \main.demo._q_prev_hs ;
 wire \main.demo._q_prev_vs ;
 wire \main.demo._q_rand_0[0] ;
 wire \main.demo._q_rand_0[10] ;
 wire \main.demo._q_rand_0[11] ;
 wire \main.demo._q_rand_0[1] ;
 wire \main.demo._q_rand_0[2] ;
 wire \main.demo._q_rand_0[3] ;
 wire \main.demo._q_rand_0[4] ;
 wire \main.demo._q_rand_0[5] ;
 wire \main.demo._q_rand_0[6] ;
 wire \main.demo._q_rand_0[7] ;
 wire \main.demo._q_rand_0[8] ;
 wire \main.demo._q_rand_0[9] ;
 wire \main.demo._q_rand_1[0] ;
 wire \main.demo._q_rand_1[10] ;
 wire \main.demo._q_rand_1[11] ;
 wire \main.demo._q_rand_1[1] ;
 wire \main.demo._q_rand_1[2] ;
 wire \main.demo._q_rand_1[3] ;
 wire \main.demo._q_rand_1[4] ;
 wire \main.demo._q_rand_1[5] ;
 wire \main.demo._q_rand_1[6] ;
 wire \main.demo._q_rand_1[7] ;
 wire \main.demo._q_rand_1[8] ;
 wire \main.demo._q_rand_1[9] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[0] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[1] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[2] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[3] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[4] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[5] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[6] ;
 wire \main.demo._t___pip_24_1_0___stage___block_3_y[7] ;
 wire \main.demo._w_vga_active ;
 wire \main.demo.vga._d_active ;
 wire \main.demo.vga._d_vblank ;
 wire \main.demo.vga._q_active_h ;
 wire \main.demo.vga._q_active_v ;
 wire \main.demo.vga._q_xcount[0] ;
 wire \main.demo.vga._q_xcount[10] ;
 wire \main.demo.vga._q_xcount[1] ;
 wire \main.demo.vga._q_xcount[2] ;
 wire \main.demo.vga._q_xcount[3] ;
 wire \main.demo.vga._q_xcount[4] ;
 wire \main.demo.vga._q_xcount[5] ;
 wire \main.demo.vga._q_xcount[6] ;
 wire \main.demo.vga._q_xcount[7] ;
 wire \main.demo.vga._q_xcount[8] ;
 wire \main.demo.vga._q_xcount[9] ;
 wire \main.demo.vga._q_ycount[0] ;
 wire \main.demo.vga._q_ycount[1] ;
 wire \main.demo.vga._q_ycount[2] ;
 wire \main.demo.vga._q_ycount[3] ;
 wire \main.demo.vga._q_ycount[4] ;
 wire \main.demo.vga._q_ycount[5] ;
 wire \main.demo.vga._q_ycount[6] ;
 wire \main.demo.vga._q_ycount[7] ;
 wire \main.demo.vga._q_ycount[8] ;
 wire rst_n_q;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_o21ai_1 _1995_ (.B1(_0006_),
    .Y(_0988_),
    .A1(\main.demo._q_modulo_0[5] ),
    .A2(_0969_));
 sg13g2_inv_1 _1996_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_o21ai_1 _1997_ (.B1(_0974_),
    .Y(_0990_),
    .A1(_0987_),
    .A2(_0989_));
 sg13g2_nand2_1 _1998_ (.Y(_0991_),
    .A(_1434_),
    .B(\main.demo._q_modulo_0[13] ));
 sg13g2_nor3_1 _1999_ (.A(_1443_),
    .B(_0980_),
    .C(_0991_),
    .Y(_0992_));
 sg13g2_nand2_1 _2000_ (.Y(_0993_),
    .A(_0990_),
    .B(_0992_));
 sg13g2_nor3_1 _2001_ (.A(_1423_),
    .B(_0993_),
    .C(net20),
    .Y(_0994_));
 sg13g2_inv_1 _2002_ (.Y(_0995_),
    .A(net20));
 sg13g2_inv_1 _2003_ (.Y(_0996_),
    .A(_0993_));
 sg13g2_a21oi_1 _2004_ (.A1(_0995_),
    .A2(_0996_),
    .Y(_0997_),
    .B1(\main.demo._q_modulo_0[14] ));
 sg13g2_nor3_1 _2005_ (.A(net22),
    .B(_0994_),
    .C(_0997_),
    .Y(_0043_));
 sg13g2_nor3_1 _2006_ (.A(_1429_),
    .B(_1423_),
    .C(_0984_),
    .Y(_0998_));
 sg13g2_o21ai_1 _2007_ (.B1(net33),
    .Y(_0999_),
    .A1(\main.demo._q_modulo_0[15] ),
    .A2(_0998_));
 sg13g2_a21oi_1 _2008_ (.A1(\main.demo._q_modulo_0[15] ),
    .A2(_0998_),
    .Y(_0044_),
    .B1(_0999_));
 sg13g2_a21oi_1 _2009_ (.A1(_0995_),
    .A2(_1491_),
    .Y(_1000_),
    .B1(_1487_));
 sg13g2_and3_1 _2010_ (.X(_1001_),
    .A(_0995_),
    .B(_1491_),
    .C(_1487_));
 sg13g2_nor3_1 _2011_ (.A(net22),
    .B(_1000_),
    .C(_1001_),
    .Y(_0045_));
 sg13g2_nor2_1 _2012_ (.A(\main.demo._q_modulo_0[2] ),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nor2b_1 _2013_ (.A(_1500_),
    .B_N(_1001_),
    .Y(_1003_));
 sg13g2_nor3_1 _2014_ (.A(net22),
    .B(_1002_),
    .C(_1003_),
    .Y(_0046_));
 sg13g2_nor2_1 _2015_ (.A(_0967_),
    .B(net20),
    .Y(_1004_));
 sg13g2_nor2_1 _2016_ (.A(\main.demo._q_modulo_0[3] ),
    .B(_1003_),
    .Y(_1005_));
 sg13g2_nor3_1 _2017_ (.A(_0982_),
    .B(_1004_),
    .C(_1005_),
    .Y(_0047_));
 sg13g2_inv_1 _2018_ (.Y(_1006_),
    .A(_1004_));
 sg13g2_o21ai_1 _2019_ (.B1(net33),
    .Y(_1007_),
    .A1(_1465_),
    .A2(_1006_));
 sg13g2_a21oi_1 _2020_ (.A1(_1465_),
    .A2(_1006_),
    .Y(_0048_),
    .B1(_1007_));
 sg13g2_xor2_1 _2021_ (.B(_0968_),
    .A(_0006_),
    .X(_1008_));
 sg13g2_o21ai_1 _2022_ (.B1(net34),
    .Y(_1009_),
    .A1(_1008_),
    .A2(net20));
 sg13g2_a21oi_1 _2023_ (.A1(_1478_),
    .A2(net20),
    .Y(_0049_),
    .B1(_1009_));
 sg13g2_nor3_1 _2024_ (.A(_0970_),
    .B(_0989_),
    .C(net20),
    .Y(_1010_));
 sg13g2_a21oi_1 _2025_ (.A1(_0995_),
    .A2(_0988_),
    .Y(_1011_),
    .B1(_1482_));
 sg13g2_nor3_1 _2026_ (.A(net22),
    .B(_1010_),
    .C(_1011_),
    .Y(_0050_));
 sg13g2_inv_1 _2027_ (.Y(_1012_),
    .A(_1461_));
 sg13g2_nand2_1 _2028_ (.Y(_1013_),
    .A(_0995_),
    .B(_0971_));
 sg13g2_o21ai_1 _2029_ (.B1(net34),
    .Y(_1014_),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_a21oi_1 _2030_ (.A1(_1012_),
    .A2(_1013_),
    .Y(_0051_),
    .B1(_1014_));
 sg13g2_o21ai_1 _2031_ (.B1(\main.demo._q_modulo_0[8] ),
    .Y(_1015_),
    .A1(_0973_),
    .A2(net20));
 sg13g2_nand3_1 _2032_ (.B(_1457_),
    .C(_0972_),
    .A(_0995_),
    .Y(_1016_));
 sg13g2_buf_1 _2033_ (.A(net31),
    .X(_1017_));
 sg13g2_a21oi_1 _2034_ (.A1(_1015_),
    .A2(_1016_),
    .Y(_0052_),
    .B1(net30));
 sg13g2_o21ai_1 _2035_ (.B1(net34),
    .Y(_1018_),
    .A1(_1449_),
    .A2(_1016_));
 sg13g2_a21oi_1 _2036_ (.A1(_1449_),
    .A2(_1016_),
    .Y(_0053_),
    .B1(_1018_));
 sg13g2_inv_1 _2037_ (.Y(_1019_),
    .A(\main.demo._q_modulo_1[0] ));
 sg13g2_and3_1 _2038_ (.X(_1020_),
    .A(_0463_),
    .B(_0464_),
    .C(_0490_));
 sg13g2_nor4_1 _2039_ (.A(_0479_),
    .B(_0477_),
    .C(_0482_),
    .D(_0487_),
    .Y(_1021_));
 sg13g2_nand2_1 _2040_ (.Y(_1022_),
    .A(_0374_),
    .B(_0466_));
 sg13g2_nor3_1 _2041_ (.A(_0471_),
    .B(_1022_),
    .C(_0474_),
    .Y(_1023_));
 sg13g2_and4_1 _2042_ (.A(_0453_),
    .B(_1020_),
    .C(_1021_),
    .D(_1023_),
    .X(_1024_));
 sg13g2_nor3_1 _2043_ (.A(_0447_),
    .B(_0416_),
    .C(_0440_),
    .Y(_1025_));
 sg13g2_nand3_1 _2044_ (.B(_0430_),
    .C(_1025_),
    .A(_0459_),
    .Y(_1026_));
 sg13g2_inv_1 _2045_ (.Y(_1027_),
    .A(_0447_));
 sg13g2_nand3_1 _2046_ (.B(_1027_),
    .C(_0415_),
    .A(_0419_),
    .Y(_1028_));
 sg13g2_o21ai_1 _2047_ (.B1(_1028_),
    .Y(_1029_),
    .A1(_0447_),
    .A2(_0449_));
 sg13g2_a21oi_1 _2048_ (.A1(_0438_),
    .A2(_1025_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_nand2_1 _2049_ (.Y(_1031_),
    .A(_1026_),
    .B(_1030_));
 sg13g2_nand3_1 _2050_ (.B(_0906_),
    .C(_1031_),
    .A(_1024_),
    .Y(_1032_));
 sg13g2_buf_1 _2051_ (.A(_1032_),
    .X(_1033_));
 sg13g2_buf_1 _2052_ (.A(_1033_),
    .X(_1034_));
 sg13g2_o21ai_1 _2053_ (.B1(net34),
    .Y(_1035_),
    .A1(_0016_),
    .A2(net19));
 sg13g2_a21oi_1 _2054_ (.A1(_1019_),
    .A2(net19),
    .Y(_0054_),
    .B1(_1035_));
 sg13g2_inv_1 _2055_ (.Y(_1036_),
    .A(\main.demo._q_modulo_1[1] ));
 sg13g2_nor4_1 _2056_ (.A(_1019_),
    .B(_1036_),
    .C(_0380_),
    .D(_0389_),
    .Y(_1037_));
 sg13g2_inv_1 _2057_ (.Y(_1038_),
    .A(_1037_));
 sg13g2_nor2_1 _2058_ (.A(_0384_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_inv_1 _2059_ (.Y(_1040_),
    .A(_1039_));
 sg13g2_nand2_1 _2060_ (.Y(_1041_),
    .A(\main.demo._q_modulo_1[6] ),
    .B(\main.demo._q_modulo_1[7] ));
 sg13g2_a21oi_1 _2061_ (.A1(_1040_),
    .A2(_0399_),
    .Y(_1042_),
    .B1(_1041_));
 sg13g2_nor2_1 _2062_ (.A(_0338_),
    .B(\main.demo._q_modulo_1[9] ),
    .Y(_1043_));
 sg13g2_nor2b_1 _2063_ (.A(_1042_),
    .B_N(_1043_),
    .Y(_1044_));
 sg13g2_nand3b_1 _2064_ (.B(_1027_),
    .C(_0906_),
    .Y(_1045_),
    .A_N(_0414_));
 sg13g2_or4_1 _2065_ (.A(_0474_),
    .B(_0471_),
    .C(_1022_),
    .D(_1045_),
    .X(_1046_));
 sg13g2_nor4_1 _2066_ (.A(_0479_),
    .B(_0477_),
    .C(_0482_),
    .D(_1046_),
    .Y(_1047_));
 sg13g2_inv_1 _2067_ (.Y(_1048_),
    .A(_0487_));
 sg13g2_and4_1 _2068_ (.A(_0464_),
    .B(_1047_),
    .C(_1048_),
    .D(_0490_),
    .X(_1049_));
 sg13g2_nor2_1 _2069_ (.A(_0419_),
    .B(_0441_),
    .Y(_1050_));
 sg13g2_nand2_1 _2070_ (.Y(_1051_),
    .A(_1050_),
    .B(_0449_));
 sg13g2_nand4_1 _2071_ (.B(_1049_),
    .C(_0463_),
    .A(_0453_),
    .Y(_1052_),
    .D(_1051_));
 sg13g2_buf_1 _2072_ (.A(_1052_),
    .X(_1053_));
 sg13g2_nor2_1 _2073_ (.A(_1044_),
    .B(_1053_),
    .Y(_1054_));
 sg13g2_o21ai_1 _2074_ (.B1(net33),
    .Y(_1055_),
    .A1(\main.demo._q_modulo_1[10] ),
    .A2(_1054_));
 sg13g2_nor3_1 _2075_ (.A(_0352_),
    .B(_1044_),
    .C(_1033_),
    .Y(_1056_));
 sg13g2_nor2_1 _2076_ (.A(_1055_),
    .B(_1056_),
    .Y(_0055_));
 sg13g2_nor4_2 _2077_ (.A(_0352_),
    .B(_0367_),
    .C(_1044_),
    .Y(_1057_),
    .D(_1053_));
 sg13g2_nor2_1 _2078_ (.A(\main.demo._q_modulo_1[11] ),
    .B(_1056_),
    .Y(_1058_));
 sg13g2_nor3_1 _2079_ (.A(net22),
    .B(_1057_),
    .C(_1058_),
    .Y(_0056_));
 sg13g2_nor2_1 _2080_ (.A(_0360_),
    .B(_1057_),
    .Y(_1059_));
 sg13g2_and3_1 _2081_ (.X(_1060_),
    .A(_1056_),
    .B(\main.demo._q_modulo_1[11] ),
    .C(_0360_));
 sg13g2_buf_1 _2082_ (.A(_1060_),
    .X(_1061_));
 sg13g2_nor3_1 _2083_ (.A(net22),
    .B(_1059_),
    .C(_1061_),
    .Y(_0057_));
 sg13g2_o21ai_1 _2084_ (.B1(net34),
    .Y(_1062_),
    .A1(_0330_),
    .A2(_1061_));
 sg13g2_a21oi_1 _2085_ (.A1(_0330_),
    .A2(_1061_),
    .Y(_0058_),
    .B1(_1062_));
 sg13g2_o21ai_1 _2086_ (.B1(_0005_),
    .Y(_1063_),
    .A1(\main.demo._q_modulo_1[5] ),
    .A2(_1040_));
 sg13g2_inv_1 _2087_ (.Y(_1064_),
    .A(_1063_));
 sg13g2_o21ai_1 _2088_ (.B1(_1043_),
    .Y(_1065_),
    .A1(_1041_),
    .A2(_1064_));
 sg13g2_nand2_1 _2089_ (.Y(_1066_),
    .A(_0360_),
    .B(_0330_));
 sg13g2_nor3_1 _2090_ (.A(_0352_),
    .B(_0367_),
    .C(_1066_),
    .Y(_1067_));
 sg13g2_nand2_1 _2091_ (.Y(_1068_),
    .A(_1065_),
    .B(_1067_));
 sg13g2_nor3_1 _2092_ (.A(_0413_),
    .B(_1068_),
    .C(net19),
    .Y(_1069_));
 sg13g2_inv_1 _2093_ (.Y(_1070_),
    .A(net19));
 sg13g2_inv_1 _2094_ (.Y(_1071_),
    .A(_1068_));
 sg13g2_a21oi_1 _2095_ (.A1(_1070_),
    .A2(_1071_),
    .Y(_1072_),
    .B1(\main.demo._q_modulo_1[14] ));
 sg13g2_nor3_1 _2096_ (.A(net22),
    .B(_1069_),
    .C(_1072_),
    .Y(_0059_));
 sg13g2_nand4_1 _2097_ (.B(_0360_),
    .C(_0330_),
    .A(_1057_),
    .Y(_1073_),
    .D(\main.demo._q_modulo_1[14] ));
 sg13g2_a21oi_1 _2098_ (.A1(_1073_),
    .A2(_1027_),
    .Y(_0060_),
    .B1(net30));
 sg13g2_nor3_1 _2099_ (.A(_1019_),
    .B(_1036_),
    .C(net19),
    .Y(_1074_));
 sg13g2_a21oi_1 _2100_ (.A1(_1070_),
    .A2(\main.demo._q_modulo_1[0] ),
    .Y(_1075_),
    .B1(\main.demo._q_modulo_1[1] ));
 sg13g2_nor3_1 _2101_ (.A(_0982_),
    .B(_1074_),
    .C(_1075_),
    .Y(_0061_));
 sg13g2_buf_1 _2102_ (.A(net31),
    .X(_1076_));
 sg13g2_nor2_1 _2103_ (.A(\main.demo._q_modulo_1[2] ),
    .B(_1074_),
    .Y(_1077_));
 sg13g2_nor2b_1 _2104_ (.A(_0380_),
    .B_N(_1074_),
    .Y(_1078_));
 sg13g2_nor3_1 _2105_ (.A(_1076_),
    .B(_1077_),
    .C(_1078_),
    .Y(_0062_));
 sg13g2_nor2_1 _2106_ (.A(_1038_),
    .B(net19),
    .Y(_1079_));
 sg13g2_nor2_1 _2107_ (.A(\main.demo._q_modulo_1[3] ),
    .B(_1078_),
    .Y(_1080_));
 sg13g2_nor3_1 _2108_ (.A(net29),
    .B(_1079_),
    .C(_1080_),
    .Y(_0063_));
 sg13g2_inv_1 _2109_ (.Y(_1081_),
    .A(_1079_));
 sg13g2_o21ai_1 _2110_ (.B1(net34),
    .Y(_1082_),
    .A1(_0384_),
    .A2(_1081_));
 sg13g2_a21oi_1 _2111_ (.A1(_0384_),
    .A2(_1081_),
    .Y(_0064_),
    .B1(_1082_));
 sg13g2_xor2_1 _2112_ (.B(_1039_),
    .A(_0005_),
    .X(_1083_));
 sg13g2_o21ai_1 _2113_ (.B1(_0907_),
    .Y(_1084_),
    .A1(_1083_),
    .A2(net19));
 sg13g2_a21oi_1 _2114_ (.A1(_0399_),
    .A2(_1034_),
    .Y(_0065_),
    .B1(_1084_));
 sg13g2_nor3_1 _2115_ (.A(_0333_),
    .B(_1064_),
    .C(_1034_),
    .Y(_1085_));
 sg13g2_a21oi_1 _2116_ (.A1(_1070_),
    .A2(_1063_),
    .Y(_1086_),
    .B1(\main.demo._q_modulo_1[6] ));
 sg13g2_nor3_1 _2117_ (.A(_1076_),
    .B(_1085_),
    .C(_1086_),
    .Y(_0066_));
 sg13g2_nor2b_1 _2118_ (.A(_1053_),
    .B_N(_1042_),
    .Y(_1087_));
 sg13g2_a21oi_1 _2119_ (.A1(_1040_),
    .A2(_0399_),
    .Y(_1088_),
    .B1(_0333_));
 sg13g2_a21oi_1 _2120_ (.A1(_1070_),
    .A2(_1088_),
    .Y(_1089_),
    .B1(\main.demo._q_modulo_1[7] ));
 sg13g2_nor3_1 _2121_ (.A(net29),
    .B(_1087_),
    .C(_1089_),
    .Y(_0067_));
 sg13g2_nor2_1 _2122_ (.A(_1042_),
    .B(net19),
    .Y(_1090_));
 sg13g2_o21ai_1 _2123_ (.B1(net34),
    .Y(_1091_),
    .A1(_0338_),
    .A2(_1090_));
 sg13g2_a21oi_1 _2124_ (.A1(_0338_),
    .A2(_1090_),
    .Y(_0068_),
    .B1(_1091_));
 sg13g2_nor3_1 _2125_ (.A(_0338_),
    .B(_1042_),
    .C(_1053_),
    .Y(_1092_));
 sg13g2_nor2_1 _2126_ (.A(\main.demo._q_modulo_1[9] ),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_nor2b_1 _2127_ (.A(_0356_),
    .B_N(_1092_),
    .Y(_1094_));
 sg13g2_nor3_1 _2128_ (.A(net29),
    .B(_1093_),
    .C(_1094_),
    .Y(_0069_));
 sg13g2_nor3_1 _2129_ (.A(\main.demo._q_pix_x[0] ),
    .B(net24),
    .C(_1576_),
    .Y(_0070_));
 sg13g2_buf_1 _2130_ (.A(net31),
    .X(_1095_));
 sg13g2_nor2_1 _2131_ (.A(net28),
    .B(_1591_),
    .Y(_0071_));
 sg13g2_nor2_1 _2132_ (.A(net28),
    .B(_1595_),
    .Y(_0072_));
 sg13g2_nor2_1 _2133_ (.A(_1095_),
    .B(_0473_),
    .Y(_0073_));
 sg13g2_nor2b_1 _2134_ (.A(net28),
    .B_N(_1631_),
    .Y(_0074_));
 sg13g2_nor2_1 _2135_ (.A(net28),
    .B(_1628_),
    .Y(_0075_));
 sg13g2_nor2_1 _2136_ (.A(net28),
    .B(_1619_),
    .Y(_0076_));
 sg13g2_nor2_1 _2137_ (.A(net28),
    .B(_1615_),
    .Y(_0077_));
 sg13g2_nor2_1 _2138_ (.A(net28),
    .B(_1639_),
    .Y(_0078_));
 sg13g2_nor2_1 _2139_ (.A(net28),
    .B(_1642_),
    .Y(_0079_));
 sg13g2_nand2_1 _2140_ (.Y(_1096_),
    .A(\main._w_demo_video_hs ),
    .B(_0908_));
 sg13g2_inv_1 _2141_ (.Y(_0080_),
    .A(_1096_));
 sg13g2_nand2_1 _2142_ (.Y(_1097_),
    .A(\main._w_demo_video_vs ),
    .B(_0908_));
 sg13g2_inv_1 _2143_ (.Y(_0081_),
    .A(_1097_));
 sg13g2_buf_1 _2144_ (.A(net31),
    .X(_1098_));
 sg13g2_nor2_1 _2145_ (.A(net27),
    .B(_1743_),
    .Y(_0082_));
 sg13g2_nor2_1 _2146_ (.A(_1098_),
    .B(_1650_),
    .Y(_0083_));
 sg13g2_nor2_1 _2147_ (.A(net27),
    .B(net11),
    .Y(_0084_));
 sg13g2_nor2_1 _2148_ (.A(net27),
    .B(_1737_),
    .Y(_0085_));
 sg13g2_nor2_1 _2149_ (.A(net27),
    .B(_1727_),
    .Y(_0086_));
 sg13g2_nor2_1 _2150_ (.A(net27),
    .B(_1704_),
    .Y(_0087_));
 sg13g2_nor2_1 _2151_ (.A(net27),
    .B(_1797_),
    .Y(_0088_));
 sg13g2_nor2_1 _2152_ (.A(_1098_),
    .B(_1806_),
    .Y(_0089_));
 sg13g2_nor2_1 _2153_ (.A(net27),
    .B(_1779_),
    .Y(_0090_));
 sg13g2_nor2_1 _2154_ (.A(net27),
    .B(_1829_),
    .Y(_0091_));
 sg13g2_buf_1 _2155_ (.A(_0911_),
    .X(_1099_));
 sg13g2_nor2_1 _2156_ (.A(net26),
    .B(_0825_),
    .Y(_0094_));
 sg13g2_nor2_1 _2157_ (.A(net26),
    .B(net14),
    .Y(_0095_));
 sg13g2_nor2_1 _2158_ (.A(net26),
    .B(_0730_),
    .Y(_0096_));
 sg13g2_nor2_1 _2159_ (.A(net26),
    .B(_0802_),
    .Y(_0097_));
 sg13g2_nor2_1 _2160_ (.A(net26),
    .B(_0775_),
    .Y(_0098_));
 sg13g2_nor2_1 _2161_ (.A(net26),
    .B(_0786_),
    .Y(_0099_));
 sg13g2_nor2_1 _2162_ (.A(_1099_),
    .B(_0617_),
    .Y(_0100_));
 sg13g2_nor2_1 _2163_ (.A(_1099_),
    .B(_0856_),
    .Y(_0101_));
 sg13g2_nor2_1 _2164_ (.A(net26),
    .B(_0838_),
    .Y(_0102_));
 sg13g2_nor2_1 _2165_ (.A(net26),
    .B(_0884_),
    .Y(_0103_));
 sg13g2_nand2_1 _2166_ (.Y(_1100_),
    .A(_0558_),
    .B(_0604_));
 sg13g2_inv_1 _2167_ (.Y(_1101_),
    .A(_1100_));
 sg13g2_nand3_1 _2168_ (.B(_0561_),
    .C(_0562_),
    .A(_0560_),
    .Y(_1102_));
 sg13g2_nor3_1 _2169_ (.A(_0555_),
    .B(\main.demo.vga._q_xcount[7] ),
    .C(_1102_),
    .Y(_1103_));
 sg13g2_a22oi_1 _2170_ (.Y(_1104_),
    .B1(\main.demo.vga._q_active_h ),
    .B2(net25),
    .A2(_1103_),
    .A1(_1101_));
 sg13g2_nor2_1 _2171_ (.A(net30),
    .B(_1104_),
    .Y(_0106_));
 sg13g2_nor2_1 _2172_ (.A(net30),
    .B(_0597_),
    .Y(_0107_));
 sg13g2_nor2_1 _2173_ (.A(\main.demo.vga._q_xcount[0] ),
    .B(_1095_),
    .Y(_0118_));
 sg13g2_nor3_1 _2174_ (.A(_0560_),
    .B(_0561_),
    .C(_0612_),
    .Y(_1105_));
 sg13g2_nand3_1 _2175_ (.B(_0605_),
    .C(_0606_),
    .A(_1101_),
    .Y(_1106_));
 sg13g2_inv_1 _2176_ (.Y(_1107_),
    .A(_1106_));
 sg13g2_a21oi_1 _2177_ (.A1(_1105_),
    .A2(_0562_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_nand2b_1 _2178_ (.Y(_1109_),
    .B(\main.demo.vga._q_xcount[10] ),
    .A_N(_1105_));
 sg13g2_a21oi_1 _2179_ (.A1(_1108_),
    .A2(_1109_),
    .Y(_0119_),
    .B1(net30));
 sg13g2_nand2_1 _2180_ (.Y(_1110_),
    .A(_0557_),
    .B(_0565_));
 sg13g2_a21oi_1 _2181_ (.A1(net25),
    .A2(_1110_),
    .Y(_0120_),
    .B1(net30));
 sg13g2_xnor2_1 _2182_ (.Y(_1111_),
    .A(_0564_),
    .B(_0565_));
 sg13g2_a21oi_1 _2183_ (.A1(net25),
    .A2(_1111_),
    .Y(_0121_),
    .B1(net30));
 sg13g2_xnor2_1 _2184_ (.Y(_1112_),
    .A(\main.demo.vga._q_xcount[3] ),
    .B(_0566_));
 sg13g2_a21oi_1 _2185_ (.A1(net25),
    .A2(_1112_),
    .Y(_0122_),
    .B1(net30));
 sg13g2_xnor2_1 _2186_ (.Y(_1113_),
    .A(_0554_),
    .B(_0568_));
 sg13g2_a21oi_1 _2187_ (.A1(net25),
    .A2(_1113_),
    .Y(_0123_),
    .B1(_1017_));
 sg13g2_xnor2_1 _2188_ (.Y(_1114_),
    .A(_0555_),
    .B(_0602_));
 sg13g2_a21oi_1 _2189_ (.A1(_1114_),
    .A2(net25),
    .Y(_0125_),
    .B1(_1017_));
 sg13g2_xnor2_1 _2190_ (.Y(_1115_),
    .A(_0561_),
    .B(_0612_));
 sg13g2_a21oi_1 _2191_ (.A1(_1115_),
    .A2(net25),
    .Y(_0127_),
    .B1(net24));
 sg13g2_a21oi_1 _2192_ (.A1(_0613_),
    .A2(\main.demo.vga._q_xcount[8] ),
    .Y(_1116_),
    .B1(\main.demo.vga._q_xcount[9] ));
 sg13g2_nor3_1 _2193_ (.A(net29),
    .B(_1105_),
    .C(_1116_),
    .Y(_0128_));
 sg13g2_nor2_1 _2194_ (.A(_0593_),
    .B(_1106_),
    .Y(_1117_));
 sg13g2_nor2_1 _2195_ (.A(_0574_),
    .B(_1106_),
    .Y(_1118_));
 sg13g2_nor2_1 _2196_ (.A(_0573_),
    .B(_1107_),
    .Y(_1119_));
 sg13g2_nor4_1 _2197_ (.A(net29),
    .B(_1117_),
    .C(_1118_),
    .D(_1119_),
    .Y(_0129_));
 sg13g2_xnor2_1 _2198_ (.Y(_1120_),
    .A(_0572_),
    .B(_1118_));
 sg13g2_inv_1 _2199_ (.Y(_1121_),
    .A(_1117_));
 sg13g2_a21oi_1 _2200_ (.A1(_1120_),
    .A2(_1121_),
    .Y(_0130_),
    .B1(net24));
 sg13g2_nor3_1 _2201_ (.A(_0585_),
    .B(_0574_),
    .C(net25),
    .Y(_1122_));
 sg13g2_nor2_1 _2202_ (.A(net31),
    .B(_1117_),
    .Y(_1123_));
 sg13g2_o21ai_1 _2203_ (.B1(_1123_),
    .Y(_1124_),
    .A1(_0580_),
    .A2(_1122_));
 sg13g2_nand2_1 _2204_ (.Y(_1125_),
    .A(_1122_),
    .B(_0580_));
 sg13g2_nor2b_1 _2205_ (.A(_1124_),
    .B_N(_1125_),
    .Y(_0131_));
 sg13g2_nand3_1 _2206_ (.B(_0572_),
    .C(_0582_),
    .A(_1118_),
    .Y(_1126_));
 sg13g2_nand2_1 _2207_ (.Y(_1127_),
    .A(_1126_),
    .B(_1123_));
 sg13g2_a21oi_1 _2208_ (.A1(_0598_),
    .A2(_1125_),
    .Y(_0132_),
    .B1(_1127_));
 sg13g2_nor4_1 _2209_ (.A(_0585_),
    .B(_0574_),
    .C(_0581_),
    .D(_0608_),
    .Y(_1128_));
 sg13g2_xnor2_1 _2210_ (.Y(_1129_),
    .A(\main.demo.vga._q_ycount[4] ),
    .B(_1128_));
 sg13g2_a21oi_1 _2211_ (.A1(_1129_),
    .A2(_1121_),
    .Y(_0133_),
    .B1(_0912_));
 sg13g2_nor2_1 _2212_ (.A(_0576_),
    .B(_1126_),
    .Y(_1130_));
 sg13g2_nand2_1 _2213_ (.Y(_1131_),
    .A(_1130_),
    .B(_0575_));
 sg13g2_inv_1 _2214_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_o21ai_1 _2215_ (.B1(_1123_),
    .Y(_1133_),
    .A1(_0575_),
    .A2(_1130_));
 sg13g2_nor2_1 _2216_ (.A(_1132_),
    .B(_1133_),
    .Y(_0134_));
 sg13g2_nor2_1 _2217_ (.A(_0599_),
    .B(_1131_),
    .Y(_1134_));
 sg13g2_nor2_1 _2218_ (.A(\main.demo.vga._q_ycount[6] ),
    .B(_1132_),
    .Y(_1135_));
 sg13g2_nor3_1 _2219_ (.A(net29),
    .B(_1134_),
    .C(_1135_),
    .Y(_0135_));
 sg13g2_nor2_1 _2220_ (.A(_0577_),
    .B(_1131_),
    .Y(_1136_));
 sg13g2_nor2_1 _2221_ (.A(\main.demo.vga._q_ycount[7] ),
    .B(_1134_),
    .Y(_1137_));
 sg13g2_nor3_1 _2222_ (.A(net29),
    .B(_1136_),
    .C(_1137_),
    .Y(_0136_));
 sg13g2_nor2_1 _2223_ (.A(_0579_),
    .B(_1136_),
    .Y(_1138_));
 sg13g2_nand2_1 _2224_ (.Y(_1139_),
    .A(_1136_),
    .B(_0579_));
 sg13g2_inv_1 _2225_ (.Y(_1140_),
    .A(_1139_));
 sg13g2_nor3_1 _2226_ (.A(net29),
    .B(_1138_),
    .C(_1140_),
    .Y(_0137_));
 sg13g2_xor2_1 _2227_ (.B(_1139_),
    .A(\main.demo.vga._d_vblank ),
    .X(_1141_));
 sg13g2_a21oi_1 _2228_ (.A1(_1141_),
    .A2(_1121_),
    .Y(_0138_),
    .B1(_0912_));
 sg13g2_nor2_1 _2229_ (.A(net21),
    .B(_1104_),
    .Y(\main.demo.vga._d_active ));
 sg13g2_buf_8 _2230_ (.A(\main.demo._q_rand_0[5] ),
    .X(_1142_));
 sg13g2_xnor2_1 _2231_ (.Y(_1143_),
    .A(\main.demo._q_rand_0[6] ),
    .B(_1142_));
 sg13g2_buf_8 _2232_ (.A(\main.demo._q_rand_0[4] ),
    .X(_1144_));
 sg13g2_nand2_2 _2233_ (.Y(_1145_),
    .A(_1144_),
    .B(_1142_));
 sg13g2_nand2_1 _2234_ (.Y(_1146_),
    .A(_1143_),
    .B(_1145_));
 sg13g2_inv_2 _2235_ (.Y(_1147_),
    .A(\main.demo._q_rand_0[6] ));
 sg13g2_nand3_1 _2236_ (.B(_1144_),
    .C(_1142_),
    .A(_1147_),
    .Y(_1148_));
 sg13g2_nand2_1 _2237_ (.Y(_1149_),
    .A(_1146_),
    .B(_1148_));
 sg13g2_buf_8 _2238_ (.A(\main.demo._q_rand_0[2] ),
    .X(_1150_));
 sg13g2_inv_2 _2239_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_buf_8 _2240_ (.A(\main.demo._q_rand_0[1] ),
    .X(_1152_));
 sg13g2_buf_1 _2241_ (.A(\main.demo._q_rand_0[0] ),
    .X(_1153_));
 sg13g2_nand2_1 _2242_ (.Y(_1154_),
    .A(_1152_),
    .B(_1153_));
 sg13g2_buf_2 _2243_ (.A(_1154_),
    .X(_1155_));
 sg13g2_nor2_1 _2244_ (.A(_1151_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_inv_1 _2245_ (.Y(_1157_),
    .A(_1156_));
 sg13g2_xnor2_1 _2246_ (.Y(_1158_),
    .A(_1156_),
    .B(_1149_));
 sg13g2_buf_8 _2247_ (.A(\main.demo._q_rand_0[3] ),
    .X(_1159_));
 sg13g2_nand2_1 _2248_ (.Y(_1160_),
    .A(_1159_),
    .B(_1144_));
 sg13g2_nor2_1 _2249_ (.A(_1142_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nand2_1 _2250_ (.Y(_1162_),
    .A(_1158_),
    .B(_1161_));
 sg13g2_o21ai_1 _2251_ (.B1(_1162_),
    .Y(_1163_),
    .A1(_1149_),
    .A2(_1157_));
 sg13g2_xnor2_1 _2252_ (.Y(_1164_),
    .A(_1161_),
    .B(_1158_));
 sg13g2_inv_2 _2253_ (.Y(_1165_),
    .A(_1153_));
 sg13g2_nand2_1 _2254_ (.Y(_1166_),
    .A(_1165_),
    .B(_1151_));
 sg13g2_nand2_1 _2255_ (.Y(_1167_),
    .A(_1153_),
    .B(_1150_));
 sg13g2_inv_1 _2256_ (.Y(_1168_),
    .A(_1167_));
 sg13g2_a21oi_1 _2257_ (.A1(_1166_),
    .A2(_1152_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_inv_4 _2258_ (.A(_1159_),
    .Y(_1170_));
 sg13g2_xor2_1 _2259_ (.B(_1150_),
    .A(_1152_),
    .X(_1171_));
 sg13g2_xnor2_1 _2260_ (.Y(_1172_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_nand2b_1 _2261_ (.Y(_1173_),
    .B(_1172_),
    .A_N(_1169_));
 sg13g2_inv_2 _2262_ (.Y(_1174_),
    .A(_1152_));
 sg13g2_nand2_1 _2263_ (.Y(_1175_),
    .A(_1174_),
    .B(_1151_));
 sg13g2_nand2_1 _2264_ (.Y(_1176_),
    .A(_1152_),
    .B(_1150_));
 sg13g2_nand2_1 _2265_ (.Y(_1177_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_nand2_1 _2266_ (.Y(_1178_),
    .A(_1177_),
    .B(_1170_));
 sg13g2_nand2_1 _2267_ (.Y(_1179_),
    .A(_1171_),
    .B(_1159_));
 sg13g2_nand2_1 _2268_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_nand2_1 _2269_ (.Y(_1181_),
    .A(_1180_),
    .B(_1169_));
 sg13g2_nand2_1 _2270_ (.Y(_1182_),
    .A(_1173_),
    .B(_1181_));
 sg13g2_xnor2_1 _2271_ (.Y(_1183_),
    .A(_1165_),
    .B(_1182_));
 sg13g2_inv_1 _2272_ (.Y(_1184_),
    .A(_1183_));
 sg13g2_nand2b_1 _2273_ (.Y(_1185_),
    .B(_1184_),
    .A_N(_1164_));
 sg13g2_buf_1 _2274_ (.A(\main.demo._q_rand_0[7] ),
    .X(_1186_));
 sg13g2_inv_2 _2275_ (.Y(_1187_),
    .A(_1142_));
 sg13g2_nand2_1 _2276_ (.Y(_1188_),
    .A(_1187_),
    .B(net39));
 sg13g2_inv_1 _2277_ (.Y(_1189_),
    .A(net39));
 sg13g2_a21oi_1 _2278_ (.A1(_1189_),
    .A2(_1142_),
    .Y(_1190_),
    .B1(_1147_));
 sg13g2_a22oi_1 _2279_ (.Y(_1191_),
    .B1(_1188_),
    .B2(_1190_),
    .A2(net39),
    .A1(_1147_));
 sg13g2_xor2_1 _2280_ (.B(_1173_),
    .A(_1191_),
    .X(_1192_));
 sg13g2_xor2_1 _2281_ (.B(_1192_),
    .A(_1148_),
    .X(_1193_));
 sg13g2_nor2_1 _2282_ (.A(_1165_),
    .B(_1182_),
    .Y(_1194_));
 sg13g2_nor2_1 _2283_ (.A(_1152_),
    .B(_1153_),
    .Y(_1195_));
 sg13g2_inv_1 _2284_ (.Y(_1196_),
    .A(_1155_));
 sg13g2_nor2_1 _2285_ (.A(_1195_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_buf_2 _2286_ (.A(_1197_),
    .X(_1198_));
 sg13g2_inv_1 _2287_ (.Y(_1199_),
    .A(_1176_));
 sg13g2_a21oi_2 _2288_ (.B1(_1199_),
    .Y(_1200_),
    .A2(_1159_),
    .A1(_1175_));
 sg13g2_xnor2_1 _2289_ (.Y(_1201_),
    .A(_1150_),
    .B(_1159_));
 sg13g2_xnor2_1 _2290_ (.Y(_1202_),
    .A(_1144_),
    .B(_1201_));
 sg13g2_nand2b_1 _2291_ (.Y(_1203_),
    .B(_1202_),
    .A_N(_1200_));
 sg13g2_inv_2 _2292_ (.Y(_1204_),
    .A(_1144_));
 sg13g2_nand2_1 _2293_ (.Y(_1205_),
    .A(_1201_),
    .B(_1204_));
 sg13g2_nand2_1 _2294_ (.Y(_1206_),
    .A(_1151_),
    .B(_1170_));
 sg13g2_nand2_2 _2295_ (.Y(_1207_),
    .A(_1150_),
    .B(_1159_));
 sg13g2_nand3_1 _2296_ (.B(_1144_),
    .C(_1207_),
    .A(_1206_),
    .Y(_1208_));
 sg13g2_nand2_2 _2297_ (.Y(_1209_),
    .A(_1205_),
    .B(_1208_));
 sg13g2_nand2_1 _2298_ (.Y(_1210_),
    .A(_1209_),
    .B(_1200_));
 sg13g2_nand2_1 _2299_ (.Y(_1211_),
    .A(_1203_),
    .B(_1210_));
 sg13g2_xnor2_1 _2300_ (.Y(_1212_),
    .A(_1198_),
    .B(_1211_));
 sg13g2_xnor2_1 _2301_ (.Y(_1213_),
    .A(_1194_),
    .B(_1212_));
 sg13g2_xor2_1 _2302_ (.B(_1213_),
    .A(_1193_),
    .X(_1214_));
 sg13g2_nand2b_1 _2303_ (.Y(_1215_),
    .B(_1214_),
    .A_N(_1185_));
 sg13g2_xnor2_1 _2304_ (.Y(_1216_),
    .A(_1193_),
    .B(_1213_));
 sg13g2_nand2_1 _2305_ (.Y(_1217_),
    .A(_1216_),
    .B(_1185_));
 sg13g2_nand2_1 _2306_ (.Y(_1218_),
    .A(_1215_),
    .B(_1217_));
 sg13g2_nand2b_1 _2307_ (.Y(_1219_),
    .B(_1218_),
    .A_N(_1163_));
 sg13g2_nand3_1 _2308_ (.B(_1217_),
    .C(_1163_),
    .A(_1215_),
    .Y(_1220_));
 sg13g2_nand2_1 _2309_ (.Y(_1221_),
    .A(_1204_),
    .B(_1187_));
 sg13g2_nand2_1 _2310_ (.Y(_1222_),
    .A(_1221_),
    .B(_1145_));
 sg13g2_xnor2_1 _2311_ (.Y(_1223_),
    .A(_1160_),
    .B(_1222_));
 sg13g2_nor2_1 _2312_ (.A(_1144_),
    .B(_1207_),
    .Y(_1224_));
 sg13g2_inv_1 _2313_ (.Y(_1225_),
    .A(_1224_));
 sg13g2_nand2_1 _2314_ (.Y(_1226_),
    .A(_1223_),
    .B(_1225_));
 sg13g2_nand2_1 _2315_ (.Y(_1227_),
    .A(_1166_),
    .B(_1167_));
 sg13g2_a21oi_1 _2316_ (.A1(_1227_),
    .A2(_1174_),
    .Y(_1228_),
    .B1(_1199_));
 sg13g2_nor2_1 _2317_ (.A(_1187_),
    .B(_1225_),
    .Y(_1229_));
 sg13g2_inv_1 _2318_ (.Y(_1230_),
    .A(_1229_));
 sg13g2_nand3_1 _2319_ (.B(_1228_),
    .C(_1230_),
    .A(_1226_),
    .Y(_1231_));
 sg13g2_buf_1 _2320_ (.A(_1231_),
    .X(_1232_));
 sg13g2_nand2_1 _2321_ (.Y(_1233_),
    .A(_1183_),
    .B(_1164_));
 sg13g2_nand3b_1 _2322_ (.B(_1185_),
    .C(_1233_),
    .Y(_1234_),
    .A_N(_1232_));
 sg13g2_xnor2_1 _2323_ (.Y(_1235_),
    .A(_1164_),
    .B(_1183_));
 sg13g2_nand2_1 _2324_ (.Y(_1236_),
    .A(_1235_),
    .B(_1232_));
 sg13g2_nand3_1 _2325_ (.B(_1236_),
    .C(_1229_),
    .A(_1234_),
    .Y(_1237_));
 sg13g2_nand2_1 _2326_ (.Y(_1238_),
    .A(_1237_),
    .B(_1234_));
 sg13g2_a21oi_1 _2327_ (.A1(_1219_),
    .A2(_1220_),
    .Y(_1239_),
    .B1(_1238_));
 sg13g2_nand2_1 _2328_ (.Y(_1240_),
    .A(_1199_),
    .B(_1170_));
 sg13g2_nor2_1 _2329_ (.A(_1204_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nand2_1 _2330_ (.Y(_1242_),
    .A(_1176_),
    .B(_1170_));
 sg13g2_a21o_1 _2331_ (.A2(_1207_),
    .A1(_1242_),
    .B1(_1204_),
    .X(_1243_));
 sg13g2_nand3_1 _2332_ (.B(_1204_),
    .C(_1207_),
    .A(_1242_),
    .Y(_1244_));
 sg13g2_nand2_1 _2333_ (.Y(_1245_),
    .A(_1243_),
    .B(_1244_));
 sg13g2_nand2_1 _2334_ (.Y(_1246_),
    .A(_1245_),
    .B(_1198_));
 sg13g2_nand2_1 _2335_ (.Y(_1247_),
    .A(_1226_),
    .B(_1230_));
 sg13g2_nand2b_1 _2336_ (.Y(_1248_),
    .B(_1247_),
    .A_N(_1228_));
 sg13g2_nand3b_1 _2337_ (.B(_1248_),
    .C(_1232_),
    .Y(_1249_),
    .A_N(_1246_));
 sg13g2_nand2_1 _2338_ (.Y(_1250_),
    .A(_1248_),
    .B(_1232_));
 sg13g2_nand2_1 _2339_ (.Y(_1251_),
    .A(_1250_),
    .B(_1246_));
 sg13g2_nand2_1 _2340_ (.Y(_1252_),
    .A(_1249_),
    .B(_1251_));
 sg13g2_xor2_1 _2341_ (.B(_1252_),
    .A(_1241_),
    .X(_1253_));
 sg13g2_inv_1 _2342_ (.Y(_1254_),
    .A(_1198_));
 sg13g2_nand3_1 _2343_ (.B(_1244_),
    .C(_1254_),
    .A(_1243_),
    .Y(_1255_));
 sg13g2_nand2_1 _2344_ (.Y(_1256_),
    .A(_1201_),
    .B(_1176_));
 sg13g2_nand2_1 _2345_ (.Y(_1257_),
    .A(_1256_),
    .B(_1240_));
 sg13g2_nor2_1 _2346_ (.A(_1165_),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_nand3_1 _2347_ (.B(_1255_),
    .C(_1258_),
    .A(_1246_),
    .Y(_1259_));
 sg13g2_nand2_1 _2348_ (.Y(_1260_),
    .A(_1253_),
    .B(_1259_));
 sg13g2_nor3_1 _2349_ (.A(_1196_),
    .B(_1195_),
    .C(_1177_),
    .Y(_1261_));
 sg13g2_inv_1 _2350_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_o21ai_1 _2351_ (.B1(_1258_),
    .Y(_1263_),
    .A1(_1174_),
    .A2(_1150_));
 sg13g2_nand2_1 _2352_ (.Y(_1264_),
    .A(_1257_),
    .B(_1165_));
 sg13g2_nor2_1 _2353_ (.A(_1155_),
    .B(_1206_),
    .Y(_1265_));
 sg13g2_inv_1 _2354_ (.Y(_1266_),
    .A(_1265_));
 sg13g2_nand3_1 _2355_ (.B(_1264_),
    .C(_1266_),
    .A(_1263_),
    .Y(_1267_));
 sg13g2_nand2_1 _2356_ (.Y(_1268_),
    .A(_1156_),
    .B(_1170_));
 sg13g2_o21ai_1 _2357_ (.B1(_1268_),
    .Y(_1269_),
    .A1(_1262_),
    .A2(_1267_));
 sg13g2_nand2_1 _2358_ (.Y(_1270_),
    .A(_1246_),
    .B(_1255_));
 sg13g2_xor2_1 _2359_ (.B(_1270_),
    .A(_1258_),
    .X(_1271_));
 sg13g2_nand2_1 _2360_ (.Y(_1272_),
    .A(_1271_),
    .B(_1266_));
 sg13g2_nor2_1 _2361_ (.A(_1266_),
    .B(_1271_),
    .Y(_1273_));
 sg13g2_a21oi_1 _2362_ (.A1(_1269_),
    .A2(_1272_),
    .Y(_1274_),
    .B1(_1273_));
 sg13g2_inv_1 _2363_ (.Y(_1275_),
    .A(_1274_));
 sg13g2_nor2_1 _2364_ (.A(_1259_),
    .B(_1253_),
    .Y(_1276_));
 sg13g2_a21oi_1 _2365_ (.A1(_1260_),
    .A2(_1275_),
    .Y(_1277_),
    .B1(_1276_));
 sg13g2_inv_1 _2366_ (.Y(_1278_),
    .A(_1277_));
 sg13g2_nand2_1 _2367_ (.Y(_1279_),
    .A(_1234_),
    .B(_1236_));
 sg13g2_nand2_1 _2368_ (.Y(_1280_),
    .A(_1279_),
    .B(_1230_));
 sg13g2_nand2_1 _2369_ (.Y(_1281_),
    .A(_1280_),
    .B(_1237_));
 sg13g2_inv_1 _2370_ (.Y(_1282_),
    .A(_1249_));
 sg13g2_a21oi_1 _2371_ (.A1(_1251_),
    .A2(_1241_),
    .Y(_1283_),
    .B1(_1282_));
 sg13g2_nand2_1 _2372_ (.Y(_1284_),
    .A(_1281_),
    .B(_1283_));
 sg13g2_nor2_1 _2373_ (.A(_1283_),
    .B(_1281_),
    .Y(_1285_));
 sg13g2_a21oi_1 _2374_ (.A1(_1278_),
    .A2(_1284_),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_nand3_1 _2375_ (.B(_1220_),
    .C(_1238_),
    .A(_1219_),
    .Y(_1287_));
 sg13g2_o21ai_1 _2376_ (.B1(_1287_),
    .Y(_1288_),
    .A1(_1239_),
    .A2(_1286_));
 sg13g2_nor2_1 _2377_ (.A(_1193_),
    .B(_1213_),
    .Y(_1289_));
 sg13g2_nand2_1 _2378_ (.Y(_1290_),
    .A(_1212_),
    .B(_1194_));
 sg13g2_nor2b_1 _2379_ (.A(_1289_),
    .B_N(_1290_),
    .Y(_1291_));
 sg13g2_nand2_1 _2380_ (.Y(_1292_),
    .A(_1211_),
    .B(_1198_));
 sg13g2_nand2_2 _2381_ (.Y(_1293_),
    .A(_1208_),
    .B(_1207_));
 sg13g2_nor2_1 _2382_ (.A(_1155_),
    .B(_1209_),
    .Y(_1294_));
 sg13g2_nand2_1 _2383_ (.Y(_1295_),
    .A(_1209_),
    .B(_1155_));
 sg13g2_nor2b_1 _2384_ (.A(_1294_),
    .B_N(_1295_),
    .Y(_1296_));
 sg13g2_xnor2_1 _2385_ (.Y(_1297_),
    .A(_1293_),
    .B(_1296_));
 sg13g2_xnor2_1 _2386_ (.Y(_1298_),
    .A(_1292_),
    .B(_1297_));
 sg13g2_nor3_1 _2387_ (.A(net39),
    .B(_1147_),
    .C(_1187_),
    .Y(_1299_));
 sg13g2_buf_2 _2388_ (.A(\main.demo._q_rand_0[8] ),
    .X(_1300_));
 sg13g2_nand2_1 _2389_ (.Y(_1301_),
    .A(_1143_),
    .B(net39));
 sg13g2_o21ai_1 _2390_ (.B1(_1301_),
    .Y(_1302_),
    .A1(_1187_),
    .A2(net39));
 sg13g2_xnor2_1 _2391_ (.Y(_1303_),
    .A(_1300_),
    .B(_1302_));
 sg13g2_xnor2_1 _2392_ (.Y(_1304_),
    .A(_1203_),
    .B(_1303_));
 sg13g2_xnor2_1 _2393_ (.Y(_1305_),
    .A(_1299_),
    .B(_1304_));
 sg13g2_xor2_1 _2394_ (.B(_1305_),
    .A(_1298_),
    .X(_1306_));
 sg13g2_nand2b_1 _2395_ (.Y(_1307_),
    .B(_1306_),
    .A_N(_1291_));
 sg13g2_xnor2_1 _2396_ (.Y(_1308_),
    .A(_1298_),
    .B(_1305_));
 sg13g2_nand2_1 _2397_ (.Y(_1309_),
    .A(_1308_),
    .B(_1291_));
 sg13g2_nand2_1 _2398_ (.Y(_1310_),
    .A(_1307_),
    .B(_1309_));
 sg13g2_nor2_1 _2399_ (.A(_1191_),
    .B(_1173_),
    .Y(_1311_));
 sg13g2_nor2b_1 _2400_ (.A(_1148_),
    .B_N(_1192_),
    .Y(_1312_));
 sg13g2_nor2_1 _2401_ (.A(_1311_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_nand2_1 _2402_ (.Y(_1314_),
    .A(_1310_),
    .B(_1313_));
 sg13g2_inv_1 _2403_ (.Y(_1315_),
    .A(_1313_));
 sg13g2_nand3_1 _2404_ (.B(_1309_),
    .C(_1315_),
    .A(_1307_),
    .Y(_1316_));
 sg13g2_inv_1 _2405_ (.Y(_1317_),
    .A(_1215_));
 sg13g2_a21oi_1 _2406_ (.A1(_1217_),
    .A2(_1163_),
    .Y(_1318_),
    .B1(_1317_));
 sg13g2_inv_1 _2407_ (.Y(_1319_),
    .A(_1318_));
 sg13g2_a21oi_1 _2408_ (.A1(_1314_),
    .A2(_1316_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nand3_1 _2409_ (.B(_1316_),
    .C(_1319_),
    .A(_1314_),
    .Y(_1321_));
 sg13g2_nor2b_1 _2410_ (.A(_1320_),
    .B_N(_1321_),
    .Y(_1322_));
 sg13g2_nand2_1 _2411_ (.Y(_1323_),
    .A(_1288_),
    .B(_1322_));
 sg13g2_nand2_1 _2412_ (.Y(_1324_),
    .A(_1323_),
    .B(_1321_));
 sg13g2_and2_1 _2413_ (.A(_1316_),
    .B(_1307_),
    .X(_1325_));
 sg13g2_nor2_1 _2414_ (.A(_1198_),
    .B(_1297_),
    .Y(_1326_));
 sg13g2_inv_1 _2415_ (.Y(_1327_),
    .A(_1326_));
 sg13g2_inv_1 _2416_ (.Y(_1328_),
    .A(_0013_));
 sg13g2_nand2_1 _2417_ (.Y(_1329_),
    .A(_1172_),
    .B(_1328_));
 sg13g2_nand2_1 _2418_ (.Y(_1330_),
    .A(_1180_),
    .B(_0013_));
 sg13g2_nand2_1 _2419_ (.Y(_1331_),
    .A(_1329_),
    .B(_1330_));
 sg13g2_xnor2_1 _2420_ (.Y(_1332_),
    .A(_1198_),
    .B(_1331_));
 sg13g2_nand2_1 _2421_ (.Y(_1333_),
    .A(_1222_),
    .B(_1147_));
 sg13g2_nand3_1 _2422_ (.B(\main.demo._q_rand_0[6] ),
    .C(_1145_),
    .A(_1221_),
    .Y(_1334_));
 sg13g2_nand2_1 _2423_ (.Y(_1335_),
    .A(_1333_),
    .B(_1334_));
 sg13g2_nor2_1 _2424_ (.A(_1155_),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_nand2_1 _2425_ (.Y(_1337_),
    .A(_1335_),
    .B(_1155_));
 sg13g2_nand2b_1 _2426_ (.Y(_1338_),
    .B(_1337_),
    .A_N(_1336_));
 sg13g2_xnor2_1 _2427_ (.Y(_1339_),
    .A(_1293_),
    .B(_1338_));
 sg13g2_xnor2_1 _2428_ (.Y(_1340_),
    .A(_1332_),
    .B(_1339_));
 sg13g2_nor2_1 _2429_ (.A(_1327_),
    .B(_1340_),
    .Y(_1341_));
 sg13g2_inv_1 _2430_ (.Y(_1342_),
    .A(_1341_));
 sg13g2_nand2_1 _2431_ (.Y(_1343_),
    .A(_1340_),
    .B(_1327_));
 sg13g2_nand2_1 _2432_ (.Y(_1344_),
    .A(_1342_),
    .B(_1343_));
 sg13g2_inv_1 _2433_ (.Y(_1345_),
    .A(_1344_));
 sg13g2_nor2_1 _2434_ (.A(_1147_),
    .B(_1188_),
    .Y(_1346_));
 sg13g2_a21oi_1 _2435_ (.A1(_1302_),
    .A2(_1300_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_nand2_1 _2436_ (.Y(_1348_),
    .A(_1142_),
    .B(net39));
 sg13g2_xnor2_1 _2437_ (.Y(_1349_),
    .A(_1300_),
    .B(\main.demo._q_rand_0[9] ));
 sg13g2_xor2_1 _2438_ (.B(_1349_),
    .A(_1348_),
    .X(_1350_));
 sg13g2_a21oi_1 _2439_ (.A1(_1295_),
    .A2(_1293_),
    .Y(_1351_),
    .B1(_1294_));
 sg13g2_xnor2_1 _2440_ (.Y(_1352_),
    .A(_1350_),
    .B(_1351_));
 sg13g2_xnor2_1 _2441_ (.Y(_1353_),
    .A(_1347_),
    .B(_1352_));
 sg13g2_inv_1 _2442_ (.Y(_1354_),
    .A(_1353_));
 sg13g2_nand2_1 _2443_ (.Y(_1355_),
    .A(_1345_),
    .B(_1354_));
 sg13g2_nand2_1 _2444_ (.Y(_1356_),
    .A(_1344_),
    .B(_1353_));
 sg13g2_nand2_1 _2445_ (.Y(_1357_),
    .A(_1355_),
    .B(_1356_));
 sg13g2_nor2_1 _2446_ (.A(_1254_),
    .B(_1211_),
    .Y(_1358_));
 sg13g2_a21oi_1 _2447_ (.A1(_1305_),
    .A2(_1298_),
    .Y(_1359_),
    .B1(_1358_));
 sg13g2_inv_1 _2448_ (.Y(_1360_),
    .A(_1359_));
 sg13g2_nand2_1 _2449_ (.Y(_1361_),
    .A(_1357_),
    .B(_1360_));
 sg13g2_nand3_1 _2450_ (.B(_1359_),
    .C(_1356_),
    .A(_1355_),
    .Y(_1362_));
 sg13g2_nand2_1 _2451_ (.Y(_1363_),
    .A(_1361_),
    .B(_1362_));
 sg13g2_nor2_1 _2452_ (.A(_1203_),
    .B(_1303_),
    .Y(_1364_));
 sg13g2_nor2b_1 _2453_ (.A(_1304_),
    .B_N(_1299_),
    .Y(_1365_));
 sg13g2_nor2_1 _2454_ (.A(_1364_),
    .B(_1365_),
    .Y(_1366_));
 sg13g2_nand2_1 _2455_ (.Y(_1367_),
    .A(_1363_),
    .B(_1366_));
 sg13g2_inv_1 _2456_ (.Y(_1368_),
    .A(_1366_));
 sg13g2_nand3_1 _2457_ (.B(_1362_),
    .C(_1368_),
    .A(_1361_),
    .Y(_1369_));
 sg13g2_nand2_1 _2458_ (.Y(_1370_),
    .A(_1367_),
    .B(_1369_));
 sg13g2_xor2_1 _2459_ (.B(_1370_),
    .A(_1325_),
    .X(_1371_));
 sg13g2_nand2_1 _2460_ (.Y(_1372_),
    .A(_1324_),
    .B(_1371_));
 sg13g2_nor2_1 _2461_ (.A(_1325_),
    .B(_1370_),
    .Y(_1373_));
 sg13g2_inv_1 _2462_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_nand2_1 _2463_ (.Y(_1375_),
    .A(_1372_),
    .B(_1374_));
 sg13g2_inv_1 _2464_ (.Y(_1376_),
    .A(_1347_));
 sg13g2_nor2b_1 _2465_ (.A(_1351_),
    .B_N(_1350_),
    .Y(_1377_));
 sg13g2_a21oi_1 _2466_ (.A1(_1352_),
    .A2(_1376_),
    .Y(_1378_),
    .B1(_1377_));
 sg13g2_a21oi_1 _2467_ (.A1(_1343_),
    .A2(_1353_),
    .Y(_1379_),
    .B1(_1341_));
 sg13g2_nor2_1 _2468_ (.A(_1348_),
    .B(_1349_),
    .Y(_1380_));
 sg13g2_a21oi_1 _2469_ (.A1(_1337_),
    .A2(_1293_),
    .Y(_1381_),
    .B1(_1336_));
 sg13g2_nand2_1 _2470_ (.Y(_1382_),
    .A(_1300_),
    .B(\main.demo._q_rand_0[9] ));
 sg13g2_nor2_1 _2471_ (.A(net39),
    .B(\main.demo._q_rand_0[9] ),
    .Y(_1383_));
 sg13g2_nand2_1 _2472_ (.Y(_1384_),
    .A(_1186_),
    .B(\main.demo._q_rand_0[9] ));
 sg13g2_inv_1 _2473_ (.Y(_1385_),
    .A(_1384_));
 sg13g2_o21ai_1 _2474_ (.B1(_1382_),
    .Y(_1386_),
    .A1(_1383_),
    .A2(_1385_));
 sg13g2_o21ai_1 _2475_ (.B1(_1386_),
    .Y(_1387_),
    .A1(_1186_),
    .A2(_1382_));
 sg13g2_xnor2_1 _2476_ (.Y(_1388_),
    .A(\main.demo._q_rand_0[10] ),
    .B(_1387_));
 sg13g2_xnor2_1 _2477_ (.Y(_1389_),
    .A(_1381_),
    .B(_1388_));
 sg13g2_xor2_1 _2478_ (.B(_1389_),
    .A(_1380_),
    .X(_1390_));
 sg13g2_nand2_2 _2479_ (.Y(_1391_),
    .A(_1334_),
    .B(_1145_));
 sg13g2_xnor2_1 _2480_ (.Y(_1392_),
    .A(_1200_),
    .B(_1335_));
 sg13g2_xor2_1 _2481_ (.B(_1392_),
    .A(_1391_),
    .X(_1393_));
 sg13g2_xor2_1 _2482_ (.B(_1393_),
    .A(_1330_),
    .X(_1394_));
 sg13g2_nand2_1 _2483_ (.Y(_1395_),
    .A(_1339_),
    .B(_1332_));
 sg13g2_o21ai_1 _2484_ (.B1(_1395_),
    .Y(_1396_),
    .A1(_1254_),
    .A2(_1331_));
 sg13g2_or2_1 _2485_ (.X(_1397_),
    .B(_1396_),
    .A(_1394_));
 sg13g2_buf_1 _2486_ (.A(_1397_),
    .X(_1398_));
 sg13g2_nand2_1 _2487_ (.Y(_1399_),
    .A(_1396_),
    .B(_1394_));
 sg13g2_nand3b_1 _2488_ (.B(_1398_),
    .C(_1399_),
    .Y(_1400_),
    .A_N(_1390_));
 sg13g2_nand2_1 _2489_ (.Y(_1401_),
    .A(_1398_),
    .B(_1399_));
 sg13g2_nand2_1 _2490_ (.Y(_1402_),
    .A(_1401_),
    .B(_1390_));
 sg13g2_nand2_1 _2491_ (.Y(_1403_),
    .A(_1400_),
    .B(_1402_));
 sg13g2_nand2b_1 _2492_ (.Y(_1404_),
    .B(_1403_),
    .A_N(_1379_));
 sg13g2_nand3_1 _2493_ (.B(_1402_),
    .C(_1379_),
    .A(_1400_),
    .Y(_1405_));
 sg13g2_nand3b_1 _2494_ (.B(_1404_),
    .C(_1405_),
    .Y(_1406_),
    .A_N(_1378_));
 sg13g2_nand2_1 _2495_ (.Y(_1407_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_nand2_1 _2496_ (.Y(_1408_),
    .A(_1407_),
    .B(_1378_));
 sg13g2_nand2_1 _2497_ (.Y(_1409_),
    .A(_1406_),
    .B(_1408_));
 sg13g2_inv_1 _2498_ (.Y(_1410_),
    .A(_1361_));
 sg13g2_a21oi_1 _2499_ (.A1(_1362_),
    .A2(_1368_),
    .Y(_1411_),
    .B1(_1410_));
 sg13g2_nand2_1 _2500_ (.Y(_1412_),
    .A(_1409_),
    .B(_1411_));
 sg13g2_inv_1 _2501_ (.Y(_1413_),
    .A(_1411_));
 sg13g2_nand3_1 _2502_ (.B(_1408_),
    .C(_1413_),
    .A(_1406_),
    .Y(_1414_));
 sg13g2_nand2_1 _2503_ (.Y(_1415_),
    .A(_1412_),
    .B(_1414_));
 sg13g2_inv_1 _2504_ (.Y(_1416_),
    .A(_1415_));
 sg13g2_nand2_2 _2505_ (.Y(_1417_),
    .A(_1375_),
    .B(_1416_));
 sg13g2_nand3_1 _2506_ (.B(_1374_),
    .C(_1415_),
    .A(_1372_),
    .Y(_1418_));
 sg13g2_xnor2_1 _2507_ (.Y(_1419_),
    .A(\main.demo._q_frame[15] ),
    .B(\main.demo._q_modulo_0[15] ));
 sg13g2_buf_1 _2508_ (.A(\main.demo._q_frame[14] ),
    .X(_1420_));
 sg13g2_inv_1 _2509_ (.Y(_1421_),
    .A(_1420_));
 sg13g2_nor2_1 _2510_ (.A(\main.demo._q_modulo_0[14] ),
    .B(_1421_),
    .Y(_1422_));
 sg13g2_inv_1 _2511_ (.Y(_1423_),
    .A(\main.demo._q_modulo_0[14] ));
 sg13g2_nor2_1 _2512_ (.A(_1420_),
    .B(_1423_),
    .Y(_1424_));
 sg13g2_nor2_1 _2513_ (.A(_1422_),
    .B(_1424_),
    .Y(_1425_));
 sg13g2_inv_1 _2514_ (.Y(_1426_),
    .A(_1425_));
 sg13g2_inv_1 _2515_ (.Y(_1427_),
    .A(\main.demo._q_frame[13] ));
 sg13g2_nor2_1 _2516_ (.A(\main.demo._q_modulo_0[13] ),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_inv_1 _2517_ (.Y(_1429_),
    .A(\main.demo._q_modulo_0[13] ));
 sg13g2_nor2_1 _2518_ (.A(\main.demo._q_frame[13] ),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_nor2_1 _2519_ (.A(_1428_),
    .B(_1430_),
    .Y(_1431_));
 sg13g2_inv_1 _2520_ (.Y(_1432_),
    .A(_1431_));
 sg13g2_buf_1 _2521_ (.A(\main.demo._q_frame[12] ),
    .X(_1433_));
 sg13g2_buf_1 _2522_ (.A(\main.demo._q_modulo_0[12] ),
    .X(_1434_));
 sg13g2_xnor2_1 _2523_ (.Y(_1435_),
    .A(_1433_),
    .B(_1434_));
 sg13g2_buf_1 _2524_ (.A(\main.demo._q_frame[11] ),
    .X(_1436_));
 sg13g2_xnor2_1 _2525_ (.Y(_1437_),
    .A(_1436_),
    .B(\main.demo._q_modulo_0[11] ));
 sg13g2_nand2_1 _2526_ (.Y(_1438_),
    .A(_1435_),
    .B(_1437_));
 sg13g2_nor3_1 _2527_ (.A(_1426_),
    .B(_1432_),
    .C(_1438_),
    .Y(_1439_));
 sg13g2_buf_1 _2528_ (.A(\main.demo._q_frame[10] ),
    .X(_1440_));
 sg13g2_inv_1 _2529_ (.Y(_1441_),
    .A(_1440_));
 sg13g2_nor2_1 _2530_ (.A(\main.demo._q_modulo_0[10] ),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_inv_1 _2531_ (.Y(_1443_),
    .A(\main.demo._q_modulo_0[10] ));
 sg13g2_nor2_1 _2532_ (.A(_1440_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_nor2_2 _2533_ (.A(_1442_),
    .B(_1444_),
    .Y(_1445_));
 sg13g2_inv_1 _2534_ (.Y(_1446_),
    .A(_1445_));
 sg13g2_inv_1 _2535_ (.Y(_1447_),
    .A(\main.demo._q_frame[9] ));
 sg13g2_nor2_1 _2536_ (.A(\main.demo._q_modulo_0[9] ),
    .B(_1447_),
    .Y(_1448_));
 sg13g2_inv_1 _2537_ (.Y(_1449_),
    .A(\main.demo._q_modulo_0[9] ));
 sg13g2_nor2_1 _2538_ (.A(\main.demo._q_frame[9] ),
    .B(_1449_),
    .Y(_1450_));
 sg13g2_nor2_1 _2539_ (.A(_1448_),
    .B(_1450_),
    .Y(_1451_));
 sg13g2_inv_1 _2540_ (.Y(_1452_),
    .A(_1451_));
 sg13g2_nor2_1 _2541_ (.A(_1446_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_buf_1 _2542_ (.A(\main.demo._q_frame[8] ),
    .X(_1454_));
 sg13g2_inv_1 _2543_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_nor2_1 _2544_ (.A(\main.demo._q_modulo_0[8] ),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_inv_1 _2545_ (.Y(_1457_),
    .A(\main.demo._q_modulo_0[8] ));
 sg13g2_nor2_1 _2546_ (.A(_1454_),
    .B(_1457_),
    .Y(_1458_));
 sg13g2_nor2_2 _2547_ (.A(_1456_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_buf_1 _2548_ (.A(\main.demo._q_frame[7] ),
    .X(_1460_));
 sg13g2_buf_1 _2549_ (.A(\main.demo._q_modulo_0[7] ),
    .X(_1461_));
 sg13g2_xnor2_1 _2550_ (.Y(_1462_),
    .A(_1460_),
    .B(_1461_));
 sg13g2_nand4_1 _2551_ (.B(_1453_),
    .C(_1459_),
    .A(_1439_),
    .Y(_1463_),
    .D(_1462_));
 sg13g2_buf_2 _2552_ (.A(\main.demo._q_frame[4] ),
    .X(_1464_));
 sg13g2_inv_1 _2553_ (.Y(_1465_),
    .A(\main.demo._q_modulo_0[4] ));
 sg13g2_nor2_1 _2554_ (.A(_1464_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_buf_2 _2555_ (.A(\main.demo._q_frame[3] ),
    .X(_1467_));
 sg13g2_inv_1 _2556_ (.Y(_1468_),
    .A(_1467_));
 sg13g2_nor2_1 _2557_ (.A(\main.demo._q_modulo_0[3] ),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_inv_1 _2558_ (.Y(_1470_),
    .A(_1469_));
 sg13g2_inv_1 _2559_ (.Y(_1471_),
    .A(_1464_));
 sg13g2_nor2_1 _2560_ (.A(\main.demo._q_modulo_0[4] ),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_inv_1 _2561_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_o21ai_1 _2562_ (.B1(_1473_),
    .Y(_1474_),
    .A1(_1466_),
    .A2(_1470_));
 sg13g2_buf_2 _2563_ (.A(\main.demo._q_frame[5] ),
    .X(_1475_));
 sg13g2_inv_1 _2564_ (.Y(_1476_),
    .A(_1475_));
 sg13g2_nor2_2 _2565_ (.A(\main.demo._q_modulo_0[5] ),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_inv_1 _2566_ (.Y(_1478_),
    .A(\main.demo._q_modulo_0[5] ));
 sg13g2_nor2_1 _2567_ (.A(_1475_),
    .B(_1478_),
    .Y(_1479_));
 sg13g2_nor2_1 _2568_ (.A(_1477_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_buf_1 _2569_ (.A(\main.demo._q_frame[6] ),
    .X(_1481_));
 sg13g2_buf_1 _2570_ (.A(\main.demo._q_modulo_0[6] ),
    .X(_1482_));
 sg13g2_xnor2_1 _2571_ (.Y(_1483_),
    .A(_1481_),
    .B(_1482_));
 sg13g2_nand2_1 _2572_ (.Y(_1484_),
    .A(_1480_),
    .B(_1483_));
 sg13g2_inv_1 _2573_ (.Y(_1485_),
    .A(_1484_));
 sg13g2_buf_2 _2574_ (.A(\main.demo._q_frame[1] ),
    .X(_1486_));
 sg13g2_buf_1 _2575_ (.A(\main.demo._q_modulo_0[1] ),
    .X(_1487_));
 sg13g2_xnor2_1 _2576_ (.Y(_1488_),
    .A(_1486_),
    .B(_1487_));
 sg13g2_buf_2 _2577_ (.A(\main.demo._q_frame[0] ),
    .X(_1489_));
 sg13g2_inv_1 _2578_ (.Y(_1490_),
    .A(_1489_));
 sg13g2_buf_1 _2579_ (.A(\main.demo._q_modulo_0[0] ),
    .X(_1491_));
 sg13g2_nand2_1 _2580_ (.Y(_1492_),
    .A(_1490_),
    .B(_1491_));
 sg13g2_inv_1 _2581_ (.Y(_1493_),
    .A(_1486_));
 sg13g2_nor2_1 _2582_ (.A(_1487_),
    .B(_1493_),
    .Y(_1494_));
 sg13g2_a21oi_1 _2583_ (.A1(_1488_),
    .A2(_1492_),
    .Y(_1495_),
    .B1(_1494_));
 sg13g2_buf_2 _2584_ (.A(\main.demo._q_frame[2] ),
    .X(_1496_));
 sg13g2_inv_1 _2585_ (.Y(_1497_),
    .A(_1496_));
 sg13g2_nor2_1 _2586_ (.A(\main.demo._q_modulo_0[2] ),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_inv_1 _2587_ (.Y(_1499_),
    .A(_1498_));
 sg13g2_inv_1 _2588_ (.Y(_1500_),
    .A(\main.demo._q_modulo_0[2] ));
 sg13g2_nor2_1 _2589_ (.A(_1496_),
    .B(_1500_),
    .Y(_1501_));
 sg13g2_a21oi_1 _2590_ (.A1(_1495_),
    .A2(_1499_),
    .Y(_1502_),
    .B1(_1501_));
 sg13g2_xnor2_1 _2591_ (.Y(_1503_),
    .A(_1467_),
    .B(\main.demo._q_modulo_0[3] ));
 sg13g2_inv_1 _2592_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_nor2_1 _2593_ (.A(_1466_),
    .B(_1472_),
    .Y(_1505_));
 sg13g2_inv_1 _2594_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_nor3_1 _2595_ (.A(_1504_),
    .B(_1506_),
    .C(_1484_),
    .Y(_1507_));
 sg13g2_inv_1 _2596_ (.Y(_1508_),
    .A(_1481_));
 sg13g2_nor2_1 _2597_ (.A(_1482_),
    .B(_1508_),
    .Y(_1509_));
 sg13g2_a21o_1 _2598_ (.A2(_1477_),
    .A1(_1483_),
    .B1(_1509_),
    .X(_1510_));
 sg13g2_a221oi_1 _2599_ (.B2(_1507_),
    .C1(_1510_),
    .B1(_1502_),
    .A1(_1474_),
    .Y(_1511_),
    .A2(_1485_));
 sg13g2_buf_1 _2600_ (.A(_1511_),
    .X(_1512_));
 sg13g2_inv_1 _2601_ (.Y(_1513_),
    .A(_1436_));
 sg13g2_nor2_1 _2602_ (.A(\main.demo._q_modulo_0[11] ),
    .B(_1513_),
    .Y(_1514_));
 sg13g2_inv_1 _2603_ (.Y(_1515_),
    .A(_1433_));
 sg13g2_nor2_1 _2604_ (.A(_1434_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_a21oi_1 _2605_ (.A1(_1435_),
    .A2(_1514_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_inv_1 _2606_ (.Y(_1518_),
    .A(_1517_));
 sg13g2_nor2_1 _2607_ (.A(_1426_),
    .B(_1432_),
    .Y(_1519_));
 sg13g2_inv_1 _2608_ (.Y(_1520_),
    .A(_1453_));
 sg13g2_inv_1 _2609_ (.Y(_1521_),
    .A(_1460_));
 sg13g2_nor2_1 _2610_ (.A(_1461_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_a21oi_1 _2611_ (.A1(_1459_),
    .A2(_1522_),
    .Y(_1523_),
    .B1(_1456_));
 sg13g2_a21oi_1 _2612_ (.A1(_1445_),
    .A2(_1448_),
    .Y(_1524_),
    .B1(_1442_));
 sg13g2_o21ai_1 _2613_ (.B1(_1524_),
    .Y(_1525_),
    .A1(_1520_),
    .A2(_1523_));
 sg13g2_nand2_1 _2614_ (.Y(_1526_),
    .A(_1425_),
    .B(_1428_));
 sg13g2_o21ai_1 _2615_ (.B1(_1526_),
    .Y(_1527_),
    .A1(_1421_),
    .A2(\main.demo._q_modulo_0[14] ));
 sg13g2_a221oi_1 _2616_ (.B2(_1439_),
    .C1(_1527_),
    .B1(_1525_),
    .A1(_1518_),
    .Y(_1528_),
    .A2(_1519_));
 sg13g2_o21ai_1 _2617_ (.B1(_1528_),
    .Y(_1529_),
    .A1(_1463_),
    .A2(_1512_));
 sg13g2_xor2_1 _2618_ (.B(_1529_),
    .A(_1419_),
    .X(_1530_));
 sg13g2_nand2_1 _2619_ (.Y(_1531_),
    .A(_1445_),
    .B(_1437_));
 sg13g2_nor2_1 _2620_ (.A(_1448_),
    .B(_1456_),
    .Y(_1532_));
 sg13g2_inv_1 _2621_ (.Y(_1533_),
    .A(_1532_));
 sg13g2_nand2_1 _2622_ (.Y(_1534_),
    .A(_1502_),
    .B(_1503_));
 sg13g2_nand2_1 _2623_ (.Y(_1535_),
    .A(_1534_),
    .B(_1470_));
 sg13g2_nand2_1 _2624_ (.Y(_1536_),
    .A(_1483_),
    .B(_1462_));
 sg13g2_nor4_1 _2625_ (.A(_1477_),
    .B(_1479_),
    .C(_1506_),
    .D(_1536_),
    .Y(_1537_));
 sg13g2_a21oi_1 _2626_ (.A1(_1480_),
    .A2(_1472_),
    .Y(_1538_),
    .B1(_1477_));
 sg13g2_a21oi_1 _2627_ (.A1(_1462_),
    .A2(_1509_),
    .Y(_1539_),
    .B1(_1522_));
 sg13g2_o21ai_1 _2628_ (.B1(_1539_),
    .Y(_1540_),
    .A1(_1536_),
    .A2(_1538_));
 sg13g2_a21oi_1 _2629_ (.A1(_1535_),
    .A2(_1537_),
    .Y(_1541_),
    .B1(_1540_));
 sg13g2_nor2b_1 _2630_ (.A(_1541_),
    .B_N(_1459_),
    .Y(_1542_));
 sg13g2_inv_1 _2631_ (.Y(_1543_),
    .A(_1450_));
 sg13g2_o21ai_1 _2632_ (.B1(_1543_),
    .Y(_1544_),
    .A1(_1533_),
    .A2(_1542_));
 sg13g2_a21oi_1 _2633_ (.A1(_1437_),
    .A2(_1442_),
    .Y(_1545_),
    .B1(_1514_));
 sg13g2_o21ai_1 _2634_ (.B1(_1545_),
    .Y(_1546_),
    .A1(_1531_),
    .A2(_1544_));
 sg13g2_xor2_1 _2635_ (.B(_1546_),
    .A(_1435_),
    .X(_1547_));
 sg13g2_nand2_1 _2636_ (.Y(_1548_),
    .A(_1535_),
    .B(_1505_));
 sg13g2_nor2_1 _2637_ (.A(_1477_),
    .B(_1472_),
    .Y(_1549_));
 sg13g2_a21oi_1 _2638_ (.A1(_1548_),
    .A2(_1549_),
    .Y(_1550_),
    .B1(_1479_));
 sg13g2_nand2_1 _2639_ (.Y(_1551_),
    .A(_1451_),
    .B(_1459_));
 sg13g2_nor2_1 _2640_ (.A(_1536_),
    .B(_1551_),
    .Y(_1552_));
 sg13g2_nand2_1 _2641_ (.Y(_1553_),
    .A(_1431_),
    .B(_1435_));
 sg13g2_nor2_1 _2642_ (.A(_1531_),
    .B(_1553_),
    .Y(_1554_));
 sg13g2_nand3_1 _2643_ (.B(_1552_),
    .C(_1554_),
    .A(_1550_),
    .Y(_1555_));
 sg13g2_inv_1 _2644_ (.Y(_1556_),
    .A(_1545_));
 sg13g2_inv_1 _2645_ (.Y(_1557_),
    .A(_1553_));
 sg13g2_nand2_1 _2646_ (.Y(_1558_),
    .A(_1533_),
    .B(_1543_));
 sg13g2_o21ai_1 _2647_ (.B1(_1558_),
    .Y(_1559_),
    .A1(_1551_),
    .A2(_1539_));
 sg13g2_a21o_1 _2648_ (.A2(_1516_),
    .A1(_1431_),
    .B1(_1428_),
    .X(_1560_));
 sg13g2_a221oi_1 _2649_ (.B2(_1554_),
    .C1(_1560_),
    .B1(_1559_),
    .A1(_1556_),
    .Y(_1561_),
    .A2(_1557_));
 sg13g2_nand2_1 _2650_ (.Y(_1562_),
    .A(_1555_),
    .B(_1561_));
 sg13g2_xnor2_1 _2651_ (.Y(_1563_),
    .A(_1426_),
    .B(_1562_));
 sg13g2_nand2_1 _2652_ (.Y(_1564_),
    .A(_1459_),
    .B(_1462_));
 sg13g2_o21ai_1 _2653_ (.B1(_1523_),
    .Y(_1565_),
    .A1(_1564_),
    .A2(_1512_));
 sg13g2_inv_1 _2654_ (.Y(_1566_),
    .A(_1524_));
 sg13g2_a21oi_1 _2655_ (.A1(_1565_),
    .A2(_1453_),
    .Y(_1567_),
    .B1(_1566_));
 sg13g2_o21ai_1 _2656_ (.B1(_1517_),
    .Y(_1568_),
    .A1(_1438_),
    .A2(_1567_));
 sg13g2_xnor2_1 _2657_ (.Y(_1569_),
    .A(_1432_),
    .B(_1568_));
 sg13g2_nor4_2 _2658_ (.A(_1530_),
    .B(_1547_),
    .C(_1563_),
    .Y(_1570_),
    .D(_1569_));
 sg13g2_xnor2_1 _2659_ (.Y(_1571_),
    .A(_1445_),
    .B(_1544_));
 sg13g2_xnor2_1 _2660_ (.Y(_1572_),
    .A(_1437_),
    .B(_1567_));
 sg13g2_nor2_1 _2661_ (.A(_1571_),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_inv_1 _2662_ (.Y(_1574_),
    .A(\main._w_demo_video_hs ));
 sg13g2_nand2_1 _2663_ (.Y(_1575_),
    .A(_1574_),
    .B(\main.demo._q_prev_hs ));
 sg13g2_inv_1 _2664_ (.Y(_1576_),
    .A(_1575_));
 sg13g2_inv_1 _2665_ (.Y(_1577_),
    .A(\main.demo._q_pix_x[2] ));
 sg13g2_nand2_1 _2666_ (.Y(_1578_),
    .A(\main.demo._q_pix_x[1] ),
    .B(\main.demo._q_pix_x[0] ));
 sg13g2_nor2_1 _2667_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nor2_1 _2668_ (.A(\main.demo._q_pix_x[3] ),
    .B(_1579_),
    .Y(_1580_));
 sg13g2_inv_1 _2669_ (.Y(_1581_),
    .A(\main.demo._q_pix_x[3] ));
 sg13g2_inv_1 _2670_ (.Y(_1582_),
    .A(_1579_));
 sg13g2_nor2_1 _2671_ (.A(_1581_),
    .B(_1582_),
    .Y(_1583_));
 sg13g2_nor3_1 _2672_ (.A(net32),
    .B(_1580_),
    .C(_1583_),
    .Y(_1584_));
 sg13g2_xnor2_1 _2673_ (.Y(_1585_),
    .A(_1504_),
    .B(_1502_));
 sg13g2_xnor2_1 _2674_ (.Y(_1586_),
    .A(_1584_),
    .B(_1585_));
 sg13g2_xnor2_1 _2675_ (.Y(_1587_),
    .A(_1491_),
    .B(_1489_));
 sg13g2_nor2_1 _2676_ (.A(\main.demo._q_pix_x[0] ),
    .B(_1576_),
    .Y(_1588_));
 sg13g2_xor2_1 _2677_ (.B(_1588_),
    .A(_1587_),
    .X(_1589_));
 sg13g2_nor2b_1 _2678_ (.A(net32),
    .B_N(_1578_),
    .Y(_1590_));
 sg13g2_o21ai_1 _2679_ (.B1(_1590_),
    .Y(_1591_),
    .A1(\main.demo._q_pix_x[1] ),
    .A2(\main.demo._q_pix_x[0] ));
 sg13g2_xor2_1 _2680_ (.B(_1488_),
    .A(_1492_),
    .X(_1592_));
 sg13g2_xor2_1 _2681_ (.B(_1592_),
    .A(_1591_),
    .X(_1593_));
 sg13g2_nand2_1 _2682_ (.Y(_1594_),
    .A(_1578_),
    .B(_1577_));
 sg13g2_nand3_1 _2683_ (.B(_1575_),
    .C(_1594_),
    .A(_1582_),
    .Y(_1595_));
 sg13g2_inv_1 _2684_ (.Y(_1596_),
    .A(_1595_));
 sg13g2_nor2_1 _2685_ (.A(_1501_),
    .B(_1498_),
    .Y(_1597_));
 sg13g2_xnor2_1 _2686_ (.Y(_1598_),
    .A(_1597_),
    .B(_1495_));
 sg13g2_xnor2_1 _2687_ (.Y(_1599_),
    .A(_1596_),
    .B(_1598_));
 sg13g2_nand4_1 _2688_ (.B(_1589_),
    .C(_1593_),
    .A(_1586_),
    .Y(_1600_),
    .D(_1599_));
 sg13g2_inv_1 _2689_ (.Y(_1601_),
    .A(\main.demo._q_pix_x[6] ));
 sg13g2_inv_1 _2690_ (.Y(_1602_),
    .A(\main.demo._q_pix_x[5] ));
 sg13g2_inv_1 _2691_ (.Y(_1603_),
    .A(\main.demo._q_pix_x[4] ));
 sg13g2_inv_1 _2692_ (.Y(_1604_),
    .A(_1583_));
 sg13g2_nor2_1 _2693_ (.A(_1603_),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_inv_1 _2694_ (.Y(_1606_),
    .A(_1605_));
 sg13g2_nor2_1 _2695_ (.A(_1602_),
    .B(_1606_),
    .Y(_1607_));
 sg13g2_inv_1 _2696_ (.Y(_1608_),
    .A(_1607_));
 sg13g2_nor2_1 _2697_ (.A(_1601_),
    .B(_1608_),
    .Y(_1609_));
 sg13g2_inv_1 _2698_ (.Y(_1610_),
    .A(_1609_));
 sg13g2_inv_1 _2699_ (.Y(_1611_),
    .A(\main.demo._q_pix_x[7] ));
 sg13g2_a21oi_1 _2700_ (.A1(_1610_),
    .A2(_1611_),
    .Y(_1612_),
    .B1(net32));
 sg13g2_nor2_1 _2701_ (.A(_1611_),
    .B(_1610_),
    .Y(_1613_));
 sg13g2_inv_1 _2702_ (.Y(_1614_),
    .A(_1613_));
 sg13g2_nand2_1 _2703_ (.Y(_1615_),
    .A(_1612_),
    .B(_1614_));
 sg13g2_xnor2_1 _2704_ (.Y(_1616_),
    .A(_1462_),
    .B(_1512_));
 sg13g2_xnor2_1 _2705_ (.Y(_1617_),
    .A(_1615_),
    .B(_1616_));
 sg13g2_a21oi_1 _2706_ (.A1(_1608_),
    .A2(_1601_),
    .Y(_1618_),
    .B1(net32));
 sg13g2_nand2_1 _2707_ (.Y(_1619_),
    .A(_1618_),
    .B(_1610_));
 sg13g2_xor2_1 _2708_ (.B(_1550_),
    .A(_1483_),
    .X(_1620_));
 sg13g2_xnor2_1 _2709_ (.Y(_1621_),
    .A(_1619_),
    .B(_1620_));
 sg13g2_inv_1 _2710_ (.Y(_1622_),
    .A(_1535_));
 sg13g2_a21oi_1 _2711_ (.A1(_1622_),
    .A2(_1473_),
    .Y(_1623_),
    .B1(_1466_));
 sg13g2_xor2_1 _2712_ (.B(_1623_),
    .A(_1480_),
    .X(_1624_));
 sg13g2_nor2_1 _2713_ (.A(\main.demo._q_pix_x[5] ),
    .B(_1605_),
    .Y(_1625_));
 sg13g2_nor3_1 _2714_ (.A(net32),
    .B(_1625_),
    .C(_1607_),
    .Y(_1626_));
 sg13g2_nand2b_1 _2715_ (.Y(_1627_),
    .B(_1626_),
    .A_N(_1624_));
 sg13g2_inv_1 _2716_ (.Y(_1628_),
    .A(_1626_));
 sg13g2_nand2_1 _2717_ (.Y(_1629_),
    .A(_1624_),
    .B(_1628_));
 sg13g2_nor2_1 _2718_ (.A(\main.demo._q_pix_x[4] ),
    .B(_1583_),
    .Y(_1630_));
 sg13g2_nor3_2 _2719_ (.A(net32),
    .B(_1630_),
    .C(_1605_),
    .Y(_1631_));
 sg13g2_xnor2_1 _2720_ (.Y(_1632_),
    .A(_1506_),
    .B(_1535_));
 sg13g2_xnor2_1 _2721_ (.Y(_1633_),
    .A(_1631_),
    .B(_1632_));
 sg13g2_nand3_1 _2722_ (.B(_1629_),
    .C(_1633_),
    .A(_1627_),
    .Y(_1634_));
 sg13g2_nor4_1 _2723_ (.A(_1600_),
    .B(_1617_),
    .C(_1621_),
    .D(_1634_),
    .Y(_1635_));
 sg13g2_xnor2_1 _2724_ (.Y(_1636_),
    .A(_1459_),
    .B(_1541_));
 sg13g2_nor2b_1 _2725_ (.A(_1614_),
    .B_N(\main.demo._q_pix_x[8] ),
    .Y(_1637_));
 sg13g2_nor2_1 _2726_ (.A(net32),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_o21ai_1 _2727_ (.B1(_1638_),
    .Y(_1639_),
    .A1(\main.demo._q_pix_x[8] ),
    .A2(_1613_));
 sg13g2_xnor2_1 _2728_ (.Y(_1640_),
    .A(_1636_),
    .B(_1639_));
 sg13g2_a21oi_1 _2729_ (.A1(_1637_),
    .A2(\main.demo._q_pix_x[9] ),
    .Y(_1641_),
    .B1(net32));
 sg13g2_o21ai_1 _2730_ (.B1(_1641_),
    .Y(_1642_),
    .A1(\main.demo._q_pix_x[9] ),
    .A2(_1637_));
 sg13g2_xnor2_1 _2731_ (.Y(_1643_),
    .A(_1452_),
    .B(_1565_));
 sg13g2_xnor2_1 _2732_ (.Y(_1644_),
    .A(_1642_),
    .B(_1643_));
 sg13g2_nor2_1 _2733_ (.A(_1640_),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_nand4_1 _2734_ (.B(_1573_),
    .C(_1635_),
    .A(_1570_),
    .Y(_1646_),
    .D(_1645_));
 sg13g2_buf_1 _2735_ (.A(_1646_),
    .X(_1647_));
 sg13g2_nand3_1 _2736_ (.B(_1418_),
    .C(_1647_),
    .A(_1417_),
    .Y(_1648_));
 sg13g2_buf_8 _2737_ (.A(_1648_),
    .X(_1649_));
 sg13g2_buf_8 _2738_ (.A(_1649_),
    .X(_1650_));
 sg13g2_nand2_1 _2739_ (.Y(_1651_),
    .A(_1406_),
    .B(_1404_));
 sg13g2_nor2b_1 _2740_ (.A(_1381_),
    .B_N(_1388_),
    .Y(_1652_));
 sg13g2_a21oi_1 _2741_ (.A1(_1389_),
    .A2(_1380_),
    .Y(_1653_),
    .B1(_1652_));
 sg13g2_inv_1 _2742_ (.Y(_1654_),
    .A(_1382_));
 sg13g2_a22oi_1 _2743_ (.Y(_1655_),
    .B1(\main.demo._q_rand_0[10] ),
    .B2(_1386_),
    .A2(_1654_),
    .A1(_1189_));
 sg13g2_xor2_1 _2744_ (.B(_1300_),
    .A(\main.demo._q_rand_0[10] ),
    .X(_1656_));
 sg13g2_xnor2_1 _2745_ (.Y(_1657_),
    .A(\main.demo._q_rand_0[11] ),
    .B(_1384_));
 sg13g2_xnor2_1 _2746_ (.Y(_1658_),
    .A(_1656_),
    .B(_1657_));
 sg13g2_inv_1 _2747_ (.Y(_1659_),
    .A(_1392_));
 sg13g2_nor2_1 _2748_ (.A(_1200_),
    .B(_1335_),
    .Y(_1660_));
 sg13g2_a21oi_1 _2749_ (.A1(_1659_),
    .A2(_1391_),
    .Y(_1661_),
    .B1(_1660_));
 sg13g2_xnor2_1 _2750_ (.Y(_1662_),
    .A(_1658_),
    .B(_1661_));
 sg13g2_xnor2_1 _2751_ (.Y(_1663_),
    .A(_1655_),
    .B(_1662_));
 sg13g2_nor2_1 _2752_ (.A(_1328_),
    .B(_1180_),
    .Y(_1664_));
 sg13g2_xnor2_1 _2753_ (.Y(_1665_),
    .A(_1152_),
    .B(_1209_));
 sg13g2_xnor2_1 _2754_ (.Y(_1666_),
    .A(_1664_),
    .B(_1665_));
 sg13g2_xnor2_1 _2755_ (.Y(_1667_),
    .A(_1189_),
    .B(_1143_));
 sg13g2_xnor2_1 _2756_ (.Y(_1668_),
    .A(_1200_),
    .B(_1667_));
 sg13g2_xnor2_1 _2757_ (.Y(_1669_),
    .A(_1391_),
    .B(_1668_));
 sg13g2_xnor2_1 _2758_ (.Y(_1670_),
    .A(_1666_),
    .B(_1669_));
 sg13g2_o21ai_1 _2759_ (.B1(_1329_),
    .Y(_1671_),
    .A1(_1330_),
    .A2(_1393_));
 sg13g2_xnor2_1 _2760_ (.Y(_1672_),
    .A(_1670_),
    .B(_1671_));
 sg13g2_xnor2_1 _2761_ (.Y(_1673_),
    .A(_1663_),
    .B(_1672_));
 sg13g2_nand3_1 _2762_ (.B(_1399_),
    .C(_1390_),
    .A(_1398_),
    .Y(_1674_));
 sg13g2_nand2_1 _2763_ (.Y(_1675_),
    .A(_1674_),
    .B(_1399_));
 sg13g2_xnor2_1 _2764_ (.Y(_1676_),
    .A(_1673_),
    .B(_1675_));
 sg13g2_xor2_1 _2765_ (.B(_1676_),
    .A(_1653_),
    .X(_1677_));
 sg13g2_xnor2_1 _2766_ (.Y(_1678_),
    .A(_1651_),
    .B(_1677_));
 sg13g2_nand3_1 _2767_ (.B(_1414_),
    .C(_1678_),
    .A(_1417_),
    .Y(_1679_));
 sg13g2_nand2_1 _2768_ (.Y(_1680_),
    .A(_1679_),
    .B(_1647_));
 sg13g2_nand2_1 _2769_ (.Y(_1681_),
    .A(_1417_),
    .B(_1414_));
 sg13g2_nand2b_1 _2770_ (.Y(_1682_),
    .B(_1681_),
    .A_N(_1678_));
 sg13g2_nor2b_2 _2771_ (.A(_1680_),
    .B_N(_1682_),
    .Y(_1683_));
 sg13g2_buf_8 _2772_ (.A(_1683_),
    .X(_1684_));
 sg13g2_nor2_1 _2773_ (.A(net16),
    .B(net12),
    .Y(_1685_));
 sg13g2_nand4_1 _2774_ (.B(_1573_),
    .C(_1635_),
    .A(_1570_),
    .Y(_1686_),
    .D(_1645_));
 sg13g2_buf_1 _2775_ (.A(_1686_),
    .X(_1687_));
 sg13g2_inv_1 _2776_ (.Y(_1688_),
    .A(_1687_));
 sg13g2_nand2_1 _2777_ (.Y(_1689_),
    .A(_1417_),
    .B(_1418_));
 sg13g2_nor2_1 _2778_ (.A(_1688_),
    .B(_1689_),
    .Y(_1690_));
 sg13g2_buf_8 _2779_ (.A(_1690_),
    .X(_1691_));
 sg13g2_nand2_1 _2780_ (.Y(_1692_),
    .A(net15),
    .B(_1464_));
 sg13g2_nand2_1 _2781_ (.Y(_1693_),
    .A(_1649_),
    .B(_1467_));
 sg13g2_nand2_1 _2782_ (.Y(_1694_),
    .A(_1692_),
    .B(_1693_));
 sg13g2_nand3_1 _2783_ (.B(_1679_),
    .C(_1647_),
    .A(_1682_),
    .Y(_1695_));
 sg13g2_buf_1 _2784_ (.A(_1695_),
    .X(_1696_));
 sg13g2_nand2_1 _2785_ (.Y(_1697_),
    .A(_1694_),
    .B(net11));
 sg13g2_nand2_1 _2786_ (.Y(_1698_),
    .A(net15),
    .B(_1481_));
 sg13g2_nand2_1 _2787_ (.Y(_1699_),
    .A(net16),
    .B(_1475_));
 sg13g2_nand2_1 _2788_ (.Y(_1700_),
    .A(_1698_),
    .B(_1699_));
 sg13g2_nand2_1 _2789_ (.Y(_1701_),
    .A(_1700_),
    .B(net12));
 sg13g2_xnor2_1 _2790_ (.Y(_1702_),
    .A(_1261_),
    .B(_1267_));
 sg13g2_xnor2_1 _2791_ (.Y(_1703_),
    .A(_1157_),
    .B(_1702_));
 sg13g2_nand2_1 _2792_ (.Y(_1704_),
    .A(_1687_),
    .B(_1703_));
 sg13g2_a21oi_2 _2793_ (.B1(_1704_),
    .Y(_1705_),
    .A2(_1701_),
    .A1(_1697_));
 sg13g2_inv_1 _2794_ (.Y(_1706_),
    .A(_1705_));
 sg13g2_nand3_1 _2795_ (.B(_1697_),
    .C(_1704_),
    .A(_1701_),
    .Y(_1707_));
 sg13g2_nand2_1 _2796_ (.Y(_1708_),
    .A(_1706_),
    .B(_1707_));
 sg13g2_nand2_1 _2797_ (.Y(_1709_),
    .A(net15),
    .B(_1476_));
 sg13g2_nand2_1 _2798_ (.Y(_1710_),
    .A(_1649_),
    .B(_1471_));
 sg13g2_nand2_1 _2799_ (.Y(_1711_),
    .A(_1709_),
    .B(_1710_));
 sg13g2_nand2_1 _2800_ (.Y(_1712_),
    .A(_1711_),
    .B(net12));
 sg13g2_nand2_1 _2801_ (.Y(_1713_),
    .A(net15),
    .B(_1468_));
 sg13g2_nand2_1 _2802_ (.Y(_1714_),
    .A(_1649_),
    .B(_1497_));
 sg13g2_nand2_1 _2803_ (.Y(_1715_),
    .A(_1713_),
    .B(_1714_));
 sg13g2_nand2_1 _2804_ (.Y(_1716_),
    .A(_1715_),
    .B(net11));
 sg13g2_nor2_1 _2805_ (.A(_1227_),
    .B(_1688_),
    .Y(_1717_));
 sg13g2_nand3_1 _2806_ (.B(_1716_),
    .C(_1717_),
    .A(_1712_),
    .Y(_1718_));
 sg13g2_nand2_1 _2807_ (.Y(_1719_),
    .A(net15),
    .B(_1475_));
 sg13g2_nand2_1 _2808_ (.Y(_1720_),
    .A(net16),
    .B(_1464_));
 sg13g2_nand2_1 _2809_ (.Y(_1721_),
    .A(_1719_),
    .B(_1720_));
 sg13g2_nand2_1 _2810_ (.Y(_1722_),
    .A(_1721_),
    .B(net12));
 sg13g2_nand2_1 _2811_ (.Y(_1723_),
    .A(net16),
    .B(_1496_));
 sg13g2_nand4_1 _2812_ (.B(_1418_),
    .C(_1467_),
    .A(_1417_),
    .Y(_1724_),
    .D(_1647_));
 sg13g2_nand2_1 _2813_ (.Y(_1725_),
    .A(_1723_),
    .B(_1724_));
 sg13g2_nand2_1 _2814_ (.Y(_1726_),
    .A(_1725_),
    .B(net11));
 sg13g2_inv_1 _2815_ (.Y(_1727_),
    .A(_1717_));
 sg13g2_nand3_1 _2816_ (.B(_1726_),
    .C(_1727_),
    .A(_1722_),
    .Y(_1728_));
 sg13g2_nand2_1 _2817_ (.Y(_1729_),
    .A(_1718_),
    .B(_1728_));
 sg13g2_nand2_1 _2818_ (.Y(_1730_),
    .A(net15),
    .B(_1496_));
 sg13g2_nand2_1 _2819_ (.Y(_1731_),
    .A(_1649_),
    .B(_1486_));
 sg13g2_nand2_1 _2820_ (.Y(_1732_),
    .A(_1730_),
    .B(_1731_));
 sg13g2_nand2_1 _2821_ (.Y(_1733_),
    .A(_1732_),
    .B(net11));
 sg13g2_nand2_1 _2822_ (.Y(_1734_),
    .A(_1694_),
    .B(_1683_));
 sg13g2_nand2_1 _2823_ (.Y(_1735_),
    .A(_1733_),
    .B(_1734_));
 sg13g2_xnor2_1 _2824_ (.Y(_1736_),
    .A(_1328_),
    .B(_1198_));
 sg13g2_nand2_1 _2825_ (.Y(_1737_),
    .A(_1647_),
    .B(_1736_));
 sg13g2_inv_1 _2826_ (.Y(_1738_),
    .A(_1737_));
 sg13g2_nand2_1 _2827_ (.Y(_1739_),
    .A(_1735_),
    .B(_1738_));
 sg13g2_nand3_1 _2828_ (.B(_1734_),
    .C(_1737_),
    .A(_1733_),
    .Y(_1740_));
 sg13g2_nand2_1 _2829_ (.Y(_1741_),
    .A(_1739_),
    .B(_1740_));
 sg13g2_nor2_1 _2830_ (.A(_1729_),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_nor2_1 _2831_ (.A(_1165_),
    .B(_1688_),
    .Y(_1743_));
 sg13g2_nor2_1 _2832_ (.A(_1493_),
    .B(net16),
    .Y(_1744_));
 sg13g2_a21oi_1 _2833_ (.A1(_1489_),
    .A2(net16),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_nand2_1 _2834_ (.Y(_1746_),
    .A(_1745_),
    .B(net11));
 sg13g2_nand2_1 _2835_ (.Y(_1747_),
    .A(_1715_),
    .B(net12));
 sg13g2_nand3b_1 _2836_ (.B(_1746_),
    .C(_1747_),
    .Y(_1748_),
    .A_N(_1743_));
 sg13g2_inv_1 _2837_ (.Y(_1749_),
    .A(_1748_));
 sg13g2_nand2_1 _2838_ (.Y(_1750_),
    .A(_1742_),
    .B(_1749_));
 sg13g2_inv_1 _2839_ (.Y(_1751_),
    .A(_1739_));
 sg13g2_inv_1 _2840_ (.Y(_1752_),
    .A(_1718_));
 sg13g2_a21oi_1 _2841_ (.A1(_1751_),
    .A2(_1728_),
    .Y(_1753_),
    .B1(_1752_));
 sg13g2_nand2_1 _2842_ (.Y(_1754_),
    .A(_1750_),
    .B(_1753_));
 sg13g2_xnor2_1 _2843_ (.Y(_1755_),
    .A(_1708_),
    .B(_1754_));
 sg13g2_inv_1 _2844_ (.Y(_1756_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[3] ));
 sg13g2_inv_1 _2845_ (.Y(_1757_),
    .A(_1740_));
 sg13g2_o21ai_1 _2846_ (.B1(_1739_),
    .Y(_1758_),
    .A1(_1757_),
    .A2(_1748_));
 sg13g2_xnor2_1 _2847_ (.Y(_1759_),
    .A(_1729_),
    .B(_1758_));
 sg13g2_inv_1 _2848_ (.Y(_1760_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[2] ));
 sg13g2_nand2_1 _2849_ (.Y(_1761_),
    .A(_1759_),
    .B(_1760_));
 sg13g2_xnor2_1 _2850_ (.Y(_1762_),
    .A(_1749_),
    .B(_1741_));
 sg13g2_inv_1 _2851_ (.Y(_1763_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[1] ));
 sg13g2_nand2_1 _2852_ (.Y(_1764_),
    .A(_1746_),
    .B(_1747_));
 sg13g2_nand2_1 _2853_ (.Y(_1765_),
    .A(_1764_),
    .B(_1743_));
 sg13g2_nand2_1 _2854_ (.Y(_1766_),
    .A(_1748_),
    .B(_1765_));
 sg13g2_xnor2_1 _2855_ (.Y(_1767_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[0] ),
    .B(_1766_));
 sg13g2_a21oi_1 _2856_ (.A1(_1762_),
    .A2(_1763_),
    .Y(_1768_),
    .B1(_1767_));
 sg13g2_nand2_1 _2857_ (.Y(_1769_),
    .A(_1761_),
    .B(_1768_));
 sg13g2_a21oi_1 _2858_ (.A1(_1755_),
    .A2(_1756_),
    .Y(_1770_),
    .B1(_1769_));
 sg13g2_nand2b_1 _2859_ (.Y(_1771_),
    .B(\main.demo._d___pip_24_1_1___stage___block_3_y[1] ),
    .A_N(_1762_));
 sg13g2_o21ai_1 _2860_ (.B1(_1771_),
    .Y(_1772_),
    .A1(_1760_),
    .A2(_1759_));
 sg13g2_nor2_1 _2861_ (.A(_1756_),
    .B(_1755_),
    .Y(_1773_));
 sg13g2_nor2_1 _2862_ (.A(_1772_),
    .B(_1773_),
    .Y(_1774_));
 sg13g2_nand2_1 _2863_ (.Y(_1775_),
    .A(_1770_),
    .B(_1774_));
 sg13g2_nor2b_1 _2864_ (.A(_1285_),
    .B_N(_1284_),
    .Y(_1776_));
 sg13g2_xnor2_1 _2865_ (.Y(_1777_),
    .A(_1278_),
    .B(_1776_));
 sg13g2_nor2_1 _2866_ (.A(_1777_),
    .B(_1688_),
    .Y(_1778_));
 sg13g2_inv_1 _2867_ (.Y(_1779_),
    .A(_1778_));
 sg13g2_nand2_1 _2868_ (.Y(_1780_),
    .A(_1649_),
    .B(_1508_));
 sg13g2_nand2_1 _2869_ (.Y(_1781_),
    .A(net15),
    .B(_1521_));
 sg13g2_nand3_1 _2870_ (.B(_1780_),
    .C(_1781_),
    .A(net11),
    .Y(_1782_));
 sg13g2_inv_1 _2871_ (.Y(_1783_),
    .A(_0002_));
 sg13g2_nor2_1 _2872_ (.A(_1783_),
    .B(net16),
    .Y(_1784_));
 sg13g2_a21oi_1 _2873_ (.A1(_0001_),
    .A2(net16),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_nand2_1 _2874_ (.Y(_1786_),
    .A(_1785_),
    .B(_1684_));
 sg13g2_nand2_1 _2875_ (.Y(_1787_),
    .A(_1782_),
    .B(_1786_));
 sg13g2_xnor2_1 _2876_ (.Y(_1788_),
    .A(_1779_),
    .B(_1787_));
 sg13g2_xnor2_1 _2877_ (.Y(_1789_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[6] ),
    .B(_1788_));
 sg13g2_a21oi_1 _2878_ (.A1(_1752_),
    .A2(_1707_),
    .Y(_1790_),
    .B1(_1705_));
 sg13g2_nand2_1 _2879_ (.Y(_1791_),
    .A(_1781_),
    .B(_1780_));
 sg13g2_nand2_1 _2880_ (.Y(_1792_),
    .A(_1791_),
    .B(_1683_));
 sg13g2_nand2_1 _2881_ (.Y(_1793_),
    .A(_1711_),
    .B(net11));
 sg13g2_nand2_1 _2882_ (.Y(_1794_),
    .A(_1792_),
    .B(_1793_));
 sg13g2_nor2b_1 _2883_ (.A(_1273_),
    .B_N(_1272_),
    .Y(_1795_));
 sg13g2_xor2_1 _2884_ (.B(_1795_),
    .A(_1269_),
    .X(_1796_));
 sg13g2_nand2_1 _2885_ (.Y(_1797_),
    .A(_1687_),
    .B(_1796_));
 sg13g2_nand2_1 _2886_ (.Y(_1798_),
    .A(_1794_),
    .B(_1797_));
 sg13g2_inv_1 _2887_ (.Y(_1799_),
    .A(_1797_));
 sg13g2_nand3_1 _2888_ (.B(_1793_),
    .C(_1799_),
    .A(_1792_),
    .Y(_1800_));
 sg13g2_nand2_1 _2889_ (.Y(_1801_),
    .A(_1798_),
    .B(_1800_));
 sg13g2_inv_2 _2890_ (.Y(_1802_),
    .A(_1801_));
 sg13g2_nor2b_1 _2891_ (.A(_1276_),
    .B_N(_1260_),
    .Y(_1803_));
 sg13g2_xnor2_1 _2892_ (.Y(_1804_),
    .A(_1275_),
    .B(_1803_));
 sg13g2_nor2_1 _2893_ (.A(_1804_),
    .B(_1688_),
    .Y(_1805_));
 sg13g2_inv_1 _2894_ (.Y(_1806_),
    .A(_1805_));
 sg13g2_inv_1 _2895_ (.Y(_1807_),
    .A(_0001_));
 sg13g2_nand2_1 _2896_ (.Y(_1808_),
    .A(net15),
    .B(_1807_));
 sg13g2_inv_1 _2897_ (.Y(_1809_),
    .A(_0000_));
 sg13g2_nand2_1 _2898_ (.Y(_1810_),
    .A(_1650_),
    .B(_1809_));
 sg13g2_nand2_1 _2899_ (.Y(_1811_),
    .A(_1808_),
    .B(_1810_));
 sg13g2_nand2_1 _2900_ (.Y(_1812_),
    .A(_1811_),
    .B(_1684_));
 sg13g2_nand2_1 _2901_ (.Y(_1813_),
    .A(_1700_),
    .B(_1696_));
 sg13g2_nand2_1 _2902_ (.Y(_1814_),
    .A(_1812_),
    .B(_1813_));
 sg13g2_xnor2_1 _2903_ (.Y(_1815_),
    .A(_1806_),
    .B(_1814_));
 sg13g2_nand2_1 _2904_ (.Y(_1816_),
    .A(_1802_),
    .B(_1815_));
 sg13g2_nor2_1 _2905_ (.A(_1790_),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_xnor2_1 _2906_ (.Y(_1818_),
    .A(_1805_),
    .B(_1814_));
 sg13g2_nand2_1 _2907_ (.Y(_1819_),
    .A(_1814_),
    .B(_1805_));
 sg13g2_o21ai_1 _2908_ (.B1(_1819_),
    .Y(_1820_),
    .A1(_1800_),
    .A2(_1818_));
 sg13g2_nor2_1 _2909_ (.A(_1817_),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_nor2_1 _2910_ (.A(_1729_),
    .B(_1708_),
    .Y(_1822_));
 sg13g2_nor2_1 _2911_ (.A(_1801_),
    .B(_1818_),
    .Y(_1823_));
 sg13g2_nand3_1 _2912_ (.B(_1822_),
    .C(_1823_),
    .A(_1758_),
    .Y(_1824_));
 sg13g2_nand2_1 _2913_ (.Y(_1825_),
    .A(_1821_),
    .B(_1824_));
 sg13g2_xnor2_1 _2914_ (.Y(_1826_),
    .A(_1789_),
    .B(_1825_));
 sg13g2_nor2b_1 _2915_ (.A(_1239_),
    .B_N(_1287_),
    .Y(_1827_));
 sg13g2_xnor2_1 _2916_ (.Y(_1828_),
    .A(_1286_),
    .B(_1827_));
 sg13g2_nand2_1 _2917_ (.Y(_1829_),
    .A(_1687_),
    .B(_1828_));
 sg13g2_xor2_1 _2918_ (.B(_1829_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[7] ),
    .X(_1830_));
 sg13g2_nor2_1 _2919_ (.A(_1783_),
    .B(_1691_),
    .Y(_1831_));
 sg13g2_a21oi_1 _2920_ (.A1(_0003_),
    .A2(_1691_),
    .Y(_1832_),
    .B1(_1831_));
 sg13g2_a21oi_1 _2921_ (.A1(_1810_),
    .A2(_1808_),
    .Y(_1833_),
    .B1(net12));
 sg13g2_a21oi_1 _2922_ (.A1(net12),
    .A2(_1832_),
    .Y(_1834_),
    .B1(_1833_));
 sg13g2_xor2_1 _2923_ (.B(_1834_),
    .A(_1830_),
    .X(_1835_));
 sg13g2_nor2b_1 _2924_ (.A(_1705_),
    .B_N(_1707_),
    .Y(_1836_));
 sg13g2_nand2_1 _2925_ (.Y(_1837_),
    .A(_1836_),
    .B(_1802_));
 sg13g2_nand2_1 _2926_ (.Y(_1838_),
    .A(_1788_),
    .B(_1815_));
 sg13g2_nor2_1 _2927_ (.A(_1837_),
    .B(_1838_),
    .Y(_1839_));
 sg13g2_nand2_1 _2928_ (.Y(_1840_),
    .A(_1754_),
    .B(_1839_));
 sg13g2_nor2_1 _2929_ (.A(_1778_),
    .B(_1787_),
    .Y(_1841_));
 sg13g2_nand2_1 _2930_ (.Y(_1842_),
    .A(_1787_),
    .B(_1778_));
 sg13g2_o21ai_1 _2931_ (.B1(_1842_),
    .Y(_1843_),
    .A1(_1819_),
    .A2(_1841_));
 sg13g2_nand2_1 _2932_ (.Y(_1844_),
    .A(_1705_),
    .B(_1798_));
 sg13g2_nand2_1 _2933_ (.Y(_1845_),
    .A(_1844_),
    .B(_1800_));
 sg13g2_nor2b_1 _2934_ (.A(_1838_),
    .B_N(_1845_),
    .Y(_1846_));
 sg13g2_nor2_1 _2935_ (.A(_1843_),
    .B(_1846_),
    .Y(_1847_));
 sg13g2_nand2_1 _2936_ (.Y(_1848_),
    .A(_1840_),
    .B(_1847_));
 sg13g2_nand2b_1 _2937_ (.Y(_1849_),
    .B(_1848_),
    .A_N(_1835_));
 sg13g2_nand3_1 _2938_ (.B(_1847_),
    .C(_1835_),
    .A(_1840_),
    .Y(_1850_));
 sg13g2_nand2_1 _2939_ (.Y(_1851_),
    .A(_1849_),
    .B(_1850_));
 sg13g2_nor2_1 _2940_ (.A(_1826_),
    .B(_1851_),
    .Y(_1852_));
 sg13g2_nand4_1 _2941_ (.B(_1749_),
    .C(_1836_),
    .A(_1742_),
    .Y(_1853_),
    .D(_1802_));
 sg13g2_nor2_1 _2942_ (.A(_1753_),
    .B(_1837_),
    .Y(_1854_));
 sg13g2_nor2_1 _2943_ (.A(_1845_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_nand2_1 _2944_ (.Y(_1856_),
    .A(_1853_),
    .B(_1855_));
 sg13g2_xnor2_1 _2945_ (.Y(_1857_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[5] ),
    .B(_1818_));
 sg13g2_nand2_1 _2946_ (.Y(_1858_),
    .A(_1856_),
    .B(_1857_));
 sg13g2_inv_1 _2947_ (.Y(_1859_),
    .A(_1857_));
 sg13g2_nand3_1 _2948_ (.B(_1855_),
    .C(_1859_),
    .A(_1853_),
    .Y(_1860_));
 sg13g2_xor2_1 _2949_ (.B(_1801_),
    .A(\main.demo._d___pip_24_1_1___stage___block_3_y[4] ),
    .X(_1861_));
 sg13g2_nand2_1 _2950_ (.Y(_1862_),
    .A(_1758_),
    .B(_1822_));
 sg13g2_nand2_1 _2951_ (.Y(_1863_),
    .A(_1862_),
    .B(_1790_));
 sg13g2_xnor2_1 _2952_ (.Y(_1864_),
    .A(_1861_),
    .B(_1863_));
 sg13g2_a21oi_1 _2953_ (.A1(_1858_),
    .A2(_1860_),
    .Y(_1865_),
    .B1(_1864_));
 sg13g2_nand2_1 _2954_ (.Y(_1866_),
    .A(_1852_),
    .B(_1865_));
 sg13g2_nor3_1 _2955_ (.A(_1685_),
    .B(_1775_),
    .C(_1866_),
    .Y(_0020_));
 sg13g2_nor3_1 _2956_ (.A(net12),
    .B(_1775_),
    .C(_1866_),
    .Y(_0021_));
 sg13g2_inv_1 _2957_ (.Y(_1867_),
    .A(_1323_));
 sg13g2_nor2_1 _2958_ (.A(_1322_),
    .B(_1288_),
    .Y(_1868_));
 sg13g2_inv_1 _2959_ (.Y(_1869_),
    .A(_0004_));
 sg13g2_nand2_1 _2960_ (.Y(_0139_),
    .A(_1647_),
    .B(_1869_));
 sg13g2_nor3_1 _2961_ (.A(_1867_),
    .B(_1868_),
    .C(_0139_),
    .Y(_0092_));
 sg13g2_xnor2_1 _2962_ (.Y(_0140_),
    .A(_1371_),
    .B(_1324_));
 sg13g2_nor2_1 _2963_ (.A(_0140_),
    .B(_0139_),
    .Y(_0093_));
 sg13g2_buf_8 _2964_ (.A(\main.demo._q_rand_1[1] ),
    .X(_0141_));
 sg13g2_buf_8 _2965_ (.A(\main.demo._q_rand_1[0] ),
    .X(_0142_));
 sg13g2_nand2_2 _2966_ (.Y(_0143_),
    .A(net38),
    .B(_0142_));
 sg13g2_buf_8 _2967_ (.A(\main.demo._q_rand_1[3] ),
    .X(_0144_));
 sg13g2_buf_1 _2968_ (.A(\main.demo._q_rand_1[2] ),
    .X(_0145_));
 sg13g2_xnor2_1 _2969_ (.Y(_0146_),
    .A(net37),
    .B(net36));
 sg13g2_xnor2_1 _2970_ (.Y(_0147_),
    .A(_0143_),
    .B(_0146_));
 sg13g2_buf_8 _2971_ (.A(\main.demo._q_rand_1[4] ),
    .X(_0148_));
 sg13g2_nand2_2 _2972_ (.Y(_0149_),
    .A(net36),
    .B(_0148_));
 sg13g2_buf_2 _2973_ (.A(\main.demo._q_rand_1[6] ),
    .X(_0150_));
 sg13g2_buf_2 _2974_ (.A(\main.demo._q_rand_1[5] ),
    .X(_0151_));
 sg13g2_xnor2_1 _2975_ (.Y(_0152_),
    .A(_0150_),
    .B(_0151_));
 sg13g2_xor2_1 _2976_ (.B(_0152_),
    .A(_0149_),
    .X(_0153_));
 sg13g2_inv_1 _2977_ (.Y(_0154_),
    .A(net36));
 sg13g2_inv_2 _2978_ (.Y(_0155_),
    .A(_0148_));
 sg13g2_nand2_1 _2979_ (.Y(_0156_),
    .A(_0154_),
    .B(_0155_));
 sg13g2_nand2_1 _2980_ (.Y(_0157_),
    .A(_0156_),
    .B(_0149_));
 sg13g2_nand2_1 _2981_ (.Y(_0158_),
    .A(net38),
    .B(net37));
 sg13g2_nand2_1 _2982_ (.Y(_0159_),
    .A(_0157_),
    .B(_0158_));
 sg13g2_nand3b_1 _2983_ (.B(_0156_),
    .C(_0149_),
    .Y(_0160_),
    .A_N(_0158_));
 sg13g2_inv_1 _2984_ (.Y(_0161_),
    .A(_0160_));
 sg13g2_a21oi_1 _2985_ (.A1(_0159_),
    .A2(_0151_),
    .Y(_0162_),
    .B1(_0161_));
 sg13g2_xnor2_1 _2986_ (.Y(_0163_),
    .A(_0153_),
    .B(_0162_));
 sg13g2_xor2_1 _2987_ (.B(_0163_),
    .A(_0147_),
    .X(_0164_));
 sg13g2_xnor2_1 _2988_ (.Y(_0165_),
    .A(net38),
    .B(net37));
 sg13g2_nand2_1 _2989_ (.Y(_0166_),
    .A(_0142_),
    .B(net36));
 sg13g2_nand2_1 _2990_ (.Y(_0167_),
    .A(_0165_),
    .B(_0166_));
 sg13g2_nor2_1 _2991_ (.A(_0166_),
    .B(_0165_),
    .Y(_0168_));
 sg13g2_a21oi_1 _2992_ (.A1(_0167_),
    .A2(_0148_),
    .Y(_0169_),
    .B1(_0168_));
 sg13g2_nand2_1 _2993_ (.Y(_0170_),
    .A(_0160_),
    .B(_0159_));
 sg13g2_xnor2_1 _2994_ (.Y(_0171_),
    .A(_0151_),
    .B(_0170_));
 sg13g2_xnor2_1 _2995_ (.Y(_0172_),
    .A(_0169_),
    .B(_0171_));
 sg13g2_inv_2 _2996_ (.Y(_0173_),
    .A(_0141_));
 sg13g2_nand2_1 _2997_ (.Y(_0174_),
    .A(_0172_),
    .B(_0173_));
 sg13g2_inv_1 _2998_ (.Y(_0175_),
    .A(_0014_));
 sg13g2_nand2_1 _2999_ (.Y(_0176_),
    .A(_0175_),
    .B(net38));
 sg13g2_nand3_1 _3000_ (.B(_0174_),
    .C(_0176_),
    .A(_0164_),
    .Y(_0177_));
 sg13g2_nand2_1 _3001_ (.Y(_0178_),
    .A(_0174_),
    .B(_0176_));
 sg13g2_inv_1 _3002_ (.Y(_0179_),
    .A(_0164_));
 sg13g2_nand2_1 _3003_ (.Y(_0180_),
    .A(_0178_),
    .B(_0179_));
 sg13g2_nand2_1 _3004_ (.Y(_0181_),
    .A(_0177_),
    .B(_0180_));
 sg13g2_inv_1 _3005_ (.Y(_0182_),
    .A(_0169_));
 sg13g2_nand2_1 _3006_ (.Y(_0183_),
    .A(_0171_),
    .B(_0182_));
 sg13g2_nand2_1 _3007_ (.Y(_0184_),
    .A(_0181_),
    .B(_0183_));
 sg13g2_inv_1 _3008_ (.Y(_0185_),
    .A(_0183_));
 sg13g2_nand3_1 _3009_ (.B(_0180_),
    .C(_0185_),
    .A(_0177_),
    .Y(_0186_));
 sg13g2_nand2_1 _3010_ (.Y(_0187_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_nand2b_1 _3011_ (.Y(_0188_),
    .B(net38),
    .A_N(_0172_));
 sg13g2_nand2_1 _3012_ (.Y(_0189_),
    .A(_0188_),
    .B(_0174_));
 sg13g2_inv_4 _3013_ (.A(_0144_),
    .Y(_0190_));
 sg13g2_nor2_1 _3014_ (.A(_0142_),
    .B(net36),
    .Y(_0191_));
 sg13g2_inv_1 _3015_ (.Y(_0192_),
    .A(_0166_));
 sg13g2_nor2_1 _3016_ (.A(_0191_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_inv_1 _3017_ (.Y(_0194_),
    .A(_0193_));
 sg13g2_nor2_1 _3018_ (.A(_0190_),
    .B(_0194_),
    .Y(_0195_));
 sg13g2_nor2b_1 _3019_ (.A(_0168_),
    .B_N(_0167_),
    .Y(_0196_));
 sg13g2_xnor2_1 _3020_ (.Y(_0197_),
    .A(_0155_),
    .B(_0196_));
 sg13g2_xnor2_1 _3021_ (.Y(_0198_),
    .A(_0195_),
    .B(_0197_));
 sg13g2_nand2_1 _3022_ (.Y(_0199_),
    .A(_0197_),
    .B(_0195_));
 sg13g2_o21ai_1 _3023_ (.B1(_0199_),
    .Y(_0200_),
    .A1(_0175_),
    .A2(_0198_));
 sg13g2_nand2b_1 _3024_ (.Y(_0201_),
    .B(_0200_),
    .A_N(_0189_));
 sg13g2_nand2_1 _3025_ (.Y(_0202_),
    .A(_0187_),
    .B(_0201_));
 sg13g2_xor2_1 _3026_ (.B(_0200_),
    .A(_0189_),
    .X(_0203_));
 sg13g2_xnor2_1 _3027_ (.Y(_0204_),
    .A(_0142_),
    .B(_0198_));
 sg13g2_inv_1 _3028_ (.Y(_0205_),
    .A(_0195_));
 sg13g2_nand2_1 _3029_ (.Y(_0206_),
    .A(_0194_),
    .B(_0190_));
 sg13g2_nor2_1 _3030_ (.A(_0173_),
    .B(_0191_),
    .Y(_0207_));
 sg13g2_a21oi_1 _3031_ (.A1(_0205_),
    .A2(_0206_),
    .Y(_0208_),
    .B1(_0207_));
 sg13g2_nand2_1 _3032_ (.Y(_0209_),
    .A(_0204_),
    .B(_0208_));
 sg13g2_nor2_1 _3033_ (.A(net38),
    .B(net36),
    .Y(_0210_));
 sg13g2_a21oi_1 _3034_ (.A1(_0207_),
    .A2(_0166_),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_inv_1 _3035_ (.Y(_0212_),
    .A(_0211_));
 sg13g2_and3_1 _3036_ (.X(_0213_),
    .A(_0205_),
    .B(_0206_),
    .C(_0207_));
 sg13g2_nor2_1 _3037_ (.A(_0208_),
    .B(_0213_),
    .Y(_0214_));
 sg13g2_nor2_1 _3038_ (.A(_0212_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor2_1 _3039_ (.A(_0208_),
    .B(_0204_),
    .Y(_0216_));
 sg13g2_a21oi_1 _3040_ (.A1(_0209_),
    .A2(_0215_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_nor2_1 _3041_ (.A(_0203_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_nor2_1 _3042_ (.A(_0201_),
    .B(_0187_),
    .Y(_0219_));
 sg13g2_a21oi_1 _3043_ (.A1(_0202_),
    .A2(_0218_),
    .Y(_0220_),
    .B1(_0219_));
 sg13g2_nor2b_1 _3044_ (.A(_0162_),
    .B_N(_0153_),
    .Y(_0221_));
 sg13g2_nor2_1 _3045_ (.A(_0149_),
    .B(_0152_),
    .Y(_0222_));
 sg13g2_inv_1 _3046_ (.Y(_0223_),
    .A(_0146_));
 sg13g2_nor2_1 _3047_ (.A(_0143_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_inv_1 _3048_ (.Y(_0225_),
    .A(_0150_));
 sg13g2_inv_1 _3049_ (.Y(_0226_),
    .A(_0151_));
 sg13g2_buf_1 _3050_ (.A(\main.demo._q_rand_1[7] ),
    .X(_0227_));
 sg13g2_xnor2_1 _3051_ (.Y(_0228_),
    .A(_0150_),
    .B(net35));
 sg13g2_o21ai_1 _3052_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_nor3_1 _3053_ (.A(net35),
    .B(_0225_),
    .C(_0226_),
    .Y(_0230_));
 sg13g2_inv_1 _3054_ (.Y(_0231_),
    .A(_0230_));
 sg13g2_nand2_1 _3055_ (.Y(_0232_),
    .A(_0229_),
    .B(_0231_));
 sg13g2_xnor2_1 _3056_ (.Y(_0233_),
    .A(_0224_),
    .B(_0232_));
 sg13g2_xor2_1 _3057_ (.B(_0233_),
    .A(_0222_),
    .X(_0234_));
 sg13g2_inv_1 _3058_ (.Y(_0235_),
    .A(_0142_));
 sg13g2_nor2_1 _3059_ (.A(_0235_),
    .B(_0146_),
    .Y(_0236_));
 sg13g2_nand2_1 _3060_ (.Y(_0237_),
    .A(net38),
    .B(_0145_));
 sg13g2_o21ai_1 _3061_ (.B1(_0237_),
    .Y(_0238_),
    .A1(_0190_),
    .A2(_0210_));
 sg13g2_xnor2_1 _3062_ (.Y(_0239_),
    .A(_0148_),
    .B(_0146_));
 sg13g2_inv_1 _3063_ (.Y(_0240_),
    .A(_0239_));
 sg13g2_nand2b_1 _3064_ (.Y(_0241_),
    .B(_0240_),
    .A_N(_0238_));
 sg13g2_nand2_2 _3065_ (.Y(_0242_),
    .A(_0239_),
    .B(_0238_));
 sg13g2_nand2_1 _3066_ (.Y(_0243_),
    .A(_0241_),
    .B(_0242_));
 sg13g2_xor2_1 _3067_ (.B(_0142_),
    .A(net38),
    .X(_0244_));
 sg13g2_inv_1 _3068_ (.Y(_0245_),
    .A(_0244_));
 sg13g2_nand2_1 _3069_ (.Y(_0246_),
    .A(_0243_),
    .B(_0245_));
 sg13g2_nand3_1 _3070_ (.B(_0242_),
    .C(_0244_),
    .A(_0241_),
    .Y(_0247_));
 sg13g2_buf_8 _3071_ (.A(_0247_),
    .X(_0248_));
 sg13g2_nand2_1 _3072_ (.Y(_0249_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_nand2b_1 _3073_ (.Y(_0250_),
    .B(_0249_),
    .A_N(_0236_));
 sg13g2_nand3_1 _3074_ (.B(_0248_),
    .C(_0236_),
    .A(_0246_),
    .Y(_0251_));
 sg13g2_nand2_1 _3075_ (.Y(_0252_),
    .A(_0250_),
    .B(_0251_));
 sg13g2_nand2b_1 _3076_ (.Y(_0253_),
    .B(_0252_),
    .A_N(_0234_));
 sg13g2_nand3_1 _3077_ (.B(_0251_),
    .C(_0234_),
    .A(_0250_),
    .Y(_0254_));
 sg13g2_nand2_1 _3078_ (.Y(_0255_),
    .A(_0253_),
    .B(_0254_));
 sg13g2_nor2_1 _3079_ (.A(_0223_),
    .B(_0245_),
    .Y(_0256_));
 sg13g2_nand2b_1 _3080_ (.Y(_0257_),
    .B(_0163_),
    .A_N(_0147_));
 sg13g2_nor2b_1 _3081_ (.A(_0256_),
    .B_N(_0257_),
    .Y(_0258_));
 sg13g2_nand2_1 _3082_ (.Y(_0259_),
    .A(_0255_),
    .B(_0258_));
 sg13g2_inv_1 _3083_ (.Y(_0260_),
    .A(_0258_));
 sg13g2_nand3_1 _3084_ (.B(_0254_),
    .C(_0260_),
    .A(_0253_),
    .Y(_0261_));
 sg13g2_nand2_1 _3085_ (.Y(_0262_),
    .A(_0259_),
    .B(_0261_));
 sg13g2_nand2b_1 _3086_ (.Y(_0263_),
    .B(_0262_),
    .A_N(_0221_));
 sg13g2_nand3_1 _3087_ (.B(_0261_),
    .C(_0221_),
    .A(_0259_),
    .Y(_0264_));
 sg13g2_nand2_1 _3088_ (.Y(_0265_),
    .A(_0186_),
    .B(_0180_));
 sg13g2_nand3_1 _3089_ (.B(_0264_),
    .C(_0265_),
    .A(_0263_),
    .Y(_0266_));
 sg13g2_nand2_1 _3090_ (.Y(_0267_),
    .A(_0220_),
    .B(_0266_));
 sg13g2_a21o_1 _3091_ (.A2(_0264_),
    .A1(_0263_),
    .B1(_0265_),
    .X(_0268_));
 sg13g2_inv_1 _3092_ (.Y(_0269_),
    .A(_0224_));
 sg13g2_nand2_1 _3093_ (.Y(_0270_),
    .A(_0233_),
    .B(_0222_));
 sg13g2_o21ai_1 _3094_ (.B1(_0270_),
    .Y(_0271_),
    .A1(_0269_),
    .A2(_0232_));
 sg13g2_inv_1 _3095_ (.Y(_0272_),
    .A(_0251_));
 sg13g2_a21oi_1 _3096_ (.A1(_0250_),
    .A2(_0234_),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_nand2_1 _3097_ (.Y(_0274_),
    .A(_0190_),
    .B(_0155_));
 sg13g2_nand2_1 _3098_ (.Y(_0275_),
    .A(net37),
    .B(_0148_));
 sg13g2_nand2_1 _3099_ (.Y(_0276_),
    .A(_0274_),
    .B(_0275_));
 sg13g2_nand2_1 _3100_ (.Y(_0277_),
    .A(_0276_),
    .B(_0226_));
 sg13g2_nand3_1 _3101_ (.B(_0151_),
    .C(_0275_),
    .A(_0274_),
    .Y(_0278_));
 sg13g2_buf_1 _3102_ (.A(_0278_),
    .X(_0279_));
 sg13g2_nand2_2 _3103_ (.Y(_0280_),
    .A(_0277_),
    .B(_0279_));
 sg13g2_nand2_1 _3104_ (.Y(_0281_),
    .A(_0280_),
    .B(_0143_));
 sg13g2_inv_1 _3105_ (.Y(_0282_),
    .A(_0143_));
 sg13g2_nand3_1 _3106_ (.B(_0279_),
    .C(_0282_),
    .A(_0277_),
    .Y(_0283_));
 sg13g2_nand2_1 _3107_ (.Y(_0284_),
    .A(net37),
    .B(net36));
 sg13g2_o21ai_1 _3108_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0155_),
    .A2(_0146_));
 sg13g2_nand3_1 _3109_ (.B(_0283_),
    .C(_0285_),
    .A(_0281_),
    .Y(_0286_));
 sg13g2_nand2_1 _3110_ (.Y(_0287_),
    .A(_0280_),
    .B(_0282_));
 sg13g2_nand3_1 _3111_ (.B(_0279_),
    .C(_0143_),
    .A(_0277_),
    .Y(_0288_));
 sg13g2_inv_1 _3112_ (.Y(_0289_),
    .A(_0285_));
 sg13g2_nand3_1 _3113_ (.B(_0288_),
    .C(_0289_),
    .A(_0287_),
    .Y(_0290_));
 sg13g2_nand2_1 _3114_ (.Y(_0291_),
    .A(_0286_),
    .B(_0290_));
 sg13g2_xnor2_1 _3115_ (.Y(_0292_),
    .A(net36),
    .B(_0244_));
 sg13g2_nand2_1 _3116_ (.Y(_0293_),
    .A(_0291_),
    .B(_0292_));
 sg13g2_inv_1 _3117_ (.Y(_0294_),
    .A(_0292_));
 sg13g2_nand3_1 _3118_ (.B(_0290_),
    .C(_0294_),
    .A(_0286_),
    .Y(_0295_));
 sg13g2_nand2_1 _3119_ (.Y(_0296_),
    .A(_0293_),
    .B(_0295_));
 sg13g2_nand2_1 _3120_ (.Y(_0297_),
    .A(_0296_),
    .B(_0248_));
 sg13g2_inv_2 _3121_ (.Y(_0298_),
    .A(_0248_));
 sg13g2_nand3_1 _3122_ (.B(_0295_),
    .C(_0298_),
    .A(_0293_),
    .Y(_0299_));
 sg13g2_buf_1 _3123_ (.A(_0299_),
    .X(_0300_));
 sg13g2_nand2_1 _3124_ (.Y(_0301_),
    .A(_0297_),
    .B(_0300_));
 sg13g2_buf_1 _3125_ (.A(\main.demo._q_rand_1[8] ),
    .X(_0302_));
 sg13g2_inv_1 _3126_ (.Y(_0303_),
    .A(_0302_));
 sg13g2_xnor2_1 _3127_ (.Y(_0304_),
    .A(_0150_),
    .B(_0302_));
 sg13g2_nand2_1 _3128_ (.Y(_0305_),
    .A(_0304_),
    .B(net35));
 sg13g2_o21ai_1 _3129_ (.B1(_0305_),
    .Y(_0306_),
    .A1(net35),
    .A2(_0303_));
 sg13g2_xnor2_1 _3130_ (.Y(_0307_),
    .A(_0306_),
    .B(_0242_));
 sg13g2_xnor2_1 _3131_ (.Y(_0308_),
    .A(_0231_),
    .B(_0307_));
 sg13g2_inv_1 _3132_ (.Y(_0309_),
    .A(_0308_));
 sg13g2_nand2_1 _3133_ (.Y(_0310_),
    .A(_0301_),
    .B(_0309_));
 sg13g2_nand3_1 _3134_ (.B(_0300_),
    .C(_0308_),
    .A(_0297_),
    .Y(_0311_));
 sg13g2_nand3b_1 _3135_ (.B(_0310_),
    .C(_0311_),
    .Y(_0312_),
    .A_N(_0273_));
 sg13g2_nand2_1 _3136_ (.Y(_0313_),
    .A(_0301_),
    .B(_0308_));
 sg13g2_nand3_1 _3137_ (.B(_0300_),
    .C(_0309_),
    .A(_0297_),
    .Y(_0314_));
 sg13g2_nand3_1 _3138_ (.B(_0314_),
    .C(_0273_),
    .A(_0313_),
    .Y(_0315_));
 sg13g2_nand2_1 _3139_ (.Y(_0316_),
    .A(_0312_),
    .B(_0315_));
 sg13g2_nand2b_1 _3140_ (.Y(_0317_),
    .B(_0316_),
    .A_N(_0271_));
 sg13g2_nand3_1 _3141_ (.B(_0315_),
    .C(_0271_),
    .A(_0312_),
    .Y(_0318_));
 sg13g2_inv_1 _3142_ (.Y(_0319_),
    .A(_0261_));
 sg13g2_a21oi_1 _3143_ (.A1(_0259_),
    .A2(_0221_),
    .Y(_0320_),
    .B1(_0319_));
 sg13g2_inv_1 _3144_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_nand3_1 _3145_ (.B(_0318_),
    .C(_0321_),
    .A(_0317_),
    .Y(_0322_));
 sg13g2_buf_1 _3146_ (.A(_0322_),
    .X(_0323_));
 sg13g2_nand2_1 _3147_ (.Y(_0324_),
    .A(_0317_),
    .B(_0318_));
 sg13g2_nand2_1 _3148_ (.Y(_0325_),
    .A(_0324_),
    .B(_0320_));
 sg13g2_a22oi_1 _3149_ (.Y(_0326_),
    .B1(_0323_),
    .B2(_0325_),
    .A2(_0268_),
    .A1(_0267_));
 sg13g2_nand2_1 _3150_ (.Y(_0327_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_nand2_1 _3151_ (.Y(_0328_),
    .A(_0325_),
    .B(_0323_));
 sg13g2_nor2_1 _3152_ (.A(_0327_),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_buf_1 _3153_ (.A(\main.demo._q_modulo_1[13] ),
    .X(_0330_));
 sg13g2_xnor2_1 _3154_ (.Y(_0331_),
    .A(_1420_),
    .B(_0330_));
 sg13g2_nor2_1 _3155_ (.A(\main.demo._q_modulo_1[6] ),
    .B(_1521_),
    .Y(_0332_));
 sg13g2_inv_1 _3156_ (.Y(_0333_),
    .A(\main.demo._q_modulo_1[6] ));
 sg13g2_nor2_1 _3157_ (.A(_1460_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_nor2_1 _3158_ (.A(_0332_),
    .B(_0334_),
    .Y(_0335_));
 sg13g2_nor2_1 _3159_ (.A(\main.demo._q_modulo_1[5] ),
    .B(_1508_),
    .Y(_0336_));
 sg13g2_a21oi_1 _3160_ (.A1(_0335_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(_0332_));
 sg13g2_buf_1 _3161_ (.A(\main.demo._q_modulo_1[8] ),
    .X(_0338_));
 sg13g2_nor2_1 _3162_ (.A(_0338_),
    .B(_1447_),
    .Y(_0339_));
 sg13g2_nor2b_1 _3163_ (.A(\main.demo._q_frame[9] ),
    .B_N(_0338_),
    .Y(_0340_));
 sg13g2_nor2_1 _3164_ (.A(_0339_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_inv_1 _3165_ (.Y(_0342_),
    .A(_0341_));
 sg13g2_nor2_1 _3166_ (.A(\main.demo._q_modulo_1[7] ),
    .B(_1455_),
    .Y(_0343_));
 sg13g2_nor2b_1 _3167_ (.A(_1454_),
    .B_N(\main.demo._q_modulo_1[7] ),
    .Y(_0344_));
 sg13g2_nor2_1 _3168_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_inv_1 _3169_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_nor2_1 _3170_ (.A(_0342_),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_inv_1 _3171_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_a21oi_1 _3172_ (.A1(_0341_),
    .A2(_0343_),
    .Y(_0349_),
    .B1(_0339_));
 sg13g2_o21ai_1 _3173_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0337_),
    .A2(_0348_));
 sg13g2_nor2_1 _3174_ (.A(\main.demo._q_modulo_1[10] ),
    .B(_1513_),
    .Y(_0351_));
 sg13g2_inv_1 _3175_ (.Y(_0352_),
    .A(\main.demo._q_modulo_1[10] ));
 sg13g2_nor2_1 _3176_ (.A(_1436_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_nor2_1 _3177_ (.A(_0351_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_nor2_1 _3178_ (.A(\main.demo._q_modulo_1[9] ),
    .B(_1441_),
    .Y(_0355_));
 sg13g2_inv_1 _3179_ (.Y(_0356_),
    .A(\main.demo._q_modulo_1[9] ));
 sg13g2_nor2_1 _3180_ (.A(_1440_),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_nor2_2 _3181_ (.A(_0355_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_nand2_1 _3182_ (.Y(_0359_),
    .A(_0354_),
    .B(_0358_));
 sg13g2_buf_1 _3183_ (.A(\main.demo._q_modulo_1[12] ),
    .X(_0360_));
 sg13g2_nor2_1 _3184_ (.A(_0360_),
    .B(_1427_),
    .Y(_0361_));
 sg13g2_inv_1 _3185_ (.Y(_0362_),
    .A(_0360_));
 sg13g2_nor2_1 _3186_ (.A(\main.demo._q_frame[13] ),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nor2_2 _3187_ (.A(_0361_),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_inv_1 _3188_ (.Y(_0365_),
    .A(_0364_));
 sg13g2_nor2_1 _3189_ (.A(\main.demo._q_modulo_1[11] ),
    .B(_1515_),
    .Y(_0366_));
 sg13g2_inv_1 _3190_ (.Y(_0367_),
    .A(\main.demo._q_modulo_1[11] ));
 sg13g2_nor2_1 _3191_ (.A(_1433_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_nor2_1 _3192_ (.A(_0366_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_inv_1 _3193_ (.Y(_0370_),
    .A(_0369_));
 sg13g2_nor2_1 _3194_ (.A(_0365_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_inv_1 _3195_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_nor2_1 _3196_ (.A(_0359_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_xnor2_1 _3197_ (.Y(_0374_),
    .A(_1496_),
    .B(\main.demo._q_modulo_1[1] ));
 sg13g2_nand2_1 _3198_ (.Y(_0375_),
    .A(_1493_),
    .B(\main.demo._q_modulo_1[0] ));
 sg13g2_nor2_1 _3199_ (.A(\main.demo._q_modulo_1[1] ),
    .B(_1497_),
    .Y(_0376_));
 sg13g2_a21oi_1 _3200_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0377_),
    .B1(_0376_));
 sg13g2_nor2_1 _3201_ (.A(\main.demo._q_modulo_1[2] ),
    .B(_1468_),
    .Y(_0378_));
 sg13g2_inv_1 _3202_ (.Y(_0379_),
    .A(_0378_));
 sg13g2_inv_1 _3203_ (.Y(_0380_),
    .A(\main.demo._q_modulo_1[2] ));
 sg13g2_nor2_1 _3204_ (.A(_1467_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_a21oi_2 _3205_ (.B1(_0381_),
    .Y(_0382_),
    .A2(_0379_),
    .A1(_0377_));
 sg13g2_nor2_2 _3206_ (.A(\main.demo._q_modulo_1[4] ),
    .B(_1476_),
    .Y(_0383_));
 sg13g2_inv_1 _3207_ (.Y(_0384_),
    .A(\main.demo._q_modulo_1[4] ));
 sg13g2_nor2_1 _3208_ (.A(_1475_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor2_2 _3209_ (.A(_0383_),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_inv_1 _3210_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_nor2_1 _3211_ (.A(\main.demo._q_modulo_1[3] ),
    .B(_1471_),
    .Y(_0388_));
 sg13g2_inv_1 _3212_ (.Y(_0389_),
    .A(\main.demo._q_modulo_1[3] ));
 sg13g2_nor2_1 _3213_ (.A(_1464_),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_nor2_1 _3214_ (.A(_0388_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_inv_1 _3215_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_nor2_1 _3216_ (.A(_0387_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_a21oi_1 _3217_ (.A1(_0386_),
    .A2(_0388_),
    .Y(_0394_),
    .B1(_0383_));
 sg13g2_inv_1 _3218_ (.Y(_0395_),
    .A(_0394_));
 sg13g2_a21oi_2 _3219_ (.B1(_0395_),
    .Y(_0396_),
    .A2(_0393_),
    .A1(_0382_));
 sg13g2_inv_1 _3220_ (.Y(_0397_),
    .A(_0396_));
 sg13g2_inv_1 _3221_ (.Y(_0398_),
    .A(_0335_));
 sg13g2_inv_1 _3222_ (.Y(_0399_),
    .A(\main.demo._q_modulo_1[5] ));
 sg13g2_nor2_1 _3223_ (.A(_1481_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_nor2_1 _3224_ (.A(_0336_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_inv_1 _3225_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_nor2_1 _3226_ (.A(_0398_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_inv_1 _3227_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_nor4_1 _3228_ (.A(_0359_),
    .B(_0372_),
    .C(_0404_),
    .D(_0348_),
    .Y(_0405_));
 sg13g2_a21oi_1 _3229_ (.A1(_0354_),
    .A2(_0355_),
    .Y(_0406_),
    .B1(_0351_));
 sg13g2_a21oi_1 _3230_ (.A1(_0364_),
    .A2(_0366_),
    .Y(_0407_),
    .B1(_0361_));
 sg13g2_o21ai_1 _3231_ (.B1(_0407_),
    .Y(_0408_),
    .A1(_0372_),
    .A2(_0406_));
 sg13g2_a221oi_1 _3232_ (.B2(_0405_),
    .C1(_0408_),
    .B1(_0397_),
    .A1(_0350_),
    .Y(_0409_),
    .A2(_0373_));
 sg13g2_xnor2_1 _3233_ (.Y(_0410_),
    .A(_0331_),
    .B(_0409_));
 sg13g2_inv_1 _3234_ (.Y(_0411_),
    .A(\main.demo._q_frame[15] ));
 sg13g2_nor2_1 _3235_ (.A(\main.demo._q_modulo_1[14] ),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_inv_1 _3236_ (.Y(_0413_),
    .A(\main.demo._q_modulo_1[14] ));
 sg13g2_nor2_1 _3237_ (.A(\main.demo._q_frame[15] ),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_nor2_1 _3238_ (.A(_0412_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_inv_1 _3239_ (.Y(_0416_),
    .A(_0415_));
 sg13g2_nand2_1 _3240_ (.Y(_0417_),
    .A(_0331_),
    .B(_0361_));
 sg13g2_o21ai_1 _3241_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_1421_),
    .A2(_0330_));
 sg13g2_buf_1 _3242_ (.A(_0418_),
    .X(_0419_));
 sg13g2_inv_1 _3243_ (.Y(_0420_),
    .A(_0390_));
 sg13g2_a21oi_1 _3244_ (.A1(_0382_),
    .A2(_0420_),
    .Y(_0421_),
    .B1(_0388_));
 sg13g2_inv_1 _3245_ (.Y(_0422_),
    .A(_0421_));
 sg13g2_nand2_1 _3246_ (.Y(_0423_),
    .A(_0345_),
    .B(_0335_));
 sg13g2_nor3_1 _3247_ (.A(_0402_),
    .B(_0387_),
    .C(_0423_),
    .Y(_0424_));
 sg13g2_inv_1 _3248_ (.Y(_0425_),
    .A(_0354_));
 sg13g2_nor2_1 _3249_ (.A(_0370_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_inv_1 _3250_ (.Y(_0427_),
    .A(_0426_));
 sg13g2_inv_1 _3251_ (.Y(_0428_),
    .A(_0358_));
 sg13g2_nor2_1 _3252_ (.A(_0428_),
    .B(_0342_),
    .Y(_0429_));
 sg13g2_nor2b_1 _3253_ (.A(_0427_),
    .B_N(_0429_),
    .Y(_0430_));
 sg13g2_nand3_1 _3254_ (.B(_0424_),
    .C(_0430_),
    .A(_0422_),
    .Y(_0431_));
 sg13g2_inv_1 _3255_ (.Y(_0432_),
    .A(_0400_));
 sg13g2_a21oi_1 _3256_ (.A1(_0432_),
    .A2(_0383_),
    .Y(_0433_),
    .B1(_0336_));
 sg13g2_a21oi_1 _3257_ (.A1(_0345_),
    .A2(_0332_),
    .Y(_0434_),
    .B1(_0343_));
 sg13g2_o21ai_1 _3258_ (.B1(_0434_),
    .Y(_0435_),
    .A1(_0423_),
    .A2(_0433_));
 sg13g2_a21oi_1 _3259_ (.A1(_0358_),
    .A2(_0339_),
    .Y(_0436_),
    .B1(_0355_));
 sg13g2_a21oi_1 _3260_ (.A1(_0369_),
    .A2(_0351_),
    .Y(_0437_),
    .B1(_0366_));
 sg13g2_o21ai_1 _3261_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0427_),
    .A2(_0436_));
 sg13g2_a21oi_1 _3262_ (.A1(_0435_),
    .A2(_0430_),
    .Y(_0439_),
    .B1(_0438_));
 sg13g2_nand2_1 _3263_ (.Y(_0440_),
    .A(_0364_),
    .B(_0331_));
 sg13g2_a21oi_2 _3264_ (.B1(_0440_),
    .Y(_0441_),
    .A2(_0439_),
    .A1(_0431_));
 sg13g2_nor3_1 _3265_ (.A(_0416_),
    .B(_0419_),
    .C(_0441_),
    .Y(_0442_));
 sg13g2_o21ai_1 _3266_ (.B1(_0416_),
    .Y(_0443_),
    .A1(_0419_),
    .A2(_0441_));
 sg13g2_nand2_1 _3267_ (.Y(_0444_),
    .A(_0431_),
    .B(_0439_));
 sg13g2_xnor2_1 _3268_ (.Y(_0445_),
    .A(_0364_),
    .B(_0444_));
 sg13g2_nand2_1 _3269_ (.Y(_0446_),
    .A(_0443_),
    .B(_0445_));
 sg13g2_buf_1 _3270_ (.A(\main.demo._q_modulo_1[15] ),
    .X(_0447_));
 sg13g2_nand2_1 _3271_ (.Y(_0448_),
    .A(_0441_),
    .B(_0415_));
 sg13g2_inv_1 _3272_ (.Y(_0449_),
    .A(_0412_));
 sg13g2_nand2b_1 _3273_ (.Y(_0450_),
    .B(_0419_),
    .A_N(_0414_));
 sg13g2_nand3_1 _3274_ (.B(_0449_),
    .C(_0450_),
    .A(_0448_),
    .Y(_0451_));
 sg13g2_xnor2_1 _3275_ (.Y(_0452_),
    .A(_0447_),
    .B(_0451_));
 sg13g2_nor4_2 _3276_ (.A(_0410_),
    .B(_0442_),
    .C(_0446_),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_o21ai_1 _3277_ (.B1(_0337_),
    .Y(_0454_),
    .A1(_0404_),
    .A2(_0396_));
 sg13g2_inv_1 _3278_ (.Y(_0455_),
    .A(_0349_));
 sg13g2_a21oi_1 _3279_ (.A1(_0454_),
    .A2(_0347_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_o21ai_1 _3280_ (.B1(_0406_),
    .Y(_0457_),
    .A1(_0359_),
    .A2(_0456_));
 sg13g2_xnor2_1 _3281_ (.Y(_0458_),
    .A(_0370_),
    .B(_0457_));
 sg13g2_a21o_1 _3282_ (.A2(_0424_),
    .A1(_0422_),
    .B1(_0435_),
    .X(_0459_));
 sg13g2_inv_1 _3283_ (.Y(_0460_),
    .A(_0436_));
 sg13g2_a21oi_1 _3284_ (.A1(_0459_),
    .A2(_0429_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_xnor2_1 _3285_ (.Y(_0462_),
    .A(_0425_),
    .B(_0461_));
 sg13g2_nor2b_1 _3286_ (.A(_0458_),
    .B_N(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _3287_ (.Y(_0464_),
    .A(_0342_),
    .B(_0459_));
 sg13g2_xor2_1 _3288_ (.B(_0464_),
    .A(_1639_),
    .X(_0465_));
 sg13g2_xnor2_1 _3289_ (.Y(_0466_),
    .A(_1486_),
    .B(\main.demo._q_modulo_1[0] ));
 sg13g2_xnor2_1 _3290_ (.Y(_0467_),
    .A(_0466_),
    .B(_1588_));
 sg13g2_xor2_1 _3291_ (.B(_0374_),
    .A(_0375_),
    .X(_0468_));
 sg13g2_xnor2_1 _3292_ (.Y(_0469_),
    .A(_1591_),
    .B(_0468_));
 sg13g2_nor2_1 _3293_ (.A(_0381_),
    .B(_0378_),
    .Y(_0470_));
 sg13g2_xnor2_1 _3294_ (.Y(_0471_),
    .A(_0470_),
    .B(_0377_));
 sg13g2_xnor2_1 _3295_ (.Y(_0472_),
    .A(_1595_),
    .B(_0471_));
 sg13g2_inv_1 _3296_ (.Y(_0473_),
    .A(_1584_));
 sg13g2_xnor2_1 _3297_ (.Y(_0474_),
    .A(_0392_),
    .B(_0382_));
 sg13g2_xnor2_1 _3298_ (.Y(_0475_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_nor4_1 _3299_ (.A(_0467_),
    .B(_0469_),
    .C(_0472_),
    .D(_0475_),
    .Y(_0476_));
 sg13g2_xnor2_1 _3300_ (.Y(_0477_),
    .A(_0386_),
    .B(_0421_));
 sg13g2_xnor2_1 _3301_ (.Y(_0478_),
    .A(_1631_),
    .B(_0477_));
 sg13g2_xnor2_1 _3302_ (.Y(_0479_),
    .A(_0402_),
    .B(_0396_));
 sg13g2_xnor2_1 _3303_ (.Y(_0480_),
    .A(_1628_),
    .B(_0479_));
 sg13g2_nand3_1 _3304_ (.B(_0478_),
    .C(_0480_),
    .A(_0476_),
    .Y(_0481_));
 sg13g2_xnor2_1 _3305_ (.Y(_0482_),
    .A(_0346_),
    .B(_0454_));
 sg13g2_xnor2_1 _3306_ (.Y(_0483_),
    .A(_1615_),
    .B(_0482_));
 sg13g2_nand2_1 _3307_ (.Y(_0484_),
    .A(_0422_),
    .B(_0386_));
 sg13g2_nor2_1 _3308_ (.A(_0336_),
    .B(_0383_),
    .Y(_0485_));
 sg13g2_a21oi_1 _3309_ (.A1(_0484_),
    .A2(_0485_),
    .Y(_0486_),
    .B1(_0400_));
 sg13g2_xnor2_1 _3310_ (.Y(_0487_),
    .A(_0398_),
    .B(_0486_));
 sg13g2_xnor2_1 _3311_ (.Y(_0488_),
    .A(_1619_),
    .B(_0487_));
 sg13g2_nor3_1 _3312_ (.A(_0481_),
    .B(_0483_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_xnor2_1 _3313_ (.Y(_0490_),
    .A(_0358_),
    .B(_0456_));
 sg13g2_xor2_1 _3314_ (.B(_0490_),
    .A(_1642_),
    .X(_0491_));
 sg13g2_and2_1 _3315_ (.A(_0489_),
    .B(_0491_),
    .X(_0492_));
 sg13g2_nand4_1 _3316_ (.B(_0463_),
    .C(_0465_),
    .A(_0453_),
    .Y(_0493_),
    .D(_0492_));
 sg13g2_buf_2 _3317_ (.A(_0493_),
    .X(_0494_));
 sg13g2_nand2_1 _3318_ (.Y(_0495_),
    .A(_0494_),
    .B(_1869_));
 sg13g2_nor3_1 _3319_ (.A(_0326_),
    .B(_0329_),
    .C(_0495_),
    .Y(_0104_));
 sg13g2_nor2b_1 _3320_ (.A(_0242_),
    .B_N(_0306_),
    .Y(_0496_));
 sg13g2_a21o_1 _3321_ (.A2(_0230_),
    .A1(_0307_),
    .B1(_0496_),
    .X(_0497_));
 sg13g2_buf_1 _3322_ (.A(_0497_),
    .X(_0498_));
 sg13g2_nand2_1 _3323_ (.Y(_0499_),
    .A(_0279_),
    .B(_0275_));
 sg13g2_inv_1 _3324_ (.Y(_0500_),
    .A(_0499_));
 sg13g2_nor2_1 _3325_ (.A(_0192_),
    .B(_0207_),
    .Y(_0501_));
 sg13g2_buf_2 _3326_ (.A(_0501_),
    .X(_0502_));
 sg13g2_xnor2_1 _3327_ (.Y(_0503_),
    .A(_0502_),
    .B(_0280_));
 sg13g2_xnor2_1 _3328_ (.Y(_0504_),
    .A(_0500_),
    .B(_0503_));
 sg13g2_nand2_1 _3329_ (.Y(_0505_),
    .A(_0291_),
    .B(_0294_));
 sg13g2_xnor2_1 _3330_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_inv_1 _3331_ (.Y(_0507_),
    .A(_0283_));
 sg13g2_a21oi_1 _3332_ (.A1(_0281_),
    .A2(_0285_),
    .Y(_0508_),
    .B1(_0507_));
 sg13g2_inv_1 _3333_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_buf_1 _3334_ (.A(\main.demo._q_rand_1[9] ),
    .X(_0510_));
 sg13g2_nand2_1 _3335_ (.Y(_0511_),
    .A(net35),
    .B(_0302_));
 sg13g2_nand2_1 _3336_ (.Y(_0512_),
    .A(_0304_),
    .B(_0511_));
 sg13g2_o21ai_1 _3337_ (.B1(_0512_),
    .Y(_0513_),
    .A1(_0150_),
    .A2(_0511_));
 sg13g2_xnor2_1 _3338_ (.Y(_0514_),
    .A(_0510_),
    .B(_0513_));
 sg13g2_inv_1 _3339_ (.Y(_0515_),
    .A(_0514_));
 sg13g2_nand2_1 _3340_ (.Y(_0516_),
    .A(_0509_),
    .B(_0515_));
 sg13g2_nand2_1 _3341_ (.Y(_0517_),
    .A(_0508_),
    .B(_0514_));
 sg13g2_nand2_1 _3342_ (.Y(_0518_),
    .A(_0516_),
    .B(_0517_));
 sg13g2_nand3_1 _3343_ (.B(_0150_),
    .C(_0227_),
    .A(_0303_),
    .Y(_0519_));
 sg13g2_inv_1 _3344_ (.Y(_0520_),
    .A(_0519_));
 sg13g2_nand2_1 _3345_ (.Y(_0521_),
    .A(_0518_),
    .B(_0520_));
 sg13g2_nand3_1 _3346_ (.B(_0519_),
    .C(_0517_),
    .A(_0516_),
    .Y(_0522_));
 sg13g2_nand2_1 _3347_ (.Y(_0523_),
    .A(_0521_),
    .B(_0522_));
 sg13g2_xnor2_1 _3348_ (.Y(_0524_),
    .A(_0506_),
    .B(_0523_));
 sg13g2_inv_1 _3349_ (.Y(_0525_),
    .A(_0300_));
 sg13g2_a21oi_1 _3350_ (.A1(_0297_),
    .A2(_0308_),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_inv_1 _3351_ (.Y(_0527_),
    .A(_0526_));
 sg13g2_nand2_1 _3352_ (.Y(_0528_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_nand2_1 _3353_ (.Y(_0529_),
    .A(_0518_),
    .B(_0519_));
 sg13g2_nand3_1 _3354_ (.B(_0520_),
    .C(_0517_),
    .A(_0516_),
    .Y(_0530_));
 sg13g2_nand2_1 _3355_ (.Y(_0531_),
    .A(_0529_),
    .B(_0530_));
 sg13g2_nand2_1 _3356_ (.Y(_0532_),
    .A(_0531_),
    .B(_0506_));
 sg13g2_inv_1 _3357_ (.Y(_0533_),
    .A(_0504_));
 sg13g2_xnor2_1 _3358_ (.Y(_0534_),
    .A(_0533_),
    .B(_0505_));
 sg13g2_nand2_1 _3359_ (.Y(_0535_),
    .A(_0523_),
    .B(_0534_));
 sg13g2_nand2_1 _3360_ (.Y(_0536_),
    .A(_0532_),
    .B(_0535_));
 sg13g2_nand2_1 _3361_ (.Y(_0537_),
    .A(_0536_),
    .B(_0526_));
 sg13g2_nand2_1 _3362_ (.Y(_0538_),
    .A(_0528_),
    .B(_0537_));
 sg13g2_xnor2_1 _3363_ (.Y(_0539_),
    .A(_0498_),
    .B(_0538_));
 sg13g2_inv_1 _3364_ (.Y(_0540_),
    .A(_0312_));
 sg13g2_a21oi_1 _3365_ (.A1(_0315_),
    .A2(_0271_),
    .Y(_0541_),
    .B1(_0540_));
 sg13g2_inv_1 _3366_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_nand2_1 _3367_ (.Y(_0543_),
    .A(_0539_),
    .B(_0542_));
 sg13g2_nand2b_1 _3368_ (.Y(_0544_),
    .B(_0538_),
    .A_N(_0498_));
 sg13g2_nand3_1 _3369_ (.B(_0537_),
    .C(_0498_),
    .A(_0528_),
    .Y(_0545_));
 sg13g2_nand2_1 _3370_ (.Y(_0546_),
    .A(_0544_),
    .B(_0545_));
 sg13g2_nand2_1 _3371_ (.Y(_0547_),
    .A(_0546_),
    .B(_0541_));
 sg13g2_nand2_1 _3372_ (.Y(_0548_),
    .A(_0543_),
    .B(_0547_));
 sg13g2_inv_1 _3373_ (.Y(_0549_),
    .A(_0325_));
 sg13g2_a21oi_1 _3374_ (.A1(_0327_),
    .A2(_0323_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_xor2_1 _3375_ (.B(_0550_),
    .A(_0548_),
    .X(_0551_));
 sg13g2_nor2_1 _3376_ (.A(_0495_),
    .B(_0551_),
    .Y(_0105_));
 sg13g2_inv_1 _3377_ (.Y(_0552_),
    .A(\main.demo.vga._q_xcount[7] ));
 sg13g2_buf_1 _3378_ (.A(\main.demo.vga._q_xcount[5] ),
    .X(_0553_));
 sg13g2_buf_1 _3379_ (.A(\main.demo.vga._q_xcount[4] ),
    .X(_0554_));
 sg13g2_buf_1 _3380_ (.A(\main.demo.vga._q_xcount[6] ),
    .X(_0555_));
 sg13g2_nand4_1 _3381_ (.B(_0553_),
    .C(_0554_),
    .A(_0552_),
    .Y(_0556_),
    .D(_0555_));
 sg13g2_or2_1 _3382_ (.X(_0557_),
    .B(\main.demo.vga._q_xcount[0] ),
    .A(\main.demo.vga._q_xcount[1] ));
 sg13g2_nor3_1 _3383_ (.A(\main.demo.vga._q_xcount[3] ),
    .B(\main.demo.vga._q_xcount[2] ),
    .C(_0557_),
    .Y(_0558_));
 sg13g2_nor2b_1 _3384_ (.A(_0556_),
    .B_N(_0558_),
    .Y(_0559_));
 sg13g2_inv_1 _3385_ (.Y(_0560_),
    .A(\main.demo.vga._q_xcount[9] ));
 sg13g2_inv_1 _3386_ (.Y(_0561_),
    .A(\main.demo.vga._q_xcount[8] ));
 sg13g2_inv_1 _3387_ (.Y(_0562_),
    .A(\main.demo.vga._q_xcount[10] ));
 sg13g2_nor3_1 _3388_ (.A(_0560_),
    .B(_0561_),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_inv_1 _3389_ (.Y(_0564_),
    .A(\main.demo.vga._q_xcount[2] ));
 sg13g2_nand2_1 _3390_ (.Y(_0565_),
    .A(\main.demo.vga._q_xcount[1] ),
    .B(\main.demo.vga._q_xcount[0] ));
 sg13g2_nor2_1 _3391_ (.A(_0564_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_and2_1 _3392_ (.A(_0566_),
    .B(\main.demo.vga._q_xcount[3] ),
    .X(_0567_));
 sg13g2_buf_1 _3393_ (.A(_0567_),
    .X(_0568_));
 sg13g2_inv_1 _3394_ (.Y(_0569_),
    .A(_0555_));
 sg13g2_nor4_1 _3395_ (.A(_0553_),
    .B(_0554_),
    .C(_0569_),
    .D(_0552_),
    .Y(_0570_));
 sg13g2_nand3_1 _3396_ (.B(_0570_),
    .C(_0563_),
    .A(_0568_),
    .Y(_0571_));
 sg13g2_a221oi_1 _3397_ (.B2(_1574_),
    .C1(_0004_),
    .B1(_0571_),
    .A1(_0559_),
    .Y(_0108_),
    .A2(_0563_));
 sg13g2_buf_1 _3398_ (.A(\main.demo.vga._q_ycount[1] ),
    .X(_0572_));
 sg13g2_buf_1 _3399_ (.A(\main.demo.vga._q_ycount[0] ),
    .X(_0573_));
 sg13g2_inv_1 _3400_ (.Y(_0574_),
    .A(_0573_));
 sg13g2_buf_1 _3401_ (.A(\main.demo.vga._q_ycount[5] ),
    .X(_0575_));
 sg13g2_inv_1 _3402_ (.Y(_0576_),
    .A(\main.demo.vga._q_ycount[4] ));
 sg13g2_nand2_1 _3403_ (.Y(_0577_),
    .A(\main.demo.vga._q_ycount[7] ),
    .B(\main.demo.vga._q_ycount[6] ));
 sg13g2_nor3_1 _3404_ (.A(_0575_),
    .B(_0576_),
    .C(_0577_),
    .Y(_0578_));
 sg13g2_buf_1 _3405_ (.A(\main.demo.vga._q_ycount[8] ),
    .X(_0579_));
 sg13g2_buf_1 _3406_ (.A(\main.demo.vga._q_ycount[2] ),
    .X(_0580_));
 sg13g2_nand2_1 _3407_ (.Y(_0581_),
    .A(\main.demo.vga._q_ycount[3] ),
    .B(_0580_));
 sg13g2_inv_1 _3408_ (.Y(_0582_),
    .A(_0581_));
 sg13g2_nand4_1 _3409_ (.B(_0579_),
    .C(\main.demo.vga._d_vblank ),
    .A(_0578_),
    .Y(_0583_),
    .D(_0582_));
 sg13g2_nor3_1 _3410_ (.A(_0572_),
    .B(_0574_),
    .C(_0583_),
    .Y(_0584_));
 sg13g2_inv_1 _3411_ (.Y(_0585_),
    .A(_0572_));
 sg13g2_nor3_1 _3412_ (.A(_0585_),
    .B(_0573_),
    .C(_0583_),
    .Y(_0586_));
 sg13g2_nor2_1 _3413_ (.A(\main._w_demo_video_vs ),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nor3_1 _3414_ (.A(_0004_),
    .B(_0584_),
    .C(_0587_),
    .Y(_0109_));
 sg13g2_nor4_1 _3415_ (.A(_0572_),
    .B(_0573_),
    .C(\main.demo.vga._q_ycount[3] ),
    .D(_0580_),
    .Y(_0588_));
 sg13g2_nor2_1 _3416_ (.A(\main.demo.vga._q_ycount[4] ),
    .B(\main.demo.vga._d_vblank ),
    .Y(_0589_));
 sg13g2_inv_1 _3417_ (.Y(_0590_),
    .A(_0575_));
 sg13g2_inv_1 _3418_ (.Y(_0591_),
    .A(_0579_));
 sg13g2_nor3_1 _3419_ (.A(_0590_),
    .B(_0591_),
    .C(_0577_),
    .Y(_0592_));
 sg13g2_nand3_1 _3420_ (.B(_0589_),
    .C(_0592_),
    .A(_0588_),
    .Y(_0593_));
 sg13g2_nor4_1 _3421_ (.A(_0575_),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(_0579_),
    .Y(_0594_));
 sg13g2_and3_1 _3422_ (.X(_0595_),
    .A(_0588_),
    .B(_0594_),
    .C(_0589_));
 sg13g2_a21oi_1 _3423_ (.A1(\main.demo.vga._q_active_v ),
    .A2(_0593_),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_buf_1 _3424_ (.A(_0596_),
    .X(_0597_));
 sg13g2_nor2_1 _3425_ (.A(_0574_),
    .B(net21),
    .Y(_0110_));
 sg13g2_nor2_1 _3426_ (.A(_0585_),
    .B(net21),
    .Y(_0111_));
 sg13g2_nor2b_1 _3427_ (.A(net21),
    .B_N(_0580_),
    .Y(_0112_));
 sg13g2_inv_1 _3428_ (.Y(_0598_),
    .A(\main.demo.vga._q_ycount[3] ));
 sg13g2_nor2_1 _3429_ (.A(_0598_),
    .B(_0597_),
    .Y(_0113_));
 sg13g2_nor2_1 _3430_ (.A(_0576_),
    .B(net21),
    .Y(_0114_));
 sg13g2_nor2_1 _3431_ (.A(_0590_),
    .B(net21),
    .Y(_0115_));
 sg13g2_inv_1 _3432_ (.Y(_0599_),
    .A(\main.demo.vga._q_ycount[6] ));
 sg13g2_nor2_1 _3433_ (.A(_0599_),
    .B(net21),
    .Y(_0116_));
 sg13g2_nor2b_1 _3434_ (.A(net21),
    .B_N(\main.demo.vga._q_ycount[7] ),
    .Y(_0117_));
 sg13g2_inv_1 _3435_ (.Y(_0600_),
    .A(_0553_));
 sg13g2_nand2_1 _3436_ (.Y(_0601_),
    .A(_0568_),
    .B(_0554_));
 sg13g2_nor2_1 _3437_ (.A(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_a21oi_1 _3438_ (.A1(_0568_),
    .A2(_0554_),
    .Y(_0603_),
    .B1(_0553_));
 sg13g2_nor2_1 _3439_ (.A(_0553_),
    .B(_0554_),
    .Y(_0604_));
 sg13g2_nor3_1 _3440_ (.A(\main.demo.vga._q_xcount[8] ),
    .B(\main.demo.vga._q_xcount[10] ),
    .C(_0560_),
    .Y(_0605_));
 sg13g2_nor2_1 _3441_ (.A(_0555_),
    .B(_0552_),
    .Y(_0606_));
 sg13g2_nand4_1 _3442_ (.B(_0604_),
    .C(_0605_),
    .A(_0558_),
    .Y(_0607_),
    .D(_0606_));
 sg13g2_buf_1 _3443_ (.A(_0607_),
    .X(_0608_));
 sg13g2_nand2_1 _3444_ (.Y(_0609_),
    .A(_0608_),
    .B(_1869_));
 sg13g2_nor3_1 _3445_ (.A(_0602_),
    .B(_0603_),
    .C(_0609_),
    .Y(_0124_));
 sg13g2_nor3_1 _3446_ (.A(_0600_),
    .B(_0569_),
    .C(_0601_),
    .Y(_0610_));
 sg13g2_nor2_1 _3447_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_nand2_1 _3448_ (.Y(_0612_),
    .A(_0610_),
    .B(\main.demo.vga._q_xcount[7] ));
 sg13g2_inv_1 _3449_ (.Y(_0613_),
    .A(_0612_));
 sg13g2_nor3_1 _3450_ (.A(_0609_),
    .B(_0611_),
    .C(_0613_),
    .Y(_0126_));
 sg13g2_nor2b_1 _3451_ (.A(_0216_),
    .B_N(_0209_),
    .Y(_0614_));
 sg13g2_inv_1 _3452_ (.Y(_0615_),
    .A(_0494_));
 sg13g2_a21oi_1 _3453_ (.A1(_0215_),
    .A2(_0614_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_o21ai_1 _3454_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0215_),
    .A2(_0614_));
 sg13g2_inv_1 _3455_ (.Y(_0618_),
    .A(_0528_));
 sg13g2_a21oi_1 _3456_ (.A1(_0537_),
    .A2(_0498_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nor2_1 _3457_ (.A(_0504_),
    .B(_0295_),
    .Y(_0620_));
 sg13g2_nand2b_1 _3458_ (.Y(_0621_),
    .B(_0532_),
    .A_N(_0620_));
 sg13g2_inv_1 _3459_ (.Y(_0622_),
    .A(_0511_));
 sg13g2_a22oi_1 _3460_ (.Y(_0623_),
    .B1(_0510_),
    .B2(_0512_),
    .A2(_0622_),
    .A1(_0225_));
 sg13g2_nand2_1 _3461_ (.Y(_0624_),
    .A(_0150_),
    .B(_0302_));
 sg13g2_xnor2_1 _3462_ (.Y(_0625_),
    .A(net35),
    .B(_0510_));
 sg13g2_nor2_1 _3463_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_nand2_1 _3464_ (.Y(_0627_),
    .A(_0625_),
    .B(_0624_));
 sg13g2_nand2b_1 _3465_ (.Y(_0628_),
    .B(_0627_),
    .A_N(_0626_));
 sg13g2_xnor2_1 _3466_ (.Y(_0629_),
    .A(\main.demo._q_rand_1[10] ),
    .B(_0628_));
 sg13g2_nand2_1 _3467_ (.Y(_0630_),
    .A(_0280_),
    .B(_0502_));
 sg13g2_nor2_1 _3468_ (.A(_0502_),
    .B(_0280_),
    .Y(_0631_));
 sg13g2_a21oi_1 _3469_ (.A1(_0630_),
    .A2(_0499_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_xnor2_1 _3470_ (.Y(_0633_),
    .A(_0629_),
    .B(_0632_));
 sg13g2_xnor2_1 _3471_ (.Y(_0634_),
    .A(_0623_),
    .B(_0633_));
 sg13g2_nor2_1 _3472_ (.A(_0294_),
    .B(_0504_),
    .Y(_0635_));
 sg13g2_xnor2_1 _3473_ (.Y(_0636_),
    .A(_0148_),
    .B(_0151_));
 sg13g2_xnor2_1 _3474_ (.Y(_0637_),
    .A(_0225_),
    .B(_0636_));
 sg13g2_xor2_1 _3475_ (.B(_0637_),
    .A(_0502_),
    .X(_0638_));
 sg13g2_nand2_1 _3476_ (.Y(_0639_),
    .A(_0638_),
    .B(_0500_));
 sg13g2_xnor2_1 _3477_ (.Y(_0640_),
    .A(_0502_),
    .B(_0637_));
 sg13g2_nand2_1 _3478_ (.Y(_0641_),
    .A(_0640_),
    .B(_0499_));
 sg13g2_nand2_1 _3479_ (.Y(_0642_),
    .A(_0639_),
    .B(_0641_));
 sg13g2_nand2_1 _3480_ (.Y(_0643_),
    .A(_0642_),
    .B(_0190_));
 sg13g2_nand3_1 _3481_ (.B(_0641_),
    .C(net37),
    .A(_0639_),
    .Y(_0644_));
 sg13g2_nand2_1 _3482_ (.Y(_0645_),
    .A(_0643_),
    .B(_0644_));
 sg13g2_nand2b_1 _3483_ (.Y(_0646_),
    .B(_0645_),
    .A_N(_0635_));
 sg13g2_nand3_1 _3484_ (.B(_0643_),
    .C(_0644_),
    .A(_0635_),
    .Y(_0647_));
 sg13g2_nand2_1 _3485_ (.Y(_0648_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_nand2b_1 _3486_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0634_));
 sg13g2_nand3_1 _3487_ (.B(_0634_),
    .C(_0647_),
    .A(_0646_),
    .Y(_0650_));
 sg13g2_nand2_1 _3488_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nand2b_1 _3489_ (.Y(_0652_),
    .B(_0651_),
    .A_N(_0621_));
 sg13g2_nand3_1 _3490_ (.B(_0650_),
    .C(_0621_),
    .A(_0649_),
    .Y(_0653_));
 sg13g2_nand2_1 _3491_ (.Y(_0654_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_nor2_1 _3492_ (.A(_0508_),
    .B(_0515_),
    .Y(_0655_));
 sg13g2_a21oi_1 _3493_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_nand2_1 _3494_ (.Y(_0657_),
    .A(_0654_),
    .B(_0656_));
 sg13g2_inv_1 _3495_ (.Y(_0658_),
    .A(_0656_));
 sg13g2_nand3_1 _3496_ (.B(_0653_),
    .C(_0658_),
    .A(_0652_),
    .Y(_0659_));
 sg13g2_nand3b_1 _3497_ (.B(_0657_),
    .C(_0659_),
    .Y(_0660_),
    .A_N(_0619_));
 sg13g2_nand2_1 _3498_ (.Y(_0661_),
    .A(_0657_),
    .B(_0659_));
 sg13g2_nand2_1 _3499_ (.Y(_0662_),
    .A(_0661_),
    .B(_0619_));
 sg13g2_nand2_1 _3500_ (.Y(_0663_),
    .A(_0660_),
    .B(_0662_));
 sg13g2_inv_1 _3501_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_inv_1 _3502_ (.Y(_0665_),
    .A(_0547_));
 sg13g2_a21oi_1 _3503_ (.A1(_0323_),
    .A2(_0543_),
    .Y(_0666_),
    .B1(_0665_));
 sg13g2_nor3_1 _3504_ (.A(_0327_),
    .B(_0548_),
    .C(_0328_),
    .Y(_0667_));
 sg13g2_nor3_1 _3505_ (.A(_0664_),
    .B(_0666_),
    .C(_0667_),
    .Y(_0668_));
 sg13g2_nor2b_1 _3506_ (.A(_0668_),
    .B_N(_0494_),
    .Y(_0669_));
 sg13g2_buf_8 _3507_ (.A(_0669_),
    .X(_0670_));
 sg13g2_o21ai_1 _3508_ (.B1(_0664_),
    .Y(_0671_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_buf_1 _3509_ (.A(_0671_),
    .X(_0672_));
 sg13g2_nand2_2 _3510_ (.Y(_0673_),
    .A(net17),
    .B(net18));
 sg13g2_buf_8 _3511_ (.A(_0673_),
    .X(_0674_));
 sg13g2_inv_1 _3512_ (.Y(_0675_),
    .A(_0010_));
 sg13g2_nand2_1 _3513_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_inv_1 _3514_ (.Y(_0677_),
    .A(_0011_));
 sg13g2_nand3_1 _3515_ (.B(_0677_),
    .C(net18),
    .A(net17),
    .Y(_0678_));
 sg13g2_nand2_1 _3516_ (.Y(_0679_),
    .A(_0676_),
    .B(_0678_));
 sg13g2_nand2_1 _3517_ (.Y(_0680_),
    .A(_0659_),
    .B(_0653_));
 sg13g2_inv_1 _3518_ (.Y(_0681_),
    .A(_0647_));
 sg13g2_inv_1 _3519_ (.Y(_0682_),
    .A(_0650_));
 sg13g2_nor2_1 _3520_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_nor2_1 _3521_ (.A(_0190_),
    .B(_0292_),
    .Y(_0684_));
 sg13g2_a21oi_1 _3522_ (.A1(_0642_),
    .A2(_0190_),
    .Y(_0685_),
    .B1(_0684_));
 sg13g2_a21oi_1 _3523_ (.A1(_0627_),
    .A2(\main.demo._q_rand_1[10] ),
    .Y(_0686_),
    .B1(_0626_));
 sg13g2_xor2_1 _3524_ (.B(_0302_),
    .A(\main.demo._q_rand_1[10] ),
    .X(_0687_));
 sg13g2_nand2_1 _3525_ (.Y(_0688_),
    .A(net35),
    .B(_0510_));
 sg13g2_xnor2_1 _3526_ (.Y(_0689_),
    .A(\main.demo._q_rand_1[11] ),
    .B(_0688_));
 sg13g2_xnor2_1 _3527_ (.Y(_0690_),
    .A(_0687_),
    .B(_0689_));
 sg13g2_xnor2_1 _3528_ (.Y(_0691_),
    .A(_0686_),
    .B(_0690_));
 sg13g2_nor2_1 _3529_ (.A(_0502_),
    .B(_0637_),
    .Y(_0692_));
 sg13g2_a21oi_1 _3530_ (.A1(_0638_),
    .A2(_0499_),
    .Y(_0693_),
    .B1(_0692_));
 sg13g2_xnor2_1 _3531_ (.Y(_0694_),
    .A(_0691_),
    .B(_0693_));
 sg13g2_xnor2_1 _3532_ (.Y(_0695_),
    .A(_0685_),
    .B(_0694_));
 sg13g2_nand2_1 _3533_ (.Y(_0696_),
    .A(_0148_),
    .B(_0151_));
 sg13g2_o21ai_1 _3534_ (.B1(_0696_),
    .Y(_0697_),
    .A1(_0225_),
    .A2(_0636_));
 sg13g2_xnor2_1 _3535_ (.Y(_0698_),
    .A(net35),
    .B(_0152_));
 sg13g2_xnor2_1 _3536_ (.Y(_0699_),
    .A(_0238_),
    .B(_0698_));
 sg13g2_xnor2_1 _3537_ (.Y(_0700_),
    .A(_0697_),
    .B(_0699_));
 sg13g2_xnor2_1 _3538_ (.Y(_0701_),
    .A(_0173_),
    .B(_0239_));
 sg13g2_nor2b_1 _3539_ (.A(_0210_),
    .B_N(_0237_),
    .Y(_0702_));
 sg13g2_o21ai_1 _3540_ (.B1(_0014_),
    .Y(_0703_),
    .A1(net37),
    .A2(_0702_));
 sg13g2_a21oi_1 _3541_ (.A1(net37),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_xnor2_1 _3542_ (.Y(_0705_),
    .A(_0701_),
    .B(_0704_));
 sg13g2_xnor2_1 _3543_ (.Y(_0706_),
    .A(_0700_),
    .B(_0705_));
 sg13g2_nand2b_1 _3544_ (.Y(_0707_),
    .B(_0706_),
    .A_N(_0695_));
 sg13g2_nand2b_1 _3545_ (.Y(_0708_),
    .B(_0695_),
    .A_N(_0706_));
 sg13g2_nand2_1 _3546_ (.Y(_0709_),
    .A(_0707_),
    .B(_0708_));
 sg13g2_or2_1 _3547_ (.X(_0710_),
    .B(_0709_),
    .A(_0683_));
 sg13g2_nand2_1 _3548_ (.Y(_0711_),
    .A(_0709_),
    .B(_0683_));
 sg13g2_nand2_1 _3549_ (.Y(_0712_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_inv_1 _3550_ (.Y(_0713_),
    .A(_0623_));
 sg13g2_nor2b_1 _3551_ (.A(_0632_),
    .B_N(_0629_),
    .Y(_0714_));
 sg13g2_a21oi_1 _3552_ (.A1(_0633_),
    .A2(_0713_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nand2_1 _3553_ (.Y(_0716_),
    .A(_0712_),
    .B(_0715_));
 sg13g2_inv_1 _3554_ (.Y(_0717_),
    .A(_0715_));
 sg13g2_nand3_1 _3555_ (.B(_0711_),
    .C(_0717_),
    .A(_0710_),
    .Y(_0718_));
 sg13g2_nand2_1 _3556_ (.Y(_0719_),
    .A(_0716_),
    .B(_0718_));
 sg13g2_xnor2_1 _3557_ (.Y(_0720_),
    .A(_0680_),
    .B(_0719_));
 sg13g2_nor2_1 _3558_ (.A(_0548_),
    .B(_0663_),
    .Y(_0721_));
 sg13g2_nand2_1 _3559_ (.Y(_0722_),
    .A(_0721_),
    .B(_0550_));
 sg13g2_nand2_1 _3560_ (.Y(_0723_),
    .A(_0660_),
    .B(_0543_));
 sg13g2_nand2_1 _3561_ (.Y(_0724_),
    .A(_0723_),
    .B(_0662_));
 sg13g2_nand2_1 _3562_ (.Y(_0725_),
    .A(_0722_),
    .B(_0724_));
 sg13g2_nand2b_1 _3563_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0720_));
 sg13g2_nand3_1 _3564_ (.B(_0720_),
    .C(_0724_),
    .A(_0722_),
    .Y(_0727_));
 sg13g2_nand3_1 _3565_ (.B(_0727_),
    .C(_0494_),
    .A(_0726_),
    .Y(_0728_));
 sg13g2_buf_2 _3566_ (.A(_0728_),
    .X(_0729_));
 sg13g2_buf_8 _3567_ (.A(_0729_),
    .X(_0730_));
 sg13g2_nand2_1 _3568_ (.Y(_0731_),
    .A(_0679_),
    .B(net10));
 sg13g2_nand2_1 _3569_ (.Y(_0732_),
    .A(net14),
    .B(_0012_));
 sg13g2_nand3_1 _3570_ (.B(_0000_),
    .C(net18),
    .A(net17),
    .Y(_0733_));
 sg13g2_nand2_1 _3571_ (.Y(_0734_),
    .A(_0727_),
    .B(_0494_));
 sg13g2_nor2b_1 _3572_ (.A(_0734_),
    .B_N(_0726_),
    .Y(_0735_));
 sg13g2_buf_1 _3573_ (.A(_0735_),
    .X(_0736_));
 sg13g2_nand3_1 _3574_ (.B(_0733_),
    .C(net13),
    .A(_0732_),
    .Y(_0737_));
 sg13g2_nand2_1 _3575_ (.Y(_0738_),
    .A(_0731_),
    .B(_0737_));
 sg13g2_nand2b_1 _3576_ (.Y(_0739_),
    .B(_0738_),
    .A_N(_0617_));
 sg13g2_nand3_1 _3577_ (.B(_0737_),
    .C(_0617_),
    .A(_0731_),
    .Y(_0740_));
 sg13g2_nand2_2 _3578_ (.Y(_0741_),
    .A(_0739_),
    .B(_0740_));
 sg13g2_xor2_1 _3579_ (.B(_0741_),
    .A(\main.demo._d___pip_24_1_2___stage___block_3_y[4] ),
    .X(_0742_));
 sg13g2_nand2b_1 _3580_ (.Y(_0743_),
    .B(_0674_),
    .A_N(_0008_));
 sg13g2_inv_1 _3581_ (.Y(_0744_),
    .A(_0009_));
 sg13g2_nand3_1 _3582_ (.B(_0744_),
    .C(net18),
    .A(net17),
    .Y(_0745_));
 sg13g2_nand3_1 _3583_ (.B(_0745_),
    .C(net13),
    .A(_0743_),
    .Y(_0746_));
 sg13g2_inv_1 _3584_ (.Y(_0747_),
    .A(_0017_));
 sg13g2_nand2_1 _3585_ (.Y(_0748_),
    .A(net14),
    .B(_0747_));
 sg13g2_inv_1 _3586_ (.Y(_0749_),
    .A(_0007_));
 sg13g2_nand3_1 _3587_ (.B(_0749_),
    .C(net18),
    .A(net17),
    .Y(_0750_));
 sg13g2_nand3_1 _3588_ (.B(_0750_),
    .C(_0730_),
    .A(_0748_),
    .Y(_0751_));
 sg13g2_nor2_1 _3589_ (.A(_0235_),
    .B(_0615_),
    .Y(_0752_));
 sg13g2_nand3_1 _3590_ (.B(_0751_),
    .C(_0752_),
    .A(_0746_),
    .Y(_0753_));
 sg13g2_buf_2 _3591_ (.A(_0753_),
    .X(_0754_));
 sg13g2_nor2_1 _3592_ (.A(_0245_),
    .B(_0615_),
    .Y(_0755_));
 sg13g2_nand2_1 _3593_ (.Y(_0756_),
    .A(_0673_),
    .B(_0744_));
 sg13g2_nand3_1 _3594_ (.B(_0675_),
    .C(_0672_),
    .A(_0670_),
    .Y(_0757_));
 sg13g2_nand2_1 _3595_ (.Y(_0758_),
    .A(_0756_),
    .B(_0757_));
 sg13g2_nand2_1 _3596_ (.Y(_0759_),
    .A(_0758_),
    .B(net13));
 sg13g2_nand2_1 _3597_ (.Y(_0760_),
    .A(_0673_),
    .B(_0007_));
 sg13g2_nand3_1 _3598_ (.B(_0008_),
    .C(_0672_),
    .A(_0670_),
    .Y(_0761_));
 sg13g2_nand3_1 _3599_ (.B(_0761_),
    .C(_0729_),
    .A(_0760_),
    .Y(_0762_));
 sg13g2_nand2_1 _3600_ (.Y(_0763_),
    .A(_0759_),
    .B(_0762_));
 sg13g2_nor2_1 _3601_ (.A(_0755_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_nand2_1 _3602_ (.Y(_0765_),
    .A(_0763_),
    .B(_0755_));
 sg13g2_o21ai_1 _3603_ (.B1(_0765_),
    .Y(_0766_),
    .A1(_0754_),
    .A2(_0764_));
 sg13g2_nand3_1 _3604_ (.B(_0745_),
    .C(net10),
    .A(_0743_),
    .Y(_0767_));
 sg13g2_nand3_1 _3605_ (.B(_0678_),
    .C(net13),
    .A(_0676_),
    .Y(_0768_));
 sg13g2_nor2_1 _3606_ (.A(_0211_),
    .B(_0615_),
    .Y(_0769_));
 sg13g2_nand3_1 _3607_ (.B(_0768_),
    .C(_0769_),
    .A(_0767_),
    .Y(_0770_));
 sg13g2_nand2_1 _3608_ (.Y(_0771_),
    .A(_0679_),
    .B(_0736_));
 sg13g2_nand2_1 _3609_ (.Y(_0772_),
    .A(net14),
    .B(_0008_));
 sg13g2_nand3_1 _3610_ (.B(_0009_),
    .C(net18),
    .A(net17),
    .Y(_0773_));
 sg13g2_nand3_1 _3611_ (.B(_0773_),
    .C(net10),
    .A(_0772_),
    .Y(_0774_));
 sg13g2_inv_1 _3612_ (.Y(_0775_),
    .A(_0769_));
 sg13g2_nand3_1 _3613_ (.B(_0774_),
    .C(_0775_),
    .A(_0771_),
    .Y(_0776_));
 sg13g2_nand2_1 _3614_ (.Y(_0777_),
    .A(_0770_),
    .B(_0776_));
 sg13g2_nand2_1 _3615_ (.Y(_0778_),
    .A(net14),
    .B(_0677_));
 sg13g2_inv_1 _3616_ (.Y(_0779_),
    .A(_0012_));
 sg13g2_nand3_1 _3617_ (.B(_0779_),
    .C(net18),
    .A(net17),
    .Y(_0780_));
 sg13g2_nand3_1 _3618_ (.B(_0780_),
    .C(net13),
    .A(_0778_),
    .Y(_0781_));
 sg13g2_nand3_1 _3619_ (.B(_0757_),
    .C(_0729_),
    .A(_0756_),
    .Y(_0782_));
 sg13g2_nand2_1 _3620_ (.Y(_0783_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_xnor2_1 _3621_ (.Y(_0784_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_nand2_1 _3622_ (.Y(_0785_),
    .A(_0494_),
    .B(_0784_));
 sg13g2_inv_1 _3623_ (.Y(_0786_),
    .A(_0785_));
 sg13g2_nand2_1 _3624_ (.Y(_0787_),
    .A(_0783_),
    .B(_0786_));
 sg13g2_nand3_1 _3625_ (.B(_0781_),
    .C(_0785_),
    .A(_0782_),
    .Y(_0788_));
 sg13g2_nand2_1 _3626_ (.Y(_0789_),
    .A(_0787_),
    .B(_0788_));
 sg13g2_nor2_1 _3627_ (.A(_0777_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_nand2_1 _3628_ (.Y(_0791_),
    .A(_0766_),
    .B(_0790_));
 sg13g2_nor2_1 _3629_ (.A(_0786_),
    .B(_0783_),
    .Y(_0792_));
 sg13g2_inv_1 _3630_ (.Y(_0793_),
    .A(_0770_));
 sg13g2_nor2_1 _3631_ (.A(_0792_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nor2b_1 _3632_ (.A(_0794_),
    .B_N(_0787_),
    .Y(_0795_));
 sg13g2_inv_1 _3633_ (.Y(_0796_),
    .A(_0795_));
 sg13g2_nand2_1 _3634_ (.Y(_0797_),
    .A(_0791_),
    .B(_0796_));
 sg13g2_nor2_1 _3635_ (.A(_0742_),
    .B(_0797_),
    .Y(_0798_));
 sg13g2_nand2_1 _3636_ (.Y(_0799_),
    .A(_0797_),
    .B(_0742_));
 sg13g2_nand2b_1 _3637_ (.Y(_0800_),
    .B(_0766_),
    .A_N(_0777_));
 sg13g2_inv_2 _3638_ (.Y(_0801_),
    .A(_0754_));
 sg13g2_inv_1 _3639_ (.Y(_0802_),
    .A(_0755_));
 sg13g2_nand3_1 _3640_ (.B(_0762_),
    .C(_0802_),
    .A(_0759_),
    .Y(_0803_));
 sg13g2_a21oi_1 _3641_ (.A1(_0759_),
    .A2(_0762_),
    .Y(_0804_),
    .B1(_0802_));
 sg13g2_a21oi_1 _3642_ (.A1(_0801_),
    .A2(_0803_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nand2_1 _3643_ (.Y(_0806_),
    .A(_0805_),
    .B(_0777_));
 sg13g2_nand2_1 _3644_ (.Y(_0807_),
    .A(_0800_),
    .B(_0806_));
 sg13g2_nand2_1 _3645_ (.Y(_0808_),
    .A(_0807_),
    .B(\main.demo._d___pip_24_1_2___stage___block_3_y[2] ));
 sg13g2_nand3b_1 _3646_ (.B(_0799_),
    .C(_0808_),
    .Y(_0809_),
    .A_N(_0798_));
 sg13g2_nand2b_1 _3647_ (.Y(_0810_),
    .B(_0789_),
    .A_N(\main.demo._d___pip_24_1_2___stage___block_3_y[3] ));
 sg13g2_nand3_1 _3648_ (.B(_0788_),
    .C(\main.demo._d___pip_24_1_2___stage___block_3_y[3] ),
    .A(_0787_),
    .Y(_0811_));
 sg13g2_nand2_1 _3649_ (.Y(_0812_),
    .A(_0810_),
    .B(_0811_));
 sg13g2_nand2_1 _3650_ (.Y(_0813_),
    .A(_0765_),
    .B(_0803_));
 sg13g2_nor2_1 _3651_ (.A(_0777_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_nand2_1 _3652_ (.Y(_0815_),
    .A(_0814_),
    .B(_0801_));
 sg13g2_a21oi_1 _3653_ (.A1(_0804_),
    .A2(_0776_),
    .Y(_0816_),
    .B1(_0793_));
 sg13g2_nand2_1 _3654_ (.Y(_0817_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_nand2b_1 _3655_ (.Y(_0818_),
    .B(_0817_),
    .A_N(_0812_));
 sg13g2_nand3_1 _3656_ (.B(_0812_),
    .C(_0816_),
    .A(_0815_),
    .Y(_0819_));
 sg13g2_nand2_1 _3657_ (.Y(_0820_),
    .A(_0818_),
    .B(_0819_));
 sg13g2_nand2_1 _3658_ (.Y(_0821_),
    .A(_0813_),
    .B(_0801_));
 sg13g2_nand3_1 _3659_ (.B(_0754_),
    .C(_0803_),
    .A(_0765_),
    .Y(_0822_));
 sg13g2_nand3_1 _3660_ (.B(_0822_),
    .C(\main.demo._d___pip_24_1_2___stage___block_3_y[1] ),
    .A(_0821_),
    .Y(_0823_));
 sg13g2_nand2_1 _3661_ (.Y(_0824_),
    .A(_0746_),
    .B(_0751_));
 sg13g2_inv_1 _3662_ (.Y(_0825_),
    .A(_0752_));
 sg13g2_nand2_1 _3663_ (.Y(_0826_),
    .A(_0824_),
    .B(_0825_));
 sg13g2_nand2_1 _3664_ (.Y(_0827_),
    .A(_0826_),
    .B(_0754_));
 sg13g2_xor2_1 _3665_ (.B(_0827_),
    .A(\main.demo._d___pip_24_1_2___stage___block_3_y[0] ),
    .X(_0828_));
 sg13g2_nand2_1 _3666_ (.Y(_0829_),
    .A(_0823_),
    .B(_0828_));
 sg13g2_nand2_1 _3667_ (.Y(_0830_),
    .A(_0821_),
    .B(_0822_));
 sg13g2_nand2b_1 _3668_ (.Y(_0831_),
    .B(_0830_),
    .A_N(\main.demo._d___pip_24_1_2___stage___block_3_y[1] ));
 sg13g2_nor2b_1 _3669_ (.A(_0829_),
    .B_N(_0831_),
    .Y(_0832_));
 sg13g2_nand3b_1 _3670_ (.B(_0800_),
    .C(_0806_),
    .Y(_0833_),
    .A_N(\main.demo._d___pip_24_1_2___stage___block_3_y[2] ));
 sg13g2_nand3_1 _3671_ (.B(_0832_),
    .C(_0833_),
    .A(_0820_),
    .Y(_0834_));
 sg13g2_nor2_1 _3672_ (.A(_0809_),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_nand2b_1 _3673_ (.Y(_0836_),
    .B(_0202_),
    .A_N(_0219_));
 sg13g2_xnor2_1 _3674_ (.Y(_0837_),
    .A(_0218_),
    .B(_0836_));
 sg13g2_nor2_1 _3675_ (.A(_0837_),
    .B(_0615_),
    .Y(_0838_));
 sg13g2_inv_2 _3676_ (.Y(_0839_),
    .A(net14));
 sg13g2_nand2_1 _3677_ (.Y(_0840_),
    .A(_0839_),
    .B(_0002_));
 sg13g2_nand2_1 _3678_ (.Y(_0841_),
    .A(net14),
    .B(_0001_));
 sg13g2_nand3_1 _3679_ (.B(net13),
    .C(_0841_),
    .A(_0840_),
    .Y(_0842_));
 sg13g2_nand3_1 _3680_ (.B(_0733_),
    .C(net10),
    .A(_0732_),
    .Y(_0843_));
 sg13g2_nand2_1 _3681_ (.Y(_0844_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_nand2b_1 _3682_ (.Y(_0845_),
    .B(_0844_),
    .A_N(_0838_));
 sg13g2_nand3_1 _3683_ (.B(_0838_),
    .C(_0843_),
    .A(_0842_),
    .Y(_0846_));
 sg13g2_nand2_1 _3684_ (.Y(_0847_),
    .A(_0845_),
    .B(_0846_));
 sg13g2_xnor2_1 _3685_ (.Y(_0848_),
    .A(\main.demo._d___pip_24_1_2___stage___block_3_y[6] ),
    .B(_0847_));
 sg13g2_nand2_1 _3686_ (.Y(_0849_),
    .A(net14),
    .B(_1809_));
 sg13g2_nand3_1 _3687_ (.B(_1807_),
    .C(net18),
    .A(net17),
    .Y(_0850_));
 sg13g2_nand3_1 _3688_ (.B(_0850_),
    .C(net13),
    .A(_0849_),
    .Y(_0851_));
 sg13g2_nand3_1 _3689_ (.B(_0780_),
    .C(net10),
    .A(_0778_),
    .Y(_0852_));
 sg13g2_nand2_1 _3690_ (.Y(_0853_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_xnor2_1 _3691_ (.Y(_0854_),
    .A(_0203_),
    .B(_0217_));
 sg13g2_nand2_1 _3692_ (.Y(_0855_),
    .A(_0494_),
    .B(_0854_));
 sg13g2_inv_1 _3693_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_nand2_1 _3694_ (.Y(_0857_),
    .A(_0853_),
    .B(_0856_));
 sg13g2_nand3_1 _3695_ (.B(_0852_),
    .C(_0855_),
    .A(_0851_),
    .Y(_0858_));
 sg13g2_nand2_1 _3696_ (.Y(_0859_),
    .A(_0857_),
    .B(_0858_));
 sg13g2_nor2_1 _3697_ (.A(_0859_),
    .B(_0741_),
    .Y(_0860_));
 sg13g2_inv_1 _3698_ (.Y(_0861_),
    .A(_0857_));
 sg13g2_a21oi_1 _3699_ (.A1(_0739_),
    .A2(_0858_),
    .Y(_0862_),
    .B1(_0861_));
 sg13g2_a21oi_1 _3700_ (.A1(_0795_),
    .A2(_0860_),
    .Y(_0863_),
    .B1(_0862_));
 sg13g2_nand3_1 _3701_ (.B(_0860_),
    .C(_0790_),
    .A(_0766_),
    .Y(_0864_));
 sg13g2_nand2_1 _3702_ (.Y(_0865_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_nand2b_1 _3703_ (.Y(_0866_),
    .B(_0865_),
    .A_N(_0848_));
 sg13g2_nand3_1 _3704_ (.B(_0864_),
    .C(_0848_),
    .A(_0863_),
    .Y(_0867_));
 sg13g2_nand2_1 _3705_ (.Y(_0868_),
    .A(_0866_),
    .B(_0867_));
 sg13g2_xor2_1 _3706_ (.B(_0859_),
    .A(\main.demo._d___pip_24_1_2___stage___block_3_y[5] ),
    .X(_0869_));
 sg13g2_nand2_1 _3707_ (.Y(_0870_),
    .A(_0792_),
    .B(_0740_));
 sg13g2_nand2_1 _3708_ (.Y(_0871_),
    .A(_0870_),
    .B(_0739_));
 sg13g2_inv_1 _3709_ (.Y(_0872_),
    .A(_0741_));
 sg13g2_xnor2_1 _3710_ (.Y(_0873_),
    .A(_0785_),
    .B(_0783_));
 sg13g2_nand2_1 _3711_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_));
 sg13g2_nor2_1 _3712_ (.A(_0816_),
    .B(_0874_),
    .Y(_0875_));
 sg13g2_nor2_1 _3713_ (.A(_0871_),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2_1 _3714_ (.A(_0789_),
    .B(_0741_),
    .Y(_0877_));
 sg13g2_nand3_1 _3715_ (.B(_0814_),
    .C(_0801_),
    .A(_0877_),
    .Y(_0878_));
 sg13g2_nand2_1 _3716_ (.Y(_0879_),
    .A(_0876_),
    .B(_0878_));
 sg13g2_xnor2_1 _3717_ (.Y(_0880_),
    .A(_0869_),
    .B(_0879_));
 sg13g2_nor2_1 _3718_ (.A(_0868_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nand2_1 _3719_ (.Y(_0882_),
    .A(_0268_),
    .B(_0266_));
 sg13g2_a21oi_1 _3720_ (.A1(_0220_),
    .A2(_0882_),
    .Y(_0883_),
    .B1(_0615_));
 sg13g2_o21ai_1 _3721_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0220_),
    .A2(_0882_));
 sg13g2_xor2_1 _3722_ (.B(_0884_),
    .A(\main.demo._d___pip_24_1_2___stage___block_3_y[7] ),
    .X(_0885_));
 sg13g2_nand2_1 _3723_ (.Y(_0886_),
    .A(_0839_),
    .B(_0003_));
 sg13g2_o21ai_1 _3724_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_1783_),
    .A2(_0839_));
 sg13g2_and3_1 _3725_ (.X(_0888_),
    .A(_0849_),
    .B(_0850_),
    .C(net10));
 sg13g2_a21oi_1 _3726_ (.A1(_0887_),
    .A2(net13),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_xnor2_1 _3727_ (.Y(_0890_),
    .A(_0885_),
    .B(_0889_));
 sg13g2_nor2_1 _3728_ (.A(_0859_),
    .B(_0847_),
    .Y(_0891_));
 sg13g2_nor2b_1 _3729_ (.A(_0874_),
    .B_N(_0891_),
    .Y(_0892_));
 sg13g2_nand2_1 _3730_ (.Y(_0893_),
    .A(_0817_),
    .B(_0892_));
 sg13g2_nand2b_1 _3731_ (.Y(_0894_),
    .B(_0846_),
    .A_N(_0858_));
 sg13g2_nand2_1 _3732_ (.Y(_0895_),
    .A(_0894_),
    .B(_0845_));
 sg13g2_a21oi_1 _3733_ (.A1(_0891_),
    .A2(_0871_),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_nand2_1 _3734_ (.Y(_0897_),
    .A(_0893_),
    .B(_0896_));
 sg13g2_xnor2_1 _3735_ (.Y(_0898_),
    .A(_0890_),
    .B(_0897_));
 sg13g2_nand4_1 _3736_ (.B(_0881_),
    .C(net10),
    .A(_0835_),
    .Y(_0899_),
    .D(_0898_));
 sg13g2_inv_1 _3737_ (.Y(_0900_),
    .A(\main.demo._q___pip_24_1_2___stage___block_3_s[1] ));
 sg13g2_inv_1 _3738_ (.Y(_0901_),
    .A(\main.demo._w_vga_active ));
 sg13g2_a21oi_1 _3739_ (.A1(_0899_),
    .A2(_0900_),
    .Y(_0018_),
    .B1(_0901_));
 sg13g2_nand2_1 _3740_ (.Y(_0902_),
    .A(net10),
    .B(_0839_));
 sg13g2_nand4_1 _3741_ (.B(_0881_),
    .C(_0898_),
    .A(_0835_),
    .Y(_0903_),
    .D(_0902_));
 sg13g2_inv_1 _3742_ (.Y(_0904_),
    .A(\main.demo._q___pip_24_1_2___stage___block_3_s[0] ));
 sg13g2_a21oi_1 _3743_ (.A1(_0903_),
    .A2(_0904_),
    .Y(_0019_),
    .B1(_0901_));
 sg13g2_nor2b_1 _3744_ (.A(\main._w_demo_video_vs ),
    .B_N(\main.demo._q_prev_vs ),
    .Y(_0905_));
 sg13g2_buf_2 _3745_ (.A(_0905_),
    .X(_0906_));
 sg13g2_buf_1 _3746_ (.A(rst_n_q),
    .X(_0907_));
 sg13g2_buf_1 _3747_ (.A(net34),
    .X(_0908_));
 sg13g2_o21ai_1 _3748_ (.B1(net33),
    .Y(_0909_),
    .A1(_1489_),
    .A2(_0906_));
 sg13g2_a21oi_1 _3749_ (.A1(_0747_),
    .A2(_0906_),
    .Y(_0022_),
    .B1(_0909_));
 sg13g2_inv_1 _3750_ (.Y(_0910_),
    .A(_0907_));
 sg13g2_buf_1 _3751_ (.A(_0910_),
    .X(_0911_));
 sg13g2_buf_1 _3752_ (.A(net31),
    .X(_0912_));
 sg13g2_inv_1 _3753_ (.Y(_0913_),
    .A(_0906_));
 sg13g2_nor3_1 _3754_ (.A(_1490_),
    .B(_1493_),
    .C(_0913_),
    .Y(_0914_));
 sg13g2_nand2_1 _3755_ (.Y(_0915_),
    .A(_0914_),
    .B(_1496_));
 sg13g2_nor2_1 _3756_ (.A(_1468_),
    .B(_0915_),
    .Y(_0916_));
 sg13g2_nand2_1 _3757_ (.Y(_0917_),
    .A(_0916_),
    .B(_1464_));
 sg13g2_nor2_1 _3758_ (.A(_1476_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_inv_1 _3759_ (.Y(_0919_),
    .A(_0918_));
 sg13g2_nor2_1 _3760_ (.A(_1508_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_inv_1 _3761_ (.Y(_0921_),
    .A(_0920_));
 sg13g2_nor2_1 _3762_ (.A(_1521_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_inv_1 _3763_ (.Y(_0923_),
    .A(_0922_));
 sg13g2_nor3_1 _3764_ (.A(_1455_),
    .B(_1447_),
    .C(_0923_),
    .Y(_0924_));
 sg13g2_nor2_1 _3765_ (.A(_1440_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nand2_1 _3766_ (.Y(_0926_),
    .A(_0924_),
    .B(_1440_));
 sg13g2_inv_1 _3767_ (.Y(_0927_),
    .A(_0926_));
 sg13g2_nor3_1 _3768_ (.A(net24),
    .B(_0925_),
    .C(_0927_),
    .Y(_0023_));
 sg13g2_nor2_1 _3769_ (.A(_1513_),
    .B(_0926_),
    .Y(_0928_));
 sg13g2_nor2_1 _3770_ (.A(_1436_),
    .B(_0927_),
    .Y(_0929_));
 sg13g2_nor3_1 _3771_ (.A(net24),
    .B(_0928_),
    .C(_0929_),
    .Y(_0024_));
 sg13g2_nor2_1 _3772_ (.A(_1433_),
    .B(_0928_),
    .Y(_0930_));
 sg13g2_nand2_1 _3773_ (.Y(_0931_),
    .A(_0928_),
    .B(_1433_));
 sg13g2_inv_1 _3774_ (.Y(_0932_),
    .A(_0931_));
 sg13g2_nor3_1 _3775_ (.A(net24),
    .B(_0930_),
    .C(_0932_),
    .Y(_0025_));
 sg13g2_nor2_1 _3776_ (.A(_1427_),
    .B(_0931_),
    .Y(_0933_));
 sg13g2_nor2_1 _3777_ (.A(\main.demo._q_frame[13] ),
    .B(_0932_),
    .Y(_0934_));
 sg13g2_nor3_1 _3778_ (.A(net24),
    .B(_0933_),
    .C(_0934_),
    .Y(_0026_));
 sg13g2_nor2_1 _3779_ (.A(_1420_),
    .B(_0933_),
    .Y(_0935_));
 sg13g2_nand2_1 _3780_ (.Y(_0936_),
    .A(_0933_),
    .B(_1420_));
 sg13g2_inv_1 _3781_ (.Y(_0937_),
    .A(_0936_));
 sg13g2_nor3_1 _3782_ (.A(net24),
    .B(_0935_),
    .C(_0937_),
    .Y(_0027_));
 sg13g2_o21ai_1 _3783_ (.B1(net33),
    .Y(_0938_),
    .A1(_0411_),
    .A2(_0936_));
 sg13g2_a21oi_1 _3784_ (.A1(_0411_),
    .A2(_0936_),
    .Y(_0028_),
    .B1(_0938_));
 sg13g2_buf_1 _3785_ (.A(net31),
    .X(_0939_));
 sg13g2_a21oi_1 _3786_ (.A1(_0906_),
    .A2(_1489_),
    .Y(_0940_),
    .B1(_1486_));
 sg13g2_nor3_1 _3787_ (.A(net23),
    .B(_0940_),
    .C(_0914_),
    .Y(_0029_));
 sg13g2_nor2_1 _3788_ (.A(_1496_),
    .B(_0914_),
    .Y(_0941_));
 sg13g2_inv_1 _3789_ (.Y(_0942_),
    .A(_0915_));
 sg13g2_nor3_1 _3790_ (.A(net23),
    .B(_0941_),
    .C(_0942_),
    .Y(_0030_));
 sg13g2_nor2_1 _3791_ (.A(_1467_),
    .B(_0942_),
    .Y(_0943_));
 sg13g2_nor3_1 _3792_ (.A(net23),
    .B(_0916_),
    .C(_0943_),
    .Y(_0031_));
 sg13g2_nor2_1 _3793_ (.A(_1464_),
    .B(_0916_),
    .Y(_0944_));
 sg13g2_inv_1 _3794_ (.Y(_0945_),
    .A(_0917_));
 sg13g2_nor3_1 _3795_ (.A(net23),
    .B(_0944_),
    .C(_0945_),
    .Y(_0032_));
 sg13g2_nor2_1 _3796_ (.A(_1475_),
    .B(_0945_),
    .Y(_0946_));
 sg13g2_nor3_1 _3797_ (.A(net23),
    .B(_0918_),
    .C(_0946_),
    .Y(_0033_));
 sg13g2_nor2_1 _3798_ (.A(_1481_),
    .B(_0918_),
    .Y(_0947_));
 sg13g2_nor3_1 _3799_ (.A(_0939_),
    .B(_0947_),
    .C(_0920_),
    .Y(_0034_));
 sg13g2_nor2_1 _3800_ (.A(_1460_),
    .B(_0920_),
    .Y(_0948_));
 sg13g2_nor3_1 _3801_ (.A(_0939_),
    .B(_0948_),
    .C(_0922_),
    .Y(_0035_));
 sg13g2_nor2_1 _3802_ (.A(_1454_),
    .B(_0922_),
    .Y(_0949_));
 sg13g2_nor2_1 _3803_ (.A(_1455_),
    .B(_0923_),
    .Y(_0950_));
 sg13g2_nor3_1 _3804_ (.A(net23),
    .B(_0949_),
    .C(_0950_),
    .Y(_0036_));
 sg13g2_nor2_1 _3805_ (.A(\main.demo._q_frame[9] ),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_nor3_1 _3806_ (.A(net23),
    .B(_0924_),
    .C(_0951_),
    .Y(_0037_));
 sg13g2_inv_1 _3807_ (.Y(_0952_),
    .A(_1491_));
 sg13g2_nor2_1 _3808_ (.A(_1616_),
    .B(_1620_),
    .Y(_0953_));
 sg13g2_inv_1 _3809_ (.Y(_0954_),
    .A(_1632_));
 sg13g2_nand3_1 _3810_ (.B(_1587_),
    .C(_0906_),
    .A(_1488_),
    .Y(_0955_));
 sg13g2_nor3_1 _3811_ (.A(_1598_),
    .B(_0955_),
    .C(_1585_),
    .Y(_0956_));
 sg13g2_nand4_1 _3812_ (.B(_1624_),
    .C(_0954_),
    .A(_0953_),
    .Y(_0957_),
    .D(_0956_));
 sg13g2_nand2_1 _3813_ (.Y(_0958_),
    .A(_1643_),
    .B(_1636_));
 sg13g2_nor2b_1 _3814_ (.A(_1426_),
    .B_N(_1419_),
    .Y(_0959_));
 sg13g2_nor2_1 _3815_ (.A(\main.demo._q_modulo_0[15] ),
    .B(_0411_),
    .Y(_0960_));
 sg13g2_a221oi_1 _3816_ (.B2(_0959_),
    .C1(_0960_),
    .B1(_1562_),
    .A1(_1422_),
    .Y(_0961_),
    .A2(_1419_));
 sg13g2_nor3_1 _3817_ (.A(_0957_),
    .B(_0958_),
    .C(_0961_),
    .Y(_0962_));
 sg13g2_nand3_1 _3818_ (.B(_1573_),
    .C(_0962_),
    .A(_1570_),
    .Y(_0963_));
 sg13g2_buf_1 _3819_ (.A(_0963_),
    .X(_0964_));
 sg13g2_buf_1 _3820_ (.A(_0964_),
    .X(_0965_));
 sg13g2_o21ai_1 _3821_ (.B1(net33),
    .Y(_0966_),
    .A1(_0015_),
    .A2(_0965_));
 sg13g2_a21oi_1 _3822_ (.A1(_0952_),
    .A2(_0965_),
    .Y(_0038_),
    .B1(_0966_));
 sg13g2_nand4_1 _3823_ (.B(_1487_),
    .C(\main.demo._q_modulo_0[2] ),
    .A(_1491_),
    .Y(_0967_),
    .D(\main.demo._q_modulo_0[3] ));
 sg13g2_nor2_1 _3824_ (.A(_1465_),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_inv_1 _3825_ (.Y(_0969_),
    .A(_0968_));
 sg13g2_inv_1 _3826_ (.Y(_0970_),
    .A(_1482_));
 sg13g2_a21oi_1 _3827_ (.A1(_0969_),
    .A2(_1478_),
    .Y(_0971_),
    .B1(_0970_));
 sg13g2_nand2_1 _3828_ (.Y(_0972_),
    .A(_0971_),
    .B(_1461_));
 sg13g2_inv_1 _3829_ (.Y(_0973_),
    .A(_0972_));
 sg13g2_nor2_1 _3830_ (.A(\main.demo._q_modulo_0[8] ),
    .B(\main.demo._q_modulo_0[9] ),
    .Y(_0974_));
 sg13g2_nor2b_1 _3831_ (.A(_0973_),
    .B_N(_0974_),
    .Y(_0975_));
 sg13g2_o21ai_1 _3832_ (.B1(_1443_),
    .Y(_0976_),
    .A1(_0975_),
    .A2(net20));
 sg13g2_nor3_1 _3833_ (.A(_1443_),
    .B(_0975_),
    .C(_0964_),
    .Y(_0977_));
 sg13g2_inv_1 _3834_ (.Y(_0978_),
    .A(_0977_));
 sg13g2_and3_1 _3835_ (.X(_0039_),
    .A(_0976_),
    .B(_0978_),
    .C(net33));
 sg13g2_nor2_1 _3836_ (.A(\main.demo._q_modulo_0[11] ),
    .B(_0977_),
    .Y(_0979_));
 sg13g2_inv_1 _3837_ (.Y(_0980_),
    .A(\main.demo._q_modulo_0[11] ));
 sg13g2_nor2_1 _3838_ (.A(_0980_),
    .B(_0978_),
    .Y(_0981_));
 sg13g2_nor3_1 _3839_ (.A(net23),
    .B(_0979_),
    .C(_0981_),
    .Y(_0040_));
 sg13g2_buf_1 _3840_ (.A(net31),
    .X(_0982_));
 sg13g2_nor2_1 _3841_ (.A(_1434_),
    .B(_0981_),
    .Y(_0983_));
 sg13g2_nand2_1 _3842_ (.Y(_0984_),
    .A(_0981_),
    .B(_1434_));
 sg13g2_inv_1 _3843_ (.Y(_0985_),
    .A(_0984_));
 sg13g2_nor3_1 _3844_ (.A(net22),
    .B(_0983_),
    .C(_0985_),
    .Y(_0041_));
 sg13g2_o21ai_1 _3845_ (.B1(net33),
    .Y(_0986_),
    .A1(_1429_),
    .A2(_0984_));
 sg13g2_a21oi_1 _3846_ (.A1(_1429_),
    .A2(_0984_),
    .Y(_0042_),
    .B1(_0986_));
 sg13g2_nand2_1 _3847_ (.Y(_0987_),
    .A(_1482_),
    .B(_1461_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \main._q_uo[2]$_SDFF_PN0__56  (.L_HI(net56));
 sg13g2_buf_1 _3850_ (.A(net40),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3851_ (.A(net41),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3852_ (.A(net42),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3853_ (.A(net43),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3854_ (.A(net44),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3855_ (.A(net45),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3856_ (.A(net46),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3857_ (.A(net47),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3858_ (.A(net48),
    .X(uio_out[0]));
 sg13g2_buf_1 _3859_ (.A(net49),
    .X(uio_out[1]));
 sg13g2_buf_1 _3860_ (.A(net50),
    .X(uio_out[2]));
 sg13g2_buf_1 _3861_ (.A(net51),
    .X(uio_out[3]));
 sg13g2_buf_1 _3862_ (.A(net52),
    .X(uio_out[4]));
 sg13g2_buf_1 _3863_ (.A(net53),
    .X(uio_out[5]));
 sg13g2_buf_1 _3864_ (.A(net54),
    .X(uio_out[6]));
 sg13g2_buf_1 _3865_ (.A(net55),
    .X(uio_out[7]));
 sg13g2_buf_1 _3866_ (.A(net4),
    .X(net2));
 sg13g2_buf_1 _3867_ (.A(net4),
    .X(net3));
 sg13g2_buf_1 _3868_ (.A(net8),
    .X(net6));
 sg13g2_buf_1 _3869_ (.A(net8),
    .X(net7));
 sg13g2_dfrbp_1 \main._q_uo[2]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net56),
    .D(_0018_),
    .Q_N(_1973_),
    .Q(net4));
 sg13g2_dfrbp_1 \main._q_uo[3]$_DFF_P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net57),
    .D(\main._w_demo_video_vs ),
    .Q_N(_1972_),
    .Q(net5));
 sg13g2_dfrbp_1 \main._q_uo[6]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net58),
    .D(_0019_),
    .Q_N(_1974_),
    .Q(net8));
 sg13g2_dfrbp_1 \main._q_uo[7]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net59),
    .D(\main._w_demo_video_hs ),
    .Q_N(_1975_),
    .Q(net9));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[0]$_DFF_P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net60),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[0] ),
    .Q_N(_1976_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[1]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net61),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[1] ),
    .Q_N(_1977_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[2]$_DFF_P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net62),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[2] ),
    .Q_N(_1978_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[3]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[3] ),
    .Q_N(_1979_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[4]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net64),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[4] ),
    .Q_N(_1980_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[5]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net65),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[5] ),
    .Q_N(_1981_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[6]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net66),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[6] ),
    .Q_N(_1982_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_1___stage___block_3_y[7]$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net67),
    .D(\main.demo._t___pip_24_1_0___stage___block_3_y[7] ),
    .Q_N(_1971_),
    .Q(\main.demo._d___pip_24_1_1___stage___block_3_y[7] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_s[0]$_SDFF_PP0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net68),
    .D(_0020_),
    .Q_N(_1970_),
    .Q(\main.demo._q___pip_24_1_2___stage___block_3_s[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_s[1]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net69),
    .D(_0021_),
    .Q_N(_1983_),
    .Q(\main.demo._q___pip_24_1_2___stage___block_3_s[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[0]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net70),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[0] ),
    .Q_N(_1984_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[1]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net71),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[1] ),
    .Q_N(_1985_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[2]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net72),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[2] ),
    .Q_N(_1986_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[3]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net73),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[3] ),
    .Q_N(_1987_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[3] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[4]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net74),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[4] ),
    .Q_N(_1988_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[4] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[5]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net75),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[5] ),
    .Q_N(_1989_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[5] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[6]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net76),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[6] ),
    .Q_N(_1990_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[6] ));
 sg13g2_dfrbp_1 \main.demo._q___pip_24_1_2___stage___block_3_y[7]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net77),
    .D(\main.demo._d___pip_24_1_1___stage___block_3_y[7] ),
    .Q_N(_1969_),
    .Q(\main.demo._d___pip_24_1_2___stage___block_3_y[7] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[0]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net78),
    .D(_0022_),
    .Q_N(_0017_),
    .Q(\main.demo._q_frame[0] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[10]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net79),
    .D(_0023_),
    .Q_N(_0003_),
    .Q(\main.demo._q_frame[10] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[11]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net80),
    .D(_0024_),
    .Q_N(_1968_),
    .Q(\main.demo._q_frame[11] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[12]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net81),
    .D(_0025_),
    .Q_N(_1967_),
    .Q(\main.demo._q_frame[12] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[13]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net82),
    .D(_0026_),
    .Q_N(_1966_),
    .Q(\main.demo._q_frame[13] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[14]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net83),
    .D(_0027_),
    .Q_N(_1965_),
    .Q(\main.demo._q_frame[14] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[15]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net84),
    .D(_0028_),
    .Q_N(_1964_),
    .Q(\main.demo._q_frame[15] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[1]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net85),
    .D(_0029_),
    .Q_N(_0007_),
    .Q(\main.demo._q_frame[1] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[2]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net86),
    .D(_0030_),
    .Q_N(_0008_),
    .Q(\main.demo._q_frame[2] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[3]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net87),
    .D(_0031_),
    .Q_N(_0009_),
    .Q(\main.demo._q_frame[3] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[4]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net88),
    .D(_0032_),
    .Q_N(_0010_),
    .Q(\main.demo._q_frame[4] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[5]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net89),
    .D(_0033_),
    .Q_N(_0011_),
    .Q(\main.demo._q_frame[5] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[6]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net90),
    .D(_0034_),
    .Q_N(_0012_),
    .Q(\main.demo._q_frame[6] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[7]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net91),
    .D(_0035_),
    .Q_N(_0000_),
    .Q(\main.demo._q_frame[7] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[8]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net92),
    .D(_0036_),
    .Q_N(_0001_),
    .Q(\main.demo._q_frame[8] ));
 sg13g2_dfrbp_1 \main.demo._q_frame[9]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net93),
    .D(_0037_),
    .Q_N(_0002_),
    .Q(\main.demo._q_frame[9] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[0]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net94),
    .D(_0038_),
    .Q_N(_0015_),
    .Q(\main.demo._q_modulo_0[0] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[10]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net95),
    .D(_0039_),
    .Q_N(_1963_),
    .Q(\main.demo._q_modulo_0[10] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[11]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net96),
    .D(_0040_),
    .Q_N(_1962_),
    .Q(\main.demo._q_modulo_0[11] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[12]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net97),
    .D(_0041_),
    .Q_N(_1961_),
    .Q(\main.demo._q_modulo_0[12] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[13]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net98),
    .D(_0042_),
    .Q_N(_1960_),
    .Q(\main.demo._q_modulo_0[13] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[14]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net99),
    .D(_0043_),
    .Q_N(_1959_),
    .Q(\main.demo._q_modulo_0[14] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[15]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net100),
    .D(_0044_),
    .Q_N(_1958_),
    .Q(\main.demo._q_modulo_0[15] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[1]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net101),
    .D(_0045_),
    .Q_N(_1957_),
    .Q(\main.demo._q_modulo_0[1] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[2]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net102),
    .D(_0046_),
    .Q_N(_1956_),
    .Q(\main.demo._q_modulo_0[2] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[3]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net103),
    .D(_0047_),
    .Q_N(_1955_),
    .Q(\main.demo._q_modulo_0[3] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[4]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net104),
    .D(_0048_),
    .Q_N(_1954_),
    .Q(\main.demo._q_modulo_0[4] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[5]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net105),
    .D(_0049_),
    .Q_N(_0006_),
    .Q(\main.demo._q_modulo_0[5] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[6]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net106),
    .D(_0050_),
    .Q_N(_1953_),
    .Q(\main.demo._q_modulo_0[6] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[7]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net107),
    .D(_0051_),
    .Q_N(_1952_),
    .Q(\main.demo._q_modulo_0[7] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[8]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net108),
    .D(_0052_),
    .Q_N(_1951_),
    .Q(\main.demo._q_modulo_0[8] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_0[9]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net109),
    .D(_0053_),
    .Q_N(_1950_),
    .Q(\main.demo._q_modulo_0[9] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[0]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net110),
    .D(_0054_),
    .Q_N(_0016_),
    .Q(\main.demo._q_modulo_1[0] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[10]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net111),
    .D(_0055_),
    .Q_N(_1949_),
    .Q(\main.demo._q_modulo_1[10] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[11]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net112),
    .D(_0056_),
    .Q_N(_1948_),
    .Q(\main.demo._q_modulo_1[11] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[12]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net113),
    .D(_0057_),
    .Q_N(_1947_),
    .Q(\main.demo._q_modulo_1[12] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[13]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net114),
    .D(_0058_),
    .Q_N(_1946_),
    .Q(\main.demo._q_modulo_1[13] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[14]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net115),
    .D(_0059_),
    .Q_N(_1945_),
    .Q(\main.demo._q_modulo_1[14] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[15]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net116),
    .D(_0060_),
    .Q_N(_1944_),
    .Q(\main.demo._q_modulo_1[15] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net117),
    .D(_0061_),
    .Q_N(_1943_),
    .Q(\main.demo._q_modulo_1[1] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[2]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net118),
    .D(_0062_),
    .Q_N(_1942_),
    .Q(\main.demo._q_modulo_1[2] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[3]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net119),
    .D(_0063_),
    .Q_N(_1941_),
    .Q(\main.demo._q_modulo_1[3] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[4]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net120),
    .D(_0064_),
    .Q_N(_1940_),
    .Q(\main.demo._q_modulo_1[4] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[5]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net121),
    .D(_0065_),
    .Q_N(_0005_),
    .Q(\main.demo._q_modulo_1[5] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[6]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net122),
    .D(_0066_),
    .Q_N(_1939_),
    .Q(\main.demo._q_modulo_1[6] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[7]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net123),
    .D(_0067_),
    .Q_N(_1938_),
    .Q(\main.demo._q_modulo_1[7] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[8]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net124),
    .D(_0068_),
    .Q_N(_1937_),
    .Q(\main.demo._q_modulo_1[8] ));
 sg13g2_dfrbp_1 \main.demo._q_modulo_1[9]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net125),
    .D(_0069_),
    .Q_N(_1936_),
    .Q(\main.demo._q_modulo_1[9] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[0]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net126),
    .D(_0070_),
    .Q_N(_1935_),
    .Q(\main.demo._q_pix_x[0] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[1]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net127),
    .D(_0071_),
    .Q_N(_1934_),
    .Q(\main.demo._q_pix_x[1] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[2]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net128),
    .D(_0072_),
    .Q_N(_1933_),
    .Q(\main.demo._q_pix_x[2] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[3]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net129),
    .D(_0073_),
    .Q_N(_1932_),
    .Q(\main.demo._q_pix_x[3] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[4]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0074_),
    .Q_N(_1931_),
    .Q(\main.demo._q_pix_x[4] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[5]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net131),
    .D(_0075_),
    .Q_N(_1930_),
    .Q(\main.demo._q_pix_x[5] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[6]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net132),
    .D(_0076_),
    .Q_N(_1929_),
    .Q(\main.demo._q_pix_x[6] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[7]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0077_),
    .Q_N(_1928_),
    .Q(\main.demo._q_pix_x[7] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[8]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net134),
    .D(_0078_),
    .Q_N(_1927_),
    .Q(\main.demo._q_pix_x[8] ));
 sg13g2_dfrbp_1 \main.demo._q_pix_x[9]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net135),
    .D(_0079_),
    .Q_N(_1926_),
    .Q(\main.demo._q_pix_x[9] ));
 sg13g2_dfrbp_1 \main.demo._q_prev_hs$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net136),
    .D(_0080_),
    .Q_N(_1925_),
    .Q(\main.demo._q_prev_hs ));
 sg13g2_dfrbp_1 \main.demo._q_prev_vs$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net137),
    .D(_0081_),
    .Q_N(_1924_),
    .Q(\main.demo._q_prev_vs ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[0]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0082_),
    .Q_N(_0013_),
    .Q(\main.demo._q_rand_0[0] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[10]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net139),
    .D(_0083_),
    .Q_N(_1923_),
    .Q(\main.demo._q_rand_0[10] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[11]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net140),
    .D(_0084_),
    .Q_N(_1922_),
    .Q(\main.demo._q_rand_0[11] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[1]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net141),
    .D(_0085_),
    .Q_N(_1921_),
    .Q(\main.demo._q_rand_0[1] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[2]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net142),
    .D(_0086_),
    .Q_N(_1920_),
    .Q(\main.demo._q_rand_0[2] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[3]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net143),
    .D(_0087_),
    .Q_N(_1919_),
    .Q(\main.demo._q_rand_0[3] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[4]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net144),
    .D(_0088_),
    .Q_N(_1918_),
    .Q(\main.demo._q_rand_0[4] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[5]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(_0089_),
    .Q_N(_1917_),
    .Q(\main.demo._q_rand_0[5] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[6]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net146),
    .D(_0090_),
    .Q_N(_1916_),
    .Q(\main.demo._q_rand_0[6] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[7]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0091_),
    .Q_N(_1915_),
    .Q(\main.demo._q_rand_0[7] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[8]$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net148),
    .D(_0092_),
    .Q_N(_1914_),
    .Q(\main.demo._q_rand_0[8] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_0[9]$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net149),
    .D(_0093_),
    .Q_N(_1913_),
    .Q(\main.demo._q_rand_0[9] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[0]$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net150),
    .D(_0094_),
    .Q_N(_0014_),
    .Q(\main.demo._q_rand_1[0] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[10]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(_0095_),
    .Q_N(_1912_),
    .Q(\main.demo._q_rand_1[10] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[11]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net152),
    .D(_0096_),
    .Q_N(_1911_),
    .Q(\main.demo._q_rand_1[11] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[1]$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net153),
    .D(_0097_),
    .Q_N(_1910_),
    .Q(\main.demo._q_rand_1[1] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[2]$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net154),
    .D(_0098_),
    .Q_N(_1909_),
    .Q(\main.demo._q_rand_1[2] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[3]$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net155),
    .D(_0099_),
    .Q_N(_1908_),
    .Q(\main.demo._q_rand_1[3] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[4]$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net156),
    .D(_0100_),
    .Q_N(_1907_),
    .Q(\main.demo._q_rand_1[4] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[5]$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net157),
    .D(_0101_),
    .Q_N(_1906_),
    .Q(\main.demo._q_rand_1[5] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[6]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net158),
    .D(_0102_),
    .Q_N(_1905_),
    .Q(\main.demo._q_rand_1[6] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[7]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net159),
    .D(_0103_),
    .Q_N(_1904_),
    .Q(\main.demo._q_rand_1[7] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[8]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net160),
    .D(_0104_),
    .Q_N(_1903_),
    .Q(\main.demo._q_rand_1[8] ));
 sg13g2_dfrbp_1 \main.demo._q_rand_1[9]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net161),
    .D(_0105_),
    .Q_N(_1991_),
    .Q(\main.demo._q_rand_1[9] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net162),
    .D(\main.demo.vga._d_active ),
    .Q_N(_1902_),
    .Q(\main.demo._w_vga_active ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active_h$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net163),
    .D(_0106_),
    .Q_N(_1901_),
    .Q(\main.demo.vga._q_active_h ));
 sg13g2_dfrbp_1 \main.demo.vga._q_active_v$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net164),
    .D(_0107_),
    .Q_N(_1900_),
    .Q(\main.demo.vga._q_active_v ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_hs$_SDFFE_PP0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net165),
    .D(_0108_),
    .Q_N(_1899_),
    .Q(\main._w_demo_video_hs ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_vs$_SDFFE_PP0N_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net166),
    .D(_0109_),
    .Q_N(_1898_),
    .Q(\main._w_demo_video_vs ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[0]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net167),
    .D(_0110_),
    .Q_N(_1897_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[1]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net168),
    .D(_0111_),
    .Q_N(_1896_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[2]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net169),
    .D(_0112_),
    .Q_N(_1895_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[3]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net170),
    .D(_0113_),
    .Q_N(_1894_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[4]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net171),
    .D(_0114_),
    .Q_N(_1893_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[5]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net172),
    .D(_0115_),
    .Q_N(_1892_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[6]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net173),
    .D(_0116_),
    .Q_N(_1891_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_vga_y[7]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net174),
    .D(_0117_),
    .Q_N(_1890_),
    .Q(\main.demo._t___pip_24_1_0___stage___block_3_y[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[0]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net175),
    .D(_0118_),
    .Q_N(_1889_),
    .Q(\main.demo.vga._q_xcount[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[10]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net176),
    .D(_0119_),
    .Q_N(_1888_),
    .Q(\main.demo.vga._q_xcount[10] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[1]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net177),
    .D(_0120_),
    .Q_N(_1887_),
    .Q(\main.demo.vga._q_xcount[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[2]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net178),
    .D(_0121_),
    .Q_N(_1886_),
    .Q(\main.demo.vga._q_xcount[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[3]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net179),
    .D(_0122_),
    .Q_N(_1885_),
    .Q(\main.demo.vga._q_xcount[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[4]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net180),
    .D(_0123_),
    .Q_N(_1884_),
    .Q(\main.demo.vga._q_xcount[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[5]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net181),
    .D(_0124_),
    .Q_N(_1883_),
    .Q(\main.demo.vga._q_xcount[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[6]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net182),
    .D(_0125_),
    .Q_N(_1882_),
    .Q(\main.demo.vga._q_xcount[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[7]$_SDFF_PP0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net183),
    .D(_0126_),
    .Q_N(_1881_),
    .Q(\main.demo.vga._q_xcount[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[8]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net184),
    .D(_0127_),
    .Q_N(_1880_),
    .Q(\main.demo.vga._q_xcount[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_xcount[9]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net185),
    .D(_0128_),
    .Q_N(_1879_),
    .Q(\main.demo.vga._q_xcount[9] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[0]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net186),
    .D(_0129_),
    .Q_N(_1878_),
    .Q(\main.demo.vga._q_ycount[0] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[1]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net187),
    .D(_0130_),
    .Q_N(_1877_),
    .Q(\main.demo.vga._q_ycount[1] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[2]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net188),
    .D(_0131_),
    .Q_N(_1876_),
    .Q(\main.demo.vga._q_ycount[2] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[3]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net189),
    .D(_0132_),
    .Q_N(_1875_),
    .Q(\main.demo.vga._q_ycount[3] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[4]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net190),
    .D(_0133_),
    .Q_N(_1874_),
    .Q(\main.demo.vga._q_ycount[4] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[5]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net191),
    .D(_0134_),
    .Q_N(_1873_),
    .Q(\main.demo.vga._q_ycount[5] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[6]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net192),
    .D(_0135_),
    .Q_N(_1872_),
    .Q(\main.demo.vga._q_ycount[6] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[7]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net193),
    .D(_0136_),
    .Q_N(_1871_),
    .Q(\main.demo.vga._q_ycount[7] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[8]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net194),
    .D(_0137_),
    .Q_N(_1870_),
    .Q(\main.demo.vga._q_ycount[8] ));
 sg13g2_dfrbp_1 \main.demo.vga._q_ycount[9]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net195),
    .D(_0138_),
    .Q_N(_1992_),
    .Q(\main.demo.vga._d_vblank ));
 sg13g2_dfrbp_1 \rst_n_q$_DFF_P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net196),
    .D(net1),
    .Q_N(_0004_),
    .Q(rst_n_q));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_0730_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_1696_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_1684_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0736_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0674_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1691_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_1650_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0670_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0672_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_1034_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0965_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0597_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0982_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0939_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0912_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0608_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1099_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1098_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1095_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1076_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1017_),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(_0911_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1576_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0908_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0907_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0227_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0145_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0144_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0141_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1186_),
    .X(net39));
 sg13g2_tielo _3850__40 (.L_LO(net40));
 sg13g2_tielo _3851__41 (.L_LO(net41));
 sg13g2_tielo _3852__42 (.L_LO(net42));
 sg13g2_tielo _3853__43 (.L_LO(net43));
 sg13g2_tielo _3854__44 (.L_LO(net44));
 sg13g2_tielo _3855__45 (.L_LO(net45));
 sg13g2_tielo _3856__46 (.L_LO(net46));
 sg13g2_tielo _3857__47 (.L_LO(net47));
 sg13g2_tielo _3858__48 (.L_LO(net48));
 sg13g2_tielo _3859__49 (.L_LO(net49));
 sg13g2_tielo _3860__50 (.L_LO(net50));
 sg13g2_tielo _3861__51 (.L_LO(net51));
 sg13g2_tielo _3862__52 (.L_LO(net52));
 sg13g2_tielo _3863__53 (.L_LO(net53));
 sg13g2_tielo _3864__54 (.L_LO(net54));
 sg13g2_tielo _3865__55 (.L_LO(net55));
 sg13g2_tiehi \main._q_uo[3]$_DFF_P__57  (.L_HI(net57));
 sg13g2_tiehi \main._q_uo[6]$_SDFF_PN0__58  (.L_HI(net58));
 sg13g2_tiehi \main._q_uo[7]$_DFF_P__59  (.L_HI(net59));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[0]$_DFF_P__60  (.L_HI(net60));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[1]$_DFF_P__61  (.L_HI(net61));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[2]$_DFF_P__62  (.L_HI(net62));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[3]$_DFF_P__63  (.L_HI(net63));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[4]$_DFF_P__64  (.L_HI(net64));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[5]$_DFF_P__65  (.L_HI(net65));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[6]$_DFF_P__66  (.L_HI(net66));
 sg13g2_tiehi \main.demo._q___pip_24_1_1___stage___block_3_y[7]$_DFF_P__67  (.L_HI(net67));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_s[0]$_SDFF_PP0__68  (.L_HI(net68));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_s[1]$_SDFF_PP0__69  (.L_HI(net69));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[0]$_DFF_P__70  (.L_HI(net70));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[1]$_DFF_P__71  (.L_HI(net71));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[2]$_DFF_P__72  (.L_HI(net72));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[3]$_DFF_P__73  (.L_HI(net73));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[4]$_DFF_P__74  (.L_HI(net74));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[5]$_DFF_P__75  (.L_HI(net75));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[6]$_DFF_P__76  (.L_HI(net76));
 sg13g2_tiehi \main.demo._q___pip_24_1_2___stage___block_3_y[7]$_DFF_P__77  (.L_HI(net77));
 sg13g2_tiehi \main.demo._q_frame[0]$_SDFFE_PN0P__78  (.L_HI(net78));
 sg13g2_tiehi \main.demo._q_frame[10]$_SDFFE_PN0P__79  (.L_HI(net79));
 sg13g2_tiehi \main.demo._q_frame[11]$_SDFFE_PN0P__80  (.L_HI(net80));
 sg13g2_tiehi \main.demo._q_frame[12]$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_tiehi \main.demo._q_frame[13]$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \main.demo._q_frame[14]$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \main.demo._q_frame[15]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \main.demo._q_frame[1]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \main.demo._q_frame[2]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \main.demo._q_frame[3]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \main.demo._q_frame[4]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \main.demo._q_frame[5]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \main.demo._q_frame[6]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \main.demo._q_frame[7]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \main.demo._q_frame[8]$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \main.demo._q_frame[9]$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \main.demo._q_modulo_0[0]$_SDFFE_PN0P__94  (.L_HI(net94));
 sg13g2_tiehi \main.demo._q_modulo_0[10]$_SDFFE_PN0P__95  (.L_HI(net95));
 sg13g2_tiehi \main.demo._q_modulo_0[11]$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \main.demo._q_modulo_0[12]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \main.demo._q_modulo_0[13]$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \main.demo._q_modulo_0[14]$_SDFFE_PN0P__99  (.L_HI(net99));
 sg13g2_tiehi \main.demo._q_modulo_0[15]$_SDFFE_PN0P__100  (.L_HI(net100));
 sg13g2_tiehi \main.demo._q_modulo_0[1]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \main.demo._q_modulo_0[2]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \main.demo._q_modulo_0[3]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \main.demo._q_modulo_0[4]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \main.demo._q_modulo_0[5]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \main.demo._q_modulo_0[6]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \main.demo._q_modulo_0[7]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \main.demo._q_modulo_0[8]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \main.demo._q_modulo_0[9]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \main.demo._q_modulo_1[0]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \main.demo._q_modulo_1[10]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \main.demo._q_modulo_1[11]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \main.demo._q_modulo_1[12]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \main.demo._q_modulo_1[13]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \main.demo._q_modulo_1[14]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \main.demo._q_modulo_1[15]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \main.demo._q_modulo_1[1]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \main.demo._q_modulo_1[2]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \main.demo._q_modulo_1[3]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \main.demo._q_modulo_1[4]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \main.demo._q_modulo_1[5]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \main.demo._q_modulo_1[6]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \main.demo._q_modulo_1[7]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \main.demo._q_modulo_1[8]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \main.demo._q_modulo_1[9]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \main.demo._q_pix_x[0]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \main.demo._q_pix_x[1]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \main.demo._q_pix_x[2]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \main.demo._q_pix_x[3]$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \main.demo._q_pix_x[4]$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \main.demo._q_pix_x[5]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \main.demo._q_pix_x[6]$_SDFF_PN0__132  (.L_HI(net132));
 sg13g2_tiehi \main.demo._q_pix_x[7]$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \main.demo._q_pix_x[8]$_SDFF_PN0__134  (.L_HI(net134));
 sg13g2_tiehi \main.demo._q_pix_x[9]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \main.demo._q_prev_hs$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \main.demo._q_prev_vs$_SDFF_PN0__137  (.L_HI(net137));
 sg13g2_tiehi \main.demo._q_rand_0[0]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_tiehi \main.demo._q_rand_0[10]$_SDFF_PN0__139  (.L_HI(net139));
 sg13g2_tiehi \main.demo._q_rand_0[11]$_SDFF_PN0__140  (.L_HI(net140));
 sg13g2_tiehi \main.demo._q_rand_0[1]$_SDFF_PN0__141  (.L_HI(net141));
 sg13g2_tiehi \main.demo._q_rand_0[2]$_SDFF_PN0__142  (.L_HI(net142));
 sg13g2_tiehi \main.demo._q_rand_0[3]$_SDFF_PN0__143  (.L_HI(net143));
 sg13g2_tiehi \main.demo._q_rand_0[4]$_SDFF_PN0__144  (.L_HI(net144));
 sg13g2_tiehi \main.demo._q_rand_0[5]$_SDFF_PN0__145  (.L_HI(net145));
 sg13g2_tiehi \main.demo._q_rand_0[6]$_SDFF_PN0__146  (.L_HI(net146));
 sg13g2_tiehi \main.demo._q_rand_0[7]$_SDFF_PN0__147  (.L_HI(net147));
 sg13g2_tiehi \main.demo._q_rand_0[8]$_SDFF_PP0__148  (.L_HI(net148));
 sg13g2_tiehi \main.demo._q_rand_0[9]$_SDFF_PP0__149  (.L_HI(net149));
 sg13g2_tiehi \main.demo._q_rand_1[0]$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \main.demo._q_rand_1[10]$_SDFF_PN0__151  (.L_HI(net151));
 sg13g2_tiehi \main.demo._q_rand_1[11]$_SDFF_PN0__152  (.L_HI(net152));
 sg13g2_tiehi \main.demo._q_rand_1[1]$_SDFF_PN0__153  (.L_HI(net153));
 sg13g2_tiehi \main.demo._q_rand_1[2]$_SDFF_PN0__154  (.L_HI(net154));
 sg13g2_tiehi \main.demo._q_rand_1[3]$_SDFF_PN0__155  (.L_HI(net155));
 sg13g2_tiehi \main.demo._q_rand_1[4]$_SDFF_PN0__156  (.L_HI(net156));
 sg13g2_tiehi \main.demo._q_rand_1[5]$_SDFF_PN0__157  (.L_HI(net157));
 sg13g2_tiehi \main.demo._q_rand_1[6]$_SDFF_PN0__158  (.L_HI(net158));
 sg13g2_tiehi \main.demo._q_rand_1[7]$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \main.demo._q_rand_1[8]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \main.demo._q_rand_1[9]$_SDFF_PP0__161  (.L_HI(net161));
 sg13g2_tiehi \main.demo.vga._q_active$_DFF_P__162  (.L_HI(net162));
 sg13g2_tiehi \main.demo.vga._q_active_h$_SDFF_PN0__163  (.L_HI(net163));
 sg13g2_tiehi \main.demo.vga._q_active_v$_SDFF_PN0__164  (.L_HI(net164));
 sg13g2_tiehi \main.demo.vga._q_vga_hs$_SDFFE_PP0N__165  (.L_HI(net165));
 sg13g2_tiehi \main.demo.vga._q_vga_vs$_SDFFE_PP0N__166  (.L_HI(net166));
 sg13g2_tiehi \main.demo.vga._q_vga_y[0]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \main.demo.vga._q_vga_y[1]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \main.demo.vga._q_vga_y[2]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \main.demo.vga._q_vga_y[3]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \main.demo.vga._q_vga_y[4]$_SDFF_PP0__171  (.L_HI(net171));
 sg13g2_tiehi \main.demo.vga._q_vga_y[5]$_SDFF_PP0__172  (.L_HI(net172));
 sg13g2_tiehi \main.demo.vga._q_vga_y[6]$_SDFF_PP0__173  (.L_HI(net173));
 sg13g2_tiehi \main.demo.vga._q_vga_y[7]$_SDFF_PP0__174  (.L_HI(net174));
 sg13g2_tiehi \main.demo.vga._q_xcount[0]$_SDFF_PN0__175  (.L_HI(net175));
 sg13g2_tiehi \main.demo.vga._q_xcount[10]$_SDFF_PN0__176  (.L_HI(net176));
 sg13g2_tiehi \main.demo.vga._q_xcount[1]$_SDFF_PN0__177  (.L_HI(net177));
 sg13g2_tiehi \main.demo.vga._q_xcount[2]$_SDFF_PN0__178  (.L_HI(net178));
 sg13g2_tiehi \main.demo.vga._q_xcount[3]$_SDFF_PN0__179  (.L_HI(net179));
 sg13g2_tiehi \main.demo.vga._q_xcount[4]$_SDFF_PN0__180  (.L_HI(net180));
 sg13g2_tiehi \main.demo.vga._q_xcount[5]$_SDFF_PP0__181  (.L_HI(net181));
 sg13g2_tiehi \main.demo.vga._q_xcount[6]$_SDFF_PN0__182  (.L_HI(net182));
 sg13g2_tiehi \main.demo.vga._q_xcount[7]$_SDFF_PP0__183  (.L_HI(net183));
 sg13g2_tiehi \main.demo.vga._q_xcount[8]$_SDFF_PN0__184  (.L_HI(net184));
 sg13g2_tiehi \main.demo.vga._q_xcount[9]$_SDFF_PN0__185  (.L_HI(net185));
 sg13g2_tiehi \main.demo.vga._q_ycount[0]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \main.demo.vga._q_ycount[1]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \main.demo.vga._q_ycount[2]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \main.demo.vga._q_ycount[3]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \main.demo.vga._q_ycount[4]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \main.demo.vga._q_ycount[5]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \main.demo.vga._q_ycount[6]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \main.demo.vga._q_ycount[7]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \main.demo.vga._q_ycount[8]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \main.demo.vga._q_ycount[9]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \rst_n_q$_DFF_P__196  (.L_HI(net196));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(net1));
 sg13g2_antennanp ANTENNA_2 (.A(net1));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_decap_4 FILLER_1_277 ();
 sg13g2_fill_2 FILLER_1_281 ();
 sg13g2_fill_2 FILLER_1_286 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_1 FILLER_1_298 ();
 sg13g2_decap_4 FILLER_1_311 ();
 sg13g2_fill_2 FILLER_1_319 ();
 sg13g2_fill_1 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_fill_2 FILLER_1_332 ();
 sg13g2_fill_1 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_4 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_256 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_312 ();
 sg13g2_fill_2 FILLER_2_320 ();
 sg13g2_fill_1 FILLER_2_332 ();
 sg13g2_fill_1 FILLER_2_338 ();
 sg13g2_decap_4 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_266 ();
 sg13g2_fill_2 FILLER_3_284 ();
 sg13g2_fill_2 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_315 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_330 ();
 sg13g2_fill_1 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_4 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_235 ();
 sg13g2_fill_1 FILLER_4_244 ();
 sg13g2_fill_2 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_285 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_349 ();
 sg13g2_fill_2 FILLER_4_376 ();
 sg13g2_fill_2 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_80 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_decap_4 FILLER_5_89 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_fill_2 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_169 ();
 sg13g2_decap_8 FILLER_5_176 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_2 FILLER_5_331 ();
 sg13g2_fill_2 FILLER_5_337 ();
 sg13g2_fill_1 FILLER_5_373 ();
 sg13g2_fill_1 FILLER_5_403 ();
 sg13g2_fill_1 FILLER_5_418 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_51 ();
 sg13g2_fill_2 FILLER_6_65 ();
 sg13g2_fill_1 FILLER_6_85 ();
 sg13g2_fill_2 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_fill_2 FILLER_6_123 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_136 ();
 sg13g2_fill_2 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_155 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_decap_8 FILLER_6_180 ();
 sg13g2_decap_8 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_4 FILLER_6_229 ();
 sg13g2_fill_2 FILLER_6_233 ();
 sg13g2_fill_1 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_1 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_fill_2 FILLER_7_10 ();
 sg13g2_fill_2 FILLER_7_15 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_43 ();
 sg13g2_fill_1 FILLER_7_101 ();
 sg13g2_fill_1 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_fill_2 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_292 ();
 sg13g2_fill_1 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_319 ();
 sg13g2_fill_2 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_fill_1 FILLER_8_19 ();
 sg13g2_fill_1 FILLER_8_26 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_fill_1 FILLER_8_37 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_1 FILLER_8_54 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_fill_1 FILLER_8_173 ();
 sg13g2_fill_2 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_254 ();
 sg13g2_fill_1 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_fill_2 FILLER_8_376 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_fill_2 FILLER_9_317 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_fill_2 FILLER_9_375 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_1 FILLER_10_22 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_fill_2 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_2 FILLER_10_333 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_fill_1 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_354 ();
 sg13g2_fill_1 FILLER_10_395 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_406 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_fill_2 FILLER_11_148 ();
 sg13g2_fill_1 FILLER_11_166 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_369 ();
 sg13g2_fill_2 FILLER_11_398 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_1 FILLER_12_8 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_246 ();
 sg13g2_fill_1 FILLER_12_412 ();
 sg13g2_fill_1 FILLER_12_420 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_fill_1 FILLER_13_90 ();
 sg13g2_fill_2 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_223 ();
 sg13g2_fill_2 FILLER_13_270 ();
 sg13g2_fill_1 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_356 ();
 sg13g2_fill_2 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_8 FILLER_13_404 ();
 sg13g2_decap_8 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_fill_1 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_95 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_115 ();
 sg13g2_fill_2 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_decap_4 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_196 ();
 sg13g2_fill_1 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_8 FILLER_18_404 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_12 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_219 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_20_409 ();
 sg13g2_decap_4 FILLER_20_413 ();
 sg13g2_fill_2 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_425 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_396 ();
 sg13g2_fill_1 FILLER_21_425 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_383 ();
 sg13g2_fill_1 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_2 FILLER_26_356 ();
 sg13g2_fill_1 FILLER_27_9 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_2 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_fill_2 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_410 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_170 ();
endmodule
