module tt_um_hpretl_spi (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire clknet_0_clk;
 wire net106;
 wire \dac.accu1[0] ;
 wire \dac.accu1[10] ;
 wire \dac.accu1[11] ;
 wire \dac.accu1[12] ;
 wire \dac.accu1[13] ;
 wire \dac.accu1[14] ;
 wire \dac.accu1[15] ;
 wire \dac.accu1[1] ;
 wire \dac.accu1[2] ;
 wire \dac.accu1[3] ;
 wire \dac.accu1[4] ;
 wire \dac.accu1[5] ;
 wire \dac.accu1[6] ;
 wire \dac.accu1[7] ;
 wire \dac.accu1[8] ;
 wire \dac.accu1[9] ;
 wire \dac.accu2[0] ;
 wire \dac.accu2[10] ;
 wire \dac.accu2[11] ;
 wire \dac.accu2[12] ;
 wire \dac.accu2[13] ;
 wire \dac.accu2[14] ;
 wire \dac.accu2[15] ;
 wire \dac.accu2[1] ;
 wire \dac.accu2[2] ;
 wire \dac.accu2[3] ;
 wire \dac.accu2[4] ;
 wire \dac.accu2[5] ;
 wire \dac.accu2[6] ;
 wire \dac.accu2[7] ;
 wire \dac.accu2[8] ;
 wire \dac.accu2[9] ;
 wire \dac.accu3[0] ;
 wire \dac.accu3[1] ;
 wire \dac.mod2_ctr[0] ;
 wire \dac.mod2_ctr[1] ;
 wire \dac.mod2_out[0] ;
 wire \dac.mod2_out[1] ;
 wire \dac.o_ds ;
 wire \dac.o_ds_n ;
 wire \reg_out_w[0] ;
 wire \reg_out_w[10] ;
 wire \reg_out_w[11] ;
 wire \reg_out_w[12] ;
 wire \reg_out_w[13] ;
 wire \reg_out_w[14] ;
 wire \reg_out_w[15] ;
 wire \reg_out_w[1] ;
 wire \reg_out_w[2] ;
 wire \reg_out_w[3] ;
 wire \reg_out_w[4] ;
 wire \reg_out_w[5] ;
 wire \reg_out_w[6] ;
 wire \reg_out_w[7] ;
 wire \reg_out_w[8] ;
 wire \reg_out_w[9] ;
 wire \sine.ctr_msb_last_r ;
 wire \sine.ctr_r[0] ;
 wire \sine.ctr_r[10] ;
 wire \sine.ctr_r[11] ;
 wire \sine.ctr_r[12] ;
 wire \sine.ctr_r[13] ;
 wire \sine.ctr_r[14] ;
 wire \sine.ctr_r[15] ;
 wire \sine.ctr_r[1] ;
 wire \sine.ctr_r[2] ;
 wire \sine.ctr_r[3] ;
 wire \sine.ctr_r[4] ;
 wire \sine.ctr_r[5] ;
 wire \sine.ctr_r[6] ;
 wire \sine.ctr_r[7] ;
 wire \sine.ctr_r[8] ;
 wire \sine.ctr_r[9] ;
 wire \sine.read_ptr_r[0] ;
 wire \sine.read_ptr_r[1] ;
 wire \sine.read_ptr_r[2] ;
 wire \sine.read_ptr_r[3] ;
 wire \sine.read_ptr_r[4] ;
 wire \sine.read_ptr_r[5] ;
 wire \spi.last_spi_clk_r ;
 wire \spi.o_check ;
 wire \spi.o_det ;
 wire \spi.o_spi_dat ;
 wire \spi.scan_r[0] ;
 wire \spi.scan_r[10] ;
 wire \spi.scan_r[11] ;
 wire \spi.scan_r[12] ;
 wire \spi.scan_r[13] ;
 wire \spi.scan_r[14] ;
 wire \spi.scan_r[1] ;
 wire \spi.scan_r[2] ;
 wire \spi.scan_r[3] ;
 wire \spi.scan_r[4] ;
 wire \spi.scan_r[5] ;
 wire \spi.scan_r[6] ;
 wire \spi.scan_r[7] ;
 wire \spi.scan_r[8] ;
 wire \spi.scan_r[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _1358_ (.A(net5),
    .X(_0532_));
 sg13g2_buf_1 _1359_ (.A(_0532_),
    .X(_0533_));
 sg13g2_nand2_1 _1360_ (.Y(_0534_),
    .A(\dac.accu3[1] ),
    .B(\dac.mod2_out[1] ));
 sg13g2_nand2_1 _1361_ (.Y(_0535_),
    .A(\dac.accu3[0] ),
    .B(\dac.mod2_out[0] ));
 sg13g2_nand2_1 _1362_ (.Y(_0536_),
    .A(_0534_),
    .B(_0535_));
 sg13g2_o21ai_1 _1363_ (.B1(_0536_),
    .Y(_0537_),
    .A1(\dac.accu3[1] ),
    .A2(\dac.mod2_out[1] ));
 sg13g2_buf_2 _1364_ (.A(\dac.accu1[15] ),
    .X(_0538_));
 sg13g2_inv_1 _1365_ (.Y(_0539_),
    .A(_0001_));
 sg13g2_buf_1 _1366_ (.A(ui_in[6]),
    .X(_0540_));
 sg13g2_inv_1 _1367_ (.Y(_0541_),
    .A(net84));
 sg13g2_buf_1 _1368_ (.A(_0541_),
    .X(_0542_));
 sg13g2_buf_1 _1369_ (.A(net64),
    .X(_0543_));
 sg13g2_buf_8 _1370_ (.A(\sine.read_ptr_r[1] ),
    .X(_0544_));
 sg13g2_buf_1 _1371_ (.A(net81),
    .X(_0545_));
 sg13g2_buf_1 _1372_ (.A(net63),
    .X(_0546_));
 sg13g2_buf_8 _1373_ (.A(\sine.read_ptr_r[0] ),
    .X(_0547_));
 sg13g2_buf_1 _1374_ (.A(net80),
    .X(_0548_));
 sg13g2_buf_1 _1375_ (.A(net62),
    .X(_0549_));
 sg13g2_buf_8 _1376_ (.A(\sine.read_ptr_r[2] ),
    .X(_0550_));
 sg13g2_buf_8 _1377_ (.A(_0550_),
    .X(_0551_));
 sg13g2_buf_1 _1378_ (.A(net61),
    .X(_0552_));
 sg13g2_buf_1 _1379_ (.A(net43),
    .X(_0553_));
 sg13g2_buf_1 _1380_ (.A(\sine.read_ptr_r[3] ),
    .X(_0554_));
 sg13g2_buf_1 _1381_ (.A(net79),
    .X(_0555_));
 sg13g2_buf_1 _1382_ (.A(_0555_),
    .X(_0556_));
 sg13g2_nor4_1 _1383_ (.A(net45),
    .B(net44),
    .C(net27),
    .D(net42),
    .Y(_0557_));
 sg13g2_buf_1 _1384_ (.A(\sine.read_ptr_r[5] ),
    .X(_0558_));
 sg13g2_inv_2 _1385_ (.Y(_0559_),
    .A(net78));
 sg13g2_buf_1 _1386_ (.A(net59),
    .X(_0560_));
 sg13g2_a21o_1 _1387_ (.A2(_0557_),
    .A1(_0002_),
    .B1(net41),
    .X(_0561_));
 sg13g2_buf_2 _1388_ (.A(ui_in[4]),
    .X(_0562_));
 sg13g2_buf_1 _1389_ (.A(_0562_),
    .X(_0563_));
 sg13g2_buf_1 _1390_ (.A(ui_in[5]),
    .X(_0564_));
 sg13g2_buf_1 _1391_ (.A(_0564_),
    .X(_0565_));
 sg13g2_buf_1 _1392_ (.A(net84),
    .X(_0566_));
 sg13g2_nand2b_1 _1393_ (.Y(_0567_),
    .B(_0566_),
    .A_N(_0565_));
 sg13g2_nor2_1 _1394_ (.A(net77),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_a22oi_1 _1395_ (.Y(_0569_),
    .B1(_0561_),
    .B2(_0568_),
    .A2(net46),
    .A1(_0539_));
 sg13g2_buf_1 _1396_ (.A(_0569_),
    .X(_0570_));
 sg13g2_inv_1 _1397_ (.Y(_0571_),
    .A(_0570_));
 sg13g2_inv_1 _1398_ (.Y(_0572_),
    .A(_0003_));
 sg13g2_nor2_2 _1399_ (.A(_0562_),
    .B(_0564_),
    .Y(_0573_));
 sg13g2_nand2_1 _1400_ (.Y(_0574_),
    .A(net84),
    .B(_0573_));
 sg13g2_buf_1 _1401_ (.A(net61),
    .X(_0575_));
 sg13g2_and2_1 _1402_ (.A(\sine.read_ptr_r[1] ),
    .B(net80),
    .X(_0576_));
 sg13g2_buf_2 _1403_ (.A(_0576_),
    .X(_0577_));
 sg13g2_buf_1 _1404_ (.A(\sine.read_ptr_r[4] ),
    .X(_0578_));
 sg13g2_nor2b_1 _1405_ (.A(_0004_),
    .B_N(_0578_),
    .Y(_0579_));
 sg13g2_o21ai_1 _1406_ (.B1(_0579_),
    .Y(_0580_),
    .A1(net40),
    .A2(_0577_));
 sg13g2_nor2_1 _1407_ (.A(net79),
    .B(net74),
    .Y(_0581_));
 sg13g2_buf_8 _1408_ (.A(_0550_),
    .X(_0582_));
 sg13g2_nand2_1 _1409_ (.Y(_0583_),
    .A(net81),
    .B(net57));
 sg13g2_a21oi_1 _1410_ (.A1(net58),
    .A2(_0583_),
    .Y(_0584_),
    .B1(net78));
 sg13g2_and2_1 _1411_ (.A(_0580_),
    .B(_0584_),
    .X(_0585_));
 sg13g2_buf_8 _1412_ (.A(net80),
    .X(_0586_));
 sg13g2_buf_1 _1413_ (.A(net56),
    .X(_0587_));
 sg13g2_nand2_1 _1414_ (.Y(_0588_),
    .A(net39),
    .B(net58));
 sg13g2_or2_1 _1415_ (.X(_0589_),
    .B(net61),
    .A(net81));
 sg13g2_o21ai_1 _1416_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net58),
    .A2(_0579_));
 sg13g2_nand2_2 _1417_ (.Y(_0591_),
    .A(_0545_),
    .B(net56));
 sg13g2_nor2_1 _1418_ (.A(_0579_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_a221oi_1 _1419_ (.B2(_0553_),
    .C1(net59),
    .B1(_0592_),
    .A1(_0588_),
    .Y(_0593_),
    .A2(_0590_));
 sg13g2_nor2_1 _1420_ (.A(_0585_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_nor2_1 _1421_ (.A(_0574_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_a21oi_2 _1422_ (.B1(_0595_),
    .Y(_0596_),
    .A2(_0572_),
    .A1(net46));
 sg13g2_inv_1 _1423_ (.Y(_0597_),
    .A(_0596_));
 sg13g2_buf_2 _1424_ (.A(\dac.accu1[4] ),
    .X(_0598_));
 sg13g2_nand2_1 _1425_ (.Y(_0599_),
    .A(net64),
    .B(_0018_));
 sg13g2_and2_1 _1426_ (.A(net79),
    .B(net74),
    .X(_0600_));
 sg13g2_buf_1 _1427_ (.A(_0600_),
    .X(_0601_));
 sg13g2_or2_1 _1428_ (.X(_0602_),
    .B(net74),
    .A(_0554_));
 sg13g2_buf_1 _1429_ (.A(_0602_),
    .X(_0603_));
 sg13g2_o21ai_1 _1430_ (.B1(_0603_),
    .Y(_0604_),
    .A1(net27),
    .A2(net38));
 sg13g2_buf_1 _1431_ (.A(net78),
    .X(_0605_));
 sg13g2_buf_1 _1432_ (.A(net81),
    .X(_0606_));
 sg13g2_nor2b_1 _1433_ (.A(net54),
    .B_N(net62),
    .Y(_0607_));
 sg13g2_and2_1 _1434_ (.A(net55),
    .B(_0607_),
    .X(_0608_));
 sg13g2_buf_8 _1435_ (.A(net74),
    .X(_0609_));
 sg13g2_or3_1 _1436_ (.A(net62),
    .B(net57),
    .C(net53),
    .X(_0610_));
 sg13g2_buf_1 _1437_ (.A(net53),
    .X(_0611_));
 sg13g2_nand2_1 _1438_ (.Y(_0612_),
    .A(net39),
    .B(net37));
 sg13g2_buf_1 _1439_ (.A(net79),
    .X(_0613_));
 sg13g2_nand3_1 _1440_ (.B(net52),
    .C(net78),
    .A(net45),
    .Y(_0614_));
 sg13g2_a21oi_1 _1441_ (.A1(_0610_),
    .A2(_0612_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_a21oi_1 _1442_ (.A1(_0604_),
    .A2(_0608_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_nor2_2 _1443_ (.A(net43),
    .B(net60),
    .Y(_0617_));
 sg13g2_o21ai_1 _1444_ (.B1(_0607_),
    .Y(_0618_),
    .A1(net55),
    .A2(_0617_));
 sg13g2_inv_2 _1445_ (.Y(_0619_),
    .A(net61));
 sg13g2_inv_1 _1446_ (.Y(_0620_),
    .A(net74));
 sg13g2_buf_1 _1447_ (.A(_0620_),
    .X(_0621_));
 sg13g2_a21oi_1 _1448_ (.A1(net36),
    .A2(net55),
    .Y(_0622_),
    .B1(net35));
 sg13g2_nor2b_1 _1449_ (.A(\sine.read_ptr_r[5] ),
    .B_N(net43),
    .Y(_0623_));
 sg13g2_nor2b_1 _1450_ (.A(net61),
    .B_N(net79),
    .Y(_0624_));
 sg13g2_buf_1 _1451_ (.A(_0624_),
    .X(_0625_));
 sg13g2_a22oi_1 _1452_ (.Y(_0626_),
    .B1(net26),
    .B2(net45),
    .A2(_0623_),
    .A1(_0577_));
 sg13g2_nor2b_1 _1453_ (.A(net39),
    .B_N(net52),
    .Y(_0627_));
 sg13g2_buf_2 _1454_ (.A(net79),
    .X(_0628_));
 sg13g2_nor2_1 _1455_ (.A(net56),
    .B(net51),
    .Y(_0629_));
 sg13g2_a22oi_1 _1456_ (.Y(_0630_),
    .B1(_0629_),
    .B2(_0623_),
    .A2(_0627_),
    .A1(net55));
 sg13g2_nand4_1 _1457_ (.B(_0622_),
    .C(_0626_),
    .A(_0618_),
    .Y(_0631_),
    .D(_0630_));
 sg13g2_nand2_1 _1458_ (.Y(_0632_),
    .A(net61),
    .B(net51));
 sg13g2_xnor2_1 _1459_ (.Y(_0633_),
    .A(net61),
    .B(net51));
 sg13g2_xor2_1 _1460_ (.B(net56),
    .A(net81),
    .X(_0634_));
 sg13g2_mux2_1 _1461_ (.A0(_0632_),
    .A1(_0633_),
    .S(_0634_),
    .X(_0635_));
 sg13g2_buf_2 _1462_ (.A(_0009_),
    .X(_0636_));
 sg13g2_or2_1 _1463_ (.X(_0637_),
    .B(net37),
    .A(net78));
 sg13g2_a21oi_1 _1464_ (.A1(_0636_),
    .A2(_0617_),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_buf_1 _1465_ (.A(net53),
    .X(_0639_));
 sg13g2_or2_1 _1466_ (.X(_0640_),
    .B(net80),
    .A(net81));
 sg13g2_buf_1 _1467_ (.A(_0640_),
    .X(_0641_));
 sg13g2_o21ai_1 _1468_ (.B1(_0591_),
    .Y(_0642_),
    .A1(net34),
    .A2(_0641_));
 sg13g2_nor2_1 _1469_ (.A(net59),
    .B(_0632_),
    .Y(_0643_));
 sg13g2_a221oi_1 _1470_ (.B2(_0643_),
    .C1(_0542_),
    .B1(_0642_),
    .A1(_0635_),
    .Y(_0644_),
    .A2(_0638_));
 sg13g2_nand3_1 _1471_ (.B(_0631_),
    .C(_0644_),
    .A(_0616_),
    .Y(_0645_));
 sg13g2_o21ai_1 _1472_ (.B1(net75),
    .Y(_0646_),
    .A1(net77),
    .A2(net76));
 sg13g2_nand3_1 _1473_ (.B(_0645_),
    .C(_0646_),
    .A(_0599_),
    .Y(_0647_));
 sg13g2_nand2b_1 _1474_ (.Y(_0648_),
    .B(net63),
    .A_N(net53));
 sg13g2_or2_1 _1475_ (.X(_0649_),
    .B(_0648_),
    .A(_0633_));
 sg13g2_nand2b_1 _1476_ (.Y(_0650_),
    .B(net63),
    .A_N(net57));
 sg13g2_buf_8 _1477_ (.A(net74),
    .X(_0651_));
 sg13g2_and2_1 _1478_ (.A(net63),
    .B(net50),
    .X(_0652_));
 sg13g2_a22oi_1 _1479_ (.Y(_0653_),
    .B1(_0652_),
    .B2(_0617_),
    .A2(_0650_),
    .A1(net38));
 sg13g2_inv_2 _1480_ (.Y(_0654_),
    .A(net56));
 sg13g2_a21o_1 _1481_ (.A2(_0653_),
    .A1(_0649_),
    .B1(net33),
    .X(_0655_));
 sg13g2_buf_1 _1482_ (.A(_0022_),
    .X(_0656_));
 sg13g2_nor4_1 _1483_ (.A(net40),
    .B(_0613_),
    .C(_0611_),
    .D(_0656_),
    .Y(_0657_));
 sg13g2_nand2b_1 _1484_ (.Y(_0658_),
    .B(net40),
    .A_N(net63));
 sg13g2_a21oi_1 _1485_ (.A1(_0587_),
    .A2(net58),
    .Y(_0659_),
    .B1(_0658_));
 sg13g2_nor3_1 _1486_ (.A(net41),
    .B(_0657_),
    .C(_0659_),
    .Y(_0660_));
 sg13g2_xnor2_1 _1487_ (.Y(_0661_),
    .A(_0547_),
    .B(_0551_));
 sg13g2_nand2b_1 _1488_ (.Y(_0662_),
    .B(net38),
    .A_N(_0661_));
 sg13g2_nand2_1 _1489_ (.Y(_0663_),
    .A(net51),
    .B(net53));
 sg13g2_nor2_2 _1490_ (.A(net80),
    .B(net61),
    .Y(_0664_));
 sg13g2_inv_2 _1491_ (.Y(_0665_),
    .A(net81));
 sg13g2_a21oi_1 _1492_ (.A1(_0663_),
    .A2(_0664_),
    .Y(_0666_),
    .B1(_0665_));
 sg13g2_and2_1 _1493_ (.A(_0547_),
    .B(_0550_),
    .X(_0667_));
 sg13g2_buf_1 _1494_ (.A(_0667_),
    .X(_0668_));
 sg13g2_a221oi_1 _1495_ (.B2(net33),
    .C1(_0546_),
    .B1(net26),
    .A1(net58),
    .Y(_0669_),
    .A2(_0668_));
 sg13g2_a21o_1 _1496_ (.A2(_0666_),
    .A1(_0662_),
    .B1(_0669_),
    .X(_0670_));
 sg13g2_buf_1 _1497_ (.A(net78),
    .X(_0671_));
 sg13g2_nand2b_1 _1498_ (.Y(_0672_),
    .B(net60),
    .A_N(net53));
 sg13g2_nand2b_2 _1499_ (.Y(_0673_),
    .B(net50),
    .A_N(_0628_));
 sg13g2_nor2b_1 _1500_ (.A(net43),
    .B_N(net63),
    .Y(_0674_));
 sg13g2_a221oi_1 _1501_ (.B2(_0673_),
    .C1(_0674_),
    .B1(_0672_),
    .A1(net40),
    .Y(_0675_),
    .A2(_0636_));
 sg13g2_nor2_1 _1502_ (.A(net49),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_a22oi_1 _1503_ (.Y(_0677_),
    .B1(_0670_),
    .B2(_0676_),
    .A2(_0660_),
    .A1(_0655_));
 sg13g2_nor2b_2 _1504_ (.A(_0562_),
    .B_N(_0564_),
    .Y(_0678_));
 sg13g2_nand3_1 _1505_ (.B(_0678_),
    .C(_0599_),
    .A(_0677_),
    .Y(_0679_));
 sg13g2_buf_1 _1506_ (.A(net54),
    .X(_0680_));
 sg13g2_nor2b_1 _1507_ (.A(net54),
    .B_N(net43),
    .Y(_0681_));
 sg13g2_a22oi_1 _1508_ (.Y(_0682_),
    .B1(_0612_),
    .B2(_0681_),
    .A2(_0664_),
    .A1(net32));
 sg13g2_nor2b_1 _1509_ (.A(net57),
    .B_N(net53),
    .Y(_0683_));
 sg13g2_buf_1 _1510_ (.A(_0008_),
    .X(_0684_));
 sg13g2_nand2b_1 _1511_ (.Y(_0685_),
    .B(net73),
    .A_N(net37));
 sg13g2_a22oi_1 _1512_ (.Y(_0686_),
    .B1(_0685_),
    .B2(net42),
    .A2(_0683_),
    .A1(net44));
 sg13g2_o21ai_1 _1513_ (.B1(_0686_),
    .Y(_0687_),
    .A1(net42),
    .A2(_0682_));
 sg13g2_nand2_1 _1514_ (.Y(_0688_),
    .A(net36),
    .B(_0577_));
 sg13g2_nor2b_1 _1515_ (.A(net56),
    .B_N(net57),
    .Y(_0689_));
 sg13g2_nor2_1 _1516_ (.A(_0663_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_a21oi_1 _1517_ (.A1(_0688_),
    .A2(_0690_),
    .Y(_0691_),
    .B1(net41));
 sg13g2_nor2b_1 _1518_ (.A(net51),
    .B_N(_0656_),
    .Y(_0692_));
 sg13g2_o21ai_1 _1519_ (.B1(net32),
    .Y(_0693_),
    .A1(net34),
    .A2(_0692_));
 sg13g2_nor2b_2 _1520_ (.A(net51),
    .B_N(net74),
    .Y(_0694_));
 sg13g2_a21oi_1 _1521_ (.A1(net44),
    .A2(_0694_),
    .Y(_0695_),
    .B1(net27));
 sg13g2_o21ai_1 _1522_ (.B1(net37),
    .Y(_0696_),
    .A1(net62),
    .A2(net52));
 sg13g2_nand2b_1 _1523_ (.Y(_0697_),
    .B(net37),
    .A_N(_0656_));
 sg13g2_o21ai_1 _1524_ (.B1(net40),
    .Y(_0698_),
    .A1(net39),
    .A2(net37));
 sg13g2_a221oi_1 _1525_ (.B2(net42),
    .C1(_0698_),
    .B1(_0697_),
    .A1(_0665_),
    .Y(_0699_),
    .A2(_0696_));
 sg13g2_a21o_1 _1526_ (.A2(_0695_),
    .A1(_0693_),
    .B1(_0699_),
    .X(_0700_));
 sg13g2_nor2_1 _1527_ (.A(net63),
    .B(net50),
    .Y(_0701_));
 sg13g2_a21oi_1 _1528_ (.A1(_0692_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(_0671_));
 sg13g2_a22oi_1 _1529_ (.Y(_0703_),
    .B1(_0700_),
    .B2(_0702_),
    .A2(_0691_),
    .A1(_0687_));
 sg13g2_inv_1 _1530_ (.Y(_0704_),
    .A(_0562_));
 sg13g2_nor2_1 _1531_ (.A(_0704_),
    .B(net76),
    .Y(_0705_));
 sg13g2_nand3b_1 _1532_ (.B(_0705_),
    .C(_0599_),
    .Y(_0706_),
    .A_N(_0703_));
 sg13g2_and3_1 _1533_ (.X(_0707_),
    .A(_0647_),
    .B(_0679_),
    .C(_0706_));
 sg13g2_nand2_1 _1534_ (.Y(_0708_),
    .A(_0598_),
    .B(_0707_));
 sg13g2_inv_2 _1535_ (.Y(_0709_),
    .A(_0598_));
 sg13g2_nand3_1 _1536_ (.B(_0679_),
    .C(_0706_),
    .A(_0647_),
    .Y(_0710_));
 sg13g2_buf_2 _1537_ (.A(_0710_),
    .X(_0711_));
 sg13g2_nand2_1 _1538_ (.Y(_0712_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_nor2b_1 _1539_ (.A(_0636_),
    .B_N(net57),
    .Y(_0713_));
 sg13g2_nor2_1 _1540_ (.A(_0663_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_a21o_1 _1541_ (.A2(net57),
    .A1(net56),
    .B1(_0609_),
    .X(_0715_));
 sg13g2_a21oi_1 _1542_ (.A1(net54),
    .A2(_0664_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_nand2b_1 _1543_ (.Y(_0717_),
    .B(net80),
    .A_N(net79));
 sg13g2_a21o_1 _1544_ (.A2(_0632_),
    .A1(_0717_),
    .B1(_0606_),
    .X(_0718_));
 sg13g2_a221oi_1 _1545_ (.B2(_0718_),
    .C1(net49),
    .B1(_0716_),
    .A1(_0688_),
    .Y(_0719_),
    .A2(_0714_));
 sg13g2_nand2b_1 _1546_ (.Y(_0720_),
    .B(net50),
    .A_N(net43));
 sg13g2_nand2b_1 _1547_ (.Y(_0721_),
    .B(_0545_),
    .A_N(net60));
 sg13g2_nor3_1 _1548_ (.A(_0587_),
    .B(_0720_),
    .C(_0721_),
    .Y(_0722_));
 sg13g2_nand2_1 _1549_ (.Y(_0723_),
    .A(net39),
    .B(_0575_));
 sg13g2_a21oi_1 _1550_ (.A1(_0673_),
    .A2(_0721_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_nor2_1 _1551_ (.A(_0722_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_and2_1 _1552_ (.A(_0550_),
    .B(net79),
    .X(_0726_));
 sg13g2_buf_1 _1553_ (.A(_0726_),
    .X(_0727_));
 sg13g2_nand2_1 _1554_ (.Y(_0728_),
    .A(net35),
    .B(_0727_));
 sg13g2_nand2b_1 _1555_ (.Y(_0729_),
    .B(net81),
    .A_N(_0586_));
 sg13g2_nor2_1 _1556_ (.A(_0694_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_nor2_1 _1557_ (.A(net45),
    .B(net26),
    .Y(_0731_));
 sg13g2_o21ai_1 _1558_ (.B1(net40),
    .Y(_0732_),
    .A1(net37),
    .A2(_0629_));
 sg13g2_nor2_1 _1559_ (.A(_0582_),
    .B(_0609_),
    .Y(_0733_));
 sg13g2_nor2b_2 _1560_ (.A(net60),
    .B_N(_0551_),
    .Y(_0734_));
 sg13g2_nor3_1 _1561_ (.A(_0591_),
    .B(_0733_),
    .C(_0734_),
    .Y(_0735_));
 sg13g2_a221oi_1 _1562_ (.B2(_0732_),
    .C1(_0735_),
    .B1(_0731_),
    .A1(_0728_),
    .Y(_0736_),
    .A2(_0730_));
 sg13g2_nand2b_1 _1563_ (.Y(_0737_),
    .B(_0552_),
    .A_N(net60));
 sg13g2_nand2_1 _1564_ (.Y(_0738_),
    .A(_0651_),
    .B(_0656_));
 sg13g2_nor2_1 _1565_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_nor2_1 _1566_ (.A(net59),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_a22oi_1 _1567_ (.Y(_0741_),
    .B1(_0736_),
    .B2(_0740_),
    .A2(_0725_),
    .A1(_0719_));
 sg13g2_nand2b_2 _1568_ (.Y(_0742_),
    .B(_0562_),
    .A_N(_0564_));
 sg13g2_nor2_1 _1569_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sg13g2_nor2_1 _1570_ (.A(_0558_),
    .B(net34),
    .Y(_0744_));
 sg13g2_nor2_1 _1571_ (.A(net55),
    .B(net35),
    .Y(_0745_));
 sg13g2_inv_1 _1572_ (.Y(_0746_),
    .A(net60));
 sg13g2_nor3_1 _1573_ (.A(_0746_),
    .B(net59),
    .C(_0589_),
    .Y(_0747_));
 sg13g2_a221oi_1 _1574_ (.B2(_0617_),
    .C1(_0747_),
    .B1(_0745_),
    .A1(_0744_),
    .Y(_0748_),
    .A2(_0727_));
 sg13g2_nor2b_2 _1575_ (.A(net57),
    .B_N(net80),
    .Y(_0749_));
 sg13g2_nor2b_1 _1576_ (.A(_0613_),
    .B_N(_0558_),
    .Y(_0750_));
 sg13g2_a22oi_1 _1577_ (.Y(_0751_),
    .B1(_0668_),
    .B2(_0750_),
    .A2(_0749_),
    .A1(net59));
 sg13g2_nor3_1 _1578_ (.A(net62),
    .B(net43),
    .C(net50),
    .Y(_0752_));
 sg13g2_and2_1 _1579_ (.A(_0550_),
    .B(net74),
    .X(_0753_));
 sg13g2_buf_1 _1580_ (.A(_0753_),
    .X(_0754_));
 sg13g2_o21ai_1 _1581_ (.B1(_0605_),
    .Y(_0755_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_buf_1 _1582_ (.A(_0665_),
    .X(_0756_));
 sg13g2_a21o_1 _1583_ (.A2(_0755_),
    .A1(_0751_),
    .B1(_0756_),
    .X(_0757_));
 sg13g2_nor2b_1 _1584_ (.A(net50),
    .B_N(\sine.read_ptr_r[5] ),
    .Y(_0758_));
 sg13g2_a21oi_1 _1585_ (.A1(_0749_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(_0623_));
 sg13g2_or2_1 _1586_ (.X(_0760_),
    .B(_0759_),
    .A(net32));
 sg13g2_and3_1 _1587_ (.X(_0761_),
    .A(_0748_),
    .B(_0757_),
    .C(_0760_));
 sg13g2_nand2_1 _1588_ (.Y(_0762_),
    .A(_0704_),
    .B(net76));
 sg13g2_inv_1 _1589_ (.Y(_0763_),
    .A(net73));
 sg13g2_a21oi_1 _1590_ (.A1(_0763_),
    .A2(_0641_),
    .Y(_0764_),
    .B1(_0673_));
 sg13g2_mux2_1 _1591_ (.A0(_0555_),
    .A1(net62),
    .S(_0582_),
    .X(_0765_));
 sg13g2_o21ai_1 _1592_ (.B1(_0605_),
    .Y(_0766_),
    .A1(_0648_),
    .A2(_0765_));
 sg13g2_a221oi_1 _1593_ (.B2(net36),
    .C1(_0746_),
    .B1(_0738_),
    .A1(_0754_),
    .Y(_0767_),
    .A2(_0729_));
 sg13g2_nand3_1 _1594_ (.B(net40),
    .C(net52),
    .A(net39),
    .Y(_0768_));
 sg13g2_a21oi_1 _1595_ (.A1(_0610_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(net45));
 sg13g2_nor4_2 _1596_ (.A(_0764_),
    .B(_0766_),
    .C(_0767_),
    .Y(_0770_),
    .D(_0769_));
 sg13g2_nor2_2 _1597_ (.A(_0544_),
    .B(net80),
    .Y(_0771_));
 sg13g2_nor2_1 _1598_ (.A(net73),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_nor2b_1 _1599_ (.A(_0586_),
    .B_N(_0544_),
    .Y(_0773_));
 sg13g2_a22oi_1 _1600_ (.Y(_0774_),
    .B1(_0727_),
    .B2(_0773_),
    .A2(_0617_),
    .A1(net45));
 sg13g2_nor2b_1 _1601_ (.A(net54),
    .B_N(net51),
    .Y(_0775_));
 sg13g2_a221oi_1 _1602_ (.B2(_0775_),
    .C1(_0694_),
    .B1(_0661_),
    .A1(net35),
    .Y(_0776_),
    .A2(_0727_));
 sg13g2_a221oi_1 _1603_ (.B2(_0776_),
    .C1(net49),
    .B1(_0774_),
    .A1(_0694_),
    .Y(_0777_),
    .A2(_0772_));
 sg13g2_o21ai_1 _1604_ (.B1(_0573_),
    .Y(_0778_),
    .A1(_0770_),
    .A2(_0777_));
 sg13g2_o21ai_1 _1605_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0761_),
    .A2(_0762_));
 sg13g2_nor3_1 _1606_ (.A(net46),
    .B(_0743_),
    .C(_0779_),
    .Y(_0780_));
 sg13g2_buf_1 _1607_ (.A(net75),
    .X(_0781_));
 sg13g2_nor2b_1 _1608_ (.A(net48),
    .B_N(_0017_),
    .Y(_0782_));
 sg13g2_o21ai_1 _1609_ (.B1(\dac.accu1[5] ),
    .Y(_0783_),
    .A1(_0780_),
    .A2(_0782_));
 sg13g2_inv_1 _1610_ (.Y(_0784_),
    .A(\dac.accu1[5] ));
 sg13g2_or3_1 _1611_ (.A(net64),
    .B(_0743_),
    .C(_0779_),
    .X(_0785_));
 sg13g2_buf_2 _1612_ (.A(_0785_),
    .X(_0786_));
 sg13g2_nand2_2 _1613_ (.Y(_0787_),
    .A(net46),
    .B(_0017_));
 sg13g2_nand3_1 _1614_ (.B(_0786_),
    .C(_0787_),
    .A(net72),
    .Y(_0788_));
 sg13g2_or2_1 _1615_ (.X(_0789_),
    .B(net73),
    .A(net52));
 sg13g2_inv_1 _1616_ (.Y(_0790_),
    .A(_0656_));
 sg13g2_nand2_1 _1617_ (.Y(_0791_),
    .A(net52),
    .B(_0790_));
 sg13g2_o21ai_1 _1618_ (.B1(_0791_),
    .Y(_0792_),
    .A1(_0634_),
    .A2(_0789_));
 sg13g2_a22oi_1 _1619_ (.Y(_0793_),
    .B1(_0683_),
    .B2(_0773_),
    .A2(_0754_),
    .A1(_0771_));
 sg13g2_a22oi_1 _1620_ (.Y(_0794_),
    .B1(_0749_),
    .B2(_0665_),
    .A2(_0620_),
    .A1(_0548_));
 sg13g2_a21o_1 _1621_ (.A2(_0794_),
    .A1(_0793_),
    .B1(_0746_),
    .X(_0795_));
 sg13g2_nand2_1 _1622_ (.Y(_0796_),
    .A(_0654_),
    .B(_0589_));
 sg13g2_o21ai_1 _1623_ (.B1(_0583_),
    .Y(_0797_),
    .A1(net54),
    .A2(_0790_));
 sg13g2_a221oi_1 _1624_ (.B2(net58),
    .C1(net55),
    .B1(_0797_),
    .A1(_0694_),
    .Y(_0798_),
    .A2(_0796_));
 sg13g2_nand2_1 _1625_ (.Y(_0799_),
    .A(net33),
    .B(_0625_));
 sg13g2_and2_1 _1626_ (.A(net78),
    .B(_0651_),
    .X(_0800_));
 sg13g2_and2_1 _1627_ (.A(net56),
    .B(net51),
    .X(_0801_));
 sg13g2_o21ai_1 _1628_ (.B1(net40),
    .Y(_0802_),
    .A1(_0692_),
    .A2(_0801_));
 sg13g2_o21ai_1 _1629_ (.B1(net54),
    .Y(_0803_),
    .A1(net52),
    .A2(_0664_));
 sg13g2_and4_1 _1630_ (.A(_0799_),
    .B(_0800_),
    .C(_0802_),
    .D(_0803_),
    .X(_0804_));
 sg13g2_a221oi_1 _1631_ (.B2(_0798_),
    .C1(_0804_),
    .B1(_0795_),
    .A1(_0758_),
    .Y(_0805_),
    .A2(_0792_));
 sg13g2_a22oi_1 _1632_ (.Y(_0806_),
    .B1(_0805_),
    .B2(_0573_),
    .A2(_0594_),
    .A1(net76));
 sg13g2_o21ai_1 _1633_ (.B1(_0650_),
    .Y(_0807_),
    .A1(net36),
    .A2(_0790_));
 sg13g2_nand3b_1 _1634_ (.B(net62),
    .C(net43),
    .Y(_0808_),
    .A_N(net63));
 sg13g2_o21ai_1 _1635_ (.B1(_0808_),
    .Y(_0809_),
    .A1(_0665_),
    .A2(_0661_));
 sg13g2_a221oi_1 _1636_ (.B2(_0694_),
    .C1(net59),
    .B1(_0809_),
    .A1(net38),
    .Y(_0810_),
    .A2(_0807_));
 sg13g2_or2_1 _1637_ (.X(_0811_),
    .B(_0656_),
    .A(net60));
 sg13g2_a22oi_1 _1638_ (.Y(_0812_),
    .B1(_0811_),
    .B2(_0674_),
    .A2(_0734_),
    .A1(net33));
 sg13g2_o21ai_1 _1639_ (.B1(_0665_),
    .Y(_0813_),
    .A1(_0668_),
    .A2(_0692_));
 sg13g2_a21o_1 _1640_ (.A2(_0813_),
    .A1(_0812_),
    .B1(net34),
    .X(_0814_));
 sg13g2_nand2b_1 _1641_ (.Y(_0815_),
    .B(net52),
    .A_N(_0548_));
 sg13g2_o21ai_1 _1642_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net45),
    .A2(_0717_));
 sg13g2_o21ai_1 _1643_ (.B1(net34),
    .Y(_0817_),
    .A1(_0665_),
    .A2(_0661_));
 sg13g2_a21o_1 _1644_ (.A2(_0816_),
    .A1(net27),
    .B1(_0817_),
    .X(_0818_));
 sg13g2_nor2b_1 _1645_ (.A(net53),
    .B_N(_0628_),
    .Y(_0819_));
 sg13g2_inv_1 _1646_ (.Y(_0820_),
    .A(_0636_));
 sg13g2_a22oi_1 _1647_ (.Y(_0821_),
    .B1(_0668_),
    .B2(_0665_),
    .A2(_0820_),
    .A1(net36));
 sg13g2_nand2_1 _1648_ (.Y(_0822_),
    .A(net45),
    .B(_0664_));
 sg13g2_nor2_1 _1649_ (.A(_0603_),
    .B(_0681_),
    .Y(_0823_));
 sg13g2_a221oi_1 _1650_ (.B2(_0823_),
    .C1(net49),
    .B1(_0822_),
    .A1(_0819_),
    .Y(_0824_),
    .A2(_0821_));
 sg13g2_a22oi_1 _1651_ (.Y(_0825_),
    .B1(_0818_),
    .B2(_0824_),
    .A2(_0814_),
    .A1(_0810_));
 sg13g2_o21ai_1 _1652_ (.B1(net77),
    .Y(_0826_),
    .A1(net76),
    .A2(_0825_));
 sg13g2_nand3_1 _1653_ (.B(_0806_),
    .C(_0826_),
    .A(net48),
    .Y(_0827_));
 sg13g2_buf_1 _1654_ (.A(_0827_),
    .X(_0828_));
 sg13g2_or2_1 _1655_ (.X(_0829_),
    .B(_0016_),
    .A(net48));
 sg13g2_buf_1 _1656_ (.A(_0829_),
    .X(_0830_));
 sg13g2_inv_1 _1657_ (.Y(_0831_),
    .A(_0015_));
 sg13g2_nor2b_1 _1658_ (.A(_0611_),
    .B_N(_0636_),
    .Y(_0832_));
 sg13g2_or2_1 _1659_ (.X(_0833_),
    .B(_0832_),
    .A(net26));
 sg13g2_nor2_1 _1660_ (.A(net37),
    .B(_0636_),
    .Y(_0834_));
 sg13g2_o21ai_1 _1661_ (.B1(_0556_),
    .Y(_0835_),
    .A1(net32),
    .A2(_0834_));
 sg13g2_nor2_1 _1662_ (.A(_0820_),
    .B(_0603_),
    .Y(_0836_));
 sg13g2_a221oi_1 _1663_ (.B2(net27),
    .C1(_0836_),
    .B1(_0835_),
    .A1(net32),
    .Y(_0837_),
    .A2(_0833_));
 sg13g2_or2_1 _1664_ (.X(_0838_),
    .B(_0837_),
    .A(net44));
 sg13g2_o21ai_1 _1665_ (.B1(net32),
    .Y(_0839_),
    .A1(net26),
    .A2(_0834_));
 sg13g2_o21ai_1 _1666_ (.B1(_0737_),
    .Y(_0840_),
    .A1(net26),
    .A2(_0832_));
 sg13g2_a21oi_1 _1667_ (.A1(_0756_),
    .A2(_0840_),
    .Y(_0841_),
    .B1(net33));
 sg13g2_o21ai_1 _1668_ (.B1(net49),
    .Y(_0842_),
    .A1(_0556_),
    .A2(_0583_));
 sg13g2_a21oi_1 _1669_ (.A1(_0839_),
    .A2(_0841_),
    .Y(_0843_),
    .B1(_0842_));
 sg13g2_xnor2_1 _1670_ (.Y(_0844_),
    .A(net60),
    .B(net50));
 sg13g2_mux2_1 _1671_ (.A0(_0723_),
    .A1(_0661_),
    .S(net31),
    .X(_0845_));
 sg13g2_xnor2_1 _1672_ (.Y(_0846_),
    .A(net31),
    .B(_0664_));
 sg13g2_nand2_1 _1673_ (.Y(_0847_),
    .A(net44),
    .B(_0636_));
 sg13g2_nand2b_1 _1674_ (.Y(_0848_),
    .B(net73),
    .A_N(net39));
 sg13g2_a21oi_1 _1675_ (.A1(_0847_),
    .A2(_0848_),
    .Y(_0849_),
    .B1(_0673_));
 sg13g2_a221oi_1 _1676_ (.B2(_0819_),
    .C1(_0849_),
    .B1(_0846_),
    .A1(_0844_),
    .Y(_0850_),
    .A2(_0845_));
 sg13g2_and2_1 _1677_ (.A(net41),
    .B(_0850_),
    .X(_0851_));
 sg13g2_a21o_1 _1678_ (.A2(_0843_),
    .A1(_0838_),
    .B1(_0851_),
    .X(_0852_));
 sg13g2_nor2_1 _1679_ (.A(_0541_),
    .B(_0742_),
    .Y(_0853_));
 sg13g2_and2_1 _1680_ (.A(net27),
    .B(net55),
    .X(_0854_));
 sg13g2_mux4_1 _1681_ (.S0(net33),
    .A0(net59),
    .A1(_0854_),
    .A2(_0800_),
    .A3(_0733_),
    .S1(net31),
    .X(_0855_));
 sg13g2_o21ai_1 _1682_ (.B1(_0746_),
    .Y(_0856_),
    .A1(_0744_),
    .A2(_0855_));
 sg13g2_and2_1 _1683_ (.A(_0606_),
    .B(net78),
    .X(_0857_));
 sg13g2_o21ai_1 _1684_ (.B1(_0672_),
    .Y(_0858_),
    .A1(net44),
    .A2(_0720_));
 sg13g2_a21o_1 _1685_ (.A2(_0717_),
    .A1(net31),
    .B1(net38),
    .X(_0859_));
 sg13g2_a221oi_1 _1686_ (.B2(net41),
    .C1(net76),
    .B1(_0859_),
    .A1(_0857_),
    .Y(_0860_),
    .A2(_0858_));
 sg13g2_and2_1 _1687_ (.A(_0565_),
    .B(_0561_),
    .X(_0861_));
 sg13g2_a21o_1 _1688_ (.A2(_0860_),
    .A1(_0856_),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_and3_1 _1689_ (.X(_0863_),
    .A(_0704_),
    .B(net75),
    .C(_0862_));
 sg13g2_a221oi_1 _1690_ (.B2(_0853_),
    .C1(_0863_),
    .B1(_0852_),
    .A1(_0543_),
    .Y(_0864_),
    .A2(_0831_));
 sg13g2_buf_2 _1691_ (.A(_0864_),
    .X(_0865_));
 sg13g2_a21o_1 _1692_ (.A2(net25),
    .A1(net21),
    .B1(_0865_),
    .X(_0866_));
 sg13g2_a221oi_1 _1693_ (.B2(_0788_),
    .C1(_0866_),
    .B1(_0783_),
    .A1(_0708_),
    .Y(_0867_),
    .A2(_0712_));
 sg13g2_inv_1 _1694_ (.Y(_0868_),
    .A(\dac.accu1[6] ));
 sg13g2_or2_1 _1695_ (.X(_0869_),
    .B(_0865_),
    .A(net71));
 sg13g2_a221oi_1 _1696_ (.B2(_0788_),
    .C1(_0869_),
    .B1(_0783_),
    .A1(_0708_),
    .Y(_0870_),
    .A2(_0712_));
 sg13g2_a22oi_1 _1697_ (.Y(_0871_),
    .B1(_0642_),
    .B2(_0643_),
    .A2(_0638_),
    .A1(_0635_));
 sg13g2_and3_1 _1698_ (.X(_0872_),
    .A(_0871_),
    .B(_0616_),
    .C(_0631_));
 sg13g2_a22oi_1 _1699_ (.Y(_0873_),
    .B1(_0872_),
    .B2(_0705_),
    .A2(_0678_),
    .A1(_0703_));
 sg13g2_nor2_1 _1700_ (.A(net50),
    .B(net73),
    .Y(_0874_));
 sg13g2_a21oi_1 _1701_ (.A1(_0575_),
    .A2(_0600_),
    .Y(_0875_),
    .B1(_0874_));
 sg13g2_nand2_1 _1702_ (.Y(_0876_),
    .A(net38),
    .B(_0674_));
 sg13g2_o21ai_1 _1703_ (.B1(_0876_),
    .Y(_0877_),
    .A1(_0641_),
    .A2(_0875_));
 sg13g2_nand2b_1 _1704_ (.Y(_0878_),
    .B(net62),
    .A_N(_0552_));
 sg13g2_nor3_1 _1705_ (.A(net54),
    .B(net39),
    .C(net73),
    .Y(_0879_));
 sg13g2_a221oi_1 _1706_ (.B2(_0878_),
    .C1(_0879_),
    .B1(_0701_),
    .A1(_0621_),
    .Y(_0880_),
    .A2(_0689_));
 sg13g2_inv_1 _1707_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_nor3_1 _1708_ (.A(net42),
    .B(_0562_),
    .C(net76),
    .Y(_0882_));
 sg13g2_a221oi_1 _1709_ (.B2(_0882_),
    .C1(_0541_),
    .B1(_0881_),
    .A1(_0573_),
    .Y(_0883_),
    .A2(_0877_));
 sg13g2_nand2_1 _1710_ (.Y(_0884_),
    .A(_0562_),
    .B(_0564_));
 sg13g2_nor4_1 _1711_ (.A(_0559_),
    .B(_0657_),
    .C(_0659_),
    .D(_0884_),
    .Y(_0885_));
 sg13g2_nor3_1 _1712_ (.A(net49),
    .B(_0675_),
    .C(_0884_),
    .Y(_0886_));
 sg13g2_a22oi_1 _1713_ (.Y(_0887_),
    .B1(_0886_),
    .B2(_0670_),
    .A2(_0885_),
    .A1(_0655_));
 sg13g2_and2_1 _1714_ (.A(_0883_),
    .B(_0887_),
    .X(_0888_));
 sg13g2_nor4_2 _1715_ (.A(net64),
    .B(_0742_),
    .C(_0770_),
    .Y(_0889_),
    .D(_0777_));
 sg13g2_nor2b_1 _1716_ (.A(_0540_),
    .B_N(_0021_),
    .Y(_0890_));
 sg13g2_nand3_1 _1717_ (.B(net84),
    .C(_0573_),
    .A(net55),
    .Y(_0891_));
 sg13g2_a21oi_1 _1718_ (.A1(net34),
    .A2(_0771_),
    .Y(_0892_),
    .B1(_0832_));
 sg13g2_nor4_1 _1719_ (.A(_0553_),
    .B(net42),
    .C(_0891_),
    .D(_0892_),
    .Y(_0893_));
 sg13g2_o21ai_1 _1720_ (.B1(_0601_),
    .Y(_0894_),
    .A1(_0668_),
    .A2(_0664_));
 sg13g2_nand2_1 _1721_ (.Y(_0895_),
    .A(net58),
    .B(_0689_));
 sg13g2_nand3_1 _1722_ (.B(_0573_),
    .C(_0857_),
    .A(net84),
    .Y(_0896_));
 sg13g2_a21oi_1 _1723_ (.A1(_0894_),
    .A2(_0895_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_a22oi_1 _1724_ (.Y(_0898_),
    .B1(_0844_),
    .B2(net36),
    .A2(_0819_),
    .A1(_0684_));
 sg13g2_mux2_1 _1725_ (.A0(_0581_),
    .A1(_0601_),
    .S(_0546_),
    .X(_0899_));
 sg13g2_nand3_1 _1726_ (.B(net84),
    .C(_0573_),
    .A(_0559_),
    .Y(_0900_));
 sg13g2_a221oi_1 _1727_ (.B2(_0549_),
    .C1(_0900_),
    .B1(_0899_),
    .A1(_0771_),
    .Y(_0901_),
    .A2(_0898_));
 sg13g2_or4_1 _1728_ (.A(_0890_),
    .B(_0893_),
    .C(_0897_),
    .D(_0901_),
    .X(_0902_));
 sg13g2_nor2_1 _1729_ (.A(_0541_),
    .B(_0884_),
    .Y(_0903_));
 sg13g2_and4_1 _1730_ (.A(_0748_),
    .B(_0757_),
    .C(_0760_),
    .D(_0903_),
    .X(_0904_));
 sg13g2_nor3_1 _1731_ (.A(_0889_),
    .B(_0902_),
    .C(_0904_),
    .Y(_0905_));
 sg13g2_buf_2 _1732_ (.A(\dac.accu1[0] ),
    .X(_0906_));
 sg13g2_inv_2 _1733_ (.Y(_0907_),
    .A(_0906_));
 sg13g2_nand2_1 _1734_ (.Y(_0908_),
    .A(net84),
    .B(_0678_));
 sg13g2_a221oi_1 _1735_ (.B2(_0740_),
    .C1(_0908_),
    .B1(_0736_),
    .A1(_0719_),
    .Y(_0909_),
    .A2(_0725_));
 sg13g2_nor2_1 _1736_ (.A(_0907_),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_nand4_1 _1737_ (.B(_0888_),
    .C(_0905_),
    .A(_0873_),
    .Y(_0911_),
    .D(_0910_));
 sg13g2_buf_2 _1738_ (.A(\dac.accu1[1] ),
    .X(_0912_));
 sg13g2_inv_1 _1739_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_nor2_1 _1740_ (.A(_0913_),
    .B(_0909_),
    .Y(_0914_));
 sg13g2_buf_1 _1741_ (.A(\reg_out_w[0] ),
    .X(_0915_));
 sg13g2_inv_2 _1742_ (.Y(_0916_),
    .A(_0915_));
 sg13g2_nor3_1 _1743_ (.A(_0916_),
    .B(net75),
    .C(_0907_),
    .Y(_0917_));
 sg13g2_o21ai_1 _1744_ (.B1(_0905_),
    .Y(_0918_),
    .A1(_0914_),
    .A2(_0917_));
 sg13g2_and4_1 _1745_ (.A(_0912_),
    .B(_0906_),
    .C(_0883_),
    .D(_0887_),
    .X(_0919_));
 sg13g2_a22oi_1 _1746_ (.Y(_0920_),
    .B1(_0919_),
    .B2(_0873_),
    .A2(_0917_),
    .A1(_0912_));
 sg13g2_nor2_1 _1747_ (.A(net44),
    .B(_0636_),
    .Y(_0921_));
 sg13g2_o21ai_1 _1748_ (.B1(net42),
    .Y(_0922_),
    .A1(_0701_),
    .A2(_0921_));
 sg13g2_a21oi_1 _1749_ (.A1(_0673_),
    .A2(_0922_),
    .Y(_0923_),
    .B1(net36));
 sg13g2_nor3_1 _1750_ (.A(net38),
    .B(_0734_),
    .C(_0729_),
    .Y(_0924_));
 sg13g2_a221oi_1 _1751_ (.B2(_0619_),
    .C1(net31),
    .B1(_0603_),
    .A1(_0639_),
    .Y(_0925_),
    .A2(_0820_));
 sg13g2_nor3_1 _1752_ (.A(net32),
    .B(net35),
    .C(_0713_),
    .Y(_0926_));
 sg13g2_nor3_1 _1753_ (.A(net33),
    .B(_0925_),
    .C(_0926_),
    .Y(_0927_));
 sg13g2_nor4_2 _1754_ (.A(_0923_),
    .B(_0900_),
    .C(_0924_),
    .Y(_0928_),
    .D(_0927_));
 sg13g2_a22oi_1 _1755_ (.Y(_0929_),
    .B1(_0859_),
    .B2(net41),
    .A2(_0858_),
    .A1(_0857_));
 sg13g2_nor2b_1 _1756_ (.A(_0929_),
    .B_N(_0853_),
    .Y(_0930_));
 sg13g2_nand2_1 _1757_ (.Y(_0931_),
    .A(_0771_),
    .B(_0734_));
 sg13g2_o21ai_1 _1758_ (.B1(_0931_),
    .Y(_0932_),
    .A1(_0591_),
    .A2(net26));
 sg13g2_o21ai_1 _1759_ (.B1(_0799_),
    .Y(_0933_),
    .A1(net35),
    .A2(_0734_));
 sg13g2_a221oi_1 _1760_ (.B2(net31),
    .C1(_0891_),
    .B1(_0933_),
    .A1(net35),
    .Y(_0934_),
    .A2(_0932_));
 sg13g2_nand3_1 _1761_ (.B(net75),
    .C(_0678_),
    .A(net41),
    .Y(_0935_));
 sg13g2_a21oi_1 _1762_ (.A1(_0002_),
    .A2(_0557_),
    .Y(_0936_),
    .B1(_0560_));
 sg13g2_a22oi_1 _1763_ (.Y(_0937_),
    .B1(_0936_),
    .B2(_0903_),
    .A2(_0019_),
    .A1(_0542_));
 sg13g2_o21ai_1 _1764_ (.B1(_0937_),
    .Y(_0938_),
    .A1(_0850_),
    .A2(_0935_));
 sg13g2_nor4_2 _1765_ (.A(_0928_),
    .B(_0930_),
    .C(_0934_),
    .Y(_0939_),
    .D(_0938_));
 sg13g2_buf_1 _1766_ (.A(\dac.accu1[3] ),
    .X(_0940_));
 sg13g2_nand2b_1 _1767_ (.Y(_0941_),
    .B(_0853_),
    .A_N(_0856_));
 sg13g2_a21o_1 _1768_ (.A2(_0834_),
    .A1(_0737_),
    .B1(net26),
    .X(_0942_));
 sg13g2_mux2_1 _1769_ (.A0(_0840_),
    .A1(_0942_),
    .S(_0680_),
    .X(_0943_));
 sg13g2_nand2_1 _1770_ (.Y(_0944_),
    .A(_0671_),
    .B(_0678_));
 sg13g2_or4_1 _1771_ (.A(_0654_),
    .B(net64),
    .C(_0943_),
    .D(_0944_),
    .X(_0945_));
 sg13g2_buf_1 _1772_ (.A(_0945_),
    .X(_0946_));
 sg13g2_or4_1 _1773_ (.A(_0549_),
    .B(net64),
    .C(_0837_),
    .D(_0944_),
    .X(_0947_));
 sg13g2_buf_1 _1774_ (.A(_0947_),
    .X(_0948_));
 sg13g2_and4_1 _1775_ (.A(net70),
    .B(_0941_),
    .C(_0946_),
    .D(_0948_),
    .X(_0949_));
 sg13g2_nor2b_1 _1776_ (.A(net75),
    .B_N(_0020_),
    .Y(_0950_));
 sg13g2_a221oi_1 _1777_ (.B2(_0594_),
    .C1(_0950_),
    .B1(_0903_),
    .A1(_0853_),
    .Y(_0951_),
    .A2(_0805_));
 sg13g2_buf_2 _1778_ (.A(_0951_),
    .X(_0952_));
 sg13g2_nor2_1 _1779_ (.A(net64),
    .B(_0762_),
    .Y(_0953_));
 sg13g2_or2_1 _1780_ (.X(_0954_),
    .B(_0874_),
    .A(_0625_));
 sg13g2_o21ai_1 _1781_ (.B1(_0878_),
    .Y(_0955_),
    .A1(_0689_),
    .A2(_0721_));
 sg13g2_nor2_1 _1782_ (.A(_0591_),
    .B(_0789_),
    .Y(_0956_));
 sg13g2_a221oi_1 _1783_ (.B2(_0639_),
    .C1(_0956_),
    .B1(_0955_),
    .A1(net31),
    .Y(_0957_),
    .A2(_0954_));
 sg13g2_nor2_1 _1784_ (.A(_0621_),
    .B(_0641_),
    .Y(_0958_));
 sg13g2_o21ai_1 _1785_ (.B1(net27),
    .Y(_0959_),
    .A1(_0819_),
    .A2(_0958_));
 sg13g2_a21o_1 _1786_ (.A2(_0959_),
    .A1(_0957_),
    .B1(net49),
    .X(_0960_));
 sg13g2_a22oi_1 _1787_ (.Y(_0961_),
    .B1(_0754_),
    .B2(_0773_),
    .A2(_0733_),
    .A1(_0680_));
 sg13g2_nand3_1 _1788_ (.B(net34),
    .C(_0661_),
    .A(net31),
    .Y(_0962_));
 sg13g2_a21oi_1 _1789_ (.A1(net58),
    .A2(_0749_),
    .Y(_0963_),
    .B1(net38));
 sg13g2_nand3_1 _1790_ (.B(_0962_),
    .C(_0963_),
    .A(_0961_),
    .Y(_0964_));
 sg13g2_a21oi_1 _1791_ (.A1(_0763_),
    .A2(_0641_),
    .Y(_0965_),
    .B1(_0663_));
 sg13g2_nor2_1 _1792_ (.A(net41),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_a21oi_1 _1793_ (.A1(_0964_),
    .A2(_0966_),
    .Y(_0967_),
    .B1(_0574_));
 sg13g2_a22oi_1 _1794_ (.Y(_0968_),
    .B1(_0960_),
    .B2(_0967_),
    .A2(_0953_),
    .A1(_0825_));
 sg13g2_buf_2 _1795_ (.A(_0968_),
    .X(_0969_));
 sg13g2_a22oi_1 _1796_ (.Y(_0970_),
    .B1(_0952_),
    .B2(_0969_),
    .A2(_0949_),
    .A1(_0939_));
 sg13g2_and4_1 _1797_ (.A(_0911_),
    .B(_0918_),
    .C(_0920_),
    .D(_0970_),
    .X(_0971_));
 sg13g2_buf_2 _1798_ (.A(\dac.accu1[2] ),
    .X(_0972_));
 sg13g2_a21oi_1 _1799_ (.A1(_0939_),
    .A2(_0949_),
    .Y(_0973_),
    .B1(_0972_));
 sg13g2_and4_1 _1800_ (.A(_0911_),
    .B(_0918_),
    .C(_0920_),
    .D(_0973_),
    .X(_0974_));
 sg13g2_inv_1 _1801_ (.Y(_0975_),
    .A(_0972_));
 sg13g2_and3_1 _1802_ (.X(_0976_),
    .A(_0941_),
    .B(_0946_),
    .C(_0948_));
 sg13g2_a21oi_1 _1803_ (.A1(_0939_),
    .A2(_0976_),
    .Y(_0977_),
    .B1(net70));
 sg13g2_a21o_1 _1804_ (.A2(_0970_),
    .A1(_0975_),
    .B1(_0977_),
    .X(_0978_));
 sg13g2_nor3_2 _1805_ (.A(_0971_),
    .B(_0974_),
    .C(_0978_),
    .Y(_0979_));
 sg13g2_o21ai_1 _1806_ (.B1(_0979_),
    .Y(_0980_),
    .A1(_0867_),
    .A2(_0870_));
 sg13g2_nand2_2 _1807_ (.Y(_0981_),
    .A(net21),
    .B(net25));
 sg13g2_nor2_1 _1808_ (.A(net71),
    .B(_0865_),
    .Y(_0982_));
 sg13g2_nand2_1 _1809_ (.Y(_0983_),
    .A(_0981_),
    .B(_0982_));
 sg13g2_a21oi_1 _1810_ (.A1(net21),
    .A2(net25),
    .Y(_0984_),
    .B1(_0865_));
 sg13g2_a22oi_1 _1811_ (.Y(_0985_),
    .B1(_0711_),
    .B2(_0598_),
    .A2(_0787_),
    .A1(_0786_));
 sg13g2_nand4_1 _1812_ (.B(_0786_),
    .C(_0787_),
    .A(_0598_),
    .Y(_0986_),
    .D(_0711_));
 sg13g2_o21ai_1 _1813_ (.B1(_0986_),
    .Y(_0987_),
    .A1(net72),
    .A2(_0985_));
 sg13g2_o21ai_1 _1814_ (.B1(_0987_),
    .Y(_0988_),
    .A1(_0984_),
    .A2(_0982_));
 sg13g2_and3_1 _1815_ (.X(_0989_),
    .A(_0980_),
    .B(_0983_),
    .C(_0988_));
 sg13g2_buf_1 _1816_ (.A(\dac.accu1[7] ),
    .X(_0990_));
 sg13g2_a221oi_1 _1817_ (.B2(_0852_),
    .C1(net46),
    .B1(_0705_),
    .A1(_0704_),
    .Y(_0991_),
    .A2(_0862_));
 sg13g2_a21oi_1 _1818_ (.A1(_0543_),
    .A2(_0015_),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_a21oi_1 _1819_ (.A1(net21),
    .A2(net25),
    .Y(_0993_),
    .B1(net71));
 sg13g2_or4_1 _1820_ (.A(_0992_),
    .B(_0979_),
    .C(_0987_),
    .D(_0993_),
    .X(_0994_));
 sg13g2_buf_2 _1821_ (.A(\dac.accu1[10] ),
    .X(_0995_));
 sg13g2_inv_1 _1822_ (.Y(_0996_),
    .A(_0995_));
 sg13g2_or2_1 _1823_ (.X(_0997_),
    .B(_0012_),
    .A(net48));
 sg13g2_nor3_1 _1824_ (.A(_0704_),
    .B(_0585_),
    .C(_0593_),
    .Y(_0998_));
 sg13g2_a221oi_1 _1825_ (.B2(_0824_),
    .C1(net77),
    .B1(_0818_),
    .A1(_0810_),
    .Y(_0999_),
    .A2(_0814_));
 sg13g2_or3_1 _1826_ (.A(_0567_),
    .B(_0998_),
    .C(_0999_),
    .X(_1000_));
 sg13g2_and2_1 _1827_ (.A(_0997_),
    .B(_1000_),
    .X(_1001_));
 sg13g2_buf_1 _1828_ (.A(_1001_),
    .X(_1002_));
 sg13g2_or2_1 _1829_ (.X(_1003_),
    .B(_0014_),
    .A(net75));
 sg13g2_buf_2 _1830_ (.A(_1003_),
    .X(_1004_));
 sg13g2_nor2_2 _1831_ (.A(net76),
    .B(net64),
    .Y(_1005_));
 sg13g2_nand2b_1 _1832_ (.Y(_1006_),
    .B(_0563_),
    .A_N(_0677_));
 sg13g2_nand2_1 _1833_ (.Y(_1007_),
    .A(_0704_),
    .B(_0703_));
 sg13g2_nand3_1 _1834_ (.B(_1006_),
    .C(_1007_),
    .A(_1005_),
    .Y(_1008_));
 sg13g2_buf_2 _1835_ (.A(_1008_),
    .X(_1009_));
 sg13g2_buf_2 _1836_ (.A(\dac.accu1[8] ),
    .X(_1010_));
 sg13g2_inv_1 _1837_ (.Y(_1011_),
    .A(_1010_));
 sg13g2_a21o_1 _1838_ (.A2(_1009_),
    .A1(_1004_),
    .B1(_1011_),
    .X(_1012_));
 sg13g2_a221oi_1 _1839_ (.B2(_0740_),
    .C1(net77),
    .B1(_0736_),
    .A1(_0719_),
    .Y(_1013_),
    .A2(_0725_));
 sg13g2_a21oi_1 _1840_ (.A1(_0563_),
    .A2(_0761_),
    .Y(_1014_),
    .B1(_1013_));
 sg13g2_nor2_1 _1841_ (.A(_0566_),
    .B(_0013_),
    .Y(_1015_));
 sg13g2_a21oi_2 _1842_ (.B1(_1015_),
    .Y(_1016_),
    .A2(_1014_),
    .A1(_1005_));
 sg13g2_buf_2 _1843_ (.A(\dac.accu1[9] ),
    .X(_1017_));
 sg13g2_inv_1 _1844_ (.Y(_1018_),
    .A(_1017_));
 sg13g2_a221oi_1 _1845_ (.B2(_1016_),
    .C1(_1018_),
    .B1(_1012_),
    .A1(_0996_),
    .Y(_1019_),
    .A2(_1002_));
 sg13g2_nand2_1 _1846_ (.Y(_1020_),
    .A(_0997_),
    .B(_1000_));
 sg13g2_inv_1 _1847_ (.Y(_1021_),
    .A(_1016_));
 sg13g2_a221oi_1 _1848_ (.B2(_1009_),
    .C1(_1011_),
    .B1(_1004_),
    .A1(_0996_),
    .Y(_1022_),
    .A2(_1002_));
 sg13g2_a22oi_1 _1849_ (.Y(_1023_),
    .B1(_1021_),
    .B2(_1022_),
    .A2(_1020_),
    .A1(_0995_));
 sg13g2_a221oi_1 _1850_ (.B2(_0560_),
    .C1(net77),
    .B1(_0850_),
    .A1(_0838_),
    .Y(_1024_),
    .A2(_0843_));
 sg13g2_a21oi_1 _1851_ (.A1(net77),
    .A2(_0936_),
    .Y(_1025_),
    .B1(_0567_));
 sg13g2_inv_1 _1852_ (.Y(_1026_),
    .A(_1025_));
 sg13g2_or2_1 _1853_ (.X(_1027_),
    .B(_0011_),
    .A(net48));
 sg13g2_o21ai_1 _1854_ (.B1(_1027_),
    .Y(_1028_),
    .A1(_1024_),
    .A2(_1026_));
 sg13g2_buf_1 _1855_ (.A(_1028_),
    .X(_1029_));
 sg13g2_inv_1 _1856_ (.Y(_1030_),
    .A(net20));
 sg13g2_nand3b_1 _1857_ (.B(_1023_),
    .C(_1030_),
    .Y(_1031_),
    .A_N(_1019_));
 sg13g2_a21oi_1 _1858_ (.A1(net69),
    .A2(_0994_),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_and4_1 _1859_ (.A(_0709_),
    .B(_0647_),
    .C(_0679_),
    .D(_0706_),
    .X(_1033_));
 sg13g2_a221oi_1 _1860_ (.B2(_1033_),
    .C1(_0780_),
    .B1(net72),
    .A1(net46),
    .Y(_1034_),
    .A2(_0017_));
 sg13g2_nor2_1 _1861_ (.A(net72),
    .B(_1033_),
    .Y(_1035_));
 sg13g2_o21ai_1 _1862_ (.B1(_0981_),
    .Y(_1036_),
    .A1(_1034_),
    .A2(_1035_));
 sg13g2_nand3_1 _1863_ (.B(_0865_),
    .C(_1036_),
    .A(net71),
    .Y(_1037_));
 sg13g2_nor3_1 _1864_ (.A(_0981_),
    .B(_1034_),
    .C(_1035_),
    .Y(_1038_));
 sg13g2_xnor2_1 _1865_ (.Y(_1039_),
    .A(_1017_),
    .B(_1016_));
 sg13g2_nand3_1 _1866_ (.B(_1004_),
    .C(_1009_),
    .A(_1011_),
    .Y(_1040_));
 sg13g2_xnor2_1 _1867_ (.Y(_1041_),
    .A(_0995_),
    .B(_1002_));
 sg13g2_nand4_1 _1868_ (.B(_1039_),
    .C(_1040_),
    .A(_1012_),
    .Y(_1042_),
    .D(_1041_));
 sg13g2_a21oi_1 _1869_ (.A1(_0865_),
    .A2(_1038_),
    .Y(_1043_),
    .B1(_1042_));
 sg13g2_nand3b_1 _1870_ (.B(_1023_),
    .C(_0010_),
    .Y(_1044_),
    .A_N(_1019_));
 sg13g2_a22oi_1 _1871_ (.Y(_1045_),
    .B1(_1044_),
    .B2(_1031_),
    .A2(_1043_),
    .A1(_1037_));
 sg13g2_a21oi_2 _1872_ (.B1(_1045_),
    .Y(_1046_),
    .A2(_1032_),
    .A1(_0989_));
 sg13g2_a21oi_1 _1873_ (.A1(net69),
    .A2(_0994_),
    .Y(_1047_),
    .B1(_1044_));
 sg13g2_a22oi_1 _1874_ (.Y(_1048_),
    .B1(_0989_),
    .B2(_1047_),
    .A2(_1030_),
    .A1(_0010_));
 sg13g2_buf_1 _1875_ (.A(_1048_),
    .X(_1049_));
 sg13g2_nor2_1 _1876_ (.A(_0781_),
    .B(_0007_),
    .Y(_1050_));
 sg13g2_a21o_1 _1877_ (.A2(_0677_),
    .A1(_0568_),
    .B1(_1050_),
    .X(_1051_));
 sg13g2_buf_2 _1878_ (.A(_1051_),
    .X(_1052_));
 sg13g2_xnor2_1 _1879_ (.Y(_1053_),
    .A(_0006_),
    .B(_1052_));
 sg13g2_buf_2 _1880_ (.A(\dac.accu1[13] ),
    .X(_1054_));
 sg13g2_or2_1 _1881_ (.X(_1055_),
    .B(_0005_),
    .A(_0781_));
 sg13g2_o21ai_1 _1882_ (.B1(_1055_),
    .Y(_1056_),
    .A1(_0574_),
    .A2(_0761_));
 sg13g2_buf_2 _1883_ (.A(_1056_),
    .X(_1057_));
 sg13g2_xor2_1 _1884_ (.B(_1057_),
    .A(_1054_),
    .X(_1058_));
 sg13g2_and2_1 _1885_ (.A(_1053_),
    .B(_1058_),
    .X(_1059_));
 sg13g2_nand4_1 _1886_ (.B(_1046_),
    .C(_1049_),
    .A(_0597_),
    .Y(_1060_),
    .D(_1059_));
 sg13g2_buf_2 _1887_ (.A(\dac.accu1[14] ),
    .X(_1061_));
 sg13g2_nand4_1 _1888_ (.B(_1046_),
    .C(_1049_),
    .A(_1061_),
    .Y(_1062_),
    .D(_1059_));
 sg13g2_inv_1 _1889_ (.Y(_1063_),
    .A(_1061_));
 sg13g2_inv_1 _1890_ (.Y(_1064_),
    .A(_1052_));
 sg13g2_nor2_1 _1891_ (.A(_0006_),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_a21o_1 _1892_ (.A2(_1065_),
    .A1(_1057_),
    .B1(_1054_),
    .X(_1066_));
 sg13g2_o21ai_1 _1893_ (.B1(_1066_),
    .Y(_1067_),
    .A1(_1057_),
    .A2(_1065_));
 sg13g2_a21oi_1 _1894_ (.A1(_1063_),
    .A2(_0596_),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_a21oi_1 _1895_ (.A1(_1061_),
    .A2(_0597_),
    .Y(_1069_),
    .B1(_1068_));
 sg13g2_nand3_1 _1896_ (.B(_1062_),
    .C(_1069_),
    .A(_1060_),
    .Y(_1070_));
 sg13g2_o21ai_1 _1897_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_0538_),
    .A2(_0571_));
 sg13g2_a21oi_1 _1898_ (.A1(_0538_),
    .A2(_0571_),
    .Y(_1072_),
    .B1(net85));
 sg13g2_a22oi_1 _1899_ (.Y(_0000_),
    .B1(_1071_),
    .B2(_1072_),
    .A2(_0537_),
    .A1(_0533_));
 sg13g2_nand2_1 _1900_ (.Y(_1073_),
    .A(_0915_),
    .B(\sine.ctr_r[0] ));
 sg13g2_buf_2 _1901_ (.A(\reg_out_w[1] ),
    .X(_1074_));
 sg13g2_xor2_1 _1902_ (.B(\sine.ctr_r[1] ),
    .A(_1074_),
    .X(_1075_));
 sg13g2_xnor2_1 _1903_ (.Y(_0031_),
    .A(_1073_),
    .B(_1075_));
 sg13g2_a21o_1 _1904_ (.A2(\sine.ctr_r[0] ),
    .A1(_0915_),
    .B1(\sine.ctr_r[1] ),
    .X(_1076_));
 sg13g2_and3_1 _1905_ (.X(_1077_),
    .A(_0915_),
    .B(\sine.ctr_r[1] ),
    .C(\sine.ctr_r[0] ));
 sg13g2_a21oi_1 _1906_ (.A1(_1074_),
    .A2(_1076_),
    .Y(_1078_),
    .B1(_1077_));
 sg13g2_buf_2 _1907_ (.A(\reg_out_w[2] ),
    .X(_1079_));
 sg13g2_xor2_1 _1908_ (.B(\sine.ctr_r[2] ),
    .A(_1079_),
    .X(_1080_));
 sg13g2_xnor2_1 _1909_ (.Y(_0032_),
    .A(_1078_),
    .B(_1080_));
 sg13g2_a221oi_1 _1910_ (.B2(_1074_),
    .C1(_1077_),
    .B1(_1076_),
    .A1(_1079_),
    .Y(_1081_),
    .A2(\sine.ctr_r[2] ));
 sg13g2_buf_1 _1911_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nor2_2 _1912_ (.A(_1079_),
    .B(\sine.ctr_r[2] ),
    .Y(_1083_));
 sg13g2_nor2_1 _1913_ (.A(_1082_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_buf_2 _1914_ (.A(\reg_out_w[3] ),
    .X(_1085_));
 sg13g2_xnor2_1 _1915_ (.Y(_1086_),
    .A(_1085_),
    .B(\sine.ctr_r[3] ));
 sg13g2_xnor2_1 _1916_ (.Y(_0033_),
    .A(_1084_),
    .B(_1086_));
 sg13g2_inv_1 _1917_ (.Y(_1087_),
    .A(\sine.ctr_r[3] ));
 sg13g2_o21ai_1 _1918_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1082_),
    .A2(_1083_));
 sg13g2_nor3_1 _1919_ (.A(_1087_),
    .B(_1082_),
    .C(_1083_),
    .Y(_1089_));
 sg13g2_a21o_1 _1920_ (.A2(_1088_),
    .A1(_1085_),
    .B1(_1089_),
    .X(_1090_));
 sg13g2_buf_2 _1921_ (.A(_1090_),
    .X(_1091_));
 sg13g2_buf_2 _1922_ (.A(\sine.ctr_r[4] ),
    .X(_1092_));
 sg13g2_xnor2_1 _1923_ (.Y(_1093_),
    .A(\reg_out_w[4] ),
    .B(_1092_));
 sg13g2_xnor2_1 _1924_ (.Y(_0034_),
    .A(_1091_),
    .B(_1093_));
 sg13g2_nor2_1 _1925_ (.A(\sine.ctr_r[3] ),
    .B(_1092_),
    .Y(_1094_));
 sg13g2_o21ai_1 _1926_ (.B1(_1094_),
    .Y(_1095_),
    .A1(_1082_),
    .A2(_1083_));
 sg13g2_nor2_1 _1927_ (.A(_1085_),
    .B(_1092_),
    .Y(_1096_));
 sg13g2_o21ai_1 _1928_ (.B1(_1096_),
    .Y(_1097_),
    .A1(_1082_),
    .A2(_1083_));
 sg13g2_nor3_1 _1929_ (.A(_1085_),
    .B(\sine.ctr_r[3] ),
    .C(_1092_),
    .Y(_1098_));
 sg13g2_nor2b_1 _1930_ (.A(_1098_),
    .B_N(\reg_out_w[4] ),
    .Y(_1099_));
 sg13g2_and3_1 _1931_ (.X(_1100_),
    .A(_1095_),
    .B(_1097_),
    .C(_1099_));
 sg13g2_buf_1 _1932_ (.A(_1100_),
    .X(_1101_));
 sg13g2_a21oi_1 _1933_ (.A1(_1092_),
    .A2(_1091_),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_buf_2 _1934_ (.A(\sine.ctr_r[5] ),
    .X(_1103_));
 sg13g2_xor2_1 _1935_ (.B(_1103_),
    .A(\reg_out_w[5] ),
    .X(_1104_));
 sg13g2_xnor2_1 _1936_ (.Y(_0035_),
    .A(_1102_),
    .B(_1104_));
 sg13g2_and2_1 _1937_ (.A(_1092_),
    .B(_1103_),
    .X(_1105_));
 sg13g2_buf_1 _1938_ (.A(_1105_),
    .X(_1106_));
 sg13g2_inv_2 _1939_ (.Y(_1107_),
    .A(\reg_out_w[5] ));
 sg13g2_and2_1 _1940_ (.A(_1095_),
    .B(_1097_),
    .X(_1108_));
 sg13g2_a221oi_1 _1941_ (.B2(_1099_),
    .C1(_1103_),
    .B1(_1108_),
    .A1(_1092_),
    .Y(_1109_),
    .A2(_1091_));
 sg13g2_buf_1 _1942_ (.A(_1109_),
    .X(_1110_));
 sg13g2_nor2_1 _1943_ (.A(_1107_),
    .B(_1110_),
    .Y(_1111_));
 sg13g2_a221oi_1 _1944_ (.B2(_1091_),
    .C1(_1111_),
    .B1(_1106_),
    .A1(_1103_),
    .Y(_1112_),
    .A2(_1101_));
 sg13g2_buf_1 _1945_ (.A(\reg_out_w[6] ),
    .X(_1113_));
 sg13g2_buf_2 _1946_ (.A(\sine.ctr_r[6] ),
    .X(_1114_));
 sg13g2_xor2_1 _1947_ (.B(_1114_),
    .A(_1113_),
    .X(_1115_));
 sg13g2_xnor2_1 _1948_ (.Y(_0036_),
    .A(_1112_),
    .B(_1115_));
 sg13g2_inv_1 _1949_ (.Y(_1116_),
    .A(_1113_));
 sg13g2_nor2b_1 _1950_ (.A(_1114_),
    .B_N(_1112_),
    .Y(_1117_));
 sg13g2_nand2b_1 _1951_ (.Y(_1118_),
    .B(_1114_),
    .A_N(_1112_));
 sg13g2_o21ai_1 _1952_ (.B1(_1118_),
    .Y(_1119_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_buf_2 _1953_ (.A(\reg_out_w[7] ),
    .X(_1120_));
 sg13g2_xnor2_1 _1954_ (.Y(_1121_),
    .A(_1120_),
    .B(\sine.ctr_r[7] ));
 sg13g2_xnor2_1 _1955_ (.Y(_0037_),
    .A(_1119_),
    .B(_1121_));
 sg13g2_buf_2 _1956_ (.A(\reg_out_w[8] ),
    .X(_1122_));
 sg13g2_xor2_1 _1957_ (.B(\sine.ctr_r[8] ),
    .A(_1122_),
    .X(_1123_));
 sg13g2_or2_1 _1958_ (.X(_1124_),
    .B(\sine.ctr_r[7] ),
    .A(_1114_));
 sg13g2_a221oi_1 _1959_ (.B2(_1091_),
    .C1(_1124_),
    .B1(_1106_),
    .A1(_1103_),
    .Y(_1125_),
    .A2(_1101_));
 sg13g2_o21ai_1 _1960_ (.B1(_1125_),
    .Y(_1126_),
    .A1(_1107_),
    .A2(_1110_));
 sg13g2_or2_1 _1961_ (.X(_1127_),
    .B(\sine.ctr_r[7] ),
    .A(_1113_));
 sg13g2_a221oi_1 _1962_ (.B2(_1091_),
    .C1(_1127_),
    .B1(_1106_),
    .A1(_1103_),
    .Y(_1128_),
    .A2(_1101_));
 sg13g2_o21ai_1 _1963_ (.B1(_1128_),
    .Y(_1129_),
    .A1(_1107_),
    .A2(_1110_));
 sg13g2_or2_1 _1964_ (.X(_1130_),
    .B(_1114_),
    .A(_1120_));
 sg13g2_a221oi_1 _1965_ (.B2(_1091_),
    .C1(_1130_),
    .B1(_1106_),
    .A1(_1103_),
    .Y(_1131_),
    .A2(_1101_));
 sg13g2_o21ai_1 _1966_ (.B1(_1131_),
    .Y(_1132_),
    .A1(_1107_),
    .A2(_1110_));
 sg13g2_or2_1 _1967_ (.X(_1133_),
    .B(_1113_),
    .A(_1120_));
 sg13g2_a221oi_1 _1968_ (.B2(_1091_),
    .C1(_1133_),
    .B1(_1106_),
    .A1(_1103_),
    .Y(_1134_),
    .A2(_1101_));
 sg13g2_o21ai_1 _1969_ (.B1(_1134_),
    .Y(_1135_),
    .A1(_1107_),
    .A2(_1110_));
 sg13g2_and4_1 _1970_ (.A(_1126_),
    .B(_1129_),
    .C(_1132_),
    .D(_1135_),
    .X(_1136_));
 sg13g2_nor2_1 _1971_ (.A(_1120_),
    .B(\sine.ctr_r[7] ),
    .Y(_1137_));
 sg13g2_nor3_1 _1972_ (.A(_1113_),
    .B(_1114_),
    .C(\sine.ctr_r[7] ),
    .Y(_1138_));
 sg13g2_nor2_1 _1973_ (.A(_1114_),
    .B(_1133_),
    .Y(_1139_));
 sg13g2_nor3_1 _1974_ (.A(_1137_),
    .B(_1138_),
    .C(_1139_),
    .Y(_1140_));
 sg13g2_nand2_1 _1975_ (.Y(_1141_),
    .A(_1136_),
    .B(_1140_));
 sg13g2_xnor2_1 _1976_ (.Y(_0038_),
    .A(_1123_),
    .B(_1141_));
 sg13g2_nand2_1 _1977_ (.Y(_1142_),
    .A(_1122_),
    .B(\sine.ctr_r[8] ));
 sg13g2_nor2_1 _1978_ (.A(_1122_),
    .B(\sine.ctr_r[8] ),
    .Y(_1143_));
 sg13g2_a21oi_2 _1979_ (.B1(_1143_),
    .Y(_1144_),
    .A2(_1142_),
    .A1(_1141_));
 sg13g2_buf_2 _1980_ (.A(\reg_out_w[9] ),
    .X(_1145_));
 sg13g2_buf_1 _1981_ (.A(\sine.ctr_r[9] ),
    .X(_1146_));
 sg13g2_xnor2_1 _1982_ (.Y(_1147_),
    .A(_1145_),
    .B(_1146_));
 sg13g2_xnor2_1 _1983_ (.Y(_0039_),
    .A(_1144_),
    .B(_1147_));
 sg13g2_a21o_1 _1984_ (.A2(_1144_),
    .A1(_1146_),
    .B1(_1145_),
    .X(_1148_));
 sg13g2_o21ai_1 _1985_ (.B1(_1148_),
    .Y(_1149_),
    .A1(_1146_),
    .A2(_1144_));
 sg13g2_buf_2 _1986_ (.A(\reg_out_w[10] ),
    .X(_1150_));
 sg13g2_xor2_1 _1987_ (.B(\sine.ctr_r[10] ),
    .A(_1150_),
    .X(_1151_));
 sg13g2_xnor2_1 _1988_ (.Y(_0025_),
    .A(_1149_),
    .B(_1151_));
 sg13g2_and2_1 _1989_ (.A(_1150_),
    .B(\sine.ctr_r[10] ),
    .X(_1152_));
 sg13g2_a21oi_1 _1990_ (.A1(_1122_),
    .A2(\sine.ctr_r[8] ),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_nand2b_1 _1991_ (.Y(_1154_),
    .B(_1153_),
    .A_N(_1146_));
 sg13g2_nand2b_1 _1992_ (.Y(_1155_),
    .B(_1153_),
    .A_N(_1145_));
 sg13g2_a22oi_1 _1993_ (.Y(_1156_),
    .B1(_1154_),
    .B2(_1155_),
    .A2(_1140_),
    .A1(_1136_));
 sg13g2_or2_1 _1994_ (.X(_1157_),
    .B(\sine.ctr_r[8] ),
    .A(_1122_));
 sg13g2_a221oi_1 _1995_ (.B2(_1150_),
    .C1(_1157_),
    .B1(\sine.ctr_r[10] ),
    .A1(_1145_),
    .Y(_1158_),
    .A2(_1146_));
 sg13g2_nor3_1 _1996_ (.A(_1145_),
    .B(_1146_),
    .C(_1152_),
    .Y(_1159_));
 sg13g2_nor2_1 _1997_ (.A(_1150_),
    .B(\sine.ctr_r[10] ),
    .Y(_1160_));
 sg13g2_nor4_2 _1998_ (.A(_1156_),
    .B(_1158_),
    .C(_1159_),
    .Y(_1161_),
    .D(_1160_));
 sg13g2_xnor2_1 _1999_ (.Y(_1162_),
    .A(\reg_out_w[11] ),
    .B(\sine.ctr_r[11] ));
 sg13g2_xnor2_1 _2000_ (.Y(_0026_),
    .A(_1161_),
    .B(_1162_));
 sg13g2_a21oi_1 _2001_ (.A1(\sine.ctr_r[11] ),
    .A2(_1161_),
    .Y(_1163_),
    .B1(\reg_out_w[11] ));
 sg13g2_nor2_1 _2002_ (.A(\sine.ctr_r[11] ),
    .B(_1161_),
    .Y(_1164_));
 sg13g2_nor2_1 _2003_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_xnor2_1 _2004_ (.Y(_1166_),
    .A(\reg_out_w[12] ),
    .B(\sine.ctr_r[12] ));
 sg13g2_xnor2_1 _2005_ (.Y(_0027_),
    .A(_1165_),
    .B(_1166_));
 sg13g2_inv_1 _2006_ (.Y(_1167_),
    .A(\reg_out_w[12] ));
 sg13g2_inv_1 _2007_ (.Y(_1168_),
    .A(\sine.ctr_r[12] ));
 sg13g2_nor2_1 _2008_ (.A(_1167_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_nand2_1 _2009_ (.Y(_1170_),
    .A(_1167_),
    .B(_1168_));
 sg13g2_o21ai_1 _2010_ (.B1(_1170_),
    .Y(_1171_),
    .A1(_1165_),
    .A2(_1169_));
 sg13g2_xor2_1 _2011_ (.B(\sine.ctr_r[13] ),
    .A(\reg_out_w[13] ),
    .X(_1172_));
 sg13g2_xnor2_1 _2012_ (.Y(_0028_),
    .A(_1171_),
    .B(_1172_));
 sg13g2_buf_2 _2013_ (.A(\reg_out_w[14] ),
    .X(_1173_));
 sg13g2_xnor2_1 _2014_ (.Y(_1174_),
    .A(_1173_),
    .B(\sine.ctr_r[14] ));
 sg13g2_inv_1 _2015_ (.Y(_1175_),
    .A(\sine.ctr_r[13] ));
 sg13g2_inv_1 _2016_ (.Y(_1176_),
    .A(\reg_out_w[13] ));
 sg13g2_or2_1 _2017_ (.X(_1177_),
    .B(_1164_),
    .A(_1163_));
 sg13g2_a221oi_1 _2018_ (.B2(_1176_),
    .C1(_1177_),
    .B1(_1175_),
    .A1(_1167_),
    .Y(_1178_),
    .A2(_1168_));
 sg13g2_nand2_1 _2019_ (.Y(_1179_),
    .A(\reg_out_w[13] ),
    .B(\sine.ctr_r[13] ));
 sg13g2_o21ai_1 _2020_ (.B1(_1169_),
    .Y(_1180_),
    .A1(\reg_out_w[13] ),
    .A2(\sine.ctr_r[13] ));
 sg13g2_nand3b_1 _2021_ (.B(_1179_),
    .C(_1180_),
    .Y(_1181_),
    .A_N(_1178_));
 sg13g2_xnor2_1 _2022_ (.Y(_0029_),
    .A(_1174_),
    .B(_1181_));
 sg13g2_xor2_1 _2023_ (.B(\sine.ctr_r[15] ),
    .A(\reg_out_w[15] ),
    .X(_1182_));
 sg13g2_or2_1 _2024_ (.X(_1183_),
    .B(\sine.ctr_r[14] ),
    .A(_1173_));
 sg13g2_and2_1 _2025_ (.A(_1173_),
    .B(\sine.ctr_r[14] ),
    .X(_1184_));
 sg13g2_a21oi_1 _2026_ (.A1(_1181_),
    .A2(_1183_),
    .Y(_1185_),
    .B1(_1184_));
 sg13g2_xnor2_1 _2027_ (.Y(_0030_),
    .A(_1182_),
    .B(_1185_));
 sg13g2_xor2_1 _2028_ (.B(\sine.ctr_r[0] ),
    .A(_0915_),
    .X(_0024_));
 sg13g2_inv_2 _2029_ (.Y(_1186_),
    .A(net5));
 sg13g2_nand2_1 _2030_ (.Y(_1187_),
    .A(_0873_),
    .B(_0888_));
 sg13g2_o21ai_1 _2031_ (.B1(_1187_),
    .Y(_1188_),
    .A1(_0916_),
    .A2(net48));
 sg13g2_xnor2_1 _2032_ (.Y(_1189_),
    .A(_0906_),
    .B(_1188_));
 sg13g2_or2_1 _2033_ (.X(_1190_),
    .B(\dac.mod2_ctr[0] ),
    .A(\dac.mod2_ctr[1] ));
 sg13g2_buf_1 _2034_ (.A(_1190_),
    .X(_1191_));
 sg13g2_buf_1 _2035_ (.A(_1191_),
    .X(_1192_));
 sg13g2_xnor2_1 _2036_ (.Y(_1193_),
    .A(\dac.accu2[0] ),
    .B(_1188_));
 sg13g2_buf_1 _2037_ (.A(_1191_),
    .X(_1194_));
 sg13g2_nand2_1 _2038_ (.Y(_1195_),
    .A(_0906_),
    .B(net29));
 sg13g2_o21ai_1 _2039_ (.B1(_1195_),
    .Y(_1196_),
    .A1(net30),
    .A2(_1193_));
 sg13g2_nor2_1 _2040_ (.A(_1186_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_a21oi_1 _2041_ (.A1(_1186_),
    .A2(_1189_),
    .Y(_0040_),
    .B1(_1197_));
 sg13g2_nand2_1 _2042_ (.Y(_1198_),
    .A(_1004_),
    .B(_1009_));
 sg13g2_a21oi_1 _2043_ (.A1(net71),
    .A2(_1036_),
    .Y(_1199_),
    .B1(_1038_));
 sg13g2_nor2_1 _2044_ (.A(_0992_),
    .B(_1199_),
    .Y(_1200_));
 sg13g2_nand2_1 _2045_ (.Y(_1201_),
    .A(net69),
    .B(_0994_));
 sg13g2_o21ai_1 _2046_ (.B1(_0989_),
    .Y(_1202_),
    .A1(_1200_),
    .A2(_1201_));
 sg13g2_buf_1 _2047_ (.A(_1202_),
    .X(_1203_));
 sg13g2_a221oi_1 _2048_ (.B2(_1017_),
    .C1(_1203_),
    .B1(_1021_),
    .A1(_1010_),
    .Y(_1204_),
    .A2(_1198_));
 sg13g2_nor2_1 _2049_ (.A(_1018_),
    .B(_1016_),
    .Y(_1205_));
 sg13g2_nand2_1 _2050_ (.Y(_1206_),
    .A(_1018_),
    .B(_1016_));
 sg13g2_o21ai_1 _2051_ (.B1(_1206_),
    .Y(_1207_),
    .A1(_1205_),
    .A2(_1040_));
 sg13g2_nor2_1 _2052_ (.A(_1204_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_xnor2_1 _2053_ (.Y(_1209_),
    .A(_1041_),
    .B(_1208_));
 sg13g2_buf_1 _2054_ (.A(net85),
    .X(_1210_));
 sg13g2_nand2_1 _2055_ (.Y(_1211_),
    .A(_0709_),
    .B(\dac.accu2[5] ));
 sg13g2_nand2b_1 _2056_ (.Y(_1212_),
    .B(_0598_),
    .A_N(\dac.accu2[5] ));
 sg13g2_a21oi_1 _2057_ (.A1(_1211_),
    .A2(_1212_),
    .Y(_1213_),
    .B1(_0782_));
 sg13g2_nand2_1 _2058_ (.Y(_1214_),
    .A(_1211_),
    .B(_1212_));
 sg13g2_a21oi_1 _2059_ (.A1(_0786_),
    .A2(_0787_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_a21o_1 _2060_ (.A2(_1213_),
    .A1(_0786_),
    .B1(_1215_),
    .X(_1216_));
 sg13g2_buf_1 _2061_ (.A(\dac.accu2[4] ),
    .X(_1217_));
 sg13g2_or4_2 _2062_ (.A(_0928_),
    .B(_0930_),
    .C(_0934_),
    .D(_0938_),
    .X(_1218_));
 sg13g2_nand3_1 _2063_ (.B(_0946_),
    .C(_0948_),
    .A(_0941_),
    .Y(_1219_));
 sg13g2_nor3_2 _2064_ (.A(\dac.accu2[3] ),
    .B(_1218_),
    .C(_1219_),
    .Y(_1220_));
 sg13g2_nand4_1 _2065_ (.B(_0941_),
    .C(_0946_),
    .A(_0972_),
    .Y(_1221_),
    .D(_0948_));
 sg13g2_inv_1 _2066_ (.Y(_1222_),
    .A(\dac.accu2[3] ));
 sg13g2_nand2_1 _2067_ (.Y(_1223_),
    .A(_0972_),
    .B(_1222_));
 sg13g2_o21ai_1 _2068_ (.B1(_1223_),
    .Y(_1224_),
    .A1(_1218_),
    .A2(_1221_));
 sg13g2_o21ai_1 _2069_ (.B1(_0711_),
    .Y(_1225_),
    .A1(_1220_),
    .A2(_1224_));
 sg13g2_nor3_1 _2070_ (.A(_0711_),
    .B(_1220_),
    .C(_1224_),
    .Y(_1226_));
 sg13g2_a21oi_1 _2071_ (.A1(_1217_),
    .A2(_1225_),
    .Y(_1227_),
    .B1(_1226_));
 sg13g2_nand2_1 _2072_ (.Y(_1228_),
    .A(_1216_),
    .B(_1227_));
 sg13g2_nor2_2 _2073_ (.A(_1218_),
    .B(_1219_),
    .Y(_1229_));
 sg13g2_xnor2_1 _2074_ (.Y(_1230_),
    .A(_0972_),
    .B(\dac.accu2[3] ));
 sg13g2_xnor2_1 _2075_ (.Y(_1231_),
    .A(_1229_),
    .B(_1230_));
 sg13g2_inv_1 _2076_ (.Y(_1232_),
    .A(\dac.accu2[2] ));
 sg13g2_nand3_1 _2077_ (.B(_0952_),
    .C(_0969_),
    .A(_1232_),
    .Y(_1233_));
 sg13g2_a21oi_1 _2078_ (.A1(_0952_),
    .A2(_0969_),
    .Y(_1234_),
    .B1(_1232_));
 sg13g2_a21oi_2 _2079_ (.B1(_1234_),
    .Y(_1235_),
    .A2(_1233_),
    .A1(_0913_));
 sg13g2_nand2b_1 _2080_ (.Y(_1236_),
    .B(_1235_),
    .A_N(_1231_));
 sg13g2_nor2_1 _2081_ (.A(_0743_),
    .B(_0779_),
    .Y(_1237_));
 sg13g2_nor2_1 _2082_ (.A(net46),
    .B(_1214_),
    .Y(_1238_));
 sg13g2_nor2_1 _2083_ (.A(_0787_),
    .B(_1214_),
    .Y(_1239_));
 sg13g2_a221oi_1 _2084_ (.B2(_0786_),
    .C1(_1239_),
    .B1(_1213_),
    .A1(_1237_),
    .Y(_1240_),
    .A2(_1238_));
 sg13g2_buf_1 _2085_ (.A(_1240_),
    .X(_1241_));
 sg13g2_nor2_1 _2086_ (.A(_1241_),
    .B(_1226_),
    .Y(_1242_));
 sg13g2_a21oi_1 _2087_ (.A1(_1241_),
    .A2(_1225_),
    .Y(_1243_),
    .B1(_1217_));
 sg13g2_o21ai_1 _2088_ (.B1(net70),
    .Y(_1244_),
    .A1(_1242_),
    .A2(_1243_));
 sg13g2_xor2_1 _2089_ (.B(\dac.accu2[2] ),
    .A(_0912_),
    .X(_1245_));
 sg13g2_a21o_1 _2090_ (.A2(_0969_),
    .A1(_0952_),
    .B1(_1245_),
    .X(_1246_));
 sg13g2_o21ai_1 _2091_ (.B1(\dac.accu2[0] ),
    .Y(_1247_),
    .A1(_0916_),
    .A2(net84));
 sg13g2_a21o_1 _2092_ (.A2(_0887_),
    .A1(_0883_),
    .B1(_1247_),
    .X(_1248_));
 sg13g2_buf_1 _2093_ (.A(_1248_),
    .X(_1249_));
 sg13g2_nor2_1 _2094_ (.A(_0742_),
    .B(_1247_),
    .Y(_1250_));
 sg13g2_nor2_1 _2095_ (.A(_0762_),
    .B(_1247_),
    .Y(_1251_));
 sg13g2_a22oi_1 _2096_ (.Y(_1252_),
    .B1(_1251_),
    .B2(_0703_),
    .A2(_1250_),
    .A1(_0872_));
 sg13g2_buf_1 _2097_ (.A(_1252_),
    .X(_1253_));
 sg13g2_nor4_2 _2098_ (.A(_0889_),
    .B(_0902_),
    .C(_0904_),
    .Y(_1254_),
    .D(_0909_));
 sg13g2_a21oi_2 _2099_ (.B1(_1254_),
    .Y(_1255_),
    .A2(_1253_),
    .A1(_1249_));
 sg13g2_nor3_1 _2100_ (.A(_0907_),
    .B(_1246_),
    .C(_1255_),
    .Y(_1256_));
 sg13g2_buf_1 _2101_ (.A(\dac.accu2[1] ),
    .X(_1257_));
 sg13g2_nor2_1 _2102_ (.A(_0907_),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_nand4_1 _2103_ (.B(_1249_),
    .C(_1253_),
    .A(_1254_),
    .Y(_1259_),
    .D(_1258_));
 sg13g2_nand4_1 _2104_ (.B(_0969_),
    .C(_1245_),
    .A(_0952_),
    .Y(_1260_),
    .D(_1258_));
 sg13g2_nand2b_1 _2105_ (.Y(_1261_),
    .B(_0906_),
    .A_N(_1257_));
 sg13g2_or2_1 _2106_ (.X(_1262_),
    .B(_1261_),
    .A(_1245_));
 sg13g2_a21o_1 _2107_ (.A2(_0969_),
    .A1(_0952_),
    .B1(_1262_),
    .X(_1263_));
 sg13g2_nand3_1 _2108_ (.B(_1260_),
    .C(_1263_),
    .A(_1259_),
    .Y(_1264_));
 sg13g2_nand3_1 _2109_ (.B(_0969_),
    .C(_1245_),
    .A(_0952_),
    .Y(_1265_));
 sg13g2_nor3_1 _2110_ (.A(_0907_),
    .B(_1255_),
    .C(_1265_),
    .Y(_1266_));
 sg13g2_nand3_1 _2111_ (.B(_1249_),
    .C(_1253_),
    .A(_1254_),
    .Y(_1267_));
 sg13g2_a221oi_1 _2112_ (.B2(_1257_),
    .C1(_1255_),
    .B1(_1267_),
    .A1(_1246_),
    .Y(_1268_),
    .A2(_1265_));
 sg13g2_or4_1 _2113_ (.A(_1256_),
    .B(_1264_),
    .C(_1266_),
    .D(_1268_),
    .X(_1269_));
 sg13g2_buf_2 _2114_ (.A(_1269_),
    .X(_1270_));
 sg13g2_nand2b_1 _2115_ (.Y(_1271_),
    .B(_1231_),
    .A_N(_1235_));
 sg13g2_nand2_1 _2116_ (.Y(_1272_),
    .A(_1270_),
    .B(_1271_));
 sg13g2_nand4_1 _2117_ (.B(_1236_),
    .C(_1244_),
    .A(_1228_),
    .Y(_1273_),
    .D(_1272_));
 sg13g2_nor2b_1 _2118_ (.A(\dac.accu2[8] ),
    .B_N(net69),
    .Y(_1274_));
 sg13g2_nor2b_1 _2119_ (.A(net69),
    .B_N(\dac.accu2[8] ),
    .Y(_1275_));
 sg13g2_or2_1 _2120_ (.X(_1276_),
    .B(_1275_),
    .A(_1274_));
 sg13g2_buf_1 _2121_ (.A(_1276_),
    .X(_1277_));
 sg13g2_nand4_1 _2122_ (.B(_1006_),
    .C(_1007_),
    .A(_1005_),
    .Y(_1278_),
    .D(_1277_));
 sg13g2_nand2b_1 _2123_ (.Y(_1279_),
    .B(_1004_),
    .A_N(_1277_));
 sg13g2_a21o_1 _2124_ (.A2(_1007_),
    .A1(_1006_),
    .B1(_1279_),
    .X(_1280_));
 sg13g2_nor2_1 _2125_ (.A(net75),
    .B(_0014_),
    .Y(_1281_));
 sg13g2_nor3_1 _2126_ (.A(_1005_),
    .B(_1281_),
    .C(_1277_),
    .Y(_1282_));
 sg13g2_a21oi_1 _2127_ (.A1(_1281_),
    .A2(_1277_),
    .Y(_1283_),
    .B1(_1282_));
 sg13g2_nand3_1 _2128_ (.B(_1280_),
    .C(_1283_),
    .A(_1278_),
    .Y(_1284_));
 sg13g2_nand2_1 _2129_ (.Y(_0116_),
    .A(net71),
    .B(\dac.accu2[7] ));
 sg13g2_o21ai_1 _2130_ (.B1(_0116_),
    .Y(_0117_),
    .A1(net48),
    .A2(_0831_));
 sg13g2_nand2b_1 _2131_ (.Y(_0118_),
    .B(\dac.accu1[6] ),
    .A_N(\dac.accu2[7] ));
 sg13g2_o21ai_1 _2132_ (.B1(_0118_),
    .Y(_0119_),
    .A1(_0991_),
    .A2(_0117_));
 sg13g2_buf_2 _2133_ (.A(_0119_),
    .X(_0120_));
 sg13g2_xor2_1 _2134_ (.B(_0120_),
    .A(_1284_),
    .X(_0121_));
 sg13g2_xnor2_1 _2135_ (.Y(_0122_),
    .A(_1010_),
    .B(\dac.accu2[9] ));
 sg13g2_nor2_1 _2136_ (.A(_0567_),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_nor2b_1 _2137_ (.A(_1015_),
    .B_N(_0122_),
    .Y(_0124_));
 sg13g2_nand4_1 _2138_ (.B(_0748_),
    .C(_0757_),
    .A(net77),
    .Y(_0125_),
    .D(_0760_));
 sg13g2_nand3b_1 _2139_ (.B(_1005_),
    .C(_0125_),
    .Y(_0126_),
    .A_N(_1013_));
 sg13g2_nor2b_1 _2140_ (.A(_0122_),
    .B_N(_1015_),
    .Y(_0127_));
 sg13g2_a221oi_1 _2141_ (.B2(_0126_),
    .C1(_0127_),
    .B1(_0124_),
    .A1(_1014_),
    .Y(_0128_),
    .A2(_0123_));
 sg13g2_buf_1 _2142_ (.A(_0128_),
    .X(_0129_));
 sg13g2_nor2_1 _2143_ (.A(_1004_),
    .B(_1275_),
    .Y(_0130_));
 sg13g2_nor2_1 _2144_ (.A(_1274_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_o21ai_1 _2145_ (.B1(_0131_),
    .Y(_0132_),
    .A1(_1009_),
    .A2(_1275_));
 sg13g2_buf_1 _2146_ (.A(_0132_),
    .X(_0133_));
 sg13g2_xnor2_1 _2147_ (.Y(_0134_),
    .A(_0129_),
    .B(_0133_));
 sg13g2_nand2_2 _2148_ (.Y(_0135_),
    .A(_0121_),
    .B(_0134_));
 sg13g2_nor3_1 _2149_ (.A(net70),
    .B(_1242_),
    .C(_1243_),
    .Y(_0136_));
 sg13g2_nand2_1 _2150_ (.Y(_0137_),
    .A(_0118_),
    .B(_0116_));
 sg13g2_xor2_1 _2151_ (.B(_0137_),
    .A(_0865_),
    .X(_0138_));
 sg13g2_buf_1 _2152_ (.A(_0138_),
    .X(_0139_));
 sg13g2_inv_1 _2153_ (.Y(_0140_),
    .A(\dac.accu2[6] ));
 sg13g2_nand2_1 _2154_ (.Y(_0141_),
    .A(\dac.accu1[5] ),
    .B(_0140_));
 sg13g2_nand3_1 _2155_ (.B(net25),
    .C(_0141_),
    .A(net21),
    .Y(_0142_));
 sg13g2_nand2_1 _2156_ (.Y(_0143_),
    .A(net72),
    .B(\dac.accu2[6] ));
 sg13g2_nand2_1 _2157_ (.Y(_0144_),
    .A(_0142_),
    .B(_0143_));
 sg13g2_xor2_1 _2158_ (.B(_0144_),
    .A(net19),
    .X(_0145_));
 sg13g2_nand2_1 _2159_ (.Y(_0146_),
    .A(_0141_),
    .B(_0143_));
 sg13g2_a21oi_1 _2160_ (.A1(net21),
    .A2(net25),
    .Y(_0147_),
    .B1(_0146_));
 sg13g2_and3_1 _2161_ (.X(_0148_),
    .A(net21),
    .B(net25),
    .C(_0146_));
 sg13g2_o21ai_1 _2162_ (.B1(_1212_),
    .Y(_0149_),
    .A1(net48),
    .A2(_0017_));
 sg13g2_nand2_1 _2163_ (.Y(_0150_),
    .A(_1211_),
    .B(_0149_));
 sg13g2_a21oi_1 _2164_ (.A1(_0709_),
    .A2(\dac.accu2[5] ),
    .Y(_0151_),
    .B1(net46));
 sg13g2_o21ai_1 _2165_ (.B1(_0151_),
    .Y(_0152_),
    .A1(_0743_),
    .A2(_0779_));
 sg13g2_and2_1 _2166_ (.A(_0150_),
    .B(_0152_),
    .X(_0153_));
 sg13g2_o21ai_1 _2167_ (.B1(_0153_),
    .Y(_0154_),
    .A1(_0147_),
    .A2(_0148_));
 sg13g2_or3_1 _2168_ (.A(_0153_),
    .B(_0147_),
    .C(_0148_),
    .X(_0155_));
 sg13g2_nand2b_1 _2169_ (.Y(_0156_),
    .B(_0711_),
    .A_N(_1217_));
 sg13g2_nand4_1 _2170_ (.B(_0647_),
    .C(_0679_),
    .A(_1217_),
    .Y(_0157_),
    .D(_0706_));
 sg13g2_o21ai_1 _2171_ (.B1(_0157_),
    .Y(_0158_),
    .A1(_1220_),
    .A2(_1224_));
 sg13g2_nand3_1 _2172_ (.B(_0156_),
    .C(_0158_),
    .A(_1241_),
    .Y(_0159_));
 sg13g2_nand3_1 _2173_ (.B(_0155_),
    .C(_0159_),
    .A(_0154_),
    .Y(_0160_));
 sg13g2_nor4_2 _2174_ (.A(_0135_),
    .B(_0136_),
    .C(_0145_),
    .Y(_0161_),
    .D(_0160_));
 sg13g2_nand4_1 _2175_ (.B(net25),
    .C(_0150_),
    .A(net21),
    .Y(_0162_),
    .D(_0152_));
 sg13g2_a22oi_1 _2176_ (.Y(_0163_),
    .B1(_0150_),
    .B2(_0152_),
    .A2(_0830_),
    .A1(_0828_));
 sg13g2_a21o_1 _2177_ (.A2(_0162_),
    .A1(_0140_),
    .B1(_0163_),
    .X(_0164_));
 sg13g2_or2_1 _2178_ (.X(_0165_),
    .B(_0163_),
    .A(net19));
 sg13g2_nor2_1 _2179_ (.A(net72),
    .B(\dac.accu2[6] ),
    .Y(_0166_));
 sg13g2_and3_1 _2180_ (.X(_0167_),
    .A(\dac.accu1[5] ),
    .B(net19),
    .C(_0162_));
 sg13g2_a221oi_1 _2181_ (.B2(_0166_),
    .C1(_0167_),
    .B1(_0165_),
    .A1(_0139_),
    .Y(_0168_),
    .A2(_0164_));
 sg13g2_nand2b_1 _2182_ (.Y(_0169_),
    .B(_0133_),
    .A_N(_0129_));
 sg13g2_a21oi_1 _2183_ (.A1(_1004_),
    .A2(_1009_),
    .Y(_0170_),
    .B1(_0129_));
 sg13g2_nor2_1 _2184_ (.A(\dac.accu2[8] ),
    .B(_0129_),
    .Y(_0171_));
 sg13g2_o21ai_1 _2185_ (.B1(_0120_),
    .Y(_0172_),
    .A1(_0170_),
    .A2(_0171_));
 sg13g2_nand3b_1 _2186_ (.B(net69),
    .C(_0120_),
    .Y(_0173_),
    .A_N(_0129_));
 sg13g2_nand3_1 _2187_ (.B(_1274_),
    .C(_0120_),
    .A(_1198_),
    .Y(_0174_));
 sg13g2_and4_1 _2188_ (.A(_0169_),
    .B(_0172_),
    .C(_0173_),
    .D(_0174_),
    .X(_0175_));
 sg13g2_o21ai_1 _2189_ (.B1(_0175_),
    .Y(_0176_),
    .A1(_0135_),
    .A2(_0168_));
 sg13g2_a21oi_1 _2190_ (.A1(_1273_),
    .A2(_0161_),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_nand2_1 _2191_ (.Y(_0178_),
    .A(\dac.accu2[9] ),
    .B(_1016_));
 sg13g2_or2_1 _2192_ (.X(_0179_),
    .B(_1016_),
    .A(\dac.accu2[9] ));
 sg13g2_nand2_1 _2193_ (.Y(_0180_),
    .A(_1011_),
    .B(_0179_));
 sg13g2_nand2_2 _2194_ (.Y(_0181_),
    .A(_0178_),
    .B(_0180_));
 sg13g2_xnor2_1 _2195_ (.Y(_0182_),
    .A(_1017_),
    .B(\dac.accu2[10] ));
 sg13g2_xnor2_1 _2196_ (.Y(_0183_),
    .A(_1002_),
    .B(_0182_));
 sg13g2_xor2_1 _2197_ (.B(_0183_),
    .A(_0181_),
    .X(_0184_));
 sg13g2_xnor2_1 _2198_ (.Y(_0185_),
    .A(_0177_),
    .B(_0184_));
 sg13g2_nand2_1 _2199_ (.Y(_0186_),
    .A(_0995_),
    .B(net29));
 sg13g2_o21ai_1 _2200_ (.B1(_0186_),
    .Y(_0187_),
    .A1(net30),
    .A2(_0185_));
 sg13g2_nand2_1 _2201_ (.Y(_0188_),
    .A(_1210_),
    .B(_0187_));
 sg13g2_o21ai_1 _2202_ (.B1(_0188_),
    .Y(_0041_),
    .A1(net82),
    .A2(_1209_));
 sg13g2_nor2b_1 _2203_ (.A(_1019_),
    .B_N(_1023_),
    .Y(_0189_));
 sg13g2_nand2b_1 _2204_ (.Y(_0190_),
    .B(_1203_),
    .A_N(_1042_));
 sg13g2_and2_1 _2205_ (.A(_0189_),
    .B(_0190_),
    .X(_0191_));
 sg13g2_xor2_1 _2206_ (.B(net20),
    .A(_0010_),
    .X(_0192_));
 sg13g2_xnor2_1 _2207_ (.Y(_0193_),
    .A(_0191_),
    .B(_0192_));
 sg13g2_nor2_1 _2208_ (.A(\dac.mod2_ctr[1] ),
    .B(\dac.mod2_ctr[0] ),
    .Y(_0194_));
 sg13g2_buf_1 _2209_ (.A(_0194_),
    .X(_0195_));
 sg13g2_nand2_1 _2210_ (.Y(_0196_),
    .A(net70),
    .B(_0157_));
 sg13g2_nand2_2 _2211_ (.Y(_0197_),
    .A(_0156_),
    .B(_0196_));
 sg13g2_nor2_1 _2212_ (.A(_1216_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_xnor2_1 _2213_ (.Y(_0199_),
    .A(net70),
    .B(_1217_));
 sg13g2_xnor2_1 _2214_ (.Y(_0200_),
    .A(_0707_),
    .B(_0199_));
 sg13g2_and2_1 _2215_ (.A(_1235_),
    .B(_0200_),
    .X(_0201_));
 sg13g2_a21o_1 _2216_ (.A2(_1270_),
    .A1(_1235_),
    .B1(_0200_),
    .X(_0202_));
 sg13g2_or2_1 _2217_ (.X(_0203_),
    .B(_1224_),
    .A(_1220_));
 sg13g2_and2_1 _2218_ (.A(_1246_),
    .B(_1265_),
    .X(_0204_));
 sg13g2_nand2_1 _2219_ (.Y(_0205_),
    .A(_1249_),
    .B(_1253_));
 sg13g2_nor2b_1 _2220_ (.A(_0906_),
    .B_N(_1257_),
    .Y(_0206_));
 sg13g2_a21oi_1 _2221_ (.A1(_0205_),
    .A2(_1261_),
    .Y(_0207_),
    .B1(_0206_));
 sg13g2_nand2b_1 _2222_ (.Y(_0208_),
    .B(_0207_),
    .A_N(_0204_));
 sg13g2_nor2_1 _2223_ (.A(_1254_),
    .B(_1235_),
    .Y(_0209_));
 sg13g2_o21ai_1 _2224_ (.B1(_0200_),
    .Y(_0210_),
    .A1(_1222_),
    .A2(_1229_));
 sg13g2_o21ai_1 _2225_ (.B1(_0972_),
    .Y(_0211_),
    .A1(_1220_),
    .A2(_0200_));
 sg13g2_a21oi_1 _2226_ (.A1(_1233_),
    .A2(_0206_),
    .Y(_0212_),
    .B1(_1234_));
 sg13g2_nand2_1 _2227_ (.Y(_0213_),
    .A(_0913_),
    .B(_0205_));
 sg13g2_inv_1 _2228_ (.Y(_0214_),
    .A(_0206_));
 sg13g2_a21oi_1 _2229_ (.A1(_1249_),
    .A2(_1253_),
    .Y(_0215_),
    .B1(_0214_));
 sg13g2_nor2_1 _2230_ (.A(_0912_),
    .B(_1258_),
    .Y(_0216_));
 sg13g2_o21ai_1 _2231_ (.B1(_1234_),
    .Y(_0217_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_o21ai_1 _2232_ (.B1(_0217_),
    .Y(_0218_),
    .A1(_0212_),
    .A2(_0213_));
 sg13g2_a221oi_1 _2233_ (.B2(_0211_),
    .C1(_0218_),
    .B1(_0210_),
    .A1(_0208_),
    .Y(_0219_),
    .A2(_0209_));
 sg13g2_a221oi_1 _2234_ (.B2(_0203_),
    .C1(_0219_),
    .B1(_0202_),
    .A1(_1270_),
    .Y(_0220_),
    .A2(_0201_));
 sg13g2_nand2_1 _2235_ (.Y(_0221_),
    .A(_0150_),
    .B(_0152_));
 sg13g2_nor2_1 _2236_ (.A(_0147_),
    .B(_0148_),
    .Y(_0222_));
 sg13g2_a22oi_1 _2237_ (.Y(_0223_),
    .B1(_0197_),
    .B2(_1216_),
    .A2(_0222_),
    .A1(_0221_));
 sg13g2_nor2_1 _2238_ (.A(_0221_),
    .B(_0222_),
    .Y(_0224_));
 sg13g2_a221oi_1 _2239_ (.B2(_0223_),
    .C1(_0224_),
    .B1(_0220_),
    .A1(_0155_),
    .Y(_0225_),
    .A2(_0198_));
 sg13g2_buf_2 _2240_ (.A(_0225_),
    .X(_0226_));
 sg13g2_nor3_1 _2241_ (.A(_0135_),
    .B(_0145_),
    .C(_0184_),
    .Y(_0227_));
 sg13g2_nand2_1 _2242_ (.Y(_0228_),
    .A(_1284_),
    .B(_0120_));
 sg13g2_nand4_1 _2243_ (.B(net19),
    .C(_0142_),
    .A(_0120_),
    .Y(_0229_),
    .D(_0143_));
 sg13g2_nand4_1 _2244_ (.B(net19),
    .C(_0142_),
    .A(_1284_),
    .Y(_0230_),
    .D(_0143_));
 sg13g2_nand3_1 _2245_ (.B(_0229_),
    .C(_0230_),
    .A(_0228_),
    .Y(_0231_));
 sg13g2_o21ai_1 _2246_ (.B1(_0183_),
    .Y(_0232_),
    .A1(_0133_),
    .A2(_0231_));
 sg13g2_nand2b_1 _2247_ (.Y(_0233_),
    .B(_0179_),
    .A_N(_0183_));
 sg13g2_a22oi_1 _2248_ (.Y(_0234_),
    .B1(_0233_),
    .B2(_1010_),
    .A2(_0183_),
    .A1(_0178_));
 sg13g2_nand2_1 _2249_ (.Y(_0235_),
    .A(_0133_),
    .B(_0231_));
 sg13g2_nor3_1 _2250_ (.A(_0133_),
    .B(_0183_),
    .C(_0231_),
    .Y(_0236_));
 sg13g2_a221oi_1 _2251_ (.B2(_0235_),
    .C1(_0236_),
    .B1(_0234_),
    .A1(_0181_),
    .Y(_0237_),
    .A2(_0232_));
 sg13g2_a21o_1 _2252_ (.A2(_0227_),
    .A1(_0226_),
    .B1(_0237_),
    .X(_0238_));
 sg13g2_nand2b_1 _2253_ (.Y(_0239_),
    .B(_1020_),
    .A_N(\dac.accu2[10] ));
 sg13g2_and2_1 _2254_ (.A(\dac.accu2[10] ),
    .B(_1002_),
    .X(_0240_));
 sg13g2_a21oi_2 _2255_ (.B1(_0240_),
    .Y(_0241_),
    .A2(_0239_),
    .A1(_1018_));
 sg13g2_buf_1 _2256_ (.A(\dac.accu2[11] ),
    .X(_0242_));
 sg13g2_xnor2_1 _2257_ (.Y(_0243_),
    .A(_0995_),
    .B(_0242_));
 sg13g2_xnor2_1 _2258_ (.Y(_0244_),
    .A(net20),
    .B(_0243_));
 sg13g2_xor2_1 _2259_ (.B(_0244_),
    .A(_0241_),
    .X(_0245_));
 sg13g2_xor2_1 _2260_ (.B(_0245_),
    .A(_0238_),
    .X(_0246_));
 sg13g2_buf_1 _2261_ (.A(\dac.accu1[11] ),
    .X(_0247_));
 sg13g2_o21ai_1 _2262_ (.B1(net85),
    .Y(_0248_),
    .A1(net67),
    .A2(net47));
 sg13g2_a21o_1 _2263_ (.A2(_0246_),
    .A1(net47),
    .B1(_0248_),
    .X(_0249_));
 sg13g2_o21ai_1 _2264_ (.B1(_0249_),
    .Y(_0042_),
    .A1(_0533_),
    .A2(_0193_));
 sg13g2_buf_2 _2265_ (.A(\dac.accu2[12] ),
    .X(_0250_));
 sg13g2_xnor2_1 _2266_ (.Y(_0251_),
    .A(_0250_),
    .B(net67));
 sg13g2_xnor2_1 _2267_ (.Y(_0252_),
    .A(_1052_),
    .B(_0251_));
 sg13g2_inv_1 _2268_ (.Y(_0253_),
    .A(_0252_));
 sg13g2_inv_1 _2269_ (.Y(_0254_),
    .A(_0242_));
 sg13g2_o21ai_1 _2270_ (.B1(_0995_),
    .Y(_0255_),
    .A1(_0254_),
    .A2(net20));
 sg13g2_o21ai_1 _2271_ (.B1(_0255_),
    .Y(_0256_),
    .A1(_0242_),
    .A2(_1030_));
 sg13g2_xnor2_1 _2272_ (.Y(_0257_),
    .A(_0253_),
    .B(_0256_));
 sg13g2_nor2b_1 _2273_ (.A(_0241_),
    .B_N(_0244_),
    .Y(_0258_));
 sg13g2_inv_1 _2274_ (.Y(_0259_),
    .A(_0135_));
 sg13g2_a22oi_1 _2275_ (.Y(_0260_),
    .B1(_0165_),
    .B2(_0140_),
    .A2(_0162_),
    .A1(_0139_));
 sg13g2_nand2_1 _2276_ (.Y(_0261_),
    .A(net19),
    .B(_0164_));
 sg13g2_o21ai_1 _2277_ (.B1(_0261_),
    .Y(_0262_),
    .A1(net72),
    .A2(_0260_));
 sg13g2_nand2b_1 _2278_ (.Y(_0263_),
    .B(_1017_),
    .A_N(_0240_));
 sg13g2_nand4_1 _2279_ (.B(_0181_),
    .C(_0239_),
    .A(_0175_),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_a221oi_1 _2280_ (.B2(_0161_),
    .C1(_0264_),
    .B1(_1273_),
    .A1(_0259_),
    .Y(_0265_),
    .A2(_0262_));
 sg13g2_nor2_1 _2281_ (.A(_0258_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_a221oi_1 _2282_ (.B2(_0180_),
    .C1(_0176_),
    .B1(_0178_),
    .A1(_1273_),
    .Y(_0267_),
    .A2(_0161_));
 sg13g2_nor2_1 _2283_ (.A(_0240_),
    .B(_0244_),
    .Y(_0268_));
 sg13g2_nor2_1 _2284_ (.A(_1017_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_and2_1 _2285_ (.A(_0239_),
    .B(_0244_),
    .X(_0270_));
 sg13g2_or2_1 _2286_ (.X(_0271_),
    .B(_0270_),
    .A(_0269_));
 sg13g2_o21ai_1 _2287_ (.B1(_0175_),
    .Y(_0272_),
    .A1(_0269_),
    .A2(_0270_));
 sg13g2_a221oi_1 _2288_ (.B2(_0161_),
    .C1(_0272_),
    .B1(_1273_),
    .A1(_0259_),
    .Y(_0273_),
    .A2(_0262_));
 sg13g2_a221oi_1 _2289_ (.B2(_0181_),
    .C1(_0273_),
    .B1(_0271_),
    .A1(_0244_),
    .Y(_0274_),
    .A2(_0267_));
 sg13g2_nand2_1 _2290_ (.Y(_0275_),
    .A(_0266_),
    .B(_0274_));
 sg13g2_xnor2_1 _2291_ (.Y(_0276_),
    .A(_0257_),
    .B(_0275_));
 sg13g2_nand2_1 _2292_ (.Y(_0277_),
    .A(net5),
    .B(net47));
 sg13g2_buf_2 _2293_ (.A(_0277_),
    .X(_0278_));
 sg13g2_buf_1 _2294_ (.A(_0278_),
    .X(_0279_));
 sg13g2_nand2_1 _2295_ (.Y(_0280_),
    .A(_1046_),
    .B(_1049_));
 sg13g2_xnor2_1 _2296_ (.Y(_0281_),
    .A(_0280_),
    .B(_1053_));
 sg13g2_and2_1 _2297_ (.A(net85),
    .B(\dac.accu1[12] ),
    .X(_0282_));
 sg13g2_a22oi_1 _2298_ (.Y(_0283_),
    .B1(_0282_),
    .B2(_1192_),
    .A2(_0281_),
    .A1(_1186_));
 sg13g2_o21ai_1 _2299_ (.B1(_0283_),
    .Y(_0043_),
    .A1(_0276_),
    .A2(net23));
 sg13g2_a21oi_1 _2300_ (.A1(_1046_),
    .A2(_1049_),
    .Y(_0284_),
    .B1(_1065_));
 sg13g2_a21oi_1 _2301_ (.A1(_0006_),
    .A2(_1064_),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_xnor2_1 _2302_ (.Y(_0286_),
    .A(_1058_),
    .B(_0285_));
 sg13g2_nand2_1 _2303_ (.Y(_0287_),
    .A(net67),
    .B(_1052_));
 sg13g2_nor2_1 _2304_ (.A(net67),
    .B(_1052_),
    .Y(_0288_));
 sg13g2_a21oi_2 _2305_ (.B1(_0288_),
    .Y(_0289_),
    .A2(_0287_),
    .A1(_0250_));
 sg13g2_xor2_1 _2306_ (.B(\dac.accu1[12] ),
    .A(\dac.accu2[13] ),
    .X(_0290_));
 sg13g2_xnor2_1 _2307_ (.Y(_0291_),
    .A(_1057_),
    .B(_0290_));
 sg13g2_inv_1 _2308_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_xnor2_1 _2309_ (.Y(_0293_),
    .A(_0289_),
    .B(_0292_));
 sg13g2_nor2_1 _2310_ (.A(_0245_),
    .B(_0257_),
    .Y(_0294_));
 sg13g2_nand4_1 _2311_ (.B(_0238_),
    .C(_0293_),
    .A(net47),
    .Y(_0295_),
    .D(_0294_));
 sg13g2_nor2_1 _2312_ (.A(_1029_),
    .B(_0241_),
    .Y(_0296_));
 sg13g2_nand2_1 _2313_ (.Y(_0297_),
    .A(_1029_),
    .B(_0241_));
 sg13g2_o21ai_1 _2314_ (.B1(_0297_),
    .Y(_0298_),
    .A1(_0242_),
    .A2(_0296_));
 sg13g2_nand2_1 _2315_ (.Y(_0299_),
    .A(_0252_),
    .B(_0297_));
 sg13g2_nor2_1 _2316_ (.A(_0996_),
    .B(_0242_),
    .Y(_0300_));
 sg13g2_nor3_1 _2317_ (.A(_0996_),
    .B(_0252_),
    .C(_0296_),
    .Y(_0301_));
 sg13g2_a221oi_1 _2318_ (.B2(_0300_),
    .C1(_0301_),
    .B1(_0299_),
    .A1(_0253_),
    .Y(_0302_),
    .A2(_0298_));
 sg13g2_nor2_1 _2319_ (.A(_1191_),
    .B(_0293_),
    .Y(_0303_));
 sg13g2_nand3b_1 _2320_ (.B(_0302_),
    .C(_0303_),
    .Y(_0304_),
    .A_N(_0238_));
 sg13g2_nor2_1 _2321_ (.A(_0293_),
    .B(_0294_),
    .Y(_0305_));
 sg13g2_mux2_1 _2322_ (.A0(_0293_),
    .A1(_0305_),
    .S(_0302_),
    .X(_0306_));
 sg13g2_o21ai_1 _2323_ (.B1(net5),
    .Y(_0307_),
    .A1(_1054_),
    .A2(net47));
 sg13g2_a21oi_1 _2324_ (.A1(_0195_),
    .A2(_0306_),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_nand3_1 _2325_ (.B(_0304_),
    .C(_0308_),
    .A(_0295_),
    .Y(_0309_));
 sg13g2_o21ai_1 _2326_ (.B1(_0309_),
    .Y(_0044_),
    .A1(net82),
    .A2(_0286_));
 sg13g2_xnor2_1 _2327_ (.Y(_0310_),
    .A(_1061_),
    .B(_0596_));
 sg13g2_inv_1 _2328_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_nor2_1 _2329_ (.A(_1059_),
    .B(_0310_),
    .Y(_0312_));
 sg13g2_nand2_1 _2330_ (.Y(_0313_),
    .A(_1067_),
    .B(_0312_));
 sg13g2_o21ai_1 _2331_ (.B1(_0313_),
    .Y(_0314_),
    .A1(_1067_),
    .A2(_0311_));
 sg13g2_nand2_1 _2332_ (.Y(_0315_),
    .A(_1067_),
    .B(_0311_));
 sg13g2_a21oi_1 _2333_ (.A1(_1046_),
    .A2(_1049_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_and4_1 _2334_ (.A(_1046_),
    .B(_1049_),
    .C(_1059_),
    .D(_0310_),
    .X(_0317_));
 sg13g2_nor3_1 _2335_ (.A(_0314_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0318_));
 sg13g2_or2_1 _2336_ (.X(_0319_),
    .B(net20),
    .A(_0254_));
 sg13g2_or2_1 _2337_ (.X(_0320_),
    .B(_1052_),
    .A(net67));
 sg13g2_and2_1 _2338_ (.A(_0254_),
    .B(net20),
    .X(_0321_));
 sg13g2_a221oi_1 _2339_ (.B2(_0291_),
    .C1(_0321_),
    .B1(_0320_),
    .A1(_0995_),
    .Y(_0322_),
    .A2(_0319_));
 sg13g2_nand2b_1 _2340_ (.Y(_0323_),
    .B(_0250_),
    .A_N(_1052_));
 sg13g2_a21oi_1 _2341_ (.A1(_0254_),
    .A2(net20),
    .Y(_0324_),
    .B1(_0323_));
 sg13g2_nand2b_1 _2342_ (.Y(_0325_),
    .B(_0250_),
    .A_N(net67));
 sg13g2_a21oi_1 _2343_ (.A1(_0254_),
    .A2(net20),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_o21ai_1 _2344_ (.B1(_0255_),
    .Y(_0327_),
    .A1(_0324_),
    .A2(_0326_));
 sg13g2_nor2b_1 _2345_ (.A(_0322_),
    .B_N(_0327_),
    .Y(_0328_));
 sg13g2_nor2b_1 _2346_ (.A(net67),
    .B_N(_0250_),
    .Y(_0329_));
 sg13g2_a21oi_1 _2347_ (.A1(net67),
    .A2(_1052_),
    .Y(_0330_),
    .B1(_0291_));
 sg13g2_a221oi_1 _2348_ (.B2(_0250_),
    .C1(_0330_),
    .B1(_0292_),
    .A1(_1064_),
    .Y(_0331_),
    .A2(_0329_));
 sg13g2_nor2b_1 _2349_ (.A(_0257_),
    .B_N(_0293_),
    .Y(_0332_));
 sg13g2_inv_1 _2350_ (.Y(_0333_),
    .A(_0332_));
 sg13g2_nor3_1 _2351_ (.A(_0258_),
    .B(_0265_),
    .C(_0333_),
    .Y(_0334_));
 sg13g2_a22oi_1 _2352_ (.Y(_0335_),
    .B1(_0334_),
    .B2(_0274_),
    .A2(_0331_),
    .A1(_0328_));
 sg13g2_nor2_1 _2353_ (.A(_1186_),
    .B(_1191_),
    .Y(_0336_));
 sg13g2_nand2_1 _2354_ (.Y(_0337_),
    .A(\dac.accu1[12] ),
    .B(_1057_));
 sg13g2_nor2_1 _2355_ (.A(\dac.accu1[12] ),
    .B(_1057_),
    .Y(_0338_));
 sg13g2_a21oi_1 _2356_ (.A1(\dac.accu2[13] ),
    .A2(_0337_),
    .Y(_0339_),
    .B1(_0338_));
 sg13g2_xor2_1 _2357_ (.B(_0596_),
    .A(\dac.accu2[14] ),
    .X(_0340_));
 sg13g2_xor2_1 _2358_ (.B(_0340_),
    .A(_1054_),
    .X(_0341_));
 sg13g2_nand2_1 _2359_ (.Y(_0342_),
    .A(_0339_),
    .B(_0341_));
 sg13g2_inv_1 _2360_ (.Y(_0343_),
    .A(_0339_));
 sg13g2_nand2b_1 _2361_ (.Y(_0344_),
    .B(_0343_),
    .A_N(_0341_));
 sg13g2_and2_1 _2362_ (.A(_0342_),
    .B(_0344_),
    .X(_0345_));
 sg13g2_and2_1 _2363_ (.A(_0336_),
    .B(_0345_),
    .X(_0346_));
 sg13g2_a22oi_1 _2364_ (.Y(_0347_),
    .B1(_0335_),
    .B2(_0346_),
    .A2(_0318_),
    .A1(_1186_));
 sg13g2_or3_1 _2365_ (.A(_0278_),
    .B(_0335_),
    .C(_0345_),
    .X(_0348_));
 sg13g2_nand3_1 _2366_ (.B(_1061_),
    .C(_1192_),
    .A(net85),
    .Y(_0349_));
 sg13g2_nand3_1 _2367_ (.B(_0348_),
    .C(_0349_),
    .A(_0347_),
    .Y(_0045_));
 sg13g2_xnor2_1 _2368_ (.Y(_0350_),
    .A(_0538_),
    .B(_0570_));
 sg13g2_xnor2_1 _2369_ (.Y(_0351_),
    .A(_1070_),
    .B(_0350_));
 sg13g2_nor2_1 _2370_ (.A(_0289_),
    .B(_0291_),
    .Y(_0352_));
 sg13g2_nor2_1 _2371_ (.A(_0352_),
    .B(_0302_),
    .Y(_0353_));
 sg13g2_nand2_1 _2372_ (.Y(_0354_),
    .A(_0332_),
    .B(_0345_));
 sg13g2_nor2_1 _2373_ (.A(_0245_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_nand3_1 _2374_ (.B(_0291_),
    .C(_0344_),
    .A(_0289_),
    .Y(_0356_));
 sg13g2_nand2_1 _2375_ (.Y(_0357_),
    .A(_0342_),
    .B(_0356_));
 sg13g2_a221oi_1 _2376_ (.B2(_0238_),
    .C1(_0357_),
    .B1(_0355_),
    .A1(_0344_),
    .Y(_0358_),
    .A2(_0353_));
 sg13g2_xor2_1 _2377_ (.B(\dac.accu2[15] ),
    .A(_1061_),
    .X(_0359_));
 sg13g2_xnor2_1 _2378_ (.Y(_0360_),
    .A(_0570_),
    .B(_0359_));
 sg13g2_nand2_1 _2379_ (.Y(_0361_),
    .A(\dac.accu2[14] ),
    .B(_0596_));
 sg13g2_nor2_1 _2380_ (.A(\dac.accu2[14] ),
    .B(_0596_),
    .Y(_0362_));
 sg13g2_a21oi_1 _2381_ (.A1(_1054_),
    .A2(_0361_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_xnor2_1 _2382_ (.Y(_0364_),
    .A(_0360_),
    .B(_0363_));
 sg13g2_xnor2_1 _2383_ (.Y(_0365_),
    .A(_0358_),
    .B(_0364_));
 sg13g2_buf_1 _2384_ (.A(_0336_),
    .X(_0366_));
 sg13g2_nor3_1 _2385_ (.A(_1186_),
    .B(_0538_),
    .C(_0195_),
    .Y(_0367_));
 sg13g2_a221oi_1 _2386_ (.B2(net24),
    .C1(_0367_),
    .B1(_0365_),
    .A1(_1186_),
    .Y(_0046_),
    .A2(_0351_));
 sg13g2_nand2_1 _2387_ (.Y(_0368_),
    .A(_0906_),
    .B(_1188_));
 sg13g2_xnor2_1 _2388_ (.Y(_0369_),
    .A(_0912_),
    .B(_1254_));
 sg13g2_xnor2_1 _2389_ (.Y(_0370_),
    .A(_0368_),
    .B(_0369_));
 sg13g2_nor2_1 _2390_ (.A(_1258_),
    .B(_0206_),
    .Y(_0371_));
 sg13g2_xnor2_1 _2391_ (.Y(_0372_),
    .A(_1254_),
    .B(_0371_));
 sg13g2_xnor2_1 _2392_ (.Y(_0373_),
    .A(_0205_),
    .B(_0372_));
 sg13g2_nand2_1 _2393_ (.Y(_0374_),
    .A(_0912_),
    .B(net29));
 sg13g2_o21ai_1 _2394_ (.B1(_0374_),
    .Y(_0375_),
    .A1(net29),
    .A2(_0373_));
 sg13g2_nand2_1 _2395_ (.Y(_0376_),
    .A(net68),
    .B(_0375_));
 sg13g2_o21ai_1 _2396_ (.B1(_0376_),
    .Y(_0047_),
    .A1(net82),
    .A2(_0370_));
 sg13g2_and3_1 _2397_ (.X(_0377_),
    .A(_0911_),
    .B(_0918_),
    .C(_0920_));
 sg13g2_nand2_1 _2398_ (.Y(_0378_),
    .A(_0952_),
    .B(_0969_));
 sg13g2_xnor2_1 _2399_ (.Y(_0379_),
    .A(_0975_),
    .B(_0378_));
 sg13g2_xnor2_1 _2400_ (.Y(_0380_),
    .A(_0377_),
    .B(_0379_));
 sg13g2_a21o_1 _2401_ (.A2(_1267_),
    .A1(_1257_),
    .B1(_1255_),
    .X(_0381_));
 sg13g2_nand2_1 _2402_ (.Y(_0382_),
    .A(_1257_),
    .B(_1255_));
 sg13g2_nand2_1 _2403_ (.Y(_0383_),
    .A(_1259_),
    .B(_0382_));
 sg13g2_a21oi_1 _2404_ (.A1(_0907_),
    .A2(_0381_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_xnor2_1 _2405_ (.Y(_0385_),
    .A(_0204_),
    .B(_0384_));
 sg13g2_nand2_1 _2406_ (.Y(_0386_),
    .A(_0975_),
    .B(_1191_));
 sg13g2_o21ai_1 _2407_ (.B1(_0386_),
    .Y(_0387_),
    .A1(net29),
    .A2(_0385_));
 sg13g2_and2_1 _2408_ (.A(net85),
    .B(_0387_),
    .X(_0388_));
 sg13g2_a21oi_1 _2409_ (.A1(_1186_),
    .A2(_0380_),
    .Y(_0048_),
    .B1(_0388_));
 sg13g2_nand2_1 _2410_ (.Y(_0389_),
    .A(_0378_),
    .B(_0377_));
 sg13g2_o21ai_1 _2411_ (.B1(_0975_),
    .Y(_0390_),
    .A1(_0378_),
    .A2(_0377_));
 sg13g2_nand2_1 _2412_ (.Y(_0391_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_xnor2_1 _2413_ (.Y(_0392_),
    .A(net70),
    .B(_1229_));
 sg13g2_xnor2_1 _2414_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_nand2_1 _2415_ (.Y(_0394_),
    .A(_1236_),
    .B(_1271_));
 sg13g2_xor2_1 _2416_ (.B(_0394_),
    .A(_1270_),
    .X(_0395_));
 sg13g2_nand2_1 _2417_ (.Y(_0396_),
    .A(net70),
    .B(net29));
 sg13g2_o21ai_1 _2418_ (.B1(_0396_),
    .Y(_0397_),
    .A1(net29),
    .A2(_0395_));
 sg13g2_nand2_1 _2419_ (.Y(_0398_),
    .A(net68),
    .B(_0397_));
 sg13g2_o21ai_1 _2420_ (.B1(_0398_),
    .Y(_0049_),
    .A1(net82),
    .A2(_0393_));
 sg13g2_inv_1 _2421_ (.Y(_0399_),
    .A(_1236_));
 sg13g2_o21ai_1 _2422_ (.B1(_1271_),
    .Y(_0400_),
    .A1(_0399_),
    .A2(_1270_));
 sg13g2_nor2_1 _2423_ (.A(_1220_),
    .B(_1224_),
    .Y(_0401_));
 sg13g2_xnor2_1 _2424_ (.Y(_0402_),
    .A(_0401_),
    .B(_0200_));
 sg13g2_xnor2_1 _2425_ (.Y(_0403_),
    .A(_0400_),
    .B(_0402_));
 sg13g2_nand2_1 _2426_ (.Y(_0404_),
    .A(_0709_),
    .B(net30));
 sg13g2_o21ai_1 _2427_ (.B1(_0404_),
    .Y(_0405_),
    .A1(net30),
    .A2(_0403_));
 sg13g2_and2_1 _2428_ (.A(_0708_),
    .B(_0712_),
    .X(_0406_));
 sg13g2_xnor2_1 _2429_ (.Y(_0407_),
    .A(_0979_),
    .B(_0406_));
 sg13g2_nor2_1 _2430_ (.A(net68),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_a21oi_1 _2431_ (.A1(net82),
    .A2(_0405_),
    .Y(_0050_),
    .B1(_0408_));
 sg13g2_xnor2_1 _2432_ (.Y(_0409_),
    .A(_1241_),
    .B(_0197_));
 sg13g2_xnor2_1 _2433_ (.Y(_0410_),
    .A(_0220_),
    .B(_0409_));
 sg13g2_nand2_1 _2434_ (.Y(_0411_),
    .A(_0784_),
    .B(net30));
 sg13g2_o21ai_1 _2435_ (.B1(_0411_),
    .Y(_0412_),
    .A1(net30),
    .A2(_0410_));
 sg13g2_and2_1 _2436_ (.A(_0783_),
    .B(_0788_),
    .X(_0413_));
 sg13g2_inv_1 _2437_ (.Y(_0414_),
    .A(_0979_));
 sg13g2_o21ai_1 _2438_ (.B1(_0711_),
    .Y(_0415_),
    .A1(_0598_),
    .A2(_0979_));
 sg13g2_o21ai_1 _2439_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0709_),
    .A2(_0414_));
 sg13g2_xnor2_1 _2440_ (.Y(_0417_),
    .A(_0413_),
    .B(_0416_));
 sg13g2_nor2_1 _2441_ (.A(net68),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_a21oi_1 _2442_ (.A1(net82),
    .A2(_0412_),
    .Y(_0051_),
    .B1(_0418_));
 sg13g2_nor2_1 _2443_ (.A(_0406_),
    .B(_0413_),
    .Y(_0419_));
 sg13g2_a21oi_1 _2444_ (.A1(_0979_),
    .A2(_0419_),
    .Y(_0420_),
    .B1(_0987_));
 sg13g2_xnor2_1 _2445_ (.Y(_0421_),
    .A(net71),
    .B(_0981_));
 sg13g2_xnor2_1 _2446_ (.Y(_0422_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_nand2_1 _2447_ (.Y(_0423_),
    .A(_0154_),
    .B(_0155_));
 sg13g2_nand2_1 _2448_ (.Y(_0424_),
    .A(_1216_),
    .B(_0197_));
 sg13g2_a21oi_1 _2449_ (.A1(_0220_),
    .A2(_0424_),
    .Y(_0425_),
    .B1(_0198_));
 sg13g2_xnor2_1 _2450_ (.Y(_0426_),
    .A(_0423_),
    .B(_0425_));
 sg13g2_nand2_1 _2451_ (.Y(_0427_),
    .A(net47),
    .B(_0426_));
 sg13g2_o21ai_1 _2452_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0868_),
    .A2(net47));
 sg13g2_mux2_1 _2453_ (.A0(_0422_),
    .A1(_0428_),
    .S(net68),
    .X(_0052_));
 sg13g2_nor2b_1 _2454_ (.A(_0981_),
    .B_N(_0420_),
    .Y(_0429_));
 sg13g2_nand2b_1 _2455_ (.Y(_0430_),
    .B(_0981_),
    .A_N(_0420_));
 sg13g2_o21ai_1 _2456_ (.B1(_0430_),
    .Y(_0431_),
    .A1(net71),
    .A2(_0429_));
 sg13g2_xnor2_1 _2457_ (.Y(_0432_),
    .A(net69),
    .B(_0865_));
 sg13g2_xnor2_1 _2458_ (.Y(_0433_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_xnor2_1 _2459_ (.Y(_0434_),
    .A(net19),
    .B(_0144_));
 sg13g2_xnor2_1 _2460_ (.Y(_0435_),
    .A(_0434_),
    .B(_0226_));
 sg13g2_nand2_1 _2461_ (.Y(_0436_),
    .A(_0990_),
    .B(_1191_));
 sg13g2_o21ai_1 _2462_ (.B1(_0436_),
    .Y(_0437_),
    .A1(net29),
    .A2(_0435_));
 sg13g2_nand2_1 _2463_ (.Y(_0438_),
    .A(net68),
    .B(_0437_));
 sg13g2_o21ai_1 _2464_ (.B1(_0438_),
    .Y(_0053_),
    .A1(net82),
    .A2(_0433_));
 sg13g2_inv_1 _2465_ (.Y(_0439_),
    .A(_0144_));
 sg13g2_nand2_1 _2466_ (.Y(_0440_),
    .A(_0439_),
    .B(_0226_));
 sg13g2_o21ai_1 _2467_ (.B1(net19),
    .Y(_0441_),
    .A1(_0439_),
    .A2(_0226_));
 sg13g2_nand2_1 _2468_ (.Y(_0442_),
    .A(_0440_),
    .B(_0441_));
 sg13g2_nor2_1 _2469_ (.A(_1194_),
    .B(_0121_),
    .Y(_0443_));
 sg13g2_and4_1 _2470_ (.A(net47),
    .B(_0121_),
    .C(_0440_),
    .D(_0441_),
    .X(_0444_));
 sg13g2_a221oi_1 _2471_ (.B2(_0443_),
    .C1(_0444_),
    .B1(_0442_),
    .A1(_1010_),
    .Y(_0445_),
    .A2(net30));
 sg13g2_and2_1 _2472_ (.A(_1012_),
    .B(_1040_),
    .X(_0446_));
 sg13g2_xor2_1 _2473_ (.B(_1203_),
    .A(_0446_),
    .X(_0447_));
 sg13g2_nor2_1 _2474_ (.A(_1210_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_a21oi_1 _2475_ (.A1(net82),
    .A2(_0445_),
    .Y(_0054_),
    .B1(_0448_));
 sg13g2_nand2_1 _2476_ (.Y(_0449_),
    .A(_1198_),
    .B(_1203_));
 sg13g2_o21ai_1 _2477_ (.B1(_1010_),
    .Y(_0450_),
    .A1(_1198_),
    .A2(_1203_));
 sg13g2_nand2_1 _2478_ (.Y(_0451_),
    .A(_0449_),
    .B(_0450_));
 sg13g2_xor2_1 _2479_ (.B(_0451_),
    .A(_1039_),
    .X(_0452_));
 sg13g2_and2_1 _2480_ (.A(_0121_),
    .B(_0434_),
    .X(_0453_));
 sg13g2_a21o_1 _2481_ (.A2(_0453_),
    .A1(_0226_),
    .B1(_0231_),
    .X(_0454_));
 sg13g2_xnor2_1 _2482_ (.Y(_0455_),
    .A(_0134_),
    .B(_0454_));
 sg13g2_nand2_1 _2483_ (.Y(_0456_),
    .A(_1017_),
    .B(_1194_));
 sg13g2_o21ai_1 _2484_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net30),
    .A2(_0455_));
 sg13g2_mux2_1 _2485_ (.A0(_0452_),
    .A1(_0457_),
    .S(net68),
    .X(_0055_));
 sg13g2_buf_1 _2486_ (.A(_0278_),
    .X(_0458_));
 sg13g2_nand2_1 _2487_ (.Y(_0459_),
    .A(\dac.accu2[0] ),
    .B(net22));
 sg13g2_o21ai_1 _2488_ (.B1(_0459_),
    .Y(_0056_),
    .A1(_0907_),
    .A2(net23));
 sg13g2_nand2_1 _2489_ (.Y(_0460_),
    .A(\dac.accu2[10] ),
    .B(_0458_));
 sg13g2_o21ai_1 _2490_ (.B1(_0460_),
    .Y(_0057_),
    .A1(_0996_),
    .A2(net23));
 sg13g2_nand2_1 _2491_ (.Y(_0461_),
    .A(_0247_),
    .B(net24));
 sg13g2_o21ai_1 _2492_ (.B1(_0461_),
    .Y(_0058_),
    .A1(_0254_),
    .A2(net24));
 sg13g2_mux2_1 _2493_ (.A0(_0250_),
    .A1(\dac.accu1[12] ),
    .S(net24),
    .X(_0059_));
 sg13g2_mux2_1 _2494_ (.A0(_1054_),
    .A1(\dac.accu2[13] ),
    .S(_0278_),
    .X(_0060_));
 sg13g2_nand2_1 _2495_ (.Y(_0462_),
    .A(\dac.accu2[14] ),
    .B(net22));
 sg13g2_o21ai_1 _2496_ (.B1(_0462_),
    .Y(_0061_),
    .A1(_1063_),
    .A2(net23));
 sg13g2_and2_1 _2497_ (.A(_0538_),
    .B(_0336_),
    .X(_0463_));
 sg13g2_a21o_1 _2498_ (.A2(_0458_),
    .A1(\dac.accu2[15] ),
    .B1(_0463_),
    .X(_0062_));
 sg13g2_nand2_1 _2499_ (.Y(_0464_),
    .A(_1257_),
    .B(net22));
 sg13g2_o21ai_1 _2500_ (.B1(_0464_),
    .Y(_0063_),
    .A1(_0913_),
    .A2(net23));
 sg13g2_nand2_1 _2501_ (.Y(_0465_),
    .A(_0972_),
    .B(net24));
 sg13g2_o21ai_1 _2502_ (.B1(_0465_),
    .Y(_0064_),
    .A1(_1232_),
    .A2(net24));
 sg13g2_inv_1 _2503_ (.Y(_0466_),
    .A(_0940_));
 sg13g2_nand2_1 _2504_ (.Y(_0467_),
    .A(\dac.accu2[3] ),
    .B(net22));
 sg13g2_o21ai_1 _2505_ (.B1(_0467_),
    .Y(_0065_),
    .A1(_0466_),
    .A2(net23));
 sg13g2_nand2_1 _2506_ (.Y(_0468_),
    .A(_1217_),
    .B(net22));
 sg13g2_o21ai_1 _2507_ (.B1(_0468_),
    .Y(_0066_),
    .A1(_0709_),
    .A2(net23));
 sg13g2_nand2_1 _2508_ (.Y(_0469_),
    .A(\dac.accu2[5] ),
    .B(net22));
 sg13g2_o21ai_1 _2509_ (.B1(_0469_),
    .Y(_0067_),
    .A1(net72),
    .A2(net23));
 sg13g2_nand2_1 _2510_ (.Y(_0470_),
    .A(\dac.accu1[6] ),
    .B(net24));
 sg13g2_o21ai_1 _2511_ (.B1(_0470_),
    .Y(_0068_),
    .A1(_0140_),
    .A2(net24));
 sg13g2_mux2_1 _2512_ (.A0(net69),
    .A1(\dac.accu2[7] ),
    .S(_0278_),
    .X(_0069_));
 sg13g2_nand2_1 _2513_ (.Y(_0471_),
    .A(\dac.accu2[8] ),
    .B(net22));
 sg13g2_o21ai_1 _2514_ (.B1(_0471_),
    .Y(_0070_),
    .A1(_1011_),
    .A2(_0279_));
 sg13g2_nand2_1 _2515_ (.Y(_0472_),
    .A(\dac.accu2[9] ),
    .B(_0278_));
 sg13g2_o21ai_1 _2516_ (.B1(_0472_),
    .Y(_0071_),
    .A1(_1018_),
    .A2(_0279_));
 sg13g2_nand2_1 _2517_ (.Y(_0473_),
    .A(net85),
    .B(\dac.mod2_out[0] ));
 sg13g2_xnor2_1 _2518_ (.Y(_0072_),
    .A(\dac.accu3[0] ),
    .B(_0473_));
 sg13g2_xnor2_1 _2519_ (.Y(_0474_),
    .A(\dac.mod2_out[1] ),
    .B(_0535_));
 sg13g2_nand2_1 _2520_ (.Y(_0475_),
    .A(_0532_),
    .B(_0474_));
 sg13g2_xnor2_1 _2521_ (.Y(_0073_),
    .A(\dac.accu3[1] ),
    .B(_0475_));
 sg13g2_mux2_1 _2522_ (.A0(\dac.mod2_ctr[0] ),
    .A1(_0023_),
    .S(net68),
    .X(_0074_));
 sg13g2_nand2_1 _2523_ (.Y(_0476_),
    .A(net85),
    .B(\dac.mod2_ctr[0] ));
 sg13g2_xnor2_1 _2524_ (.Y(_0075_),
    .A(\dac.mod2_ctr[1] ),
    .B(_0476_));
 sg13g2_nand2_1 _2525_ (.Y(_0477_),
    .A(_0360_),
    .B(_0363_));
 sg13g2_nand2b_1 _2526_ (.Y(_0478_),
    .B(_0362_),
    .A_N(_0360_));
 sg13g2_nand3b_1 _2527_ (.B(_0327_),
    .C(_0331_),
    .Y(_0479_),
    .A_N(_0322_));
 sg13g2_nand2b_1 _2528_ (.Y(_0480_),
    .B(_0339_),
    .A_N(_0479_));
 sg13g2_a21oi_1 _2529_ (.A1(_0479_),
    .A2(_0343_),
    .Y(_0481_),
    .B1(_0340_));
 sg13g2_a21oi_1 _2530_ (.A1(\dac.accu2[14] ),
    .A2(_0596_),
    .Y(_0482_),
    .B1(_0360_));
 sg13g2_o21ai_1 _2531_ (.B1(_1054_),
    .Y(_0483_),
    .A1(_0481_),
    .A2(_0482_));
 sg13g2_nand2_1 _2532_ (.Y(_0484_),
    .A(_0479_),
    .B(_0343_));
 sg13g2_nand3b_1 _2533_ (.B(_0340_),
    .C(_0484_),
    .Y(_0485_),
    .A_N(_1054_));
 sg13g2_nand4_1 _2534_ (.B(_0480_),
    .C(_0483_),
    .A(_0478_),
    .Y(_0486_),
    .D(_0485_));
 sg13g2_nand3_1 _2535_ (.B(_0345_),
    .C(_0477_),
    .A(_0332_),
    .Y(_0487_));
 sg13g2_nor3_1 _2536_ (.A(_0258_),
    .B(_0265_),
    .C(_0487_),
    .Y(_0488_));
 sg13g2_a22oi_1 _2537_ (.Y(_0489_),
    .B1(_0488_),
    .B2(_0274_),
    .A2(_0486_),
    .A1(_0477_));
 sg13g2_a21o_1 _2538_ (.A2(_0570_),
    .A1(\dac.accu2[15] ),
    .B1(_1063_),
    .X(_0490_));
 sg13g2_o21ai_1 _2539_ (.B1(_0490_),
    .Y(_0491_),
    .A1(\dac.accu2[15] ),
    .A2(_0570_));
 sg13g2_xnor2_1 _2540_ (.Y(_0492_),
    .A(_0538_),
    .B(_0491_));
 sg13g2_xnor2_1 _2541_ (.Y(_0493_),
    .A(_0489_),
    .B(_0492_));
 sg13g2_nand2_1 _2542_ (.Y(_0494_),
    .A(\dac.mod2_out[0] ),
    .B(_0278_));
 sg13g2_o21ai_1 _2543_ (.B1(_0494_),
    .Y(_0076_),
    .A1(net22),
    .A2(_0493_));
 sg13g2_nand2_1 _2544_ (.Y(_0495_),
    .A(_0538_),
    .B(_0366_));
 sg13g2_nand2_1 _2545_ (.Y(_0496_),
    .A(_0366_),
    .B(_0491_));
 sg13g2_a21oi_1 _2546_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(_0489_));
 sg13g2_a22oi_1 _2547_ (.Y(_0498_),
    .B1(_0463_),
    .B2(_0491_),
    .A2(_0278_),
    .A1(\dac.mod2_out[1] ));
 sg13g2_nand2b_1 _2548_ (.Y(_0077_),
    .B(_0498_),
    .A_N(_0497_));
 sg13g2_nor2b_1 _2549_ (.A(\sine.ctr_r[15] ),
    .B_N(\sine.ctr_msb_last_r ),
    .Y(_0499_));
 sg13g2_buf_2 _2550_ (.A(_0499_),
    .X(_0500_));
 sg13g2_nand2_1 _2551_ (.Y(_0501_),
    .A(_0656_),
    .B(_0500_));
 sg13g2_o21ai_1 _2552_ (.B1(_0501_),
    .Y(_0078_),
    .A1(net33),
    .A2(_0500_));
 sg13g2_nand2_1 _2553_ (.Y(_0502_),
    .A(net44),
    .B(_0500_));
 sg13g2_xnor2_1 _2554_ (.Y(_0079_),
    .A(net32),
    .B(_0502_));
 sg13g2_xnor2_1 _2555_ (.Y(_0503_),
    .A(net73),
    .B(_0577_));
 sg13g2_nand2_1 _2556_ (.Y(_0504_),
    .A(_0500_),
    .B(_0503_));
 sg13g2_o21ai_1 _2557_ (.B1(_0504_),
    .Y(_0080_),
    .A1(net36),
    .A2(_0500_));
 sg13g2_nand3_1 _2558_ (.B(_0577_),
    .C(_0500_),
    .A(net27),
    .Y(_0505_));
 sg13g2_xnor2_1 _2559_ (.Y(_0081_),
    .A(net42),
    .B(_0505_));
 sg13g2_and3_1 _2560_ (.X(_0506_),
    .A(_0577_),
    .B(_0727_),
    .C(_0500_));
 sg13g2_xnor2_1 _2561_ (.Y(_0082_),
    .A(net35),
    .B(_0506_));
 sg13g2_nand2_1 _2562_ (.Y(_0507_),
    .A(net34),
    .B(_0506_));
 sg13g2_xnor2_1 _2563_ (.Y(_0083_),
    .A(net49),
    .B(_0507_));
 sg13g2_buf_2 _2564_ (.A(ui_in[2]),
    .X(_0508_));
 sg13g2_buf_1 _2565_ (.A(_0508_),
    .X(_0509_));
 sg13g2_nand2_1 _2566_ (.Y(_0510_),
    .A(net66),
    .B(\spi.scan_r[0] ));
 sg13g2_o21ai_1 _2567_ (.B1(_0510_),
    .Y(_0084_),
    .A1(_0916_),
    .A2(_0509_));
 sg13g2_inv_1 _2568_ (.Y(_0511_),
    .A(_1150_));
 sg13g2_nand2_1 _2569_ (.Y(_0512_),
    .A(net66),
    .B(\spi.scan_r[10] ));
 sg13g2_o21ai_1 _2570_ (.B1(_0512_),
    .Y(_0085_),
    .A1(_0511_),
    .A2(net66));
 sg13g2_buf_1 _2571_ (.A(_0508_),
    .X(_0513_));
 sg13g2_mux2_1 _2572_ (.A0(\reg_out_w[11] ),
    .A1(\spi.scan_r[11] ),
    .S(net65),
    .X(_0086_));
 sg13g2_nand2_1 _2573_ (.Y(_0514_),
    .A(net65),
    .B(\spi.scan_r[12] ));
 sg13g2_o21ai_1 _2574_ (.B1(_0514_),
    .Y(_0087_),
    .A1(_1167_),
    .A2(net66));
 sg13g2_nand2_1 _2575_ (.Y(_0515_),
    .A(net65),
    .B(\spi.scan_r[13] ));
 sg13g2_o21ai_1 _2576_ (.B1(_0515_),
    .Y(_0088_),
    .A1(_1176_),
    .A2(net66));
 sg13g2_mux2_1 _2577_ (.A0(_1173_),
    .A1(\spi.scan_r[14] ),
    .S(net65),
    .X(_0089_));
 sg13g2_mux2_1 _2578_ (.A0(\reg_out_w[15] ),
    .A1(\spi.o_spi_dat ),
    .S(net65),
    .X(_0090_));
 sg13g2_mux2_1 _2579_ (.A0(_1074_),
    .A1(\spi.scan_r[1] ),
    .S(net65),
    .X(_0091_));
 sg13g2_mux2_1 _2580_ (.A0(_1079_),
    .A1(\spi.scan_r[2] ),
    .S(net65),
    .X(_0092_));
 sg13g2_mux2_1 _2581_ (.A0(_1085_),
    .A1(\spi.scan_r[3] ),
    .S(_0508_),
    .X(_0093_));
 sg13g2_mux2_1 _2582_ (.A0(\reg_out_w[4] ),
    .A1(\spi.scan_r[4] ),
    .S(_0508_),
    .X(_0094_));
 sg13g2_nand2_1 _2583_ (.Y(_0516_),
    .A(_0513_),
    .B(\spi.scan_r[5] ));
 sg13g2_o21ai_1 _2584_ (.B1(_0516_),
    .Y(_0095_),
    .A1(_1107_),
    .A2(net66));
 sg13g2_nand2_1 _2585_ (.Y(_0517_),
    .A(_0513_),
    .B(\spi.scan_r[6] ));
 sg13g2_o21ai_1 _2586_ (.B1(_0517_),
    .Y(_0096_),
    .A1(_1116_),
    .A2(net66));
 sg13g2_mux2_1 _2587_ (.A0(_1120_),
    .A1(\spi.scan_r[7] ),
    .S(_0508_),
    .X(_0097_));
 sg13g2_inv_1 _2588_ (.Y(_0518_),
    .A(_1122_));
 sg13g2_nand2_1 _2589_ (.Y(_0519_),
    .A(net65),
    .B(\spi.scan_r[8] ));
 sg13g2_o21ai_1 _2590_ (.B1(_0519_),
    .Y(_0098_),
    .A1(_0518_),
    .A2(net66));
 sg13g2_mux2_1 _2591_ (.A0(_1145_),
    .A1(\spi.scan_r[9] ),
    .S(_0508_),
    .X(_0099_));
 sg13g2_inv_1 _2592_ (.Y(_0520_),
    .A(net2));
 sg13g2_nor3_1 _2593_ (.A(_0520_),
    .B(_0508_),
    .C(\spi.last_spi_clk_r ),
    .Y(_0521_));
 sg13g2_buf_2 _2594_ (.A(_0521_),
    .X(_0522_));
 sg13g2_buf_1 _2595_ (.A(_0522_),
    .X(_0523_));
 sg13g2_mux2_1 _2596_ (.A0(\spi.scan_r[0] ),
    .A1(net3),
    .S(net28),
    .X(_0100_));
 sg13g2_mux2_1 _2597_ (.A0(\spi.scan_r[10] ),
    .A1(\spi.scan_r[9] ),
    .S(net28),
    .X(_0101_));
 sg13g2_mux2_1 _2598_ (.A0(\spi.scan_r[11] ),
    .A1(\spi.scan_r[10] ),
    .S(net28),
    .X(_0102_));
 sg13g2_mux2_1 _2599_ (.A0(\spi.scan_r[12] ),
    .A1(\spi.scan_r[11] ),
    .S(net28),
    .X(_0103_));
 sg13g2_mux2_1 _2600_ (.A0(\spi.scan_r[13] ),
    .A1(\spi.scan_r[12] ),
    .S(net28),
    .X(_0104_));
 sg13g2_mux2_1 _2601_ (.A0(\spi.scan_r[14] ),
    .A1(\spi.scan_r[13] ),
    .S(net28),
    .X(_0105_));
 sg13g2_mux2_1 _2602_ (.A0(\spi.o_spi_dat ),
    .A1(\spi.scan_r[14] ),
    .S(net28),
    .X(_0106_));
 sg13g2_mux2_1 _2603_ (.A0(\spi.scan_r[1] ),
    .A1(\spi.scan_r[0] ),
    .S(net28),
    .X(_0107_));
 sg13g2_mux2_1 _2604_ (.A0(\spi.scan_r[2] ),
    .A1(\spi.scan_r[1] ),
    .S(_0523_),
    .X(_0108_));
 sg13g2_mux2_1 _2605_ (.A0(\spi.scan_r[3] ),
    .A1(\spi.scan_r[2] ),
    .S(_0523_),
    .X(_0109_));
 sg13g2_mux2_1 _2606_ (.A0(\spi.scan_r[4] ),
    .A1(\spi.scan_r[3] ),
    .S(_0522_),
    .X(_0110_));
 sg13g2_mux2_1 _2607_ (.A0(\spi.scan_r[5] ),
    .A1(\spi.scan_r[4] ),
    .S(_0522_),
    .X(_0111_));
 sg13g2_mux2_1 _2608_ (.A0(\spi.scan_r[6] ),
    .A1(\spi.scan_r[5] ),
    .S(_0522_),
    .X(_0112_));
 sg13g2_mux2_1 _2609_ (.A0(\spi.scan_r[7] ),
    .A1(\spi.scan_r[6] ),
    .S(_0522_),
    .X(_0113_));
 sg13g2_mux2_1 _2610_ (.A0(\spi.scan_r[8] ),
    .A1(\spi.scan_r[7] ),
    .S(_0522_),
    .X(_0114_));
 sg13g2_mux2_1 _2611_ (.A0(\spi.scan_r[9] ),
    .A1(\spi.scan_r[8] ),
    .S(_0522_),
    .X(_0115_));
 sg13g2_xor2_1 _2612_ (.B(net3),
    .A(_0509_),
    .X(\spi.o_check ));
 sg13g2_nand4_1 _2613_ (.B(_1145_),
    .C(_0511_),
    .A(_0518_),
    .Y(_0524_),
    .D(_1173_));
 sg13g2_nand4_1 _2614_ (.B(_1176_),
    .C(_1167_),
    .A(\reg_out_w[11] ),
    .Y(_0525_),
    .D(\reg_out_w[15] ));
 sg13g2_nand4_1 _2615_ (.B(_0916_),
    .C(_1085_),
    .A(_1074_),
    .Y(_0526_),
    .D(_1113_));
 sg13g2_nand4_1 _2616_ (.B(\reg_out_w[5] ),
    .C(\reg_out_w[4] ),
    .A(_1079_),
    .Y(_0527_),
    .D(_1120_));
 sg13g2_nor4_1 _2617_ (.A(_0524_),
    .B(_0525_),
    .C(_0526_),
    .D(_0527_),
    .Y(\spi.o_det ));
 sg13g2_buf_1 _2618_ (.A(net4),
    .X(_0528_));
 sg13g2_nand2_1 _2619_ (.Y(_0529_),
    .A(_1122_),
    .B(net83));
 sg13g2_o21ai_1 _2620_ (.B1(_0529_),
    .Y(net6),
    .A1(_0916_),
    .A2(_0528_));
 sg13g2_mux2_1 _2621_ (.A0(_1074_),
    .A1(_1145_),
    .S(net83),
    .X(net7));
 sg13g2_mux2_1 _2622_ (.A0(_1079_),
    .A1(_1150_),
    .S(_0528_),
    .X(net8));
 sg13g2_mux2_1 _2623_ (.A0(_1085_),
    .A1(\reg_out_w[11] ),
    .S(net83),
    .X(net9));
 sg13g2_mux2_1 _2624_ (.A0(\reg_out_w[4] ),
    .A1(\reg_out_w[12] ),
    .S(net83),
    .X(net10));
 sg13g2_nand2_1 _2625_ (.Y(_0530_),
    .A(\reg_out_w[13] ),
    .B(net83));
 sg13g2_o21ai_1 _2626_ (.B1(_0530_),
    .Y(net11),
    .A1(_1107_),
    .A2(net83));
 sg13g2_nand2_1 _2627_ (.Y(_0531_),
    .A(_1173_),
    .B(net83));
 sg13g2_o21ai_1 _2628_ (.B1(_0531_),
    .Y(net12),
    .A1(_1116_),
    .A2(net83));
 sg13g2_mux2_1 _2629_ (.A0(_1120_),
    .A1(\reg_out_w[15] ),
    .S(net4),
    .X(net13));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2632__106 (.L_HI(net106));
 sg13g2_buf_1 _2632_ (.A(net106),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2633_ (.A(net107),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2634_ (.A(net108),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2635_ (.A(net109),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2636_ (.A(net110),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2637_ (.A(net111),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2638_ (.A(net112),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2639_ (.A(net113),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2640_ (.A(\spi.o_spi_dat ),
    .X(net14));
 sg13g2_buf_1 _2641_ (.A(\spi.o_det ),
    .X(net15));
 sg13g2_buf_1 _2642_ (.A(\spi.o_check ),
    .X(net16));
 sg13g2_buf_1 _2643_ (.A(net103),
    .X(uo_out[3]));
 sg13g2_buf_1 _2644_ (.A(net104),
    .X(uo_out[4]));
 sg13g2_buf_1 _2645_ (.A(net105),
    .X(uo_out[5]));
 sg13g2_buf_1 _2646_ (.A(\dac.o_ds_n ),
    .X(net17));
 sg13g2_buf_1 _2647_ (.A(\dac.o_ds ),
    .X(net18));
 sg13g2_dfrbp_1 \dac.accu1[0]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net95),
    .D(_0040_),
    .Q_N(_1338_),
    .Q(\dac.accu1[0] ));
 sg13g2_dfrbp_1 \dac.accu1[10]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0041_),
    .Q_N(_1337_),
    .Q(\dac.accu1[10] ));
 sg13g2_dfrbp_1 \dac.accu1[11]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net99),
    .D(_0042_),
    .Q_N(_0010_),
    .Q(\dac.accu1[11] ));
 sg13g2_dfrbp_1 \dac.accu1[12]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0043_),
    .Q_N(_0006_),
    .Q(\dac.accu1[12] ));
 sg13g2_dfrbp_1 \dac.accu1[13]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net99),
    .D(_0044_),
    .Q_N(_1336_),
    .Q(\dac.accu1[13] ));
 sg13g2_dfrbp_1 \dac.accu1[14]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net97),
    .D(_0045_),
    .Q_N(_1335_),
    .Q(\dac.accu1[14] ));
 sg13g2_dfrbp_1 \dac.accu1[15]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0046_),
    .Q_N(_1334_),
    .Q(\dac.accu1[15] ));
 sg13g2_dfrbp_1 \dac.accu1[1]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0047_),
    .Q_N(_1333_),
    .Q(\dac.accu1[1] ));
 sg13g2_dfrbp_1 \dac.accu1[2]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net95),
    .D(_0048_),
    .Q_N(_1332_),
    .Q(\dac.accu1[2] ));
 sg13g2_dfrbp_1 \dac.accu1[3]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0049_),
    .Q_N(_1331_),
    .Q(\dac.accu1[3] ));
 sg13g2_dfrbp_1 \dac.accu1[4]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0050_),
    .Q_N(_1330_),
    .Q(\dac.accu1[4] ));
 sg13g2_dfrbp_1 \dac.accu1[5]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net96),
    .D(_0051_),
    .Q_N(_1329_),
    .Q(\dac.accu1[5] ));
 sg13g2_dfrbp_1 \dac.accu1[6]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net96),
    .D(_0052_),
    .Q_N(_1328_),
    .Q(\dac.accu1[6] ));
 sg13g2_dfrbp_1 \dac.accu1[7]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net96),
    .D(_0053_),
    .Q_N(_1327_),
    .Q(\dac.accu1[7] ));
 sg13g2_dfrbp_1 \dac.accu1[8]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net96),
    .D(_0054_),
    .Q_N(_1326_),
    .Q(\dac.accu1[8] ));
 sg13g2_dfrbp_1 \dac.accu1[9]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0055_),
    .Q_N(_1325_),
    .Q(\dac.accu1[9] ));
 sg13g2_dfrbp_1 \dac.accu2[0]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net86),
    .D(_0056_),
    .Q_N(_1324_),
    .Q(\dac.accu2[0] ));
 sg13g2_dfrbp_1 \dac.accu2[10]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net99),
    .D(_0057_),
    .Q_N(_1323_),
    .Q(\dac.accu2[10] ));
 sg13g2_dfrbp_1 \dac.accu2[11]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0058_),
    .Q_N(_1322_),
    .Q(\dac.accu2[11] ));
 sg13g2_dfrbp_1 \dac.accu2[12]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0059_),
    .Q_N(_1321_),
    .Q(\dac.accu2[12] ));
 sg13g2_dfrbp_1 \dac.accu2[13]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0060_),
    .Q_N(_1320_),
    .Q(\dac.accu2[13] ));
 sg13g2_dfrbp_1 \dac.accu2[14]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0061_),
    .Q_N(_1319_),
    .Q(\dac.accu2[14] ));
 sg13g2_dfrbp_1 \dac.accu2[15]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0062_),
    .Q_N(_1318_),
    .Q(\dac.accu2[15] ));
 sg13g2_dfrbp_1 \dac.accu2[1]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net94),
    .D(_0063_),
    .Q_N(_1317_),
    .Q(\dac.accu2[1] ));
 sg13g2_dfrbp_1 \dac.accu2[2]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net95),
    .D(_0064_),
    .Q_N(_1316_),
    .Q(\dac.accu2[2] ));
 sg13g2_dfrbp_1 \dac.accu2[3]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0065_),
    .Q_N(_1315_),
    .Q(\dac.accu2[3] ));
 sg13g2_dfrbp_1 \dac.accu2[4]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net95),
    .D(_0066_),
    .Q_N(_1314_),
    .Q(\dac.accu2[4] ));
 sg13g2_dfrbp_1 \dac.accu2[5]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net102),
    .D(_0067_),
    .Q_N(_1313_),
    .Q(\dac.accu2[5] ));
 sg13g2_dfrbp_1 \dac.accu2[6]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net96),
    .D(_0068_),
    .Q_N(_1312_),
    .Q(\dac.accu2[6] ));
 sg13g2_dfrbp_1 \dac.accu2[7]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0069_),
    .Q_N(_1311_),
    .Q(\dac.accu2[7] ));
 sg13g2_dfrbp_1 \dac.accu2[8]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(_0070_),
    .Q_N(_1310_),
    .Q(\dac.accu2[8] ));
 sg13g2_dfrbp_1 \dac.accu2[9]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(_0071_),
    .Q_N(_1309_),
    .Q(\dac.accu2[9] ));
 sg13g2_dfrbp_1 \dac.accu3[0]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0072_),
    .Q_N(_1308_),
    .Q(\dac.accu3[0] ));
 sg13g2_dfrbp_1 \dac.accu3[1]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net100),
    .D(_0073_),
    .Q_N(_1307_),
    .Q(\dac.accu3[1] ));
 sg13g2_dfrbp_1 \dac.mod2_ctr[0]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0074_),
    .Q_N(_0023_),
    .Q(\dac.mod2_ctr[0] ));
 sg13g2_dfrbp_1 \dac.mod2_ctr[1]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net97),
    .D(_0075_),
    .Q_N(_1306_),
    .Q(\dac.mod2_ctr[1] ));
 sg13g2_dfrbp_1 \dac.mod2_out[0]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net100),
    .D(_0076_),
    .Q_N(_1305_),
    .Q(\dac.mod2_out[0] ));
 sg13g2_dfrbp_1 \dac.mod2_out[1]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net98),
    .D(_0077_),
    .Q_N(_1339_),
    .Q(\dac.mod2_out[1] ));
 sg13g2_dfrbp_1 \dac.o_ds$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net92),
    .D(_0000_),
    .Q_N(\dac.o_ds_n ),
    .Q(\dac.o_ds ));
 sg13g2_dfrbp_1 \sine.ctr_msb_last_r$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net86),
    .D(\sine.ctr_r[15] ),
    .Q_N(_1340_),
    .Q(\sine.ctr_msb_last_r ));
 sg13g2_dfrbp_1 \sine.ctr_r[0]$_DFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net98),
    .D(_0024_),
    .Q_N(_1341_),
    .Q(\sine.ctr_r[0] ));
 sg13g2_dfrbp_1 \sine.ctr_r[10]$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0025_),
    .Q_N(_1342_),
    .Q(\sine.ctr_r[10] ));
 sg13g2_dfrbp_1 \sine.ctr_r[11]$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0026_),
    .Q_N(_1343_),
    .Q(\sine.ctr_r[11] ));
 sg13g2_dfrbp_1 \sine.ctr_r[12]$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0027_),
    .Q_N(_1344_),
    .Q(\sine.ctr_r[12] ));
 sg13g2_dfrbp_1 \sine.ctr_r[13]$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0028_),
    .Q_N(_1345_),
    .Q(\sine.ctr_r[13] ));
 sg13g2_dfrbp_1 \sine.ctr_r[14]$_DFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net87),
    .D(_0029_),
    .Q_N(_1346_),
    .Q(\sine.ctr_r[14] ));
 sg13g2_dfrbp_1 \sine.ctr_r[15]$_DFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0030_),
    .Q_N(_1347_),
    .Q(\sine.ctr_r[15] ));
 sg13g2_dfrbp_1 \sine.ctr_r[1]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net93),
    .D(_0031_),
    .Q_N(_1348_),
    .Q(\sine.ctr_r[1] ));
 sg13g2_dfrbp_1 \sine.ctr_r[2]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net92),
    .D(_0032_),
    .Q_N(_1349_),
    .Q(\sine.ctr_r[2] ));
 sg13g2_dfrbp_1 \sine.ctr_r[3]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net92),
    .D(_0033_),
    .Q_N(_1350_),
    .Q(\sine.ctr_r[3] ));
 sg13g2_dfrbp_1 \sine.ctr_r[4]$_DFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0034_),
    .Q_N(_1351_),
    .Q(\sine.ctr_r[4] ));
 sg13g2_dfrbp_1 \sine.ctr_r[5]$_DFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0035_),
    .Q_N(_1352_),
    .Q(\sine.ctr_r[5] ));
 sg13g2_dfrbp_1 \sine.ctr_r[6]$_DFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0036_),
    .Q_N(_1353_),
    .Q(\sine.ctr_r[6] ));
 sg13g2_dfrbp_1 \sine.ctr_r[7]$_DFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net89),
    .D(_0037_),
    .Q_N(_1354_),
    .Q(\sine.ctr_r[7] ));
 sg13g2_dfrbp_1 \sine.ctr_r[8]$_DFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net87),
    .D(_0038_),
    .Q_N(_1355_),
    .Q(\sine.ctr_r[8] ));
 sg13g2_dfrbp_1 \sine.ctr_r[9]$_DFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(_0039_),
    .Q_N(_1304_),
    .Q(\sine.ctr_r[9] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[0]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0078_),
    .Q_N(_0022_),
    .Q(\sine.read_ptr_r[0] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[1]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0079_),
    .Q_N(_0009_),
    .Q(\sine.read_ptr_r[1] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[2]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0080_),
    .Q_N(_0008_),
    .Q(\sine.read_ptr_r[2] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[3]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0081_),
    .Q_N(_0004_),
    .Q(\sine.read_ptr_r[3] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[4]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0082_),
    .Q_N(_0002_),
    .Q(\sine.read_ptr_r[4] ));
 sg13g2_dfrbp_1 \sine.read_ptr_r[5]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0083_),
    .Q_N(_1303_),
    .Q(\sine.read_ptr_r[5] ));
 sg13g2_dfrbp_1 \spi.data_r[0]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net98),
    .D(_0084_),
    .Q_N(_1302_),
    .Q(\reg_out_w[0] ));
 sg13g2_dfrbp_1 \spi.data_r[10]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net90),
    .D(_0085_),
    .Q_N(_0012_),
    .Q(\reg_out_w[10] ));
 sg13g2_dfrbp_1 \spi.data_r[11]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net90),
    .D(_0086_),
    .Q_N(_0011_),
    .Q(\reg_out_w[11] ));
 sg13g2_dfrbp_1 \spi.data_r[12]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net90),
    .D(_0087_),
    .Q_N(_0007_),
    .Q(\reg_out_w[12] ));
 sg13g2_dfrbp_1 \spi.data_r[13]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0088_),
    .Q_N(_0005_),
    .Q(\reg_out_w[13] ));
 sg13g2_dfrbp_1 \spi.data_r[14]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net94),
    .D(_0089_),
    .Q_N(_0003_),
    .Q(\reg_out_w[14] ));
 sg13g2_dfrbp_1 \spi.data_r[15]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0090_),
    .Q_N(_0001_),
    .Q(\reg_out_w[15] ));
 sg13g2_dfrbp_1 \spi.data_r[1]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net90),
    .D(_0091_),
    .Q_N(_0021_),
    .Q(\reg_out_w[1] ));
 sg13g2_dfrbp_1 \spi.data_r[2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net91),
    .D(_0092_),
    .Q_N(_0020_),
    .Q(\reg_out_w[2] ));
 sg13g2_dfrbp_1 \spi.data_r[3]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0093_),
    .Q_N(_0019_),
    .Q(\reg_out_w[3] ));
 sg13g2_dfrbp_1 \spi.data_r[4]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net93),
    .D(_0094_),
    .Q_N(_0018_),
    .Q(\reg_out_w[4] ));
 sg13g2_dfrbp_1 \spi.data_r[5]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net92),
    .D(_0095_),
    .Q_N(_0017_),
    .Q(\reg_out_w[5] ));
 sg13g2_dfrbp_1 \spi.data_r[6]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net92),
    .D(_0096_),
    .Q_N(_0016_),
    .Q(\reg_out_w[6] ));
 sg13g2_dfrbp_1 \spi.data_r[7]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net98),
    .D(_0097_),
    .Q_N(_0015_),
    .Q(\reg_out_w[7] ));
 sg13g2_dfrbp_1 \spi.data_r[8]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net90),
    .D(_0098_),
    .Q_N(_0014_),
    .Q(\reg_out_w[8] ));
 sg13g2_dfrbp_1 \spi.data_r[9]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net91),
    .D(_0099_),
    .Q_N(_0013_),
    .Q(\reg_out_w[9] ));
 sg13g2_dfrbp_1 \spi.last_spi_clk_r$_DFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(net2),
    .Q_N(_1301_),
    .Q(\spi.last_spi_clk_r ));
 sg13g2_dfrbp_1 \spi.scan_r[0]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0100_),
    .Q_N(_1300_),
    .Q(\spi.scan_r[0] ));
 sg13g2_dfrbp_1 \spi.scan_r[10]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net87),
    .D(_0101_),
    .Q_N(_1299_),
    .Q(\spi.scan_r[10] ));
 sg13g2_dfrbp_1 \spi.scan_r[11]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net88),
    .D(_0102_),
    .Q_N(_1298_),
    .Q(\spi.scan_r[11] ));
 sg13g2_dfrbp_1 \spi.scan_r[12]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net88),
    .D(_0103_),
    .Q_N(_1297_),
    .Q(\spi.scan_r[12] ));
 sg13g2_dfrbp_1 \spi.scan_r[13]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net88),
    .D(_0104_),
    .Q_N(_1296_),
    .Q(\spi.scan_r[13] ));
 sg13g2_dfrbp_1 \spi.scan_r[14]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net88),
    .D(_0105_),
    .Q_N(_1295_),
    .Q(\spi.scan_r[14] ));
 sg13g2_dfrbp_1 \spi.scan_r[15]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0106_),
    .Q_N(_1294_),
    .Q(\spi.o_spi_dat ));
 sg13g2_dfrbp_1 \spi.scan_r[1]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net97),
    .D(_0107_),
    .Q_N(_1293_),
    .Q(\spi.scan_r[1] ));
 sg13g2_dfrbp_1 \spi.scan_r[2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net91),
    .D(_0108_),
    .Q_N(_1292_),
    .Q(\spi.scan_r[2] ));
 sg13g2_dfrbp_1 \spi.scan_r[3]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net91),
    .D(_0109_),
    .Q_N(_1291_),
    .Q(\spi.scan_r[3] ));
 sg13g2_dfrbp_1 \spi.scan_r[4]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net92),
    .D(_0110_),
    .Q_N(_1290_),
    .Q(\spi.scan_r[4] ));
 sg13g2_dfrbp_1 \spi.scan_r[5]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net92),
    .D(_0111_),
    .Q_N(_1289_),
    .Q(\spi.scan_r[5] ));
 sg13g2_dfrbp_1 \spi.scan_r[6]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(_0112_),
    .Q_N(_1288_),
    .Q(\spi.scan_r[6] ));
 sg13g2_dfrbp_1 \spi.scan_r[7]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net92),
    .D(_0113_),
    .Q_N(_1287_),
    .Q(\spi.scan_r[7] ));
 sg13g2_dfrbp_1 \spi.scan_r[8]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net94),
    .D(_0114_),
    .Q_N(_1286_),
    .Q(\spi.scan_r[8] ));
 sg13g2_dfrbp_1 \spi.scan_r[9]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net88),
    .D(_0115_),
    .Q_N(_1285_),
    .Q(\spi.scan_r[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_0139_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1029_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0828_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0458_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0279_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0366_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0830_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0625_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0553_),
    .X(net27));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(_0523_));
 sg13g2_buf_2 fanout29 (.A(_1194_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1192_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0756_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0680_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0654_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0639_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0621_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0619_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0611_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0601_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0587_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0575_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0560_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0556_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0552_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0549_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0546_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0543_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0195_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0781_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0671_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0651_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0628_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0613_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0609_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0606_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0605_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0586_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0582_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0581_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0559_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0555_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0551_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0548_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0545_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0542_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0513_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0509_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0247_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1210_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0990_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0940_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0868_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0784_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0684_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0578_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0566_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0565_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0563_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0558_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0554_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0547_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0544_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0533_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0528_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0540_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0532_),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net94));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(net89));
 sg13g2_buf_2 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net94));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net93));
 sg13g2_buf_2 fanout91 (.A(net93),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net93));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net1),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(net102));
 sg13g2_buf_2 fanout96 (.A(net102),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net101));
 sg13g2_buf_2 fanout98 (.A(net101),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net101));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(net1),
    .X(net102));
 sg13g2_tielo _2643__103 (.L_LO(net103));
 sg13g2_tielo _2644__104 (.L_LO(net104));
 sg13g2_tielo _2645__105 (.L_LO(net105));
 sg13g2_tiehi _2633__107 (.L_HI(net107));
 sg13g2_tiehi _2634__108 (.L_HI(net108));
 sg13g2_tiehi _2635__109 (.L_HI(net109));
 sg13g2_tiehi _2636__110 (.L_HI(net110));
 sg13g2_tiehi _2637__111 (.L_HI(net111));
 sg13g2_tiehi _2638__112 (.L_HI(net112));
 sg13g2_tiehi _2639__113 (.L_HI(net113));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_4 FILLER_0_259 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_fill_2 FILLER_1_86 ();
 sg13g2_fill_1 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_128 ();
 sg13g2_decap_8 FILLER_1_135 ();
 sg13g2_decap_8 FILLER_1_142 ();
 sg13g2_fill_2 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_decap_8 FILLER_1_167 ();
 sg13g2_decap_8 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_181 ();
 sg13g2_decap_8 FILLER_1_188 ();
 sg13g2_decap_8 FILLER_1_195 ();
 sg13g2_decap_8 FILLER_1_202 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_252 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_275 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_299 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_decap_8 FILLER_1_313 ();
 sg13g2_decap_8 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_341 ();
 sg13g2_decap_8 FILLER_1_348 ();
 sg13g2_decap_8 FILLER_1_355 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_8 FILLER_1_404 ();
 sg13g2_decap_8 FILLER_1_411 ();
 sg13g2_decap_8 FILLER_1_418 ();
 sg13g2_decap_4 FILLER_1_425 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_25 ();
 sg13g2_fill_2 FILLER_2_65 ();
 sg13g2_fill_1 FILLER_2_67 ();
 sg13g2_decap_4 FILLER_2_94 ();
 sg13g2_decap_4 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_4 FILLER_2_140 ();
 sg13g2_fill_2 FILLER_2_144 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_decap_8 FILLER_2_173 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_fill_2 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_2 FILLER_2_244 ();
 sg13g2_fill_1 FILLER_2_246 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_fill_1 FILLER_2_271 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_330 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_24 ();
 sg13g2_decap_8 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_38 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_fill_1 FILLER_3_56 ();
 sg13g2_decap_4 FILLER_3_62 ();
 sg13g2_fill_1 FILLER_3_66 ();
 sg13g2_fill_2 FILLER_3_72 ();
 sg13g2_fill_1 FILLER_3_79 ();
 sg13g2_fill_2 FILLER_3_89 ();
 sg13g2_fill_1 FILLER_3_102 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_118 ();
 sg13g2_decap_4 FILLER_3_129 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_144 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_2 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_171 ();
 sg13g2_decap_8 FILLER_3_178 ();
 sg13g2_decap_8 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_192 ();
 sg13g2_decap_8 FILLER_3_199 ();
 sg13g2_decap_4 FILLER_3_206 ();
 sg13g2_fill_2 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_271 ();
 sg13g2_fill_1 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_303 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_4 FILLER_3_317 ();
 sg13g2_decap_4 FILLER_3_329 ();
 sg13g2_fill_2 FILLER_3_333 ();
 sg13g2_fill_2 FILLER_3_353 ();
 sg13g2_fill_1 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_19 ();
 sg13g2_fill_1 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_27 ();
 sg13g2_fill_1 FILLER_4_34 ();
 sg13g2_fill_1 FILLER_4_43 ();
 sg13g2_decap_4 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_61 ();
 sg13g2_decap_4 FILLER_4_90 ();
 sg13g2_fill_1 FILLER_4_99 ();
 sg13g2_fill_2 FILLER_4_104 ();
 sg13g2_decap_4 FILLER_4_111 ();
 sg13g2_fill_2 FILLER_4_135 ();
 sg13g2_fill_2 FILLER_4_142 ();
 sg13g2_fill_1 FILLER_4_149 ();
 sg13g2_fill_2 FILLER_4_155 ();
 sg13g2_fill_1 FILLER_4_157 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_4 FILLER_4_196 ();
 sg13g2_fill_2 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_fill_2 FILLER_4_247 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_fill_1 FILLER_4_291 ();
 sg13g2_decap_4 FILLER_4_300 ();
 sg13g2_decap_4 FILLER_4_313 ();
 sg13g2_decap_4 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_fill_1 FILLER_4_360 ();
 sg13g2_fill_2 FILLER_4_366 ();
 sg13g2_fill_2 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_2 FILLER_5_36 ();
 sg13g2_fill_2 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_92 ();
 sg13g2_decap_4 FILLER_5_99 ();
 sg13g2_fill_1 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_132 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_169 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_198 ();
 sg13g2_fill_2 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_4 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_fill_1 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_290 ();
 sg13g2_decap_4 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_fill_2 FILLER_5_366 ();
 sg13g2_decap_4 FILLER_5_376 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_16 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_1 FILLER_6_37 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_fill_2 FILLER_6_58 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_fill_2 FILLER_6_66 ();
 sg13g2_fill_1 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_92 ();
 sg13g2_fill_2 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_106 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_fill_2 FILLER_6_132 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_2 FILLER_6_148 ();
 sg13g2_fill_1 FILLER_6_150 ();
 sg13g2_fill_2 FILLER_6_156 ();
 sg13g2_decap_4 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_167 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_fill_2 FILLER_6_187 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_195 ();
 sg13g2_decap_8 FILLER_6_202 ();
 sg13g2_decap_8 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_fill_2 FILLER_6_262 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_4 FILLER_6_374 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_16 ();
 sg13g2_fill_1 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_50 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_decap_4 FILLER_7_82 ();
 sg13g2_fill_1 FILLER_7_105 ();
 sg13g2_fill_2 FILLER_7_111 ();
 sg13g2_fill_1 FILLER_7_117 ();
 sg13g2_fill_1 FILLER_7_123 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_decap_4 FILLER_7_158 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_decap_4 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_298 ();
 sg13g2_decap_4 FILLER_7_303 ();
 sg13g2_fill_2 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_344 ();
 sg13g2_fill_1 FILLER_7_346 ();
 sg13g2_decap_4 FILLER_7_354 ();
 sg13g2_decap_4 FILLER_7_374 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_decap_4 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_11 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_23 ();
 sg13g2_fill_1 FILLER_8_34 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_decap_4 FILLER_8_57 ();
 sg13g2_fill_1 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_93 ();
 sg13g2_fill_2 FILLER_8_100 ();
 sg13g2_fill_2 FILLER_8_108 ();
 sg13g2_fill_1 FILLER_8_110 ();
 sg13g2_fill_2 FILLER_8_128 ();
 sg13g2_fill_1 FILLER_8_130 ();
 sg13g2_decap_4 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_fill_1 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_4 FILLER_8_280 ();
 sg13g2_fill_2 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_decap_4 FILLER_8_331 ();
 sg13g2_fill_2 FILLER_8_335 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_2 FILLER_8_356 ();
 sg13g2_fill_1 FILLER_8_366 ();
 sg13g2_fill_2 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_2 FILLER_9_61 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_fill_2 FILLER_9_106 ();
 sg13g2_decap_4 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_160 ();
 sg13g2_fill_1 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_decap_4 FILLER_9_176 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_decap_4 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_4 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_fill_2 FILLER_9_279 ();
 sg13g2_fill_2 FILLER_9_292 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_4 FILLER_9_335 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_20 ();
 sg13g2_fill_1 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_45 ();
 sg13g2_decap_4 FILLER_10_51 ();
 sg13g2_decap_4 FILLER_10_62 ();
 sg13g2_fill_2 FILLER_10_66 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_99 ();
 sg13g2_fill_1 FILLER_10_111 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_2 FILLER_10_138 ();
 sg13g2_decap_4 FILLER_10_174 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_fill_1 FILLER_10_246 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_296 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_343 ();
 sg13g2_decap_4 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_decap_4 FILLER_10_396 ();
 sg13g2_fill_2 FILLER_10_400 ();
 sg13g2_decap_4 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_decap_4 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_64 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_decap_8 FILLER_11_97 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_116 ();
 sg13g2_decap_4 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_4 FILLER_11_177 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_fill_2 FILLER_11_219 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_4 FILLER_11_248 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_decap_4 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_decap_4 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_decap_4 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_fill_2 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_425 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_33 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_decap_4 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_decap_4 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_153 ();
 sg13g2_fill_1 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_4 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_decap_8 FILLER_12_232 ();
 sg13g2_decap_8 FILLER_12_239 ();
 sg13g2_decap_4 FILLER_12_246 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_decap_4 FILLER_12_288 ();
 sg13g2_decap_4 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_4 FILLER_12_366 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_1 FILLER_12_384 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_4 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_72 ();
 sg13g2_decap_4 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_decap_4 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_decap_8 FILLER_13_156 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_decap_8 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_177 ();
 sg13g2_decap_4 FILLER_13_184 ();
 sg13g2_fill_2 FILLER_13_202 ();
 sg13g2_decap_4 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_240 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_decap_4 FILLER_13_290 ();
 sg13g2_decap_4 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_334 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_344 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_fill_2 FILLER_13_375 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_1 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_9 ();
 sg13g2_fill_2 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_60 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_decap_4 FILLER_14_130 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_decap_4 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_4 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_4 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_4 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_decap_4 FILLER_14_283 ();
 sg13g2_decap_4 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_fill_2 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_34 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_fill_2 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_decap_4 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_159 ();
 sg13g2_decap_8 FILLER_15_166 ();
 sg13g2_decap_8 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_218 ();
 sg13g2_decap_4 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_317 ();
 sg13g2_decap_4 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_fill_1 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_15_409 ();
 sg13g2_decap_8 FILLER_15_416 ();
 sg13g2_decap_8 FILLER_15_423 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_decap_4 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_265 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_370 ();
 sg13g2_decap_4 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_34 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_fill_2 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_59 ();
 sg13g2_decap_8 FILLER_17_66 ();
 sg13g2_decap_4 FILLER_17_73 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_2 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_125 ();
 sg13g2_decap_8 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_fill_1 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_2 FILLER_17_396 ();
 sg13g2_fill_2 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_62 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_decap_8 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_121 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_decap_4 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_decap_4 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_389 ();
 sg13g2_fill_2 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_31 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_decap_8 FILLER_19_45 ();
 sg13g2_decap_4 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_61 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_decap_8 FILLER_19_75 ();
 sg13g2_decap_8 FILLER_19_82 ();
 sg13g2_decap_8 FILLER_19_89 ();
 sg13g2_decap_8 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_103 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_decap_4 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_271 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_decap_4 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_4 FILLER_19_366 ();
 sg13g2_fill_2 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_387 ();
 sg13g2_fill_2 FILLER_19_397 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_31 ();
 sg13g2_decap_4 FILLER_20_38 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_54 ();
 sg13g2_decap_8 FILLER_20_61 ();
 sg13g2_decap_4 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_111 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_4 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_4 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_4 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_fill_2 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_36 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_decap_8 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_85 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_4 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_193 ();
 sg13g2_decap_4 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_decap_4 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_fill_2 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_57 ();
 sg13g2_decap_8 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_8 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_4 FILLER_22_258 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_decap_4 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_4 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_decap_4 FILLER_22_374 ();
 sg13g2_fill_1 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_decap_8 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_4 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_decap_4 FILLER_23_213 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_decap_4 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_4 FILLER_23_378 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_4 FILLER_23_395 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_39 ();
 sg13g2_fill_2 FILLER_24_55 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_decap_8 FILLER_24_65 ();
 sg13g2_decap_4 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_decap_8 FILLER_24_80 ();
 sg13g2_decap_4 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_8 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_4 FILLER_24_381 ();
 sg13g2_fill_1 FILLER_24_385 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_219 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_decap_4 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_fill_1 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_75 ();
 sg13g2_decap_8 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_4 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_decap_4 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_4 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_356 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_373 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_29 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_111 ();
 sg13g2_decap_4 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_decap_4 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_4 FILLER_27_368 ();
 sg13g2_fill_2 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_fill_2 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_28_34 ();
 sg13g2_decap_8 FILLER_28_44 ();
 sg13g2_decap_4 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_90 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_decap_4 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_198 ();
 sg13g2_decap_4 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_4 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_decap_4 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_4 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_fill_2 FILLER_28_410 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_decap_8 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_50 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_decap_8 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_82 ();
 sg13g2_decap_4 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_357 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_4 FILLER_29_385 ();
 sg13g2_fill_1 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_4 FILLER_29_409 ();
 sg13g2_fill_2 FILLER_29_413 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_decap_8 FILLER_30_44 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_decap_8 FILLER_30_88 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_decap_4 FILLER_31_39 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_decap_8 FILLER_31_65 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_4 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_401 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_fill_1 FILLER_31_409 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_decap_4 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_212 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_decap_4 FILLER_32_283 ();
 sg13g2_decap_4 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_decap_4 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_decap_4 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_4 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_decap_8 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_4 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_decap_8 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_decap_4 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_2 FILLER_33_404 ();
 sg13g2_decap_8 FILLER_33_414 ();
 sg13g2_decap_8 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_decap_4 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_decap_4 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_251 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_4 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_34_423 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_decap_8 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_120 ();
 sg13g2_decap_4 FILLER_35_127 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_decap_4 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_decap_4 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_decap_4 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_decap_4 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_decap_4 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_decap_4 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_decap_4 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_1 FILLER_36_351 ();
 sg13g2_decap_4 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_59 ();
 sg13g2_fill_2 FILLER_37_69 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_2 FILLER_37_80 ();
 sg13g2_fill_1 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_decap_4 FILLER_37_250 ();
 sg13g2_decap_8 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_203 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_226 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_decap_4 FILLER_38_352 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_4 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_384 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
