module tt_um_dvxf_dj8v (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DJ8.ACC[0] ;
 wire \DJ8.ACC[1] ;
 wire \DJ8.ACC[2] ;
 wire \DJ8.ACC[3] ;
 wire \DJ8.ACC[4] ;
 wire \DJ8.ACC[5] ;
 wire \DJ8.ACC[6] ;
 wire \DJ8.ACC[7] ;
 wire \DJ8.ALU.c_in ;
 wire \DJ8.ALU.opalu[0] ;
 wire \DJ8.ALU.opalu[1] ;
 wire \DJ8.ALU.opalu[2] ;
 wire \DJ8.EF[0] ;
 wire \DJ8.EF[10] ;
 wire \DJ8.EF[11] ;
 wire \DJ8.EF[12] ;
 wire \DJ8.EF[13] ;
 wire \DJ8.EF[14] ;
 wire \DJ8.EF[15] ;
 wire \DJ8.EF[1] ;
 wire \DJ8.EF[2] ;
 wire \DJ8.EF[3] ;
 wire \DJ8.EF[4] ;
 wire \DJ8.EF[5] ;
 wire \DJ8.EF[6] ;
 wire \DJ8.EF[7] ;
 wire \DJ8.EF[8] ;
 wire \DJ8.EF[9] ;
 wire \DJ8.GH[0] ;
 wire \DJ8.GH[10] ;
 wire \DJ8.GH[11] ;
 wire \DJ8.GH[12] ;
 wire \DJ8.GH[13] ;
 wire \DJ8.GH[14] ;
 wire \DJ8.GH[15] ;
 wire \DJ8.GH[1] ;
 wire \DJ8.GH[2] ;
 wire \DJ8.GH[3] ;
 wire \DJ8.GH[4] ;
 wire \DJ8.GH[5] ;
 wire \DJ8.GH[6] ;
 wire \DJ8.GH[7] ;
 wire \DJ8.GH[8] ;
 wire \DJ8.GH[9] ;
 wire \DJ8.REGS.regs[1][0] ;
 wire \DJ8.REGS.regs[1][1] ;
 wire \DJ8.REGS.regs[1][2] ;
 wire \DJ8.REGS.regs[1][3] ;
 wire \DJ8.REGS.regs[1][4] ;
 wire \DJ8.REGS.regs[1][5] ;
 wire \DJ8.REGS.regs[1][6] ;
 wire \DJ8.REGS.regs[1][7] ;
 wire \DJ8.REGS.regs[2][0] ;
 wire \DJ8.REGS.regs[2][1] ;
 wire \DJ8.REGS.regs[2][2] ;
 wire \DJ8.REGS.regs[2][3] ;
 wire \DJ8.REGS.regs[2][4] ;
 wire \DJ8.REGS.regs[2][5] ;
 wire \DJ8.REGS.regs[2][6] ;
 wire \DJ8.REGS.regs[2][7] ;
 wire \DJ8.REGS.regs[3][0] ;
 wire \DJ8.REGS.regs[3][1] ;
 wire \DJ8.REGS.regs[3][2] ;
 wire \DJ8.REGS.regs[3][3] ;
 wire \DJ8.REGS.regs[3][4] ;
 wire \DJ8.REGS.regs[3][5] ;
 wire \DJ8.REGS.regs[3][6] ;
 wire \DJ8.REGS.regs[3][7] ;
 wire \DJ8.REGS.write_addr[0] ;
 wire \DJ8.REGS.write_addr[1] ;
 wire \DJ8.REGS.write_addr[2] ;
 wire \DJ8.flag_Z ;
 wire \DJ8.ir[0] ;
 wire \DJ8.ir[14] ;
 wire \DJ8.ir[15] ;
 wire \DJ8.ir[1] ;
 wire \DJ8.ir[2] ;
 wire \DJ8.ir[3] ;
 wire \DJ8.ir[4] ;
 wire \DJ8.ir[5] ;
 wire \DJ8.ir[6] ;
 wire \DJ8.ir[7] ;
 wire \DJ8.pc[0] ;
 wire \DJ8.pc[10] ;
 wire \DJ8.pc[11] ;
 wire \DJ8.pc[12] ;
 wire \DJ8.pc[13] ;
 wire \DJ8.pc[14] ;
 wire \DJ8.pc[1] ;
 wire \DJ8.pc[2] ;
 wire \DJ8.pc[3] ;
 wire \DJ8.pc[4] ;
 wire \DJ8.pc[5] ;
 wire \DJ8.pc[6] ;
 wire \DJ8.pc[7] ;
 wire \DJ8.pc[8] ;
 wire \DJ8.pc[9] ;
 wire \DJ8.state[0] ;
 wire \DJ8.state[1] ;
 wire \DJ8.state[2] ;
 wire \DJ8.state[3] ;
 wire \DJ8.we ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire clknet_0_clk;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire net113;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][0]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0043_),
    .Q_N(_1190_),
    .Q(\DJ8.ACC[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][1]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0044_),
    .Q_N(_0020_),
    .Q(\DJ8.ACC[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][2]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0045_),
    .Q_N(_0022_),
    .Q(\DJ8.ACC[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][3]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(_0046_),
    .Q_N(_0024_),
    .Q(\DJ8.ACC[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][4]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0047_),
    .Q_N(_0025_),
    .Q(\DJ8.ACC[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][5]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(_0048_),
    .Q_N(_0027_),
    .Q(\DJ8.ACC[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][6]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0049_),
    .Q_N(_0029_),
    .Q(\DJ8.ACC[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][7]$_DFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net90),
    .D(_0050_),
    .Q_N(\DJ8.ACC[7] ),
    .Q(_0031_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][0]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(_0051_),
    .Q_N(_1189_),
    .Q(\DJ8.REGS.regs[1][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][1]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net86),
    .D(_0052_),
    .Q_N(_1188_),
    .Q(\DJ8.REGS.regs[1][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][2]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0053_),
    .Q_N(_1187_),
    .Q(\DJ8.REGS.regs[1][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][3]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0054_),
    .Q_N(_1186_),
    .Q(\DJ8.REGS.regs[1][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][4]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net88),
    .D(_0055_),
    .Q_N(_1185_),
    .Q(\DJ8.REGS.regs[1][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][5]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0056_),
    .Q_N(_1184_),
    .Q(\DJ8.REGS.regs[1][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][6]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0057_),
    .Q_N(_1183_),
    .Q(\DJ8.REGS.regs[1][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][7]$_DFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net89),
    .D(_0058_),
    .Q_N(\DJ8.REGS.regs[1][7] ),
    .Q(_0032_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][0]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net88),
    .D(_0059_),
    .Q_N(_1182_),
    .Q(\DJ8.REGS.regs[2][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][1]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0060_),
    .Q_N(_1181_),
    .Q(\DJ8.REGS.regs[2][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][2]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net86),
    .D(_0061_),
    .Q_N(_1180_),
    .Q(\DJ8.REGS.regs[2][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][3]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0062_),
    .Q_N(_1179_),
    .Q(\DJ8.REGS.regs[2][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][4]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net86),
    .D(_0063_),
    .Q_N(_1178_),
    .Q(\DJ8.REGS.regs[2][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][5]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net87),
    .D(_0064_),
    .Q_N(_1177_),
    .Q(\DJ8.REGS.regs[2][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][6]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net89),
    .D(_0065_),
    .Q_N(_1176_),
    .Q(\DJ8.REGS.regs[2][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][7]$_DFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net87),
    .D(_0066_),
    .Q_N(\DJ8.REGS.regs[2][7] ),
    .Q(_0033_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][0]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0067_),
    .Q_N(_1175_),
    .Q(\DJ8.REGS.regs[3][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][1]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net86),
    .D(_0068_),
    .Q_N(_1174_),
    .Q(\DJ8.REGS.regs[3][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][2]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net87),
    .D(_0069_),
    .Q_N(_1173_),
    .Q(\DJ8.REGS.regs[3][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][3]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0070_),
    .Q_N(_1172_),
    .Q(\DJ8.REGS.regs[3][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][4]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net87),
    .D(_0071_),
    .Q_N(_1171_),
    .Q(\DJ8.REGS.regs[3][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][5]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0072_),
    .Q_N(_1170_),
    .Q(\DJ8.REGS.regs[3][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][6]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net88),
    .D(_0073_),
    .Q_N(_1169_),
    .Q(\DJ8.REGS.regs[3][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][7]$_DFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0074_),
    .Q_N(\DJ8.REGS.regs[3][7] ),
    .Q(_0034_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][0]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net94),
    .D(_0075_),
    .Q_N(_1168_),
    .Q(\DJ8.EF[8] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][1]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net93),
    .D(_0076_),
    .Q_N(_1167_),
    .Q(\DJ8.EF[9] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][2]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net93),
    .D(_0077_),
    .Q_N(_1166_),
    .Q(\DJ8.EF[10] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][3]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0078_),
    .Q_N(_1165_),
    .Q(\DJ8.EF[11] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][4]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net96),
    .D(_0079_),
    .Q_N(_1164_),
    .Q(\DJ8.EF[12] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][5]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net93),
    .D(_0080_),
    .Q_N(_1163_),
    .Q(\DJ8.EF[13] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][6]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net93),
    .D(_0081_),
    .Q_N(_1162_),
    .Q(\DJ8.EF[14] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][7]$_DFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0082_),
    .Q_N(\DJ8.EF[15] ),
    .Q(_0035_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][0]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net97),
    .D(_0083_),
    .Q_N(_1161_),
    .Q(\DJ8.EF[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][1]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0084_),
    .Q_N(_0008_),
    .Q(\DJ8.EF[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][2]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(_0085_),
    .Q_N(_0011_),
    .Q(\DJ8.EF[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][3]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0086_),
    .Q_N(_0014_),
    .Q(\DJ8.EF[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][4]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(_0087_),
    .Q_N(_0017_),
    .Q(\DJ8.EF[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][5]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0088_),
    .Q_N(_1160_),
    .Q(\DJ8.EF[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][6]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0089_),
    .Q_N(_1159_),
    .Q(\DJ8.EF[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][7]$_DFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0090_),
    .Q_N(\DJ8.EF[7] ),
    .Q(_0036_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][0]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0091_),
    .Q_N(_1158_),
    .Q(\DJ8.GH[8] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][1]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net95),
    .D(_0092_),
    .Q_N(_1157_),
    .Q(\DJ8.GH[9] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][2]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net95),
    .D(_0093_),
    .Q_N(_1156_),
    .Q(\DJ8.GH[10] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][3]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net95),
    .D(_0094_),
    .Q_N(_1155_),
    .Q(\DJ8.GH[11] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][4]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(_0095_),
    .Q_N(_1154_),
    .Q(\DJ8.GH[12] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][5]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net95),
    .D(_0096_),
    .Q_N(_1153_),
    .Q(\DJ8.GH[13] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][6]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(_0097_),
    .Q_N(_1152_),
    .Q(\DJ8.GH[14] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][7]$_DFFE_PN1P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(_0098_),
    .Q_N(\DJ8.GH[15] ),
    .Q(_0037_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][0]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net94),
    .D(_0099_),
    .Q_N(_1151_),
    .Q(\DJ8.GH[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][1]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0100_),
    .Q_N(_0007_),
    .Q(\DJ8.GH[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][2]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0101_),
    .Q_N(_0010_),
    .Q(\DJ8.GH[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][3]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0102_),
    .Q_N(_0013_),
    .Q(\DJ8.GH[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][4]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0103_),
    .Q_N(_0016_),
    .Q(\DJ8.GH[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][5]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net96),
    .D(_0104_),
    .Q_N(_1150_),
    .Q(\DJ8.GH[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][6]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net96),
    .D(_0105_),
    .Q_N(_1149_),
    .Q(\DJ8.GH[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][7]$_DFFE_PN1P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net96),
    .D(_0106_),
    .Q_N(\DJ8.GH[7] ),
    .Q(_0038_));
 sg13g2_dfrbp_1 \DJ8.flag_C$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net91),
    .D(_0107_),
    .Q_N(_1148_),
    .Q(\DJ8.ALU.c_in ));
 sg13g2_dfrbp_1 \DJ8.flag_Z$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net91),
    .D(_0108_),
    .Q_N(_1147_),
    .Q(\DJ8.flag_Z ));
 sg13g2_dfrbp_1 \DJ8.ir[0]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0109_),
    .Q_N(_1146_),
    .Q(\DJ8.ir[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[10]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0110_),
    .Q_N(_0002_),
    .Q(\DJ8.REGS.write_addr[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[11]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net103),
    .D(_0111_),
    .Q_N(_1145_),
    .Q(\DJ8.ALU.opalu[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[12]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net103),
    .D(_0112_),
    .Q_N(_1144_),
    .Q(\DJ8.ALU.opalu[1] ));
 sg13g2_dfrbp_1 \DJ8.ir[13]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0113_),
    .Q_N(_0018_),
    .Q(\DJ8.ALU.opalu[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[14]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0114_),
    .Q_N(_1143_),
    .Q(\DJ8.ir[14] ));
 sg13g2_dfrbp_1 \DJ8.ir[15]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0115_),
    .Q_N(_1142_),
    .Q(\DJ8.ir[15] ));
 sg13g2_dfrbp_1 \DJ8.ir[1]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0116_),
    .Q_N(_0019_),
    .Q(\DJ8.ir[1] ));
 sg13g2_dfrbp_1 \DJ8.ir[2]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0117_),
    .Q_N(_0021_),
    .Q(\DJ8.ir[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[3]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0118_),
    .Q_N(_0023_),
    .Q(\DJ8.ir[3] ));
 sg13g2_dfrbp_1 \DJ8.ir[4]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0119_),
    .Q_N(_0005_),
    .Q(\DJ8.ir[4] ));
 sg13g2_dfrbp_1 \DJ8.ir[5]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net91),
    .D(_0120_),
    .Q_N(_0026_),
    .Q(\DJ8.ir[5] ));
 sg13g2_dfrbp_1 \DJ8.ir[6]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net91),
    .D(_0121_),
    .Q_N(_0028_),
    .Q(\DJ8.ir[6] ));
 sg13g2_dfrbp_1 \DJ8.ir[7]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net97),
    .D(_0122_),
    .Q_N(_0003_),
    .Q(\DJ8.ir[7] ));
 sg13g2_dfrbp_1 \DJ8.ir[8]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net99),
    .D(_0123_),
    .Q_N(_1141_),
    .Q(\DJ8.REGS.write_addr[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[9]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0124_),
    .Q_N(_1140_),
    .Q(\DJ8.REGS.write_addr[1] ));
 sg13g2_dfrbp_1 \DJ8.pc[0]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0125_),
    .Q_N(_0006_),
    .Q(\DJ8.pc[0] ));
 sg13g2_dfrbp_1 \DJ8.pc[10]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net100),
    .D(_0126_),
    .Q_N(_1139_),
    .Q(\DJ8.pc[10] ));
 sg13g2_dfrbp_1 \DJ8.pc[11]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net100),
    .D(_0127_),
    .Q_N(_1138_),
    .Q(\DJ8.pc[11] ));
 sg13g2_dfrbp_1 \DJ8.pc[12]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(_0128_),
    .Q_N(_1137_),
    .Q(\DJ8.pc[12] ));
 sg13g2_dfrbp_1 \DJ8.pc[13]$_DFFE_PN1P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net96),
    .D(_0129_),
    .Q_N(\DJ8.pc[13] ),
    .Q(_0039_));
 sg13g2_dfrbp_1 \DJ8.pc[14]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net96),
    .D(_0130_),
    .Q_N(_0004_),
    .Q(\DJ8.pc[14] ));
 sg13g2_dfrbp_1 \DJ8.pc[1]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0131_),
    .Q_N(_0009_),
    .Q(\DJ8.pc[1] ));
 sg13g2_dfrbp_1 \DJ8.pc[2]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0132_),
    .Q_N(_0012_),
    .Q(\DJ8.pc[2] ));
 sg13g2_dfrbp_1 \DJ8.pc[3]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net102),
    .D(_0133_),
    .Q_N(_0015_),
    .Q(\DJ8.pc[3] ));
 sg13g2_dfrbp_1 \DJ8.pc[4]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net97),
    .D(_0134_),
    .Q_N(_1136_),
    .Q(\DJ8.pc[4] ));
 sg13g2_dfrbp_1 \DJ8.pc[5]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net97),
    .D(_0135_),
    .Q_N(_1135_),
    .Q(\DJ8.pc[5] ));
 sg13g2_dfrbp_1 \DJ8.pc[6]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0136_),
    .Q_N(_1134_),
    .Q(\DJ8.pc[6] ));
 sg13g2_dfrbp_1 \DJ8.pc[7]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net101),
    .D(_0137_),
    .Q_N(_1133_),
    .Q(\DJ8.pc[7] ));
 sg13g2_dfrbp_1 \DJ8.pc[8]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net98),
    .D(_0138_),
    .Q_N(_1132_),
    .Q(\DJ8.pc[8] ));
 sg13g2_dfrbp_1 \DJ8.pc[9]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net98),
    .D(_0139_),
    .Q_N(_1131_),
    .Q(\DJ8.pc[9] ));
 sg13g2_dfrbp_1 \DJ8.state[0]$_DFF_PN1_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(_0041_),
    .Q_N(\DJ8.state[0] ),
    .Q(_1192_));
 sg13g2_dfrbp_1 \DJ8.state[1]$_DFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net101),
    .D(\DJ8.state[2] ),
    .Q_N(_0001_),
    .Q(\DJ8.state[1] ));
 sg13g2_dfrbp_1 \DJ8.state[2]$_DFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(\DJ8.state[0] ),
    .Q_N(_1191_),
    .Q(\DJ8.state[2] ));
 sg13g2_dfrbp_1 \DJ8.state[3]$_DFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net101),
    .D(_0000_),
    .Q_N(_0030_),
    .Q(\DJ8.state[3] ));
 sg13g2_dfrbp_1 \DJ8.we$_DFFE_NN1P_  (.CLK(net113),
    .RESET_B(net102),
    .D(_0140_),
    .Q_N(\DJ8.we ),
    .Q(_0040_));
 sg13g2_buf_2 _1194_ (.A(\DJ8.ir[0] ),
    .X(_0407_));
 sg13g2_buf_8 _1195_ (.A(\DJ8.ir[14] ),
    .X(_0408_));
 sg13g2_buf_8 _1196_ (.A(\DJ8.ir[15] ),
    .X(_0409_));
 sg13g2_nor2b_1 _1197_ (.A(net85),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_nand2_2 _1198_ (.Y(_0411_),
    .A(_0407_),
    .B(_0410_));
 sg13g2_nor2_1 _1199_ (.A(_0001_),
    .B(_0411_),
    .Y(_0000_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1201_ (.A(_0018_),
    .X(_0412_));
 sg13g2_inv_2 _1202_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_buf_1 _1203_ (.A(\DJ8.ALU.opalu[1] ),
    .X(_0414_));
 sg13g2_buf_1 _1204_ (.A(\DJ8.ALU.opalu[0] ),
    .X(_0415_));
 sg13g2_inv_1 _1205_ (.Y(_0416_),
    .A(net84));
 sg13g2_nand2_1 _1206_ (.Y(_0417_),
    .A(_0414_),
    .B(_0416_));
 sg13g2_nor2_1 _1207_ (.A(_0413_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_buf_1 _1208_ (.A(_0418_),
    .X(_0419_));
 sg13g2_buf_2 _1209_ (.A(_0012_),
    .X(_0420_));
 sg13g2_nor2_2 _1210_ (.A(_0420_),
    .B(_0015_),
    .Y(_0421_));
 sg13g2_buf_2 _1211_ (.A(_0009_),
    .X(_0422_));
 sg13g2_buf_1 _1212_ (.A(_0015_),
    .X(_0423_));
 sg13g2_nand2_1 _1213_ (.Y(_0424_),
    .A(_0420_),
    .B(net83));
 sg13g2_nor2_1 _1214_ (.A(_0422_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_buf_1 _1215_ (.A(_0006_),
    .X(_0426_));
 sg13g2_o21ai_1 _1216_ (.B1(net82),
    .Y(_0427_),
    .A1(_0421_),
    .A2(_0425_));
 sg13g2_nor2b_1 _1217_ (.A(_0420_),
    .B_N(_0015_),
    .Y(_0428_));
 sg13g2_nor2_1 _1218_ (.A(net82),
    .B(_0422_),
    .Y(_0429_));
 sg13g2_buf_2 _1219_ (.A(\DJ8.state[2] ),
    .X(_0430_));
 sg13g2_nand2b_1 _1220_ (.Y(_0431_),
    .B(_0409_),
    .A_N(\DJ8.ir[14] ));
 sg13g2_nor2_2 _1221_ (.A(_0407_),
    .B(\DJ8.ir[1] ),
    .Y(_0432_));
 sg13g2_nor4_2 _1222_ (.A(_0430_),
    .B(\DJ8.state[0] ),
    .C(_0431_),
    .Y(_0433_),
    .D(_0432_));
 sg13g2_buf_8 _1223_ (.A(_0433_),
    .X(_0434_));
 sg13g2_a21oi_1 _1224_ (.A1(_0428_),
    .A2(_0429_),
    .Y(_0435_),
    .B1(net63));
 sg13g2_buf_2 _1225_ (.A(\DJ8.ir[4] ),
    .X(_0436_));
 sg13g2_buf_8 _1226_ (.A(_0436_),
    .X(_0437_));
 sg13g2_buf_1 _1227_ (.A(net75),
    .X(_0438_));
 sg13g2_buf_1 _1228_ (.A(net68),
    .X(_0439_));
 sg13g2_buf_2 _1229_ (.A(_0014_),
    .X(_0440_));
 sg13g2_buf_1 _1230_ (.A(_0008_),
    .X(_0441_));
 sg13g2_nor2b_1 _1231_ (.A(_0440_),
    .B_N(_0441_),
    .Y(_0442_));
 sg13g2_buf_2 _1232_ (.A(_0007_),
    .X(_0443_));
 sg13g2_nor2b_1 _1233_ (.A(_0438_),
    .B_N(_0443_),
    .Y(_0444_));
 sg13g2_buf_2 _1234_ (.A(_0013_),
    .X(_0445_));
 sg13g2_inv_1 _1235_ (.Y(_0446_),
    .A(_0445_));
 sg13g2_a22oi_1 _1236_ (.Y(_0447_),
    .B1(_0444_),
    .B2(_0446_),
    .A2(_0442_),
    .A1(net62));
 sg13g2_buf_2 _1237_ (.A(_0016_),
    .X(_0448_));
 sg13g2_inv_1 _1238_ (.Y(_0449_),
    .A(_0448_));
 sg13g2_buf_2 _1239_ (.A(_0010_),
    .X(_0450_));
 sg13g2_or2_1 _1240_ (.X(_0451_),
    .B(_0450_),
    .A(net68));
 sg13g2_buf_1 _1241_ (.A(_0011_),
    .X(_0452_));
 sg13g2_buf_2 _1242_ (.A(_0017_),
    .X(_0453_));
 sg13g2_nand3b_1 _1243_ (.B(_0453_),
    .C(net62),
    .Y(_0454_),
    .A_N(_0452_));
 sg13g2_o21ai_1 _1244_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0449_),
    .A2(_0451_));
 sg13g2_nor2b_1 _1245_ (.A(_0441_),
    .B_N(_0440_),
    .Y(_0456_));
 sg13g2_nand2_1 _1246_ (.Y(_0457_),
    .A(net62),
    .B(_0456_));
 sg13g2_nor2b_1 _1247_ (.A(_0443_),
    .B_N(_0445_),
    .Y(_0458_));
 sg13g2_nand2b_1 _1248_ (.Y(_0459_),
    .B(_0458_),
    .A_N(net62));
 sg13g2_nand4_1 _1249_ (.B(_0455_),
    .C(_0457_),
    .A(_0447_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_mux2_1 _1250_ (.A0(_0443_),
    .A1(_0441_),
    .S(_0436_),
    .X(_0461_));
 sg13g2_buf_1 _1251_ (.A(_0461_),
    .X(_0462_));
 sg13g2_nor2_1 _1252_ (.A(_0440_),
    .B(_0453_),
    .Y(_0463_));
 sg13g2_nor3_1 _1253_ (.A(_0436_),
    .B(_0445_),
    .C(_0448_),
    .Y(_0464_));
 sg13g2_a21o_1 _1254_ (.A2(_0463_),
    .A1(net75),
    .B1(_0464_),
    .X(_0465_));
 sg13g2_buf_1 _1255_ (.A(_0465_),
    .X(_0466_));
 sg13g2_or4_1 _1256_ (.A(_0430_),
    .B(\DJ8.state[0] ),
    .C(_0431_),
    .D(_0432_),
    .X(_0467_));
 sg13g2_buf_1 _1257_ (.A(_0467_),
    .X(_0468_));
 sg13g2_a21oi_1 _1258_ (.A1(_0462_),
    .A2(_0466_),
    .Y(_0469_),
    .B1(net61));
 sg13g2_mux2_1 _1259_ (.A0(\DJ8.GH[0] ),
    .A1(\DJ8.EF[0] ),
    .S(_0436_),
    .X(_0470_));
 sg13g2_nor4_2 _1260_ (.A(_0430_),
    .B(_0431_),
    .C(_0432_),
    .Y(_0471_),
    .D(_0470_));
 sg13g2_or2_1 _1261_ (.X(_0472_),
    .B(_0471_),
    .A(\DJ8.state[0] ));
 sg13g2_buf_2 _1262_ (.A(_0472_),
    .X(_0473_));
 sg13g2_a221oi_1 _1263_ (.B2(_0469_),
    .C1(_0473_),
    .B1(_0460_),
    .A1(_0427_),
    .Y(_0474_),
    .A2(_0435_));
 sg13g2_inv_1 _1264_ (.Y(_0475_),
    .A(_0420_));
 sg13g2_nand2_1 _1265_ (.Y(_0476_),
    .A(_0475_),
    .B(net83));
 sg13g2_nand2b_1 _1266_ (.Y(_0477_),
    .B(_0448_),
    .A_N(_0445_));
 sg13g2_nand2b_1 _1267_ (.Y(_0478_),
    .B(_0453_),
    .A_N(_0440_));
 sg13g2_mux2_1 _1268_ (.A0(_0477_),
    .A1(_0478_),
    .S(net68),
    .X(_0479_));
 sg13g2_mux2_1 _1269_ (.A0(_0476_),
    .A1(_0479_),
    .S(net63),
    .X(_0480_));
 sg13g2_nor3_1 _1270_ (.A(_0430_),
    .B(_0432_),
    .C(_0470_),
    .Y(_0481_));
 sg13g2_buf_1 _1271_ (.A(\DJ8.state[0] ),
    .X(_0482_));
 sg13g2_inv_1 _1272_ (.Y(_0483_),
    .A(net81));
 sg13g2_mux2_1 _1273_ (.A0(_0450_),
    .A1(_0452_),
    .S(net75),
    .X(_0484_));
 sg13g2_and3_1 _1274_ (.X(_0485_),
    .A(_0483_),
    .B(_0410_),
    .C(_0484_));
 sg13g2_inv_1 _1275_ (.Y(_0486_),
    .A(_0422_));
 sg13g2_nor2_1 _1276_ (.A(_0483_),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_a21oi_1 _1277_ (.A1(_0481_),
    .A2(_0485_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_inv_1 _1278_ (.Y(_0489_),
    .A(_0004_));
 sg13g2_nor2b_1 _1279_ (.A(_0436_),
    .B_N(\DJ8.GH[15] ),
    .Y(_0490_));
 sg13g2_a21o_1 _1280_ (.A2(net75),
    .A1(\DJ8.EF[15] ),
    .B1(_0490_),
    .X(_0491_));
 sg13g2_mux2_1 _1281_ (.A0(_0489_),
    .A1(_0491_),
    .S(_0433_),
    .X(_0492_));
 sg13g2_buf_1 _1282_ (.A(_0492_),
    .X(_0493_));
 sg13g2_o21ai_1 _1283_ (.B1(net53),
    .Y(_0494_),
    .A1(_0480_),
    .A2(_0488_));
 sg13g2_inv_1 _1284_ (.Y(_0495_),
    .A(net3));
 sg13g2_a21oi_1 _1285_ (.A1(\DJ8.EF[15] ),
    .A2(net75),
    .Y(_0496_),
    .B1(_0490_));
 sg13g2_mux2_1 _1286_ (.A0(_0004_),
    .A1(_0496_),
    .S(_0433_),
    .X(_0497_));
 sg13g2_buf_8 _1287_ (.A(_0497_),
    .X(_0498_));
 sg13g2_buf_8 _1288_ (.A(_0498_),
    .X(_0499_));
 sg13g2_buf_1 _1289_ (.A(_0408_),
    .X(_0500_));
 sg13g2_inv_1 _1290_ (.Y(_0501_),
    .A(net74));
 sg13g2_nand2_2 _1291_ (.Y(_0502_),
    .A(net67),
    .B(\DJ8.ir[1] ));
 sg13g2_a21oi_1 _1292_ (.A1(_0495_),
    .A2(net42),
    .Y(_0503_),
    .B1(_0502_));
 sg13g2_o21ai_1 _1293_ (.B1(_0503_),
    .Y(_0504_),
    .A1(_0474_),
    .A2(_0494_));
 sg13g2_buf_2 _1294_ (.A(\DJ8.ir[6] ),
    .X(_0505_));
 sg13g2_mux2_1 _1295_ (.A0(_0505_),
    .A1(\DJ8.REGS.write_addr[1] ),
    .S(net85),
    .X(_0506_));
 sg13g2_buf_2 _1296_ (.A(_0506_),
    .X(_0507_));
 sg13g2_buf_1 _1297_ (.A(_0507_),
    .X(_0508_));
 sg13g2_mux2_1 _1298_ (.A0(_0003_),
    .A1(_0002_),
    .S(net85),
    .X(_0509_));
 sg13g2_buf_2 _1299_ (.A(_0509_),
    .X(_0510_));
 sg13g2_nor2b_1 _1300_ (.A(net60),
    .B_N(_0510_),
    .Y(_0511_));
 sg13g2_buf_2 _1301_ (.A(\DJ8.ir[5] ),
    .X(_0512_));
 sg13g2_mux2_1 _1302_ (.A0(_0512_),
    .A1(\DJ8.REGS.write_addr[0] ),
    .S(net85),
    .X(_0513_));
 sg13g2_buf_2 _1303_ (.A(_0513_),
    .X(_0514_));
 sg13g2_buf_8 _1304_ (.A(_0514_),
    .X(_0515_));
 sg13g2_nor2_1 _1305_ (.A(\DJ8.ACC[1] ),
    .B(net59),
    .Y(_0516_));
 sg13g2_nand2_1 _1306_ (.Y(_0517_),
    .A(_0511_),
    .B(_0516_));
 sg13g2_nand2b_1 _1307_ (.Y(_0518_),
    .B(_0510_),
    .A_N(_0507_));
 sg13g2_nand2_1 _1308_ (.Y(_0519_),
    .A(net85),
    .B(_0002_));
 sg13g2_nand2b_1 _1309_ (.Y(_0520_),
    .B(_0003_),
    .A_N(net85));
 sg13g2_nand4_1 _1310_ (.B(_0519_),
    .C(_0520_),
    .A(\DJ8.GH[9] ),
    .Y(_0521_),
    .D(net60));
 sg13g2_buf_2 _1311_ (.A(_0515_),
    .X(_0522_));
 sg13g2_a21oi_1 _1312_ (.A1(_0518_),
    .A2(_0521_),
    .Y(_0523_),
    .B1(net52));
 sg13g2_buf_1 _1313_ (.A(_0507_),
    .X(_0524_));
 sg13g2_inv_1 _1314_ (.Y(_0525_),
    .A(\DJ8.EF[9] ));
 sg13g2_inv_1 _1315_ (.Y(_0526_),
    .A(\DJ8.EF[1] ));
 sg13g2_mux2_1 _1316_ (.A0(_0525_),
    .A1(_0526_),
    .S(net59),
    .X(_0527_));
 sg13g2_nand3_1 _1317_ (.B(net60),
    .C(_0522_),
    .A(\DJ8.GH[1] ),
    .Y(_0528_));
 sg13g2_o21ai_1 _1318_ (.B1(_0528_),
    .Y(_0529_),
    .A1(net58),
    .A2(_0527_));
 sg13g2_and2_1 _1319_ (.A(_0519_),
    .B(_0520_),
    .X(_0530_));
 sg13g2_buf_1 _1320_ (.A(_0530_),
    .X(_0531_));
 sg13g2_inv_1 _1321_ (.Y(_0532_),
    .A(\DJ8.REGS.regs[2][1] ));
 sg13g2_inv_1 _1322_ (.Y(_0533_),
    .A(\DJ8.REGS.regs[3][1] ));
 sg13g2_mux2_1 _1323_ (.A0(_0532_),
    .A1(_0533_),
    .S(net59),
    .X(_0534_));
 sg13g2_buf_1 _1324_ (.A(_0510_),
    .X(_0535_));
 sg13g2_o21ai_1 _1325_ (.B1(net57),
    .Y(_0536_),
    .A1(\DJ8.REGS.regs[1][1] ),
    .A2(net60));
 sg13g2_a221oi_1 _1326_ (.B2(net58),
    .C1(_0536_),
    .B1(_0534_),
    .A1(_0511_),
    .Y(_0537_),
    .A2(_0516_));
 sg13g2_a221oi_1 _1327_ (.B2(_0531_),
    .C1(_0537_),
    .B1(_0529_),
    .A1(_0517_),
    .Y(_0538_),
    .A2(_0523_));
 sg13g2_buf_1 _1328_ (.A(_0502_),
    .X(_0539_));
 sg13g2_nand2b_2 _1329_ (.Y(_0540_),
    .B(net51),
    .A_N(_0538_));
 sg13g2_nand2_2 _1330_ (.Y(_0541_),
    .A(_0504_),
    .B(_0540_));
 sg13g2_and2_1 _1331_ (.A(_0500_),
    .B(_0019_),
    .X(_0542_));
 sg13g2_a21oi_2 _1332_ (.B1(_0542_),
    .Y(_0543_),
    .A2(_0020_),
    .A1(net67));
 sg13g2_nor2_2 _1333_ (.A(_0541_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a21o_1 _1334_ (.A2(_0020_),
    .A1(net67),
    .B1(_0542_),
    .X(_0545_));
 sg13g2_buf_1 _1335_ (.A(_0545_),
    .X(_0546_));
 sg13g2_a21oi_2 _1336_ (.B1(_0546_),
    .Y(_0547_),
    .A2(_0540_),
    .A1(_0504_));
 sg13g2_nor2_2 _1337_ (.A(_0544_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_and2_1 _1338_ (.A(_0500_),
    .B(_0407_),
    .X(_0549_));
 sg13g2_a21oi_2 _1339_ (.B1(_0549_),
    .Y(_0550_),
    .A2(\DJ8.ACC[0] ),
    .A1(net67));
 sg13g2_nor2b_1 _1340_ (.A(net68),
    .B_N(_0450_),
    .Y(_0551_));
 sg13g2_and2_1 _1341_ (.A(_0437_),
    .B(_0452_),
    .X(_0552_));
 sg13g2_nor2_1 _1342_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_mux2_1 _1343_ (.A0(_0486_),
    .A1(_0553_),
    .S(net63),
    .X(_0554_));
 sg13g2_xnor2_1 _1344_ (.Y(_0555_),
    .A(_0473_),
    .B(_0554_));
 sg13g2_inv_1 _1345_ (.Y(_0556_),
    .A(net82));
 sg13g2_inv_1 _1346_ (.Y(_0557_),
    .A(_0462_));
 sg13g2_mux2_1 _1347_ (.A0(_0556_),
    .A1(_0557_),
    .S(net63),
    .X(_0558_));
 sg13g2_buf_1 _1348_ (.A(net61),
    .X(_0559_));
 sg13g2_nand2b_1 _1349_ (.Y(_0560_),
    .B(_0445_),
    .A_N(_0448_));
 sg13g2_nand2b_1 _1350_ (.Y(_0561_),
    .B(_0440_),
    .A_N(_0453_));
 sg13g2_mux2_1 _1351_ (.A0(_0560_),
    .A1(_0561_),
    .S(net68),
    .X(_0562_));
 sg13g2_nor2_1 _1352_ (.A(net50),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_buf_1 _1353_ (.A(net63),
    .X(_0564_));
 sg13g2_nand2b_1 _1354_ (.Y(_0565_),
    .B(_0420_),
    .A_N(net83));
 sg13g2_nor2_1 _1355_ (.A(net49),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nor4_1 _1356_ (.A(_0498_),
    .B(_0558_),
    .C(_0563_),
    .D(_0566_),
    .Y(_0567_));
 sg13g2_nor4_1 _1357_ (.A(net42),
    .B(_0480_),
    .C(_0554_),
    .D(_0558_),
    .Y(_0568_));
 sg13g2_a21oi_2 _1358_ (.B1(_0568_),
    .Y(_0569_),
    .A2(_0567_),
    .A1(_0555_));
 sg13g2_nor4_1 _1359_ (.A(_0004_),
    .B(net82),
    .C(net83),
    .D(net63),
    .Y(_0570_));
 sg13g2_mux2_1 _1360_ (.A0(_0448_),
    .A1(_0453_),
    .S(net75),
    .X(_0571_));
 sg13g2_buf_2 _1361_ (.A(_0571_),
    .X(_0572_));
 sg13g2_nor4_1 _1362_ (.A(net61),
    .B(_0496_),
    .C(_0462_),
    .D(_0572_),
    .Y(_0573_));
 sg13g2_or2_1 _1363_ (.X(_0574_),
    .B(_0573_),
    .A(_0570_));
 sg13g2_mux2_1 _1364_ (.A0(_0445_),
    .A1(_0440_),
    .S(_0437_),
    .X(_0575_));
 sg13g2_nor2b_1 _1365_ (.A(_0484_),
    .B_N(_0575_),
    .Y(_0576_));
 sg13g2_nor2_1 _1366_ (.A(_0422_),
    .B(_0475_),
    .Y(_0577_));
 sg13g2_mux2_1 _1367_ (.A0(_0576_),
    .A1(_0577_),
    .S(net61),
    .X(_0578_));
 sg13g2_inv_1 _1368_ (.Y(_0579_),
    .A(_0575_));
 sg13g2_mux2_1 _1369_ (.A0(_0475_),
    .A1(_0579_),
    .S(_0433_),
    .X(_0580_));
 sg13g2_mux2_1 _1370_ (.A0(_0578_),
    .A1(_0580_),
    .S(_0473_),
    .X(_0581_));
 sg13g2_a221oi_1 _1371_ (.B2(_0581_),
    .C1(_0502_),
    .B1(_0574_),
    .A1(net2),
    .Y(_0582_),
    .A2(net42));
 sg13g2_buf_1 _1372_ (.A(_0582_),
    .X(_0583_));
 sg13g2_nor2b_1 _1373_ (.A(_0408_),
    .B_N(\DJ8.ir[1] ),
    .Y(_0584_));
 sg13g2_buf_1 _1374_ (.A(_0584_),
    .X(_0585_));
 sg13g2_mux4_1 _1375_ (.S0(_0510_),
    .A0(\DJ8.EF[8] ),
    .A1(\DJ8.ACC[0] ),
    .A2(\DJ8.EF[0] ),
    .A3(\DJ8.REGS.regs[1][0] ),
    .S1(net59),
    .X(_0586_));
 sg13g2_mux4_1 _1376_ (.S0(_0510_),
    .A0(\DJ8.GH[8] ),
    .A1(\DJ8.REGS.regs[2][0] ),
    .A2(\DJ8.GH[0] ),
    .A3(\DJ8.REGS.regs[3][0] ),
    .S1(net59),
    .X(_0587_));
 sg13g2_mux2_1 _1377_ (.A0(_0586_),
    .A1(_0587_),
    .S(_0508_),
    .X(_0588_));
 sg13g2_buf_1 _1378_ (.A(_0588_),
    .X(_0589_));
 sg13g2_nor2_1 _1379_ (.A(_0585_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_a21oi_2 _1380_ (.B1(_0590_),
    .Y(_0591_),
    .A2(_0583_),
    .A1(_0569_));
 sg13g2_nand2_1 _1381_ (.Y(_0592_),
    .A(_0550_),
    .B(_0591_));
 sg13g2_buf_1 _1382_ (.A(\DJ8.ALU.c_in ),
    .X(_0593_));
 sg13g2_inv_1 _1383_ (.Y(_0594_),
    .A(_0593_));
 sg13g2_o21ai_1 _1384_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0550_),
    .A2(_0591_));
 sg13g2_nand2_1 _1385_ (.Y(_0596_),
    .A(_0592_),
    .B(_0595_));
 sg13g2_xnor2_1 _1386_ (.Y(_0597_),
    .A(_0548_),
    .B(_0596_));
 sg13g2_a21o_1 _1387_ (.A2(\DJ8.ACC[0] ),
    .A1(net67),
    .B1(_0549_),
    .X(_0598_));
 sg13g2_buf_2 _1388_ (.A(_0598_),
    .X(_0599_));
 sg13g2_nand2_1 _1389_ (.Y(_0600_),
    .A(_0599_),
    .B(_0591_));
 sg13g2_o21ai_1 _1390_ (.B1(net80),
    .Y(_0601_),
    .A1(_0599_),
    .A2(_0591_));
 sg13g2_nand2_1 _1391_ (.Y(_0602_),
    .A(_0600_),
    .B(_0601_));
 sg13g2_xor2_1 _1392_ (.B(_0602_),
    .A(_0548_),
    .X(_0603_));
 sg13g2_buf_1 _1393_ (.A(_0416_),
    .X(_0604_));
 sg13g2_nor3_1 _1394_ (.A(_0414_),
    .B(net66),
    .C(_0413_),
    .Y(_0605_));
 sg13g2_buf_1 _1395_ (.A(_0605_),
    .X(_0606_));
 sg13g2_nor2_1 _1396_ (.A(_0414_),
    .B(net84),
    .Y(_0607_));
 sg13g2_and2_1 _1397_ (.A(_0547_),
    .B(_0607_),
    .X(_0608_));
 sg13g2_buf_1 _1398_ (.A(\DJ8.ALU.opalu[2] ),
    .X(_0609_));
 sg13g2_o21ai_1 _1399_ (.B1(net79),
    .Y(_0610_),
    .A1(_0544_),
    .A2(_0608_));
 sg13g2_inv_1 _1400_ (.Y(_0611_),
    .A(_0414_));
 sg13g2_nor2_1 _1401_ (.A(_0611_),
    .B(net84),
    .Y(_0612_));
 sg13g2_inv_1 _1402_ (.Y(_0613_),
    .A(net79));
 sg13g2_o21ai_1 _1403_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_0612_),
    .A2(_0606_));
 sg13g2_buf_1 _1404_ (.A(_0412_),
    .X(_0615_));
 sg13g2_nor2_1 _1405_ (.A(net73),
    .B(_0546_),
    .Y(_0616_));
 sg13g2_a21oi_1 _1406_ (.A1(net73),
    .A2(_0541_),
    .Y(_0617_),
    .B1(_0616_));
 sg13g2_nor2_1 _1407_ (.A(net84),
    .B(_0547_),
    .Y(_0618_));
 sg13g2_buf_1 _1408_ (.A(_0414_),
    .X(_0619_));
 sg13g2_o21ai_1 _1409_ (.B1(net72),
    .Y(_0620_),
    .A1(_0617_),
    .A2(_0618_));
 sg13g2_and3_1 _1410_ (.X(_0621_),
    .A(_0610_),
    .B(_0614_),
    .C(_0620_));
 sg13g2_a221oi_1 _1411_ (.B2(net48),
    .C1(_0621_),
    .B1(_0603_),
    .A1(net54),
    .Y(_0622_),
    .A2(_0597_));
 sg13g2_buf_1 _1412_ (.A(_0611_),
    .X(_0623_));
 sg13g2_nor2_2 _1413_ (.A(net66),
    .B(_0413_),
    .Y(_0624_));
 sg13g2_nor2_1 _1414_ (.A(\DJ8.ALU.opalu[2] ),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_nand2_1 _1415_ (.Y(_0626_),
    .A(net65),
    .B(_0625_));
 sg13g2_xnor2_1 _1416_ (.Y(_0627_),
    .A(_0548_),
    .B(_0600_));
 sg13g2_nor2_1 _1417_ (.A(net41),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_buf_1 _1418_ (.A(net67),
    .X(_0629_));
 sg13g2_xor2_1 _1419_ (.B(\DJ8.ir[3] ),
    .A(\DJ8.ir[2] ),
    .X(_0630_));
 sg13g2_and2_1 _1420_ (.A(net56),
    .B(_0630_),
    .X(_0631_));
 sg13g2_buf_1 _1421_ (.A(_0631_),
    .X(_0632_));
 sg13g2_o21ai_1 _1422_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_0622_),
    .A2(_0628_));
 sg13g2_a21oi_1 _1423_ (.A1(net80),
    .A2(_0599_),
    .Y(_0634_),
    .B1(net84));
 sg13g2_nor2_1 _1424_ (.A(net66),
    .B(_0550_),
    .Y(_0635_));
 sg13g2_nand2_1 _1425_ (.Y(_0636_),
    .A(net80),
    .B(_0635_));
 sg13g2_o21ai_1 _1426_ (.B1(_0636_),
    .Y(_0637_),
    .A1(net65),
    .A2(_0634_));
 sg13g2_nor2_1 _1427_ (.A(_0414_),
    .B(net66),
    .Y(_0638_));
 sg13g2_a21oi_1 _1428_ (.A1(net72),
    .A2(_0599_),
    .Y(_0639_),
    .B1(_0638_));
 sg13g2_nand2_1 _1429_ (.Y(_0640_),
    .A(net73),
    .B(_0594_));
 sg13g2_o21ai_1 _1430_ (.B1(_0640_),
    .Y(_0641_),
    .A1(net72),
    .A2(_0624_));
 sg13g2_a221oi_1 _1431_ (.B2(_0550_),
    .C1(_0632_),
    .B1(_0641_),
    .A1(net72),
    .Y(_0642_),
    .A2(_0635_));
 sg13g2_o21ai_1 _1432_ (.B1(_0642_),
    .Y(_0643_),
    .A1(_0613_),
    .A2(_0639_));
 sg13g2_a21oi_1 _1433_ (.A1(net73),
    .A2(_0637_),
    .Y(_0644_),
    .B1(_0643_));
 sg13g2_o21ai_1 _1434_ (.B1(net80),
    .Y(_0645_),
    .A1(net48),
    .A2(net54));
 sg13g2_nor2_1 _1435_ (.A(_0599_),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_o21ai_1 _1436_ (.B1(net65),
    .Y(_0647_),
    .A1(net79),
    .A2(_0594_));
 sg13g2_a221oi_1 _1437_ (.B2(_0624_),
    .C1(_0550_),
    .B1(_0647_),
    .A1(_0612_),
    .Y(_0648_),
    .A2(_0640_));
 sg13g2_nor4_1 _1438_ (.A(_0632_),
    .B(_0591_),
    .C(_0646_),
    .D(_0648_),
    .Y(_0649_));
 sg13g2_a21oi_1 _1439_ (.A1(_0591_),
    .A2(_0644_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_and2_1 _1440_ (.A(_0633_),
    .B(_0650_),
    .X(_0651_));
 sg13g2_buf_2 _1441_ (.A(_0651_),
    .X(_0652_));
 sg13g2_buf_1 _1442_ (.A(\DJ8.REGS.write_addr[0] ),
    .X(_0653_));
 sg13g2_buf_1 _1443_ (.A(\DJ8.REGS.write_addr[1] ),
    .X(_0654_));
 sg13g2_nand2_2 _1444_ (.Y(_0655_),
    .A(_0409_),
    .B(\DJ8.state[1] ));
 sg13g2_a21oi_1 _1445_ (.A1(_0629_),
    .A2(_0407_),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_nand2b_1 _1446_ (.Y(_0657_),
    .B(_0656_),
    .A_N(\DJ8.REGS.write_addr[2] ));
 sg13g2_buf_2 _1447_ (.A(_0657_),
    .X(_0658_));
 sg13g2_nor3_2 _1448_ (.A(net78),
    .B(net77),
    .C(_0658_),
    .Y(_0659_));
 sg13g2_mux2_1 _1449_ (.A0(\DJ8.ACC[0] ),
    .A1(_0652_),
    .S(_0659_),
    .X(_0043_));
 sg13g2_buf_1 _1450_ (.A(_0659_),
    .X(_0660_));
 sg13g2_buf_1 _1451_ (.A(_0632_),
    .X(_0661_));
 sg13g2_nand2_1 _1452_ (.Y(_0662_),
    .A(net74),
    .B(_0021_));
 sg13g2_nand2b_1 _1453_ (.Y(_0663_),
    .B(_0022_),
    .A_N(net74));
 sg13g2_and2_1 _1454_ (.A(_0662_),
    .B(_0663_),
    .X(_0664_));
 sg13g2_buf_1 _1455_ (.A(_0664_),
    .X(_0665_));
 sg13g2_nor2_1 _1456_ (.A(_0441_),
    .B(_0452_),
    .Y(_0666_));
 sg13g2_nor3_1 _1457_ (.A(net75),
    .B(_0443_),
    .C(_0450_),
    .Y(_0667_));
 sg13g2_a21o_1 _1458_ (.A2(_0666_),
    .A1(net75),
    .B1(_0667_),
    .X(_0668_));
 sg13g2_and2_1 _1459_ (.A(_0456_),
    .B(_0552_),
    .X(_0669_));
 sg13g2_a221oi_1 _1460_ (.B2(_0466_),
    .C1(_0669_),
    .B1(_0668_),
    .A1(_0458_),
    .Y(_0670_),
    .A2(_0551_));
 sg13g2_nand2_1 _1461_ (.Y(_0671_),
    .A(_0486_),
    .B(_0421_));
 sg13g2_nand2_1 _1462_ (.Y(_0672_),
    .A(_0422_),
    .B(_0420_));
 sg13g2_a21o_1 _1463_ (.A2(_0672_),
    .A1(_0671_),
    .B1(_0426_),
    .X(_0673_));
 sg13g2_mux2_1 _1464_ (.A0(_0670_),
    .A1(_0673_),
    .S(net61),
    .X(_0674_));
 sg13g2_nor2_2 _1465_ (.A(_0482_),
    .B(_0471_),
    .Y(_0675_));
 sg13g2_nor2_1 _1466_ (.A(_0498_),
    .B(_0675_),
    .Y(_0676_));
 sg13g2_nor2_1 _1467_ (.A(_0498_),
    .B(_0473_),
    .Y(_0677_));
 sg13g2_xor2_1 _1468_ (.B(_0450_),
    .A(_0443_),
    .X(_0678_));
 sg13g2_xor2_1 _1469_ (.B(_0452_),
    .A(_0441_),
    .X(_0679_));
 sg13g2_mux2_1 _1470_ (.A0(_0678_),
    .A1(_0679_),
    .S(net68),
    .X(_0680_));
 sg13g2_nand2_1 _1471_ (.Y(_0681_),
    .A(_0466_),
    .B(_0680_));
 sg13g2_xor2_1 _1472_ (.B(_0422_),
    .A(_0006_),
    .X(_0682_));
 sg13g2_nand2_1 _1473_ (.Y(_0683_),
    .A(_0421_),
    .B(_0682_));
 sg13g2_mux2_1 _1474_ (.A0(_0681_),
    .A1(_0683_),
    .S(net61),
    .X(_0684_));
 sg13g2_o21ai_1 _1475_ (.B1(_0585_),
    .Y(_0685_),
    .A1(net4),
    .A2(net53));
 sg13g2_a221oi_1 _1476_ (.B2(_0684_),
    .C1(_0685_),
    .B1(_0677_),
    .A1(_0674_),
    .Y(_0686_),
    .A2(_0676_));
 sg13g2_nor2_1 _1477_ (.A(_0507_),
    .B(_0514_),
    .Y(_0687_));
 sg13g2_nor2b_1 _1478_ (.A(_0507_),
    .B_N(net59),
    .Y(_0688_));
 sg13g2_a221oi_1 _1479_ (.B2(\DJ8.EF[2] ),
    .C1(_0510_),
    .B1(_0688_),
    .A1(\DJ8.EF[10] ),
    .Y(_0689_),
    .A2(_0687_));
 sg13g2_inv_1 _1480_ (.Y(_0690_),
    .A(_0450_));
 sg13g2_mux2_1 _1481_ (.A0(\DJ8.GH[10] ),
    .A1(_0690_),
    .S(_0515_),
    .X(_0691_));
 sg13g2_nand2_1 _1482_ (.Y(_0692_),
    .A(net60),
    .B(_0691_));
 sg13g2_mux4_1 _1483_ (.S0(_0514_),
    .A0(\DJ8.ACC[2] ),
    .A1(\DJ8.REGS.regs[1][2] ),
    .A2(\DJ8.REGS.regs[2][2] ),
    .A3(\DJ8.REGS.regs[3][2] ),
    .S1(_0507_),
    .X(_0693_));
 sg13g2_nor2_1 _1484_ (.A(_0531_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_a21oi_2 _1485_ (.B1(_0694_),
    .Y(_0695_),
    .A2(_0692_),
    .A1(_0689_));
 sg13g2_and2_1 _1486_ (.A(_0502_),
    .B(_0695_),
    .X(_0696_));
 sg13g2_or3_1 _1487_ (.A(_0665_),
    .B(_0686_),
    .C(_0696_),
    .X(_0697_));
 sg13g2_buf_2 _1488_ (.A(_0697_),
    .X(_0698_));
 sg13g2_o21ai_1 _1489_ (.B1(_0665_),
    .Y(_0699_),
    .A1(_0686_),
    .A2(_0696_));
 sg13g2_nand2_2 _1490_ (.Y(_0700_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_buf_1 _1491_ (.A(_0585_),
    .X(_0701_));
 sg13g2_o21ai_1 _1492_ (.B1(_0550_),
    .Y(_0702_),
    .A1(net55),
    .A2(_0589_));
 sg13g2_o21ai_1 _1493_ (.B1(_0594_),
    .Y(_0703_),
    .A1(net55),
    .A2(_0589_));
 sg13g2_a22oi_1 _1494_ (.Y(_0704_),
    .B1(_0702_),
    .B2(_0703_),
    .A2(_0583_),
    .A1(_0569_));
 sg13g2_o21ai_1 _1495_ (.B1(_0543_),
    .Y(_0705_),
    .A1(net80),
    .A2(_0599_));
 sg13g2_or2_1 _1496_ (.X(_0706_),
    .B(_0705_),
    .A(_0704_));
 sg13g2_nand2_1 _1497_ (.Y(_0707_),
    .A(_0546_),
    .B(_0550_));
 sg13g2_or2_1 _1498_ (.X(_0708_),
    .B(_0707_),
    .A(_0590_));
 sg13g2_a21oi_1 _1499_ (.A1(_0569_),
    .A2(_0583_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_or3_1 _1500_ (.A(net80),
    .B(_0543_),
    .C(_0590_),
    .X(_0710_));
 sg13g2_a21oi_1 _1501_ (.A1(_0569_),
    .A2(_0583_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_nor2_1 _1502_ (.A(net80),
    .B(_0707_),
    .Y(_0712_));
 sg13g2_or4_1 _1503_ (.A(_0541_),
    .B(_0709_),
    .C(_0711_),
    .D(_0712_),
    .X(_0713_));
 sg13g2_nand2_1 _1504_ (.Y(_0714_),
    .A(_0706_),
    .B(_0713_));
 sg13g2_xnor2_1 _1505_ (.Y(_0715_),
    .A(_0700_),
    .B(_0714_));
 sg13g2_nand2_1 _1506_ (.Y(_0716_),
    .A(net54),
    .B(_0715_));
 sg13g2_nand2_2 _1507_ (.Y(_0717_),
    .A(net65),
    .B(_0624_));
 sg13g2_a21oi_1 _1508_ (.A1(_0600_),
    .A2(_0601_),
    .Y(_0718_),
    .B1(_0544_));
 sg13g2_nor4_1 _1509_ (.A(_0547_),
    .B(_0717_),
    .C(_0700_),
    .D(_0718_),
    .Y(_0719_));
 sg13g2_and3_1 _1510_ (.X(_0720_),
    .A(net48),
    .B(_0700_),
    .C(_0718_));
 sg13g2_nand2_1 _1511_ (.Y(_0721_),
    .A(net65),
    .B(net66));
 sg13g2_o21ai_1 _1512_ (.B1(_0698_),
    .Y(_0722_),
    .A1(_0721_),
    .A2(_0699_));
 sg13g2_a21oi_1 _1513_ (.A1(_0417_),
    .A2(_0717_),
    .Y(_0723_),
    .B1(\DJ8.ALU.opalu[2] ));
 sg13g2_a21o_1 _1514_ (.A2(_0722_),
    .A1(_0609_),
    .B1(_0723_),
    .X(_0724_));
 sg13g2_nand2_1 _1515_ (.Y(_0725_),
    .A(net66),
    .B(_0699_));
 sg13g2_or2_1 _1516_ (.X(_0726_),
    .B(_0696_),
    .A(_0686_));
 sg13g2_buf_1 _1517_ (.A(_0726_),
    .X(_0727_));
 sg13g2_mux2_1 _1518_ (.A0(_0665_),
    .A1(_0727_),
    .S(net73),
    .X(_0728_));
 sg13g2_a21oi_1 _1519_ (.A1(_0725_),
    .A2(_0728_),
    .Y(_0729_),
    .B1(net65));
 sg13g2_nand3_1 _1520_ (.B(_0606_),
    .C(_0700_),
    .A(_0547_),
    .Y(_0730_));
 sg13g2_o21ai_1 _1521_ (.B1(_0730_),
    .Y(_0731_),
    .A1(_0724_),
    .A2(_0729_));
 sg13g2_nor3_1 _1522_ (.A(_0719_),
    .B(_0720_),
    .C(_0731_),
    .Y(_0732_));
 sg13g2_a22oi_1 _1523_ (.Y(_0733_),
    .B1(_0574_),
    .B2(_0581_),
    .A2(net42),
    .A1(net2));
 sg13g2_nand4_1 _1524_ (.B(_0546_),
    .C(_0569_),
    .A(net55),
    .Y(_0734_),
    .D(_0733_));
 sg13g2_nor3_1 _1525_ (.A(_0585_),
    .B(_0543_),
    .C(_0589_),
    .Y(_0735_));
 sg13g2_a221oi_1 _1526_ (.B2(_0550_),
    .C1(_0735_),
    .B1(_0546_),
    .A1(_0504_),
    .Y(_0736_),
    .A2(_0540_));
 sg13g2_nand3b_1 _1527_ (.B(_0543_),
    .C(_0599_),
    .Y(_0737_),
    .A_N(_0590_));
 sg13g2_a21oi_1 _1528_ (.A1(_0569_),
    .A2(_0583_),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_a21oi_1 _1529_ (.A1(_0734_),
    .A2(_0736_),
    .Y(_0739_),
    .B1(_0738_));
 sg13g2_xnor2_1 _1530_ (.Y(_0740_),
    .A(_0700_),
    .B(_0739_));
 sg13g2_nor3_2 _1531_ (.A(net79),
    .B(net72),
    .C(_0624_),
    .Y(_0741_));
 sg13g2_a22oi_1 _1532_ (.Y(_0742_),
    .B1(_0740_),
    .B2(_0741_),
    .A2(_0732_),
    .A1(_0716_));
 sg13g2_nor3_1 _1533_ (.A(net37),
    .B(_0622_),
    .C(_0628_),
    .Y(_0743_));
 sg13g2_a21oi_2 _1534_ (.B1(_0743_),
    .Y(_0744_),
    .A2(_0742_),
    .A1(net37));
 sg13g2_nor2_1 _1535_ (.A(\DJ8.ACC[1] ),
    .B(net30),
    .Y(_0745_));
 sg13g2_a21oi_1 _1536_ (.A1(net30),
    .A2(_0744_),
    .Y(_0044_),
    .B1(_0745_));
 sg13g2_nand2_1 _1537_ (.Y(_0746_),
    .A(net56),
    .B(_0630_));
 sg13g2_xnor2_1 _1538_ (.Y(_0747_),
    .A(_0445_),
    .B(_0448_));
 sg13g2_xnor2_1 _1539_ (.Y(_0748_),
    .A(_0440_),
    .B(_0453_));
 sg13g2_mux2_1 _1540_ (.A0(_0747_),
    .A1(_0748_),
    .S(net62),
    .X(_0749_));
 sg13g2_nand3_1 _1541_ (.B(_0668_),
    .C(_0749_),
    .A(_0434_),
    .Y(_0750_));
 sg13g2_nand4_1 _1542_ (.B(_0476_),
    .C(_0429_),
    .A(net61),
    .Y(_0751_),
    .D(_0565_));
 sg13g2_a21oi_1 _1543_ (.A1(_0750_),
    .A2(_0751_),
    .Y(_0752_),
    .B1(_0473_));
 sg13g2_and2_1 _1544_ (.A(_0462_),
    .B(_0572_),
    .X(_0753_));
 sg13g2_nor3_1 _1545_ (.A(_0468_),
    .B(_0484_),
    .C(_0753_),
    .Y(_0754_));
 sg13g2_nor2b_1 _1546_ (.A(net83),
    .B_N(_0420_),
    .Y(_0755_));
 sg13g2_and2_1 _1547_ (.A(_0006_),
    .B(_0422_),
    .X(_0756_));
 sg13g2_a22oi_1 _1548_ (.Y(_0757_),
    .B1(_0756_),
    .B2(_0428_),
    .A2(_0755_),
    .A1(_0422_));
 sg13g2_nand2_1 _1549_ (.Y(_0758_),
    .A(_0006_),
    .B(net83));
 sg13g2_nand2_1 _1550_ (.Y(_0759_),
    .A(_0486_),
    .B(_0758_));
 sg13g2_a21oi_1 _1551_ (.A1(_0757_),
    .A2(_0759_),
    .Y(_0760_),
    .B1(_0434_));
 sg13g2_nand2b_1 _1552_ (.Y(_0761_),
    .B(_0450_),
    .A_N(net68));
 sg13g2_nand2_1 _1553_ (.Y(_0762_),
    .A(net68),
    .B(_0452_));
 sg13g2_nor2b_1 _1554_ (.A(_0445_),
    .B_N(_0448_),
    .Y(_0763_));
 sg13g2_and2_1 _1555_ (.A(_0438_),
    .B(_0453_),
    .X(_0764_));
 sg13g2_a22oi_1 _1556_ (.Y(_0765_),
    .B1(_0764_),
    .B2(_0442_),
    .A2(_0763_),
    .A1(_0444_));
 sg13g2_a221oi_1 _1557_ (.B2(_0765_),
    .C1(net61),
    .B1(_0562_),
    .A1(_0761_),
    .Y(_0766_),
    .A2(_0762_));
 sg13g2_nor4_2 _1558_ (.A(_0675_),
    .B(_0754_),
    .C(_0760_),
    .Y(_0767_),
    .D(_0766_));
 sg13g2_nor2_1 _1559_ (.A(_0502_),
    .B(_0498_),
    .Y(_0768_));
 sg13g2_o21ai_1 _1560_ (.B1(_0768_),
    .Y(_0769_),
    .A1(_0752_),
    .A2(_0767_));
 sg13g2_nand2b_1 _1561_ (.Y(_0770_),
    .B(net52),
    .A_N(\DJ8.REGS.regs[1][3] ));
 sg13g2_a22oi_1 _1562_ (.Y(_0771_),
    .B1(_0511_),
    .B2(_0770_),
    .A2(_0687_),
    .A1(\DJ8.EF[11] ));
 sg13g2_and2_1 _1563_ (.A(net60),
    .B(net59),
    .X(_0772_));
 sg13g2_nand3_1 _1564_ (.B(net57),
    .C(_0772_),
    .A(\DJ8.REGS.regs[3][3] ),
    .Y(_0773_));
 sg13g2_nor2b_1 _1565_ (.A(net85),
    .B_N(_0512_),
    .Y(_0774_));
 sg13g2_a21oi_2 _1566_ (.B1(_0774_),
    .Y(_0775_),
    .A2(net78),
    .A1(net85));
 sg13g2_mux2_1 _1567_ (.A0(\DJ8.GH[11] ),
    .A1(\DJ8.REGS.regs[2][3] ),
    .S(_0510_),
    .X(_0776_));
 sg13g2_nand3_1 _1568_ (.B(_0775_),
    .C(_0776_),
    .A(net58),
    .Y(_0777_));
 sg13g2_mux2_1 _1569_ (.A0(\DJ8.EF[3] ),
    .A1(_0446_),
    .S(_0507_),
    .X(_0778_));
 sg13g2_nand3_1 _1570_ (.B(net52),
    .C(_0778_),
    .A(_0531_),
    .Y(_0779_));
 sg13g2_nand4_1 _1571_ (.B(_0773_),
    .C(_0777_),
    .A(_0771_),
    .Y(_0780_),
    .D(_0779_));
 sg13g2_inv_1 _1572_ (.Y(_0781_),
    .A(\DJ8.ACC[3] ));
 sg13g2_nor2_1 _1573_ (.A(net52),
    .B(_0518_),
    .Y(_0782_));
 sg13g2_a21oi_1 _1574_ (.A1(_0781_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0585_));
 sg13g2_and2_1 _1575_ (.A(net5),
    .B(_0585_),
    .X(_0784_));
 sg13g2_a22oi_1 _1576_ (.Y(_0785_),
    .B1(_0784_),
    .B2(net42),
    .A2(_0783_),
    .A1(_0780_));
 sg13g2_buf_1 _1577_ (.A(net74),
    .X(_0786_));
 sg13g2_and2_1 _1578_ (.A(net64),
    .B(_0023_),
    .X(_0787_));
 sg13g2_a21o_1 _1579_ (.A2(_0024_),
    .A1(net56),
    .B1(_0787_),
    .X(_0788_));
 sg13g2_a21oi_1 _1580_ (.A1(_0769_),
    .A2(_0785_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_nand2_2 _1581_ (.Y(_0790_),
    .A(_0769_),
    .B(_0785_));
 sg13g2_a21oi_2 _1582_ (.B1(_0787_),
    .Y(_0791_),
    .A2(_0024_),
    .A1(net56));
 sg13g2_nor2_1 _1583_ (.A(_0790_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_a21o_1 _1584_ (.A2(_0789_),
    .A1(_0607_),
    .B1(_0792_),
    .X(_0793_));
 sg13g2_mux2_1 _1585_ (.A0(_0790_),
    .A1(_0791_),
    .S(_0413_),
    .X(_0794_));
 sg13g2_o21ai_1 _1586_ (.B1(_0794_),
    .Y(_0795_),
    .A1(net84),
    .A2(_0789_));
 sg13g2_a22oi_1 _1587_ (.Y(_0796_),
    .B1(_0795_),
    .B2(net72),
    .A2(_0793_),
    .A1(net79));
 sg13g2_xnor2_1 _1588_ (.Y(_0797_),
    .A(_0790_),
    .B(_0788_));
 sg13g2_o21ai_1 _1589_ (.B1(_0541_),
    .Y(_0798_),
    .A1(_0704_),
    .A2(_0705_));
 sg13g2_inv_1 _1590_ (.Y(_0799_),
    .A(net4));
 sg13g2_mux4_1 _1591_ (.S0(net50),
    .A0(_0681_),
    .A1(_0683_),
    .A2(_0670_),
    .A3(_0673_),
    .S1(_0473_),
    .X(_0800_));
 sg13g2_mux2_1 _1592_ (.A0(_0799_),
    .A1(_0800_),
    .S(net53),
    .X(_0801_));
 sg13g2_nor2_1 _1593_ (.A(net55),
    .B(_0695_),
    .Y(_0802_));
 sg13g2_a221oi_1 _1594_ (.B2(net55),
    .C1(_0802_),
    .B1(_0801_),
    .A1(_0662_),
    .Y(_0803_),
    .A2(_0663_));
 sg13g2_nor4_1 _1595_ (.A(_0803_),
    .B(_0709_),
    .C(_0711_),
    .D(_0712_),
    .Y(_0804_));
 sg13g2_nand2_2 _1596_ (.Y(_0805_),
    .A(_0662_),
    .B(_0663_));
 sg13g2_nor2_1 _1597_ (.A(_0805_),
    .B(_0727_),
    .Y(_0806_));
 sg13g2_a21oi_1 _1598_ (.A1(_0798_),
    .A2(_0804_),
    .Y(_0807_),
    .B1(_0806_));
 sg13g2_xnor2_1 _1599_ (.Y(_0808_),
    .A(_0797_),
    .B(_0807_));
 sg13g2_a22oi_1 _1600_ (.Y(_0809_),
    .B1(_0808_),
    .B2(_0419_),
    .A2(_0796_),
    .A1(_0614_));
 sg13g2_nor2_1 _1601_ (.A(_0665_),
    .B(_0727_),
    .Y(_0810_));
 sg13g2_a221oi_1 _1602_ (.B2(_0736_),
    .C1(_0738_),
    .B1(_0734_),
    .A1(_0665_),
    .Y(_0811_),
    .A2(_0727_));
 sg13g2_o21ai_1 _1603_ (.B1(_0797_),
    .Y(_0812_),
    .A1(_0810_),
    .A2(_0811_));
 sg13g2_or3_1 _1604_ (.A(_0810_),
    .B(_0797_),
    .C(_0811_),
    .X(_0813_));
 sg13g2_xnor2_1 _1605_ (.Y(_0814_),
    .A(_0599_),
    .B(_0591_));
 sg13g2_nand3_1 _1606_ (.B(_0698_),
    .C(_0699_),
    .A(net80),
    .Y(_0815_));
 sg13g2_or4_1 _1607_ (.A(_0544_),
    .B(_0547_),
    .C(_0814_),
    .D(_0815_),
    .X(_0816_));
 sg13g2_a21oi_2 _1608_ (.B1(_0816_),
    .Y(_0817_),
    .A2(_0813_),
    .A1(_0812_));
 sg13g2_nand3_1 _1609_ (.B(_0813_),
    .C(_0816_),
    .A(_0812_),
    .Y(_0818_));
 sg13g2_nand3b_1 _1610_ (.B(_0818_),
    .C(net48),
    .Y(_0819_),
    .A_N(_0817_));
 sg13g2_nand2_1 _1611_ (.Y(_0820_),
    .A(_0812_),
    .B(_0813_));
 sg13g2_o21ai_1 _1612_ (.B1(_0632_),
    .Y(_0821_),
    .A1(net41),
    .A2(_0820_));
 sg13g2_a21oi_1 _1613_ (.A1(_0809_),
    .A2(_0819_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_a21oi_1 _1614_ (.A1(_0746_),
    .A2(_0742_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_nor2_1 _1615_ (.A(\DJ8.ACC[2] ),
    .B(net30),
    .Y(_0824_));
 sg13g2_a21oi_1 _1616_ (.A1(net30),
    .A2(net26),
    .Y(_0045_),
    .B1(_0824_));
 sg13g2_and2_1 _1617_ (.A(_0786_),
    .B(_0005_),
    .X(_0825_));
 sg13g2_a21o_1 _1618_ (.A2(_0025_),
    .A1(net56),
    .B1(_0825_),
    .X(_0826_));
 sg13g2_buf_2 _1619_ (.A(_0826_),
    .X(_0827_));
 sg13g2_nor2_1 _1620_ (.A(net49),
    .B(_0671_),
    .Y(_0828_));
 sg13g2_and3_1 _1621_ (.X(_0829_),
    .A(net49),
    .B(_0466_),
    .C(_0553_));
 sg13g2_o21ai_1 _1622_ (.B1(_0675_),
    .Y(_0830_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_and2_1 _1623_ (.A(_0426_),
    .B(net83),
    .X(_0831_));
 sg13g2_mux2_1 _1624_ (.A0(_0831_),
    .A1(_0753_),
    .S(_0564_),
    .X(_0832_));
 sg13g2_o21ai_1 _1625_ (.B1(_0578_),
    .Y(_0833_),
    .A1(_0473_),
    .A2(_0832_));
 sg13g2_nand2b_1 _1626_ (.Y(_0834_),
    .B(_0462_),
    .A_N(_0572_));
 sg13g2_a21oi_1 _1627_ (.A1(_0471_),
    .A2(_0834_),
    .Y(_0835_),
    .B1(_0482_));
 sg13g2_nor3_1 _1628_ (.A(_0483_),
    .B(_0556_),
    .C(_0423_),
    .Y(_0836_));
 sg13g2_or3_1 _1629_ (.A(_0580_),
    .B(_0835_),
    .C(_0836_),
    .X(_0837_));
 sg13g2_nand4_1 _1630_ (.B(_0830_),
    .C(_0833_),
    .A(_0768_),
    .Y(_0838_),
    .D(_0837_));
 sg13g2_mux4_1 _1631_ (.S0(net59),
    .A0(\DJ8.EF[12] ),
    .A1(\DJ8.EF[4] ),
    .A2(\DJ8.GH[12] ),
    .A3(_0449_),
    .S1(_0508_),
    .X(_0839_));
 sg13g2_nand2b_1 _1632_ (.Y(_0840_),
    .B(_0531_),
    .A_N(_0839_));
 sg13g2_inv_1 _1633_ (.Y(_0841_),
    .A(\DJ8.REGS.regs[1][4] ));
 sg13g2_o21ai_1 _1634_ (.B1(_0510_),
    .Y(_0842_),
    .A1(_0841_),
    .A2(net60));
 sg13g2_nor2b_1 _1635_ (.A(\DJ8.REGS.regs[2][4] ),
    .B_N(\DJ8.REGS.write_addr[1] ),
    .Y(_0843_));
 sg13g2_nand2b_1 _1636_ (.Y(_0844_),
    .B(net74),
    .A_N(\DJ8.REGS.write_addr[0] ));
 sg13g2_nand4_1 _1637_ (.B(\DJ8.REGS.write_addr[0] ),
    .C(net77),
    .A(net74),
    .Y(_0845_),
    .D(\DJ8.REGS.regs[3][4] ));
 sg13g2_o21ai_1 _1638_ (.B1(_0845_),
    .Y(_0846_),
    .A1(_0843_),
    .A2(_0844_));
 sg13g2_nor2b_1 _1639_ (.A(\DJ8.REGS.regs[2][4] ),
    .B_N(_0505_),
    .Y(_0847_));
 sg13g2_nor3_1 _1640_ (.A(net74),
    .B(_0512_),
    .C(_0847_),
    .Y(_0848_));
 sg13g2_and3_1 _1641_ (.X(_0849_),
    .A(_0505_),
    .B(\DJ8.REGS.regs[3][4] ),
    .C(_0774_));
 sg13g2_or4_1 _1642_ (.A(_0842_),
    .B(_0846_),
    .C(_0848_),
    .D(_0849_),
    .X(_0850_));
 sg13g2_nand3_1 _1643_ (.B(_0535_),
    .C(_0687_),
    .A(_0025_),
    .Y(_0851_));
 sg13g2_nand3_1 _1644_ (.B(_0850_),
    .C(_0851_),
    .A(_0840_),
    .Y(_0852_));
 sg13g2_nor2_1 _1645_ (.A(net6),
    .B(_0502_),
    .Y(_0853_));
 sg13g2_a22oi_1 _1646_ (.Y(_0854_),
    .B1(_0853_),
    .B2(_0499_),
    .A2(_0852_),
    .A1(net51));
 sg13g2_nand2_1 _1647_ (.Y(_0855_),
    .A(_0838_),
    .B(_0854_));
 sg13g2_xnor2_1 _1648_ (.Y(_0856_),
    .A(_0827_),
    .B(_0855_));
 sg13g2_nand3_1 _1649_ (.B(_0734_),
    .C(_0736_),
    .A(_0698_),
    .Y(_0857_));
 sg13g2_nor2_1 _1650_ (.A(net55),
    .B(_0805_),
    .Y(_0858_));
 sg13g2_nor2_1 _1651_ (.A(_0502_),
    .B(_0805_),
    .Y(_0859_));
 sg13g2_o21ai_1 _1652_ (.B1(_0859_),
    .Y(_0860_),
    .A1(net4),
    .A2(net53));
 sg13g2_a221oi_1 _1653_ (.B2(_0684_),
    .C1(_0860_),
    .B1(_0677_),
    .A1(_0674_),
    .Y(_0861_),
    .A2(_0676_));
 sg13g2_a21o_1 _1654_ (.A2(_0858_),
    .A1(_0695_),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_a221oi_1 _1655_ (.B2(_0791_),
    .C1(_0862_),
    .B1(_0790_),
    .A1(_0698_),
    .Y(_0863_),
    .A2(_0738_));
 sg13g2_a21o_1 _1656_ (.A2(_0863_),
    .A1(_0857_),
    .B1(_0792_),
    .X(_0864_));
 sg13g2_xor2_1 _1657_ (.B(_0864_),
    .A(_0856_),
    .X(_0865_));
 sg13g2_nor2_1 _1658_ (.A(net41),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_nand2_1 _1659_ (.Y(_0867_),
    .A(_0817_),
    .B(_0865_));
 sg13g2_a21oi_1 _1660_ (.A1(_0769_),
    .A2(_0785_),
    .Y(_0868_),
    .B1(_0791_));
 sg13g2_or2_1 _1661_ (.X(_0869_),
    .B(_0868_),
    .A(_0803_));
 sg13g2_a21o_1 _1662_ (.A2(_0713_),
    .A1(_0706_),
    .B1(_0869_),
    .X(_0870_));
 sg13g2_nand3_1 _1663_ (.B(_0785_),
    .C(_0791_),
    .A(_0769_),
    .Y(_0871_));
 sg13g2_or3_1 _1664_ (.A(_0805_),
    .B(_0686_),
    .C(_0696_),
    .X(_0872_));
 sg13g2_or2_1 _1665_ (.X(_0873_),
    .B(_0868_),
    .A(_0872_));
 sg13g2_and2_1 _1666_ (.A(_0871_),
    .B(_0873_),
    .X(_0874_));
 sg13g2_nand2_1 _1667_ (.Y(_0875_),
    .A(_0870_),
    .B(_0874_));
 sg13g2_xnor2_1 _1668_ (.Y(_0876_),
    .A(_0856_),
    .B(_0875_));
 sg13g2_a21oi_1 _1669_ (.A1(net56),
    .A2(_0025_),
    .Y(_0877_),
    .B1(_0825_));
 sg13g2_and2_1 _1670_ (.A(_0838_),
    .B(_0854_),
    .X(_0878_));
 sg13g2_buf_2 _1671_ (.A(_0878_),
    .X(_0879_));
 sg13g2_nand2_1 _1672_ (.Y(_0880_),
    .A(_0877_),
    .B(_0879_));
 sg13g2_nand2_1 _1673_ (.Y(_0881_),
    .A(_0827_),
    .B(_0855_));
 sg13g2_o21ai_1 _1674_ (.B1(_0881_),
    .Y(_0882_),
    .A1(_0721_),
    .A2(_0880_));
 sg13g2_nor2_1 _1675_ (.A(_0615_),
    .B(_0827_),
    .Y(_0883_));
 sg13g2_a21oi_1 _1676_ (.A1(_0615_),
    .A2(_0879_),
    .Y(_0884_),
    .B1(_0883_));
 sg13g2_a21o_1 _1677_ (.A2(_0880_),
    .A1(net66),
    .B1(_0884_),
    .X(_0885_));
 sg13g2_a221oi_1 _1678_ (.B2(net72),
    .C1(_0723_),
    .B1(_0885_),
    .A1(net79),
    .Y(_0886_),
    .A2(_0882_));
 sg13g2_a221oi_1 _1679_ (.B2(net54),
    .C1(_0886_),
    .B1(_0876_),
    .A1(net48),
    .Y(_0887_),
    .A2(_0867_));
 sg13g2_or3_1 _1680_ (.A(_0817_),
    .B(_0865_),
    .C(_0886_),
    .X(_0888_));
 sg13g2_a21oi_1 _1681_ (.A1(net54),
    .A2(_0876_),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_nor3_1 _1682_ (.A(_0866_),
    .B(_0887_),
    .C(_0889_),
    .Y(_0890_));
 sg13g2_o21ai_1 _1683_ (.B1(_0746_),
    .Y(_0891_),
    .A1(net41),
    .A2(_0820_));
 sg13g2_a21oi_1 _1684_ (.A1(_0809_),
    .A2(_0819_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_a21oi_2 _1685_ (.B1(_0892_),
    .Y(_0893_),
    .A2(_0890_),
    .A1(_0661_));
 sg13g2_nor2_1 _1686_ (.A(\DJ8.ACC[3] ),
    .B(_0660_),
    .Y(_0894_));
 sg13g2_a21oi_1 _1687_ (.A1(net30),
    .A2(_0893_),
    .Y(_0046_),
    .B1(_0894_));
 sg13g2_nand3_1 _1688_ (.B(_0785_),
    .C(_0788_),
    .A(_0769_),
    .Y(_0895_));
 sg13g2_nand2_1 _1689_ (.Y(_0896_),
    .A(_0895_),
    .B(_0877_));
 sg13g2_a21oi_1 _1690_ (.A1(_0857_),
    .A2(_0863_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_nand3_1 _1691_ (.B(_0895_),
    .C(_0879_),
    .A(_0698_),
    .Y(_0898_));
 sg13g2_o21ai_1 _1692_ (.B1(_0879_),
    .Y(_0899_),
    .A1(_0789_),
    .A2(_0877_));
 sg13g2_o21ai_1 _1693_ (.B1(_0899_),
    .Y(_0900_),
    .A1(_0811_),
    .A2(_0898_));
 sg13g2_a22oi_1 _1694_ (.Y(_0901_),
    .B1(_0552_),
    .B2(_0456_),
    .A2(_0551_),
    .A1(_0458_));
 sg13g2_nor2_1 _1695_ (.A(net50),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_nor3_1 _1696_ (.A(net82),
    .B(net49),
    .C(_0672_),
    .Y(_0903_));
 sg13g2_o21ai_1 _1697_ (.B1(_0675_),
    .Y(_0904_),
    .A1(_0902_),
    .A2(_0903_));
 sg13g2_buf_1 _1698_ (.A(net49),
    .X(_0905_));
 sg13g2_a21oi_1 _1699_ (.A1(net82),
    .A2(_0475_),
    .Y(_0906_),
    .B1(net49));
 sg13g2_a21o_1 _1700_ (.A2(_0447_),
    .A1(net40),
    .B1(_0906_),
    .X(_0907_));
 sg13g2_mux2_1 _1701_ (.A0(_0423_),
    .A1(_0572_),
    .S(net49),
    .X(_0908_));
 sg13g2_a21o_1 _1702_ (.A2(_0907_),
    .A1(_0904_),
    .B1(_0908_),
    .X(_0909_));
 sg13g2_buf_1 _1703_ (.A(_0909_),
    .X(_0910_));
 sg13g2_mux2_1 _1704_ (.A0(_0421_),
    .A1(_0466_),
    .S(net63),
    .X(_0911_));
 sg13g2_nor2_1 _1705_ (.A(_0557_),
    .B(_0553_),
    .Y(_0912_));
 sg13g2_nand2_1 _1706_ (.Y(_0913_),
    .A(_0572_),
    .B(_0575_));
 sg13g2_mux2_1 _1707_ (.A0(_0424_),
    .A1(_0913_),
    .S(net63),
    .X(_0914_));
 sg13g2_mux4_1 _1708_ (.S0(net49),
    .A0(_0756_),
    .A1(_0912_),
    .A2(_0429_),
    .A3(_0668_),
    .S1(_0914_),
    .X(_0915_));
 sg13g2_o21ai_1 _1709_ (.B1(_0473_),
    .Y(_0916_),
    .A1(_0911_),
    .A2(_0915_));
 sg13g2_and2_1 _1710_ (.A(net64),
    .B(_0026_),
    .X(_0917_));
 sg13g2_a21o_1 _1711_ (.A2(_0027_),
    .A1(_0501_),
    .B1(_0917_),
    .X(_0918_));
 sg13g2_buf_2 _1712_ (.A(_0918_),
    .X(_0919_));
 sg13g2_nor2_1 _1713_ (.A(net51),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nand2_1 _1714_ (.Y(_0921_),
    .A(net53),
    .B(_0920_));
 sg13g2_a21o_1 _1715_ (.A2(_0916_),
    .A1(_0910_),
    .B1(_0921_),
    .X(_0922_));
 sg13g2_mux2_1 _1716_ (.A0(\DJ8.EF[13] ),
    .A1(\DJ8.GH[13] ),
    .S(net58),
    .X(_0923_));
 sg13g2_a22oi_1 _1717_ (.Y(_0924_),
    .B1(_0923_),
    .B2(_0775_),
    .A2(_0688_),
    .A1(\DJ8.EF[5] ));
 sg13g2_mux2_1 _1718_ (.A0(\DJ8.ACC[5] ),
    .A1(\DJ8.REGS.regs[2][5] ),
    .S(net58),
    .X(_0925_));
 sg13g2_a221oi_1 _1719_ (.B2(_0775_),
    .C1(_0531_),
    .B1(_0925_),
    .A1(\DJ8.REGS.regs[3][5] ),
    .Y(_0926_),
    .A2(_0772_));
 sg13g2_a21o_1 _1720_ (.A2(_0924_),
    .A1(_0531_),
    .B1(_0926_),
    .X(_0927_));
 sg13g2_nor2b_1 _1721_ (.A(net57),
    .B_N(net58),
    .Y(_0928_));
 sg13g2_a22oi_1 _1722_ (.Y(_0929_),
    .B1(_0928_),
    .B2(\DJ8.GH[5] ),
    .A2(_0511_),
    .A1(\DJ8.REGS.regs[1][5] ));
 sg13g2_or2_1 _1723_ (.X(_0930_),
    .B(_0929_),
    .A(_0775_));
 sg13g2_nand2_1 _1724_ (.Y(_0931_),
    .A(_0927_),
    .B(_0930_));
 sg13g2_nor2_1 _1725_ (.A(net55),
    .B(_0919_),
    .Y(_0932_));
 sg13g2_a21oi_2 _1726_ (.B1(_0917_),
    .Y(_0933_),
    .A2(_0027_),
    .A1(net56));
 sg13g2_and3_1 _1727_ (.X(_0934_),
    .A(net7),
    .B(_0701_),
    .C(_0933_));
 sg13g2_buf_1 _1728_ (.A(_0499_),
    .X(_0935_));
 sg13g2_a22oi_1 _1729_ (.Y(_0936_),
    .B1(_0934_),
    .B2(net36),
    .A2(_0932_),
    .A1(_0931_));
 sg13g2_nor3_1 _1730_ (.A(net51),
    .B(net36),
    .C(_0933_),
    .Y(_0937_));
 sg13g2_nand3_1 _1731_ (.B(_0916_),
    .C(_0937_),
    .A(_0910_),
    .Y(_0938_));
 sg13g2_and2_1 _1732_ (.A(_0927_),
    .B(_0930_),
    .X(_0939_));
 sg13g2_nor2_1 _1733_ (.A(_0701_),
    .B(_0933_),
    .Y(_0940_));
 sg13g2_nor3_1 _1734_ (.A(net7),
    .B(net51),
    .C(_0933_),
    .Y(_0941_));
 sg13g2_a22oi_1 _1735_ (.Y(_0942_),
    .B1(_0941_),
    .B2(net36),
    .A2(_0940_),
    .A1(_0939_));
 sg13g2_and4_1 _1736_ (.A(_0922_),
    .B(_0936_),
    .C(_0938_),
    .D(_0942_),
    .X(_0943_));
 sg13g2_buf_2 _1737_ (.A(_0943_),
    .X(_0944_));
 sg13g2_o21ai_1 _1738_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0897_),
    .A2(_0900_));
 sg13g2_or3_1 _1739_ (.A(_0944_),
    .B(_0897_),
    .C(_0900_),
    .X(_0946_));
 sg13g2_nand2_1 _1740_ (.Y(_0947_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_nand4_1 _1741_ (.B(_0936_),
    .C(_0938_),
    .A(_0922_),
    .Y(_0948_),
    .D(_0942_));
 sg13g2_buf_1 _1742_ (.A(_0948_),
    .X(_0949_));
 sg13g2_nor2_1 _1743_ (.A(net84),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_o21ai_1 _1744_ (.B1(net65),
    .Y(_0951_),
    .A1(_0625_),
    .A2(_0950_));
 sg13g2_nand3_1 _1745_ (.B(_0910_),
    .C(_0916_),
    .A(_0768_),
    .Y(_0952_));
 sg13g2_nor2_1 _1746_ (.A(net7),
    .B(net51),
    .Y(_0953_));
 sg13g2_a22oi_1 _1747_ (.Y(_0954_),
    .B1(_0953_),
    .B2(net36),
    .A2(_0939_),
    .A1(_0539_));
 sg13g2_nand2_1 _1748_ (.Y(_0955_),
    .A(_0952_),
    .B(_0954_));
 sg13g2_a21oi_1 _1749_ (.A1(net72),
    .A2(_0933_),
    .Y(_0956_),
    .B1(_0638_));
 sg13g2_nand2_1 _1750_ (.Y(_0957_),
    .A(_0638_),
    .B(_0933_));
 sg13g2_o21ai_1 _1751_ (.B1(_0957_),
    .Y(_0958_),
    .A1(_0955_),
    .A2(_0956_));
 sg13g2_nor2_1 _1752_ (.A(_0623_),
    .B(net66),
    .Y(_0959_));
 sg13g2_nand3_1 _1753_ (.B(_0952_),
    .C(_0954_),
    .A(net73),
    .Y(_0960_));
 sg13g2_o21ai_1 _1754_ (.B1(_0960_),
    .Y(_0961_),
    .A1(net73),
    .A2(_0919_));
 sg13g2_a22oi_1 _1755_ (.Y(_0962_),
    .B1(_0959_),
    .B2(_0961_),
    .A2(_0958_),
    .A1(net79));
 sg13g2_nor2_2 _1756_ (.A(_0827_),
    .B(_0879_),
    .Y(_0963_));
 sg13g2_xnor2_1 _1757_ (.Y(_0964_),
    .A(_0949_),
    .B(_0963_));
 sg13g2_nand4_1 _1758_ (.B(_0870_),
    .C(_0874_),
    .A(_0419_),
    .Y(_0965_),
    .D(_0964_));
 sg13g2_and3_1 _1759_ (.X(_0966_),
    .A(_0951_),
    .B(_0962_),
    .C(_0965_));
 sg13g2_nand2_2 _1760_ (.Y(_0967_),
    .A(_0412_),
    .B(_0612_));
 sg13g2_nor2_1 _1761_ (.A(_0967_),
    .B(_0856_),
    .Y(_0968_));
 sg13g2_nand2_1 _1762_ (.Y(_0969_),
    .A(_0418_),
    .B(_0856_));
 sg13g2_nor2_1 _1763_ (.A(_0964_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_a22oi_1 _1764_ (.Y(_0971_),
    .B1(_0970_),
    .B2(_0875_),
    .A2(_0968_),
    .A1(_0964_));
 sg13g2_and4_1 _1765_ (.A(_0867_),
    .B(_0947_),
    .C(_0966_),
    .D(_0971_),
    .X(_0972_));
 sg13g2_and2_1 _1766_ (.A(_0945_),
    .B(_0946_),
    .X(_0973_));
 sg13g2_nor2_1 _1767_ (.A(net41),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_a21o_1 _1768_ (.A2(_0879_),
    .A1(_0827_),
    .B1(_0868_),
    .X(_0975_));
 sg13g2_a221oi_1 _1769_ (.B2(_0713_),
    .C1(_0975_),
    .B1(_0706_),
    .A1(_0805_),
    .Y(_0976_),
    .A2(_0727_));
 sg13g2_a21o_1 _1770_ (.A2(_0879_),
    .A1(_0827_),
    .B1(_0871_),
    .X(_0977_));
 sg13g2_o21ai_1 _1771_ (.B1(_0977_),
    .Y(_0978_),
    .A1(_0872_),
    .A2(_0975_));
 sg13g2_nor3_2 _1772_ (.A(_0963_),
    .B(_0976_),
    .C(_0978_),
    .Y(_0979_));
 sg13g2_xnor2_1 _1773_ (.Y(_0980_),
    .A(_0944_),
    .B(_0979_));
 sg13g2_nand4_1 _1774_ (.B(_0865_),
    .C(_0945_),
    .A(_0817_),
    .Y(_0981_),
    .D(_0946_));
 sg13g2_nand2_1 _1775_ (.Y(_0982_),
    .A(_0951_),
    .B(_0962_));
 sg13g2_a221oi_1 _1776_ (.B2(net48),
    .C1(_0982_),
    .B1(_0981_),
    .A1(net54),
    .Y(_0983_),
    .A2(_0980_));
 sg13g2_nor3_1 _1777_ (.A(_0972_),
    .B(_0974_),
    .C(_0983_),
    .Y(_0984_));
 sg13g2_nor4_1 _1778_ (.A(net37),
    .B(_0866_),
    .C(_0887_),
    .D(_0889_),
    .Y(_0985_));
 sg13g2_a21oi_2 _1779_ (.B1(_0985_),
    .Y(_0986_),
    .A2(_0984_),
    .A1(net37));
 sg13g2_nor2_1 _1780_ (.A(\DJ8.ACC[4] ),
    .B(_0659_),
    .Y(_0987_));
 sg13g2_a21oi_1 _1781_ (.A1(net30),
    .A2(_0986_),
    .Y(_0047_),
    .B1(_0987_));
 sg13g2_mux2_1 _1782_ (.A0(_0029_),
    .A1(_0028_),
    .S(net64),
    .X(_0988_));
 sg13g2_buf_2 _1783_ (.A(_0988_),
    .X(_0989_));
 sg13g2_nand2_1 _1784_ (.Y(_0990_),
    .A(net40),
    .B(_0575_));
 sg13g2_o21ai_1 _1785_ (.B1(_0990_),
    .Y(_0991_),
    .A1(_0475_),
    .A2(_0905_));
 sg13g2_a21o_1 _1786_ (.A2(_0485_),
    .A1(_0481_),
    .B1(_0487_),
    .X(_0992_));
 sg13g2_nor2_1 _1787_ (.A(net62),
    .B(_0443_),
    .Y(_0993_));
 sg13g2_a221oi_1 _1788_ (.B2(_0690_),
    .C1(net81),
    .B1(_0993_),
    .A1(_0439_),
    .Y(_0994_),
    .A2(_0666_));
 sg13g2_nor2_1 _1789_ (.A(_0483_),
    .B(_0429_),
    .Y(_0995_));
 sg13g2_a21oi_1 _1790_ (.A1(_0471_),
    .A2(_0994_),
    .Y(_0996_),
    .B1(_0995_));
 sg13g2_mux2_1 _1791_ (.A0(_0992_),
    .A1(_0996_),
    .S(_0908_),
    .X(_0997_));
 sg13g2_mux4_1 _1792_ (.S0(_0572_),
    .A0(_0458_),
    .A1(_0443_),
    .A2(_0456_),
    .A3(_0441_),
    .S1(_0439_),
    .X(_0998_));
 sg13g2_o21ai_1 _1793_ (.B1(_0758_),
    .Y(_0999_),
    .A1(net82),
    .A2(_0565_));
 sg13g2_mux2_1 _1794_ (.A0(_0998_),
    .A1(_0999_),
    .S(_0559_),
    .X(_1000_));
 sg13g2_a21oi_1 _1795_ (.A1(_0992_),
    .A2(_1000_),
    .Y(_1001_),
    .B1(net42));
 sg13g2_o21ai_1 _1796_ (.B1(_1001_),
    .Y(_1002_),
    .A1(_0991_),
    .A2(_0997_));
 sg13g2_nand2b_1 _1797_ (.Y(_1003_),
    .B(net42),
    .A_N(net8));
 sg13g2_and2_1 _1798_ (.A(net55),
    .B(_1003_),
    .X(_1004_));
 sg13g2_inv_1 _1799_ (.Y(_1005_),
    .A(\DJ8.GH[14] ));
 sg13g2_nor3_1 _1800_ (.A(_1005_),
    .B(net57),
    .C(net52),
    .Y(_1006_));
 sg13g2_and3_1 _1801_ (.X(_1007_),
    .A(\DJ8.REGS.regs[3][6] ),
    .B(net57),
    .C(net52));
 sg13g2_o21ai_1 _1802_ (.B1(net58),
    .Y(_1008_),
    .A1(_1006_),
    .A2(_1007_));
 sg13g2_mux2_1 _1803_ (.A0(\DJ8.EF[6] ),
    .A1(\DJ8.GH[6] ),
    .S(_0524_),
    .X(_1009_));
 sg13g2_nand3_1 _1804_ (.B(net52),
    .C(_1009_),
    .A(_0531_),
    .Y(_1010_));
 sg13g2_nand2_1 _1805_ (.Y(_1011_),
    .A(_0002_),
    .B(\DJ8.REGS.regs[1][6] ));
 sg13g2_nand2b_1 _1806_ (.Y(_1012_),
    .B(net64),
    .A_N(_0654_));
 sg13g2_a21oi_1 _1807_ (.A1(net78),
    .A2(_1011_),
    .Y(_1013_),
    .B1(_1012_));
 sg13g2_nand2_1 _1808_ (.Y(_1014_),
    .A(_0003_),
    .B(\DJ8.REGS.regs[1][6] ));
 sg13g2_or2_1 _1809_ (.X(_1015_),
    .B(_0505_),
    .A(net74));
 sg13g2_a21oi_1 _1810_ (.A1(_0512_),
    .A2(_1014_),
    .Y(_1016_),
    .B1(_1015_));
 sg13g2_or2_1 _1811_ (.X(_1017_),
    .B(_0535_),
    .A(\DJ8.EF[14] ));
 sg13g2_o21ai_1 _1812_ (.B1(_1017_),
    .Y(_1018_),
    .A1(_1013_),
    .A2(_1016_));
 sg13g2_nand4_1 _1813_ (.B(net57),
    .C(net58),
    .A(\DJ8.REGS.regs[2][6] ),
    .Y(_1019_),
    .D(_0775_));
 sg13g2_nand4_1 _1814_ (.B(_1010_),
    .C(_1018_),
    .A(_1008_),
    .Y(_1020_),
    .D(_1019_));
 sg13g2_nand2b_1 _1815_ (.Y(_1021_),
    .B(_0782_),
    .A_N(\DJ8.ACC[6] ));
 sg13g2_and3_1 _1816_ (.X(_1022_),
    .A(net51),
    .B(_1020_),
    .C(_1021_));
 sg13g2_a21oi_2 _1817_ (.B1(_1022_),
    .Y(_1023_),
    .A2(_1004_),
    .A1(_1002_));
 sg13g2_xnor2_1 _1818_ (.Y(_1024_),
    .A(_0989_),
    .B(_1023_));
 sg13g2_nand4_1 _1819_ (.B(_0910_),
    .C(_0916_),
    .A(net53),
    .Y(_1025_),
    .D(_0920_));
 sg13g2_nor3_1 _1820_ (.A(net7),
    .B(_0539_),
    .C(_0919_),
    .Y(_1026_));
 sg13g2_a22oi_1 _1821_ (.Y(_1027_),
    .B1(_1026_),
    .B2(net36),
    .A2(_0932_),
    .A1(_0939_));
 sg13g2_and2_1 _1822_ (.A(_1025_),
    .B(_1027_),
    .X(_1028_));
 sg13g2_buf_1 _1823_ (.A(_1028_),
    .X(_1029_));
 sg13g2_xor2_1 _1824_ (.B(_1029_),
    .A(_1024_),
    .X(_1030_));
 sg13g2_nor3_1 _1825_ (.A(_0967_),
    .B(_0944_),
    .C(_1030_),
    .Y(_1031_));
 sg13g2_xnor2_1 _1826_ (.Y(_1032_),
    .A(_1024_),
    .B(_1029_));
 sg13g2_nor3_1 _1827_ (.A(_0967_),
    .B(_0963_),
    .C(_1032_),
    .Y(_1033_));
 sg13g2_nor2_1 _1828_ (.A(_0976_),
    .B(_0978_),
    .Y(_1034_));
 sg13g2_mux2_1 _1829_ (.A0(_1031_),
    .A1(_1033_),
    .S(_1034_),
    .X(_1035_));
 sg13g2_inv_1 _1830_ (.Y(_1036_),
    .A(_0989_));
 sg13g2_a21o_1 _1831_ (.A2(_1004_),
    .A1(_1002_),
    .B1(_1022_),
    .X(_1037_));
 sg13g2_buf_2 _1832_ (.A(_1037_),
    .X(_1038_));
 sg13g2_nor2_1 _1833_ (.A(_1036_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_nor3_1 _1834_ (.A(_0721_),
    .B(_0989_),
    .C(_1023_),
    .Y(_1040_));
 sg13g2_o21ai_1 _1835_ (.B1(_0609_),
    .Y(_1041_),
    .A1(_1039_),
    .A2(_1040_));
 sg13g2_a21oi_1 _1836_ (.A1(_1036_),
    .A2(_1038_),
    .Y(_1042_),
    .B1(net84));
 sg13g2_nand2_1 _1837_ (.Y(_1043_),
    .A(_0413_),
    .B(_0989_));
 sg13g2_o21ai_1 _1838_ (.B1(_1043_),
    .Y(_1044_),
    .A1(_0413_),
    .A2(_1038_));
 sg13g2_o21ai_1 _1839_ (.B1(_0619_),
    .Y(_1045_),
    .A1(_1042_),
    .A2(_1044_));
 sg13g2_nand3_1 _1840_ (.B(_1041_),
    .C(_1045_),
    .A(_0614_),
    .Y(_1046_));
 sg13g2_nand3_1 _1841_ (.B(_0944_),
    .C(_1030_),
    .A(net54),
    .Y(_1047_));
 sg13g2_nand4_1 _1842_ (.B(_0949_),
    .C(_0963_),
    .A(net54),
    .Y(_1048_),
    .D(_1032_));
 sg13g2_nand3_1 _1843_ (.B(_1047_),
    .C(_1048_),
    .A(_1046_),
    .Y(_1049_));
 sg13g2_o21ai_1 _1844_ (.B1(net41),
    .Y(_1050_),
    .A1(_1035_),
    .A2(_1049_));
 sg13g2_and3_1 _1845_ (.X(_1051_),
    .A(net41),
    .B(_0817_),
    .C(_0865_));
 sg13g2_a221oi_1 _1846_ (.B2(_0863_),
    .C1(_0792_),
    .B1(_0857_),
    .A1(_0827_),
    .Y(_1052_),
    .A2(_0855_));
 sg13g2_o21ai_1 _1847_ (.B1(_0880_),
    .Y(_1053_),
    .A1(_0919_),
    .A2(_0955_));
 sg13g2_nand2_1 _1848_ (.Y(_1054_),
    .A(_0919_),
    .B(_0955_));
 sg13g2_o21ai_1 _1849_ (.B1(_1054_),
    .Y(_1055_),
    .A1(_1052_),
    .A2(_1053_));
 sg13g2_xor2_1 _1850_ (.B(_1055_),
    .A(_1024_),
    .X(_1056_));
 sg13g2_a21oi_1 _1851_ (.A1(_0973_),
    .A2(_1051_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_xnor2_1 _1852_ (.Y(_1058_),
    .A(_1024_),
    .B(_1055_));
 sg13g2_o21ai_1 _1853_ (.B1(net48),
    .Y(_1059_),
    .A1(_0981_),
    .A2(_1058_));
 sg13g2_nor2_1 _1854_ (.A(_1035_),
    .B(_1049_),
    .Y(_1060_));
 sg13g2_a22oi_1 _1855_ (.Y(_1061_),
    .B1(_1059_),
    .B2(_1060_),
    .A2(_1057_),
    .A1(_1050_));
 sg13g2_nor4_1 _1856_ (.A(net37),
    .B(_0972_),
    .C(_0974_),
    .D(_0983_),
    .Y(_1062_));
 sg13g2_a21oi_2 _1857_ (.B1(_1062_),
    .Y(_1063_),
    .A2(_1061_),
    .A1(net37));
 sg13g2_nor2_1 _1858_ (.A(\DJ8.ACC[5] ),
    .B(_0659_),
    .Y(_1064_));
 sg13g2_a21oi_1 _1859_ (.A1(_0660_),
    .A2(_1063_),
    .Y(_0048_),
    .B1(_1064_));
 sg13g2_nand2_1 _1860_ (.Y(_1065_),
    .A(_1036_),
    .B(_1038_));
 sg13g2_a21oi_1 _1861_ (.A1(_0919_),
    .A2(_0955_),
    .Y(_1066_),
    .B1(_1039_));
 sg13g2_o21ai_1 _1862_ (.B1(_1066_),
    .Y(_1067_),
    .A1(_1052_),
    .A2(_1053_));
 sg13g2_and2_1 _1863_ (.A(_1065_),
    .B(_1067_),
    .X(_1068_));
 sg13g2_buf_1 _1864_ (.A(_1068_),
    .X(_1069_));
 sg13g2_inv_1 _1865_ (.Y(_1070_),
    .A(\DJ8.ACC[7] ));
 sg13g2_mux2_1 _1866_ (.A0(_0003_),
    .A1(_1070_),
    .S(net56),
    .X(_1071_));
 sg13g2_buf_1 _1867_ (.A(_1071_),
    .X(_1072_));
 sg13g2_inv_1 _1868_ (.Y(_1073_),
    .A(\DJ8.REGS.regs[2][7] ));
 sg13g2_a21oi_1 _1869_ (.A1(_0505_),
    .A2(_1073_),
    .Y(_1074_),
    .B1(_0512_));
 sg13g2_mux2_1 _1870_ (.A0(\DJ8.REGS.regs[1][7] ),
    .A1(\DJ8.REGS.regs[3][7] ),
    .S(net60),
    .X(_1075_));
 sg13g2_nor2b_1 _1871_ (.A(\DJ8.REGS.regs[2][7] ),
    .B_N(net77),
    .Y(_1076_));
 sg13g2_nor3_1 _1872_ (.A(net67),
    .B(net78),
    .C(_1076_),
    .Y(_1077_));
 sg13g2_a221oi_1 _1873_ (.B2(net52),
    .C1(_1077_),
    .B1(_1075_),
    .A1(net67),
    .Y(_1078_),
    .A2(_1074_));
 sg13g2_mux4_1 _1874_ (.S0(_0522_),
    .A0(\DJ8.EF[15] ),
    .A1(\DJ8.EF[7] ),
    .A2(\DJ8.GH[15] ),
    .A3(\DJ8.GH[7] ),
    .S1(_0524_),
    .X(_1079_));
 sg13g2_nor2_1 _1875_ (.A(net57),
    .B(_1079_),
    .Y(_1080_));
 sg13g2_a221oi_1 _1876_ (.B2(net57),
    .C1(_1080_),
    .B1(_1078_),
    .A1(_1070_),
    .Y(_1081_),
    .A2(_0782_));
 sg13g2_nor2_1 _1877_ (.A(_0585_),
    .B(_1081_),
    .Y(_1082_));
 sg13g2_nand2_1 _1878_ (.Y(_1083_),
    .A(_0462_),
    .B(_0572_));
 sg13g2_mux2_1 _1879_ (.A0(_0758_),
    .A1(_1083_),
    .S(_0564_),
    .X(_1084_));
 sg13g2_o21ai_1 _1880_ (.B1(_1084_),
    .Y(_1085_),
    .A1(_0554_),
    .A2(_0911_));
 sg13g2_a221oi_1 _1881_ (.B2(_1085_),
    .C1(net51),
    .B1(_0676_),
    .A1(net9),
    .Y(_1086_),
    .A2(net42));
 sg13g2_or3_1 _1882_ (.A(_1072_),
    .B(_1082_),
    .C(_1086_),
    .X(_1087_));
 sg13g2_buf_1 _1883_ (.A(_1087_),
    .X(_1088_));
 sg13g2_o21ai_1 _1884_ (.B1(_1072_),
    .Y(_1089_),
    .A1(_1082_),
    .A2(_1086_));
 sg13g2_and2_1 _1885_ (.A(_1088_),
    .B(_1089_),
    .X(_1090_));
 sg13g2_buf_1 _1886_ (.A(_1090_),
    .X(_1091_));
 sg13g2_nor2_1 _1887_ (.A(net41),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_nor2b_1 _1888_ (.A(_1029_),
    .B_N(_1024_),
    .Y(_1093_));
 sg13g2_nor2_1 _1889_ (.A(_0967_),
    .B(_1091_),
    .Y(_1094_));
 sg13g2_a21oi_1 _1890_ (.A1(_1025_),
    .A2(_1027_),
    .Y(_1095_),
    .B1(_1038_));
 sg13g2_nor2_1 _1891_ (.A(_0967_),
    .B(_0989_),
    .Y(_1096_));
 sg13g2_and3_1 _1892_ (.X(_1097_),
    .A(_1088_),
    .B(_1089_),
    .C(_1096_));
 sg13g2_nand2_1 _1893_ (.Y(_1098_),
    .A(_0418_),
    .B(_0989_));
 sg13g2_a21oi_1 _1894_ (.A1(_1088_),
    .A2(_1089_),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_nand3_1 _1895_ (.B(_1025_),
    .C(_1027_),
    .A(_1038_),
    .Y(_1100_));
 sg13g2_a22oi_1 _1896_ (.Y(_1101_),
    .B1(_1099_),
    .B2(_1100_),
    .A2(_1097_),
    .A1(_1095_));
 sg13g2_nand2_1 _1897_ (.Y(_1102_),
    .A(_1088_),
    .B(_1089_));
 sg13g2_nand3_1 _1898_ (.B(_1102_),
    .C(_1096_),
    .A(_1038_),
    .Y(_1103_));
 sg13g2_a21oi_1 _1899_ (.A1(_1101_),
    .A2(_1103_),
    .Y(_1104_),
    .B1(_0944_));
 sg13g2_or3_1 _1900_ (.A(_0963_),
    .B(_0976_),
    .C(_0978_),
    .X(_1105_));
 sg13g2_o21ai_1 _1901_ (.B1(_1089_),
    .Y(_1106_),
    .A1(_0721_),
    .A2(_1088_));
 sg13g2_nor2_1 _1902_ (.A(_1082_),
    .B(_1086_),
    .Y(_1107_));
 sg13g2_nor2_1 _1903_ (.A(_0412_),
    .B(_1072_),
    .Y(_1108_));
 sg13g2_a21oi_1 _1904_ (.A1(net73),
    .A2(_1107_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_a21o_1 _1905_ (.A2(_1088_),
    .A1(_0604_),
    .B1(_1109_),
    .X(_1110_));
 sg13g2_a221oi_1 _1906_ (.B2(_0619_),
    .C1(_0723_),
    .B1(_1110_),
    .A1(net79),
    .Y(_1111_),
    .A2(_1106_));
 sg13g2_a221oi_1 _1907_ (.B2(_1105_),
    .C1(_1111_),
    .B1(_1104_),
    .A1(_1093_),
    .Y(_1112_),
    .A2(_1094_));
 sg13g2_nand2_1 _1908_ (.Y(_1113_),
    .A(_0949_),
    .B(_1032_));
 sg13g2_nand2_1 _1909_ (.Y(_1114_),
    .A(_1036_),
    .B(_1023_));
 sg13g2_or2_1 _1910_ (.X(_1115_),
    .B(_1095_),
    .A(_1036_));
 sg13g2_and2_1 _1911_ (.A(_1091_),
    .B(_1100_),
    .X(_1116_));
 sg13g2_a221oi_1 _1912_ (.B2(_1116_),
    .C1(_0967_),
    .B1(_1115_),
    .A1(_1102_),
    .Y(_1117_),
    .A2(_1114_));
 sg13g2_o21ai_1 _1913_ (.B1(_1117_),
    .Y(_1118_),
    .A1(_0979_),
    .A2(_1113_));
 sg13g2_nand2_1 _1914_ (.Y(_1119_),
    .A(_0741_),
    .B(_1091_));
 sg13g2_a21oi_1 _1915_ (.A1(_1065_),
    .A2(_1067_),
    .Y(_1120_),
    .B1(_1119_));
 sg13g2_a221oi_1 _1916_ (.B2(_1118_),
    .C1(_1120_),
    .B1(_1112_),
    .A1(_1069_),
    .Y(_1121_),
    .A2(_1092_));
 sg13g2_and4_1 _1917_ (.A(_0817_),
    .B(_0865_),
    .C(_0945_),
    .D(_0946_),
    .X(_1122_));
 sg13g2_nand4_1 _1918_ (.B(_1065_),
    .C(_1091_),
    .A(net48),
    .Y(_1123_),
    .D(_1067_));
 sg13g2_a21oi_1 _1919_ (.A1(_1122_),
    .A2(_1056_),
    .Y(_1124_),
    .B1(_1123_));
 sg13g2_nor4_1 _1920_ (.A(_0717_),
    .B(_0981_),
    .C(_1058_),
    .D(_1091_),
    .Y(_1125_));
 sg13g2_nor3_1 _1921_ (.A(_0717_),
    .B(_1091_),
    .C(_1069_),
    .Y(_1126_));
 sg13g2_or4_1 _1922_ (.A(_1121_),
    .B(_1124_),
    .C(_1125_),
    .D(_1126_),
    .X(_1127_));
 sg13g2_a221oi_1 _1923_ (.B2(_1060_),
    .C1(net37),
    .B1(_1059_),
    .A1(_1050_),
    .Y(_1128_),
    .A2(_1057_));
 sg13g2_a21oi_2 _1924_ (.B1(_1128_),
    .Y(_1129_),
    .A2(_1127_),
    .A1(net37));
 sg13g2_nor2_1 _1925_ (.A(\DJ8.ACC[6] ),
    .B(_0659_),
    .Y(_1130_));
 sg13g2_a21oi_1 _1926_ (.A1(net30),
    .A2(_1129_),
    .Y(_0049_),
    .B1(_1130_));
 sg13g2_inv_1 _1927_ (.Y(_0141_),
    .A(\DJ8.ir[2] ));
 sg13g2_nor3_1 _1928_ (.A(net64),
    .B(_0141_),
    .C(\DJ8.ir[3] ),
    .Y(_0142_));
 sg13g2_nor2b_1 _1929_ (.A(_0142_),
    .B_N(_1127_),
    .Y(_0143_));
 sg13g2_buf_2 _1930_ (.A(_0143_),
    .X(_0144_));
 sg13g2_nor2_1 _1931_ (.A(_0031_),
    .B(_0659_),
    .Y(_0145_));
 sg13g2_a21oi_1 _1932_ (.A1(net30),
    .A2(_0144_),
    .Y(_0050_),
    .B1(_0145_));
 sg13g2_nand2b_1 _1933_ (.Y(_0146_),
    .B(net78),
    .A_N(net77));
 sg13g2_nor2_2 _1934_ (.A(_0658_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_mux2_1 _1935_ (.A0(\DJ8.REGS.regs[1][0] ),
    .A1(_0652_),
    .S(_0147_),
    .X(_0051_));
 sg13g2_buf_1 _1936_ (.A(_0147_),
    .X(_0148_));
 sg13g2_nor2_1 _1937_ (.A(\DJ8.REGS.regs[1][1] ),
    .B(net29),
    .Y(_0149_));
 sg13g2_a21oi_1 _1938_ (.A1(_0744_),
    .A2(net29),
    .Y(_0052_),
    .B1(_0149_));
 sg13g2_nor2_1 _1939_ (.A(\DJ8.REGS.regs[1][2] ),
    .B(net29),
    .Y(_0150_));
 sg13g2_a21oi_1 _1940_ (.A1(net26),
    .A2(net29),
    .Y(_0053_),
    .B1(_0150_));
 sg13g2_nor2_1 _1941_ (.A(\DJ8.REGS.regs[1][3] ),
    .B(_0148_),
    .Y(_0151_));
 sg13g2_a21oi_1 _1942_ (.A1(_0893_),
    .A2(net29),
    .Y(_0054_),
    .B1(_0151_));
 sg13g2_nor2_1 _1943_ (.A(\DJ8.REGS.regs[1][4] ),
    .B(_0147_),
    .Y(_0152_));
 sg13g2_a21oi_1 _1944_ (.A1(_0986_),
    .A2(net29),
    .Y(_0055_),
    .B1(_0152_));
 sg13g2_nor2_1 _1945_ (.A(\DJ8.REGS.regs[1][5] ),
    .B(_0147_),
    .Y(_0153_));
 sg13g2_a21oi_1 _1946_ (.A1(_1063_),
    .A2(net29),
    .Y(_0056_),
    .B1(_0153_));
 sg13g2_nor2_1 _1947_ (.A(\DJ8.REGS.regs[1][6] ),
    .B(_0147_),
    .Y(_0154_));
 sg13g2_a21oi_1 _1948_ (.A1(_1129_),
    .A2(net29),
    .Y(_0057_),
    .B1(_0154_));
 sg13g2_nor2_1 _1949_ (.A(_0032_),
    .B(_0147_),
    .Y(_0155_));
 sg13g2_a21oi_1 _1950_ (.A1(_0144_),
    .A2(_0148_),
    .Y(_0058_),
    .B1(_0155_));
 sg13g2_nand2b_1 _1951_ (.Y(_0156_),
    .B(net77),
    .A_N(net78));
 sg13g2_nor2_2 _1952_ (.A(_0658_),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_mux2_1 _1953_ (.A0(\DJ8.REGS.regs[2][0] ),
    .A1(_0652_),
    .S(_0157_),
    .X(_0059_));
 sg13g2_buf_1 _1954_ (.A(_0157_),
    .X(_0158_));
 sg13g2_nor2_1 _1955_ (.A(\DJ8.REGS.regs[2][1] ),
    .B(net28),
    .Y(_0159_));
 sg13g2_a21oi_1 _1956_ (.A1(_0744_),
    .A2(net28),
    .Y(_0060_),
    .B1(_0159_));
 sg13g2_nor2_1 _1957_ (.A(\DJ8.REGS.regs[2][2] ),
    .B(net28),
    .Y(_0160_));
 sg13g2_a21oi_1 _1958_ (.A1(net26),
    .A2(net28),
    .Y(_0061_),
    .B1(_0160_));
 sg13g2_nor2_1 _1959_ (.A(\DJ8.REGS.regs[2][3] ),
    .B(_0158_),
    .Y(_0161_));
 sg13g2_a21oi_1 _1960_ (.A1(_0893_),
    .A2(net28),
    .Y(_0062_),
    .B1(_0161_));
 sg13g2_nor2_1 _1961_ (.A(\DJ8.REGS.regs[2][4] ),
    .B(_0157_),
    .Y(_0162_));
 sg13g2_a21oi_1 _1962_ (.A1(_0986_),
    .A2(net28),
    .Y(_0063_),
    .B1(_0162_));
 sg13g2_nor2_1 _1963_ (.A(\DJ8.REGS.regs[2][5] ),
    .B(_0157_),
    .Y(_0163_));
 sg13g2_a21oi_1 _1964_ (.A1(_1063_),
    .A2(net28),
    .Y(_0064_),
    .B1(_0163_));
 sg13g2_nor2_1 _1965_ (.A(\DJ8.REGS.regs[2][6] ),
    .B(_0157_),
    .Y(_0164_));
 sg13g2_a21oi_1 _1966_ (.A1(_1129_),
    .A2(_0158_),
    .Y(_0065_),
    .B1(_0164_));
 sg13g2_nor2_1 _1967_ (.A(_0033_),
    .B(_0157_),
    .Y(_0165_));
 sg13g2_a21oi_1 _1968_ (.A1(_0144_),
    .A2(net28),
    .Y(_0066_),
    .B1(_0165_));
 sg13g2_nand2_1 _1969_ (.Y(_0166_),
    .A(net78),
    .B(net77));
 sg13g2_nor2_2 _1970_ (.A(_0658_),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_mux2_1 _1971_ (.A0(\DJ8.REGS.regs[3][0] ),
    .A1(_0652_),
    .S(_0167_),
    .X(_0067_));
 sg13g2_buf_1 _1972_ (.A(_0167_),
    .X(_0168_));
 sg13g2_nor2_1 _1973_ (.A(\DJ8.REGS.regs[3][1] ),
    .B(net27),
    .Y(_0169_));
 sg13g2_a21oi_1 _1974_ (.A1(_0744_),
    .A2(net27),
    .Y(_0068_),
    .B1(_0169_));
 sg13g2_nor2_1 _1975_ (.A(\DJ8.REGS.regs[3][2] ),
    .B(net27),
    .Y(_0170_));
 sg13g2_a21oi_1 _1976_ (.A1(net26),
    .A2(net27),
    .Y(_0069_),
    .B1(_0170_));
 sg13g2_nor2_1 _1977_ (.A(\DJ8.REGS.regs[3][3] ),
    .B(net27),
    .Y(_0171_));
 sg13g2_a21oi_1 _1978_ (.A1(_0893_),
    .A2(net27),
    .Y(_0070_),
    .B1(_0171_));
 sg13g2_nor2_1 _1979_ (.A(\DJ8.REGS.regs[3][4] ),
    .B(_0167_),
    .Y(_0172_));
 sg13g2_a21oi_1 _1980_ (.A1(_0986_),
    .A2(_0168_),
    .Y(_0071_),
    .B1(_0172_));
 sg13g2_nor2_1 _1981_ (.A(\DJ8.REGS.regs[3][5] ),
    .B(_0167_),
    .Y(_0173_));
 sg13g2_a21oi_1 _1982_ (.A1(_1063_),
    .A2(_0168_),
    .Y(_0072_),
    .B1(_0173_));
 sg13g2_nor2_1 _1983_ (.A(\DJ8.REGS.regs[3][6] ),
    .B(_0167_),
    .Y(_0174_));
 sg13g2_a21oi_1 _1984_ (.A1(_1129_),
    .A2(net27),
    .Y(_0073_),
    .B1(_0174_));
 sg13g2_nor2_1 _1985_ (.A(_0034_),
    .B(_0167_),
    .Y(_0175_));
 sg13g2_a21oi_1 _1986_ (.A1(_0144_),
    .A2(net27),
    .Y(_0074_),
    .B1(_0175_));
 sg13g2_nand2b_2 _1987_ (.Y(_0176_),
    .B(_0656_),
    .A_N(_0002_));
 sg13g2_nor3_2 _1988_ (.A(net78),
    .B(net77),
    .C(_0176_),
    .Y(_0177_));
 sg13g2_mux2_1 _1989_ (.A0(\DJ8.EF[8] ),
    .A1(_0652_),
    .S(_0177_),
    .X(_0075_));
 sg13g2_buf_1 _1990_ (.A(_0177_),
    .X(_0178_));
 sg13g2_nor2_1 _1991_ (.A(\DJ8.EF[9] ),
    .B(net34),
    .Y(_0179_));
 sg13g2_a21oi_1 _1992_ (.A1(_0744_),
    .A2(net34),
    .Y(_0076_),
    .B1(_0179_));
 sg13g2_nor2_1 _1993_ (.A(\DJ8.EF[10] ),
    .B(net34),
    .Y(_0180_));
 sg13g2_a21oi_1 _1994_ (.A1(net26),
    .A2(net34),
    .Y(_0077_),
    .B1(_0180_));
 sg13g2_nor2_1 _1995_ (.A(\DJ8.EF[11] ),
    .B(net34),
    .Y(_0181_));
 sg13g2_a21oi_1 _1996_ (.A1(_0893_),
    .A2(net34),
    .Y(_0078_),
    .B1(_0181_));
 sg13g2_nor2_1 _1997_ (.A(\DJ8.EF[12] ),
    .B(_0177_),
    .Y(_0182_));
 sg13g2_a21oi_1 _1998_ (.A1(_0986_),
    .A2(net34),
    .Y(_0079_),
    .B1(_0182_));
 sg13g2_nor2_1 _1999_ (.A(\DJ8.EF[13] ),
    .B(_0177_),
    .Y(_0183_));
 sg13g2_a21oi_1 _2000_ (.A1(_1063_),
    .A2(net34),
    .Y(_0080_),
    .B1(_0183_));
 sg13g2_nor2_1 _2001_ (.A(\DJ8.EF[14] ),
    .B(_0177_),
    .Y(_0184_));
 sg13g2_a21oi_1 _2002_ (.A1(_1129_),
    .A2(_0178_),
    .Y(_0081_),
    .B1(_0184_));
 sg13g2_nor2_1 _2003_ (.A(_0035_),
    .B(_0177_),
    .Y(_0185_));
 sg13g2_a21oi_1 _2004_ (.A1(_0144_),
    .A2(_0178_),
    .Y(_0082_),
    .B1(_0185_));
 sg13g2_nor2_2 _2005_ (.A(_0146_),
    .B(_0176_),
    .Y(_0186_));
 sg13g2_mux2_1 _2006_ (.A0(\DJ8.EF[0] ),
    .A1(_0652_),
    .S(_0186_),
    .X(_0083_));
 sg13g2_buf_1 _2007_ (.A(_0186_),
    .X(_0187_));
 sg13g2_nor2_1 _2008_ (.A(\DJ8.EF[1] ),
    .B(net33),
    .Y(_0188_));
 sg13g2_a21oi_1 _2009_ (.A1(_0744_),
    .A2(net33),
    .Y(_0084_),
    .B1(_0188_));
 sg13g2_nor2_1 _2010_ (.A(\DJ8.EF[2] ),
    .B(net33),
    .Y(_0189_));
 sg13g2_a21oi_1 _2011_ (.A1(net26),
    .A2(net33),
    .Y(_0085_),
    .B1(_0189_));
 sg13g2_nor2_1 _2012_ (.A(\DJ8.EF[3] ),
    .B(net33),
    .Y(_0190_));
 sg13g2_a21oi_1 _2013_ (.A1(_0893_),
    .A2(_0187_),
    .Y(_0086_),
    .B1(_0190_));
 sg13g2_nor2_1 _2014_ (.A(\DJ8.EF[4] ),
    .B(_0186_),
    .Y(_0191_));
 sg13g2_a21oi_1 _2015_ (.A1(_0986_),
    .A2(_0187_),
    .Y(_0087_),
    .B1(_0191_));
 sg13g2_nor2_1 _2016_ (.A(\DJ8.EF[5] ),
    .B(_0186_),
    .Y(_0192_));
 sg13g2_a21oi_1 _2017_ (.A1(_1063_),
    .A2(net33),
    .Y(_0088_),
    .B1(_0192_));
 sg13g2_nor2_1 _2018_ (.A(\DJ8.EF[6] ),
    .B(_0186_),
    .Y(_0193_));
 sg13g2_a21oi_1 _2019_ (.A1(_1129_),
    .A2(net33),
    .Y(_0089_),
    .B1(_0193_));
 sg13g2_nor2_1 _2020_ (.A(_0036_),
    .B(_0186_),
    .Y(_0194_));
 sg13g2_a21oi_1 _2021_ (.A1(_0144_),
    .A2(net33),
    .Y(_0090_),
    .B1(_0194_));
 sg13g2_nor2_2 _2022_ (.A(_0156_),
    .B(_0176_),
    .Y(_0195_));
 sg13g2_mux2_1 _2023_ (.A0(\DJ8.GH[8] ),
    .A1(_0652_),
    .S(_0195_),
    .X(_0091_));
 sg13g2_buf_1 _2024_ (.A(_0195_),
    .X(_0196_));
 sg13g2_nor2_1 _2025_ (.A(\DJ8.GH[9] ),
    .B(net32),
    .Y(_0197_));
 sg13g2_a21oi_1 _2026_ (.A1(_0744_),
    .A2(net32),
    .Y(_0092_),
    .B1(_0197_));
 sg13g2_nor2_1 _2027_ (.A(\DJ8.GH[10] ),
    .B(net32),
    .Y(_0198_));
 sg13g2_a21oi_1 _2028_ (.A1(net26),
    .A2(_0196_),
    .Y(_0093_),
    .B1(_0198_));
 sg13g2_nor2_1 _2029_ (.A(\DJ8.GH[11] ),
    .B(net32),
    .Y(_0199_));
 sg13g2_a21oi_1 _2030_ (.A1(_0893_),
    .A2(_0196_),
    .Y(_0094_),
    .B1(_0199_));
 sg13g2_nor2_1 _2031_ (.A(\DJ8.GH[12] ),
    .B(_0195_),
    .Y(_0200_));
 sg13g2_a21oi_1 _2032_ (.A1(_0986_),
    .A2(net32),
    .Y(_0095_),
    .B1(_0200_));
 sg13g2_nor2_1 _2033_ (.A(\DJ8.GH[13] ),
    .B(_0195_),
    .Y(_0201_));
 sg13g2_a21oi_1 _2034_ (.A1(_1063_),
    .A2(net32),
    .Y(_0096_),
    .B1(_0201_));
 sg13g2_nor2_1 _2035_ (.A(\DJ8.GH[14] ),
    .B(_0195_),
    .Y(_0202_));
 sg13g2_a21oi_1 _2036_ (.A1(_1129_),
    .A2(net32),
    .Y(_0097_),
    .B1(_0202_));
 sg13g2_nor2_1 _2037_ (.A(_0037_),
    .B(_0195_),
    .Y(_0203_));
 sg13g2_a21oi_1 _2038_ (.A1(_0144_),
    .A2(net32),
    .Y(_0098_),
    .B1(_0203_));
 sg13g2_nor2_2 _2039_ (.A(_0166_),
    .B(_0176_),
    .Y(_0204_));
 sg13g2_mux2_1 _2040_ (.A0(\DJ8.GH[0] ),
    .A1(_0652_),
    .S(_0204_),
    .X(_0099_));
 sg13g2_buf_1 _2041_ (.A(_0204_),
    .X(_0205_));
 sg13g2_nor2_1 _2042_ (.A(\DJ8.GH[1] ),
    .B(net31),
    .Y(_0206_));
 sg13g2_a21oi_1 _2043_ (.A1(_0744_),
    .A2(net31),
    .Y(_0100_),
    .B1(_0206_));
 sg13g2_nor2_1 _2044_ (.A(\DJ8.GH[2] ),
    .B(net31),
    .Y(_0207_));
 sg13g2_a21oi_1 _2045_ (.A1(_0823_),
    .A2(net31),
    .Y(_0101_),
    .B1(_0207_));
 sg13g2_nor2_1 _2046_ (.A(\DJ8.GH[3] ),
    .B(net31),
    .Y(_0208_));
 sg13g2_a21oi_1 _2047_ (.A1(_0893_),
    .A2(_0205_),
    .Y(_0102_),
    .B1(_0208_));
 sg13g2_nor2_1 _2048_ (.A(\DJ8.GH[4] ),
    .B(_0204_),
    .Y(_0209_));
 sg13g2_a21oi_1 _2049_ (.A1(_0986_),
    .A2(_0205_),
    .Y(_0103_),
    .B1(_0209_));
 sg13g2_nor2_1 _2050_ (.A(\DJ8.GH[5] ),
    .B(_0204_),
    .Y(_0210_));
 sg13g2_a21oi_1 _2051_ (.A1(_1063_),
    .A2(net31),
    .Y(_0104_),
    .B1(_0210_));
 sg13g2_nor2_1 _2052_ (.A(\DJ8.GH[6] ),
    .B(_0204_),
    .Y(_0211_));
 sg13g2_a21oi_1 _2053_ (.A1(_1129_),
    .A2(net31),
    .Y(_0105_),
    .B1(_0211_));
 sg13g2_nor2_1 _2054_ (.A(_0038_),
    .B(_0204_),
    .Y(_0212_));
 sg13g2_a21oi_1 _2055_ (.A1(_0144_),
    .A2(net31),
    .Y(_0106_),
    .B1(_0212_));
 sg13g2_a21oi_1 _2056_ (.A1(_1072_),
    .A2(_1107_),
    .Y(_0213_),
    .B1(_0967_));
 sg13g2_o21ai_1 _2057_ (.B1(_1029_),
    .Y(_0214_),
    .A1(_0944_),
    .A2(_0979_));
 sg13g2_a21oi_1 _2058_ (.A1(_1023_),
    .A2(_0214_),
    .Y(_0215_),
    .B1(_1036_));
 sg13g2_a21oi_1 _2059_ (.A1(_0949_),
    .A2(_1105_),
    .Y(_0216_),
    .B1(_1100_));
 sg13g2_nand2b_1 _2060_ (.Y(_0217_),
    .B(net64),
    .A_N(_0003_));
 sg13g2_o21ai_1 _2061_ (.B1(_0217_),
    .Y(_0218_),
    .A1(net64),
    .A2(_1070_));
 sg13g2_inv_1 _2062_ (.Y(_0219_),
    .A(_1107_));
 sg13g2_nand2_1 _2063_ (.Y(_0220_),
    .A(_0218_),
    .B(_0219_));
 sg13g2_o21ai_1 _2064_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_o21ai_1 _2065_ (.B1(_1072_),
    .Y(_0222_),
    .A1(_0219_),
    .A2(_1069_));
 sg13g2_nand2_1 _2066_ (.Y(_0223_),
    .A(_0219_),
    .B(_1069_));
 sg13g2_nor3_1 _2067_ (.A(_0741_),
    .B(_0981_),
    .C(_1058_),
    .Y(_0224_));
 sg13g2_a21o_1 _2068_ (.A2(_0223_),
    .A1(_0222_),
    .B1(_0224_),
    .X(_0225_));
 sg13g2_nor2_1 _2069_ (.A(_0218_),
    .B(_1107_),
    .Y(_0226_));
 sg13g2_a22oi_1 _2070_ (.Y(_0227_),
    .B1(_0226_),
    .B2(_1069_),
    .A2(_0626_),
    .A1(_0717_));
 sg13g2_a221oi_1 _2071_ (.B2(_0227_),
    .C1(_0655_),
    .B1(_0225_),
    .A1(_0213_),
    .Y(_0228_),
    .A2(_0221_));
 sg13g2_a21oi_1 _2072_ (.A1(_0594_),
    .A2(_0655_),
    .Y(_0107_),
    .B1(_0228_));
 sg13g2_or3_1 _2073_ (.A(_0866_),
    .B(_0887_),
    .C(_0889_),
    .X(_0229_));
 sg13g2_a221oi_1 _2074_ (.B2(_0661_),
    .C1(_0743_),
    .B1(_0742_),
    .A1(_0633_),
    .Y(_0230_),
    .A2(_0650_));
 sg13g2_nor2_1 _2075_ (.A(_0655_),
    .B(_0892_),
    .Y(_0231_));
 sg13g2_nand4_1 _2076_ (.B(_0229_),
    .C(_0230_),
    .A(net26),
    .Y(_0232_),
    .D(_0231_));
 sg13g2_or3_1 _2077_ (.A(_0984_),
    .B(_1061_),
    .C(_1127_),
    .X(_0233_));
 sg13g2_nand2_1 _2078_ (.Y(_0234_),
    .A(\DJ8.flag_Z ),
    .B(_0655_));
 sg13g2_o21ai_1 _2079_ (.B1(_0234_),
    .Y(_0108_),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_buf_1 _2080_ (.A(_0430_),
    .X(_0235_));
 sg13g2_and2_1 _2081_ (.A(_0569_),
    .B(_0733_),
    .X(_0236_));
 sg13g2_nor2_1 _2082_ (.A(_0407_),
    .B(net71),
    .Y(_0237_));
 sg13g2_a21oi_1 _2083_ (.A1(_0235_),
    .A2(_0236_),
    .Y(_0109_),
    .B1(_0237_));
 sg13g2_buf_1 _2084_ (.A(net81),
    .X(_0238_));
 sg13g2_nor2_1 _2085_ (.A(\DJ8.REGS.write_addr[2] ),
    .B(net81),
    .Y(_0239_));
 sg13g2_a21oi_1 _2086_ (.A1(net70),
    .A2(_0801_),
    .Y(_0110_),
    .B1(_0239_));
 sg13g2_nand2_1 _2087_ (.Y(_0240_),
    .A(net5),
    .B(_0935_));
 sg13g2_nand2_1 _2088_ (.Y(_0241_),
    .A(_0493_),
    .B(_0767_));
 sg13g2_a21o_1 _2089_ (.A2(_0241_),
    .A1(_0240_),
    .B1(_0483_),
    .X(_0242_));
 sg13g2_o21ai_1 _2090_ (.B1(_0242_),
    .Y(_0111_),
    .A1(_0238_),
    .A2(_0604_));
 sg13g2_nand3_1 _2091_ (.B(_0833_),
    .C(_0837_),
    .A(_0830_),
    .Y(_0243_));
 sg13g2_mux2_1 _2092_ (.A0(net6),
    .A1(_0243_),
    .S(net53),
    .X(_0244_));
 sg13g2_nand2_1 _2093_ (.Y(_0245_),
    .A(_0238_),
    .B(_0244_));
 sg13g2_o21ai_1 _2094_ (.B1(_0245_),
    .Y(_0112_),
    .A1(_0623_),
    .A2(net70));
 sg13g2_a21oi_1 _2095_ (.A1(_0910_),
    .A2(_0916_),
    .Y(_0246_),
    .B1(_0935_));
 sg13g2_a21o_1 _2096_ (.A2(net36),
    .A1(net7),
    .B1(_0246_),
    .X(_0247_));
 sg13g2_nand2_1 _2097_ (.Y(_0248_),
    .A(net70),
    .B(_0247_));
 sg13g2_o21ai_1 _2098_ (.B1(_0248_),
    .Y(_0113_),
    .A1(_0613_),
    .A2(net70));
 sg13g2_and2_1 _2099_ (.A(_1002_),
    .B(_1003_),
    .X(_0249_));
 sg13g2_nand2_1 _2100_ (.Y(_0250_),
    .A(net70),
    .B(_0249_));
 sg13g2_o21ai_1 _2101_ (.B1(_0250_),
    .Y(_0114_),
    .A1(_0629_),
    .A2(net70));
 sg13g2_a22oi_1 _2102_ (.Y(_0251_),
    .B1(_0676_),
    .B2(_1085_),
    .A2(net36),
    .A1(net9));
 sg13g2_nor2_1 _2103_ (.A(_0409_),
    .B(net81),
    .Y(_0252_));
 sg13g2_a21oi_1 _2104_ (.A1(net70),
    .A2(_0251_),
    .Y(_0115_),
    .B1(_0252_));
 sg13g2_nor2_1 _2105_ (.A(_0474_),
    .B(_0494_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2106_ (.A1(_0495_),
    .A2(net36),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_mux2_1 _2107_ (.A0(\DJ8.ir[1] ),
    .A1(_0254_),
    .S(net71),
    .X(_0116_));
 sg13g2_nor2_1 _2108_ (.A(net71),
    .B(\DJ8.ir[2] ),
    .Y(_0255_));
 sg13g2_a21oi_1 _2109_ (.A1(net71),
    .A2(_0801_),
    .Y(_0117_),
    .B1(_0255_));
 sg13g2_o21ai_1 _2110_ (.B1(net53),
    .Y(_0256_),
    .A1(_0752_),
    .A2(_0767_));
 sg13g2_nand2_1 _2111_ (.Y(_0257_),
    .A(_0240_),
    .B(_0256_));
 sg13g2_mux2_1 _2112_ (.A0(\DJ8.ir[3] ),
    .A1(_0257_),
    .S(net71),
    .X(_0118_));
 sg13g2_buf_1 _2113_ (.A(net62),
    .X(_0258_));
 sg13g2_buf_1 _2114_ (.A(_0258_),
    .X(_0259_));
 sg13g2_mux2_1 _2115_ (.A0(net39),
    .A1(_0244_),
    .S(net71),
    .X(_0119_));
 sg13g2_mux2_1 _2116_ (.A0(_0512_),
    .A1(_0247_),
    .S(net71),
    .X(_0120_));
 sg13g2_mux2_1 _2117_ (.A0(_0505_),
    .A1(_0249_),
    .S(net71),
    .X(_0121_));
 sg13g2_nor2_1 _2118_ (.A(_0430_),
    .B(\DJ8.ir[7] ),
    .Y(_0260_));
 sg13g2_a21oi_1 _2119_ (.A1(_0235_),
    .A2(_0251_),
    .Y(_0122_),
    .B1(_0260_));
 sg13g2_nor2_1 _2120_ (.A(_0653_),
    .B(net81),
    .Y(_0261_));
 sg13g2_a21oi_1 _2121_ (.A1(net70),
    .A2(_0236_),
    .Y(_0123_),
    .B1(_0261_));
 sg13g2_mux2_1 _2122_ (.A0(net77),
    .A1(_0254_),
    .S(net81),
    .X(_0124_));
 sg13g2_nand2b_1 _2123_ (.Y(_0262_),
    .B(net64),
    .A_N(_0409_));
 sg13g2_buf_1 _2124_ (.A(_0262_),
    .X(_0263_));
 sg13g2_mux2_1 _2125_ (.A0(\DJ8.GH[1] ),
    .A1(net82),
    .S(net46),
    .X(_0264_));
 sg13g2_mux2_1 _2126_ (.A0(_0613_),
    .A1(net65),
    .S(\DJ8.flag_Z ),
    .X(_0265_));
 sg13g2_or3_1 _2127_ (.A(_0786_),
    .B(_0409_),
    .C(_0265_),
    .X(_0266_));
 sg13g2_buf_2 _2128_ (.A(_0266_),
    .X(_0267_));
 sg13g2_buf_1 _2129_ (.A(_0267_),
    .X(_0268_));
 sg13g2_mux2_1 _2130_ (.A0(_0407_),
    .A1(_0264_),
    .S(net35),
    .X(_0269_));
 sg13g2_buf_1 _2131_ (.A(\DJ8.state[1] ),
    .X(_0270_));
 sg13g2_buf_1 _2132_ (.A(net76),
    .X(_0271_));
 sg13g2_mux2_1 _2133_ (.A0(\DJ8.pc[0] ),
    .A1(_0269_),
    .S(net69),
    .X(_0125_));
 sg13g2_inv_1 _2134_ (.Y(_0272_),
    .A(\DJ8.pc[10] ));
 sg13g2_buf_1 _2135_ (.A(_0262_),
    .X(_0273_));
 sg13g2_inv_1 _2136_ (.Y(_0274_),
    .A(\DJ8.pc[7] ));
 sg13g2_buf_2 _2137_ (.A(\DJ8.pc[4] ),
    .X(_0275_));
 sg13g2_inv_1 _2138_ (.Y(_0276_),
    .A(\DJ8.pc[3] ));
 sg13g2_nand3_1 _2139_ (.B(\DJ8.pc[0] ),
    .C(\DJ8.pc[2] ),
    .A(\DJ8.pc[1] ),
    .Y(_0277_));
 sg13g2_nor2_2 _2140_ (.A(_0276_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_nand4_1 _2141_ (.B(\DJ8.pc[5] ),
    .C(\DJ8.pc[6] ),
    .A(_0275_),
    .Y(_0279_),
    .D(_0278_));
 sg13g2_nor2_1 _2142_ (.A(_0274_),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_nand3_1 _2143_ (.B(\DJ8.pc[9] ),
    .C(_0280_),
    .A(\DJ8.pc[8] ),
    .Y(_0281_));
 sg13g2_xnor2_1 _2144_ (.Y(_0282_),
    .A(_0272_),
    .B(_0281_));
 sg13g2_nor2_1 _2145_ (.A(\DJ8.GH[11] ),
    .B(net46),
    .Y(_0283_));
 sg13g2_a21oi_1 _2146_ (.A1(net45),
    .A2(_0282_),
    .Y(_0284_),
    .B1(_0283_));
 sg13g2_mux2_1 _2147_ (.A0(\DJ8.REGS.write_addr[2] ),
    .A1(_0284_),
    .S(_0267_),
    .X(_0285_));
 sg13g2_nand2_1 _2148_ (.Y(_0286_),
    .A(net69),
    .B(_0285_));
 sg13g2_o21ai_1 _2149_ (.B1(_0286_),
    .Y(_0126_),
    .A1(net69),
    .A2(_0272_));
 sg13g2_inv_1 _2150_ (.Y(_0287_),
    .A(\DJ8.GH[12] ));
 sg13g2_buf_1 _2151_ (.A(_0262_),
    .X(_0288_));
 sg13g2_o21ai_1 _2152_ (.B1(_0267_),
    .Y(_0289_),
    .A1(_0287_),
    .A2(net44));
 sg13g2_nor2b_1 _2153_ (.A(\DJ8.pc[11] ),
    .B_N(\DJ8.state[1] ),
    .Y(_0290_));
 sg13g2_nor2_1 _2154_ (.A(_0272_),
    .B(_0281_),
    .Y(_0291_));
 sg13g2_mux2_1 _2155_ (.A0(\DJ8.pc[11] ),
    .A1(_0290_),
    .S(_0291_),
    .X(_0292_));
 sg13g2_a22oi_1 _2156_ (.Y(_0293_),
    .B1(_0292_),
    .B2(_0288_),
    .A2(_0289_),
    .A1(_0270_));
 sg13g2_nor2_1 _2157_ (.A(_0415_),
    .B(net35),
    .Y(_0294_));
 sg13g2_nand2b_1 _2158_ (.Y(_0295_),
    .B(\DJ8.pc[11] ),
    .A_N(net76));
 sg13g2_o21ai_1 _2159_ (.B1(_0295_),
    .Y(_0127_),
    .A1(_0293_),
    .A2(_0294_));
 sg13g2_inv_1 _2160_ (.Y(_0296_),
    .A(\DJ8.pc[12] ));
 sg13g2_inv_1 _2161_ (.Y(_0297_),
    .A(net45));
 sg13g2_and2_1 _2162_ (.A(\DJ8.pc[11] ),
    .B(_0291_),
    .X(_0298_));
 sg13g2_and2_1 _2163_ (.A(\DJ8.state[1] ),
    .B(_0267_),
    .X(_0299_));
 sg13g2_buf_1 _2164_ (.A(_0299_),
    .X(_0300_));
 sg13g2_o21ai_1 _2165_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_and2_1 _2166_ (.A(\DJ8.pc[12] ),
    .B(_0298_),
    .X(_0302_));
 sg13g2_buf_1 _2167_ (.A(_0302_),
    .X(_0303_));
 sg13g2_nand2_1 _2168_ (.Y(_0304_),
    .A(net44),
    .B(_0303_));
 sg13g2_o21ai_1 _2169_ (.B1(_0304_),
    .Y(_0305_),
    .A1(\DJ8.GH[13] ),
    .A2(net44));
 sg13g2_a22oi_1 _2170_ (.Y(_0128_),
    .B1(_0305_),
    .B2(_0300_),
    .A2(_0301_),
    .A1(_0296_));
 sg13g2_xnor2_1 _2171_ (.Y(_0306_),
    .A(\DJ8.pc[13] ),
    .B(_0303_));
 sg13g2_nor2_1 _2172_ (.A(\DJ8.GH[14] ),
    .B(net44),
    .Y(_0307_));
 sg13g2_a21oi_1 _2173_ (.A1(net44),
    .A2(_0306_),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_nor2_1 _2174_ (.A(_0039_),
    .B(_0300_),
    .Y(_0309_));
 sg13g2_a21oi_1 _2175_ (.A1(_0300_),
    .A2(_0308_),
    .Y(_0129_),
    .B1(_0309_));
 sg13g2_nand4_1 _2176_ (.B(\DJ8.pc[14] ),
    .C(net44),
    .A(\DJ8.pc[13] ),
    .Y(_0310_),
    .D(_0303_));
 sg13g2_o21ai_1 _2177_ (.B1(_0310_),
    .Y(_0311_),
    .A1(\DJ8.GH[15] ),
    .A2(net44));
 sg13g2_a21o_1 _2178_ (.A2(_0303_),
    .A1(\DJ8.pc[13] ),
    .B1(_0297_),
    .X(_0312_));
 sg13g2_a21oi_1 _2179_ (.A1(_0300_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(\DJ8.pc[14] ));
 sg13g2_a21oi_1 _2180_ (.A1(_0300_),
    .A2(_0311_),
    .Y(_0130_),
    .B1(_0313_));
 sg13g2_xnor2_1 _2181_ (.Y(_0314_),
    .A(\DJ8.pc[1] ),
    .B(\DJ8.pc[0] ));
 sg13g2_nor2_1 _2182_ (.A(\DJ8.GH[2] ),
    .B(_0273_),
    .Y(_0315_));
 sg13g2_a21oi_1 _2183_ (.A1(_0288_),
    .A2(_0314_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_mux2_1 _2184_ (.A0(\DJ8.ir[1] ),
    .A1(_0316_),
    .S(net35),
    .X(_0317_));
 sg13g2_mux2_1 _2185_ (.A0(\DJ8.pc[1] ),
    .A1(_0317_),
    .S(net69),
    .X(_0131_));
 sg13g2_nand2_1 _2186_ (.Y(_0318_),
    .A(\DJ8.pc[1] ),
    .B(\DJ8.pc[0] ));
 sg13g2_xor2_1 _2187_ (.B(_0318_),
    .A(\DJ8.pc[2] ),
    .X(_0319_));
 sg13g2_nor2_1 _2188_ (.A(\DJ8.GH[3] ),
    .B(_0263_),
    .Y(_0320_));
 sg13g2_a21oi_1 _2189_ (.A1(_0273_),
    .A2(_0319_),
    .Y(_0321_),
    .B1(_0320_));
 sg13g2_nand2_1 _2190_ (.Y(_0322_),
    .A(_0268_),
    .B(_0321_));
 sg13g2_o21ai_1 _2191_ (.B1(_0322_),
    .Y(_0323_),
    .A1(_0141_),
    .A2(_0268_));
 sg13g2_mux2_1 _2192_ (.A0(\DJ8.pc[2] ),
    .A1(_0323_),
    .S(net69),
    .X(_0132_));
 sg13g2_xnor2_1 _2193_ (.Y(_0324_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_nor2_1 _2194_ (.A(\DJ8.GH[4] ),
    .B(_0263_),
    .Y(_0325_));
 sg13g2_a21oi_1 _2195_ (.A1(net45),
    .A2(_0324_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_mux2_1 _2196_ (.A0(\DJ8.ir[3] ),
    .A1(_0326_),
    .S(_0267_),
    .X(_0327_));
 sg13g2_nand2_1 _2197_ (.Y(_0328_),
    .A(_0271_),
    .B(_0327_));
 sg13g2_o21ai_1 _2198_ (.B1(_0328_),
    .Y(_0133_),
    .A1(_0271_),
    .A2(_0276_));
 sg13g2_xnor2_1 _2199_ (.Y(_0329_),
    .A(_0275_),
    .B(_0278_));
 sg13g2_nor2_1 _2200_ (.A(\DJ8.GH[5] ),
    .B(net46),
    .Y(_0330_));
 sg13g2_a21oi_1 _2201_ (.A1(net44),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_mux2_1 _2202_ (.A0(net39),
    .A1(_0331_),
    .S(net35),
    .X(_0332_));
 sg13g2_mux2_1 _2203_ (.A0(_0275_),
    .A1(_0332_),
    .S(net76),
    .X(_0134_));
 sg13g2_nand2_1 _2204_ (.Y(_0333_),
    .A(_0275_),
    .B(_0278_));
 sg13g2_xor2_1 _2205_ (.B(_0333_),
    .A(\DJ8.pc[5] ),
    .X(_0334_));
 sg13g2_nor2_1 _2206_ (.A(\DJ8.GH[6] ),
    .B(net46),
    .Y(_0335_));
 sg13g2_a21oi_1 _2207_ (.A1(net45),
    .A2(_0334_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_mux2_1 _2208_ (.A0(_0512_),
    .A1(_0336_),
    .S(net35),
    .X(_0337_));
 sg13g2_mux2_1 _2209_ (.A0(\DJ8.pc[5] ),
    .A1(_0337_),
    .S(net76),
    .X(_0135_));
 sg13g2_nand3_1 _2210_ (.B(\DJ8.pc[5] ),
    .C(_0278_),
    .A(_0275_),
    .Y(_0338_));
 sg13g2_xor2_1 _2211_ (.B(_0338_),
    .A(\DJ8.pc[6] ),
    .X(_0339_));
 sg13g2_nor2_1 _2212_ (.A(\DJ8.GH[7] ),
    .B(net46),
    .Y(_0340_));
 sg13g2_a21oi_1 _2213_ (.A1(net45),
    .A2(_0339_),
    .Y(_0341_),
    .B1(_0340_));
 sg13g2_mux2_1 _2214_ (.A0(_0505_),
    .A1(_0341_),
    .S(net35),
    .X(_0342_));
 sg13g2_mux2_1 _2215_ (.A0(\DJ8.pc[6] ),
    .A1(_0342_),
    .S(net76),
    .X(_0136_));
 sg13g2_xnor2_1 _2216_ (.Y(_0343_),
    .A(_0274_),
    .B(_0279_));
 sg13g2_nor2_1 _2217_ (.A(\DJ8.GH[8] ),
    .B(net46),
    .Y(_0344_));
 sg13g2_a21oi_1 _2218_ (.A1(net45),
    .A2(_0343_),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_mux2_1 _2219_ (.A0(\DJ8.ir[7] ),
    .A1(_0345_),
    .S(_0267_),
    .X(_0346_));
 sg13g2_nand2_1 _2220_ (.Y(_0347_),
    .A(net69),
    .B(_0346_));
 sg13g2_o21ai_1 _2221_ (.B1(_0347_),
    .Y(_0137_),
    .A1(net69),
    .A2(_0274_));
 sg13g2_xnor2_1 _2222_ (.Y(_0348_),
    .A(\DJ8.pc[8] ),
    .B(_0280_));
 sg13g2_nor2_1 _2223_ (.A(\DJ8.GH[9] ),
    .B(net46),
    .Y(_0349_));
 sg13g2_a21oi_1 _2224_ (.A1(net45),
    .A2(_0348_),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_mux2_1 _2225_ (.A0(_0653_),
    .A1(_0350_),
    .S(net35),
    .X(_0351_));
 sg13g2_mux2_1 _2226_ (.A0(\DJ8.pc[8] ),
    .A1(_0351_),
    .S(net76),
    .X(_0138_));
 sg13g2_nand2_1 _2227_ (.Y(_0352_),
    .A(\DJ8.pc[8] ),
    .B(_0280_));
 sg13g2_xor2_1 _2228_ (.B(_0352_),
    .A(\DJ8.pc[9] ),
    .X(_0353_));
 sg13g2_nor2_1 _2229_ (.A(\DJ8.GH[10] ),
    .B(net46),
    .Y(_0354_));
 sg13g2_a21oi_1 _2230_ (.A1(net45),
    .A2(_0353_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_mux2_1 _2231_ (.A0(_0654_),
    .A1(_0355_),
    .S(net35),
    .X(_0356_));
 sg13g2_mux2_1 _2232_ (.A0(\DJ8.pc[9] ),
    .A1(_0356_),
    .S(net76),
    .X(_0139_));
 sg13g2_inv_1 _2233_ (.Y(_0357_),
    .A(\DJ8.state[3] ));
 sg13g2_nand3_1 _2234_ (.B(_0270_),
    .C(_0410_),
    .A(_0407_),
    .Y(_0358_));
 sg13g2_o21ai_1 _2235_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0357_),
    .A2(net76));
 sg13g2_mux2_1 _2236_ (.A0(_0040_),
    .A1(_0030_),
    .S(_0359_),
    .X(_0140_));
 sg13g2_a21oi_1 _2237_ (.A1(net69),
    .A2(_0411_),
    .Y(_0041_),
    .B1(\DJ8.state[3] ));
 sg13g2_nor3_2 _2238_ (.A(_0430_),
    .B(net81),
    .C(_0411_),
    .Y(_0360_));
 sg13g2_buf_1 _2239_ (.A(_0360_),
    .X(_0361_));
 sg13g2_nand2_1 _2240_ (.Y(_0362_),
    .A(_0589_),
    .B(net43));
 sg13g2_o21ai_1 _2241_ (.B1(_0675_),
    .Y(_0363_),
    .A1(_0430_),
    .A2(_0411_));
 sg13g2_nand2_1 _2242_ (.Y(net10),
    .A(_0362_),
    .B(_0363_));
 sg13g2_nor2_1 _2243_ (.A(_0558_),
    .B(net43),
    .Y(_0364_));
 sg13g2_a21oi_1 _2244_ (.A1(_0538_),
    .A2(net43),
    .Y(net11),
    .B1(_0364_));
 sg13g2_mux2_1 _2245_ (.A0(_0554_),
    .A1(_0695_),
    .S(_0360_),
    .X(net12));
 sg13g2_nand2_1 _2246_ (.Y(_0365_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_nand3_1 _2247_ (.B(_0365_),
    .C(_0360_),
    .A(_0780_),
    .Y(_0366_));
 sg13g2_o21ai_1 _2248_ (.B1(_0366_),
    .Y(net13),
    .A1(_0991_),
    .A2(net43));
 sg13g2_and2_1 _2249_ (.A(_0905_),
    .B(_0572_),
    .X(_0367_));
 sg13g2_a21oi_1 _2250_ (.A1(net83),
    .A2(_0559_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_nor2_1 _2251_ (.A(_0368_),
    .B(_0361_),
    .Y(_0369_));
 sg13g2_a21oi_1 _2252_ (.A1(_0852_),
    .A2(_0361_),
    .Y(net14),
    .B1(_0369_));
 sg13g2_buf_1 _2253_ (.A(net50),
    .X(_0370_));
 sg13g2_nor2b_1 _2254_ (.A(net47),
    .B_N(\DJ8.GH[5] ),
    .Y(_0371_));
 sg13g2_a21oi_1 _2255_ (.A1(net47),
    .A2(\DJ8.EF[5] ),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nor2_1 _2256_ (.A(net50),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_a21oi_1 _2257_ (.A1(_0275_),
    .A2(net38),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_nand2_1 _2258_ (.Y(_0375_),
    .A(_0931_),
    .B(net43));
 sg13g2_o21ai_1 _2259_ (.B1(_0375_),
    .Y(net15),
    .A1(net43),
    .A2(_0374_));
 sg13g2_nor2b_1 _2260_ (.A(net47),
    .B_N(\DJ8.GH[6] ),
    .Y(_0376_));
 sg13g2_a21oi_1 _2261_ (.A1(net47),
    .A2(\DJ8.EF[6] ),
    .Y(_0377_),
    .B1(_0376_));
 sg13g2_nor2_1 _2262_ (.A(net50),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_a21oi_1 _2263_ (.A1(\DJ8.pc[5] ),
    .A2(net38),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_and2_1 _2264_ (.A(_1020_),
    .B(_1021_),
    .X(_0380_));
 sg13g2_nand2_1 _2265_ (.Y(_0381_),
    .A(_0380_),
    .B(_0360_));
 sg13g2_o21ai_1 _2266_ (.B1(_0381_),
    .Y(net16),
    .A1(net43),
    .A2(_0379_));
 sg13g2_nor2b_1 _2267_ (.A(net62),
    .B_N(\DJ8.GH[7] ),
    .Y(_0382_));
 sg13g2_a21oi_1 _2268_ (.A1(net47),
    .A2(\DJ8.EF[7] ),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_nor2_1 _2269_ (.A(net50),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_a21oi_1 _2270_ (.A1(\DJ8.pc[6] ),
    .A2(net50),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_nand2_1 _2271_ (.Y(_0386_),
    .A(_1081_),
    .B(_0360_));
 sg13g2_o21ai_1 _2272_ (.B1(_0386_),
    .Y(net17),
    .A1(net43),
    .A2(_0385_));
 sg13g2_inv_1 _2273_ (.Y(_0387_),
    .A(\DJ8.GH[8] ));
 sg13g2_nand2_1 _2274_ (.Y(_0388_),
    .A(\DJ8.EF[8] ),
    .B(_0258_));
 sg13g2_o21ai_1 _2275_ (.B1(_0388_),
    .Y(_0389_),
    .A1(_0387_),
    .A2(net39));
 sg13g2_nand2_1 _2276_ (.Y(_0390_),
    .A(net40),
    .B(_0389_));
 sg13g2_o21ai_1 _2277_ (.B1(_0390_),
    .Y(net18),
    .A1(_0274_),
    .A2(net40));
 sg13g2_nor2b_1 _2278_ (.A(net39),
    .B_N(\DJ8.GH[9] ),
    .Y(_0391_));
 sg13g2_a21oi_1 _2279_ (.A1(net39),
    .A2(\DJ8.EF[9] ),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_nand2_1 _2280_ (.Y(_0393_),
    .A(\DJ8.pc[8] ),
    .B(_0370_));
 sg13g2_o21ai_1 _2281_ (.B1(_0393_),
    .Y(net19),
    .A1(_0370_),
    .A2(_0392_));
 sg13g2_nor2b_1 _2282_ (.A(net39),
    .B_N(\DJ8.GH[10] ),
    .Y(_0394_));
 sg13g2_a21oi_1 _2283_ (.A1(net39),
    .A2(\DJ8.EF[10] ),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_nand2_1 _2284_ (.Y(_0396_),
    .A(\DJ8.pc[9] ),
    .B(net38));
 sg13g2_o21ai_1 _2285_ (.B1(_0396_),
    .Y(net20),
    .A1(net38),
    .A2(_0395_));
 sg13g2_mux2_1 _2286_ (.A0(\DJ8.GH[11] ),
    .A1(\DJ8.EF[11] ),
    .S(net47),
    .X(_0397_));
 sg13g2_nand2_1 _2287_ (.Y(_0398_),
    .A(net40),
    .B(_0397_));
 sg13g2_o21ai_1 _2288_ (.B1(_0398_),
    .Y(net21),
    .A1(_0272_),
    .A2(net40));
 sg13g2_nor2_1 _2289_ (.A(_0259_),
    .B(_0287_),
    .Y(_0399_));
 sg13g2_a21oi_1 _2290_ (.A1(_0259_),
    .A2(\DJ8.EF[12] ),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_nand2_1 _2291_ (.Y(_0401_),
    .A(\DJ8.pc[11] ),
    .B(net38));
 sg13g2_o21ai_1 _2292_ (.B1(_0401_),
    .Y(net22),
    .A1(net38),
    .A2(_0400_));
 sg13g2_mux2_1 _2293_ (.A0(\DJ8.GH[13] ),
    .A1(\DJ8.EF[13] ),
    .S(net47),
    .X(_0402_));
 sg13g2_nand2_1 _2294_ (.Y(_0403_),
    .A(net40),
    .B(_0402_));
 sg13g2_o21ai_1 _2295_ (.B1(_0403_),
    .Y(net23),
    .A1(_0296_),
    .A2(net40));
 sg13g2_nor2_1 _2296_ (.A(net47),
    .B(_1005_),
    .Y(_0404_));
 sg13g2_a21oi_1 _2297_ (.A1(net39),
    .A2(\DJ8.EF[14] ),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_nand2_1 _2298_ (.Y(_0406_),
    .A(\DJ8.pc[13] ),
    .B(net38));
 sg13g2_o21ai_1 _2299_ (.B1(_0406_),
    .Y(net24),
    .A1(net38),
    .A2(_0405_));
 sg13g2_inv_1 _1200__1 (.Y(net113),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_1 _2301_ (.A(net105),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2302_ (.A(net106),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2303_ (.A(net107),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2304_ (.A(net108),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2305_ (.A(net109),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2306_ (.A(net110),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2307_ (.A(net111),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2308_ (.A(net112),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2309_ (.A(\DJ8.we ),
    .X(net25));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout26 (.A(_0823_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0168_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0158_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0148_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0660_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0205_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0196_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0187_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0178_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0268_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0935_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0661_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0370_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0259_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0905_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0626_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0499_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0361_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0288_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0273_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0263_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0258_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0606_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0564_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0559_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0539_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0522_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0493_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0419_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0701_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0629_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0535_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0524_),
    .X(net58));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(_0515_));
 sg13g2_buf_2 fanout60 (.A(_0508_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0468_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0439_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0434_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0786_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0623_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0604_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0501_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0438_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0271_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0238_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0235_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0619_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0615_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0500_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0437_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0270_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0654_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0653_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0609_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0593_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0482_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0426_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0423_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0415_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0408_),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net89));
 sg13g2_buf_2 fanout87 (.A(net89),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net89));
 sg13g2_buf_2 fanout89 (.A(net104),
    .X(net89));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net92));
 sg13g2_buf_2 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net104),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net98));
 sg13g2_buf_2 fanout94 (.A(net98),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(net96));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net98));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net98));
 sg13g2_buf_2 fanout98 (.A(net104),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net103));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net101));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net103));
 sg13g2_buf_2 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net1),
    .X(net104));
 sg13g2_tiehi _2301__105 (.L_HI(net105));
 sg13g2_tiehi _2302__106 (.L_HI(net106));
 sg13g2_tiehi _2303__107 (.L_HI(net107));
 sg13g2_tiehi _2304__108 (.L_HI(net108));
 sg13g2_tiehi _2305__109 (.L_HI(net109));
 sg13g2_tiehi _2306__110 (.L_HI(net110));
 sg13g2_tiehi _2307__111 (.L_HI(net111));
 sg13g2_tiehi _2308__112 (.L_HI(net112));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_fill_1 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_fill_2 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_4 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_4 FILLER_2_286 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_330 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_4 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_fill_1 FILLER_2_375 ();
 sg13g2_fill_2 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_4 FILLER_2_402 ();
 sg13g2_fill_1 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_416 ();
 sg13g2_decap_8 FILLER_2_423 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_284 ();
 sg13g2_fill_2 FILLER_3_331 ();
 sg13g2_decap_4 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_fill_2 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_388 ();
 sg13g2_fill_1 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_fill_2 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_251 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_fill_1 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_4 FILLER_4_289 ();
 sg13g2_fill_2 FILLER_4_293 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_decap_4 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_359 ();
 sg13g2_fill_1 FILLER_4_369 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_1 FILLER_4_414 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_2 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_4 FILLER_5_284 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_4 FILLER_5_334 ();
 sg13g2_decap_4 FILLER_5_349 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_fill_2 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_388 ();
 sg13g2_fill_1 FILLER_5_394 ();
 sg13g2_decap_4 FILLER_5_398 ();
 sg13g2_fill_2 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_320 ();
 sg13g2_fill_2 FILLER_6_343 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_352 ();
 sg13g2_fill_1 FILLER_6_357 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_fill_2 FILLER_6_387 ();
 sg13g2_fill_2 FILLER_6_394 ();
 sg13g2_fill_2 FILLER_6_405 ();
 sg13g2_fill_2 FILLER_6_411 ();
 sg13g2_fill_1 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_decap_4 FILLER_7_155 ();
 sg13g2_fill_2 FILLER_7_159 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_decap_4 FILLER_7_231 ();
 sg13g2_fill_1 FILLER_7_235 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_decap_4 FILLER_7_298 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_decap_4 FILLER_7_319 ();
 sg13g2_decap_4 FILLER_7_331 ();
 sg13g2_fill_1 FILLER_7_335 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_decap_4 FILLER_7_364 ();
 sg13g2_fill_2 FILLER_7_368 ();
 sg13g2_decap_4 FILLER_7_374 ();
 sg13g2_fill_1 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_8 FILLER_7_419 ();
 sg13g2_decap_4 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_38 ();
 sg13g2_fill_2 FILLER_8_45 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_decap_8 FILLER_8_52 ();
 sg13g2_fill_2 FILLER_8_59 ();
 sg13g2_fill_1 FILLER_8_61 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_151 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_199 ();
 sg13g2_fill_2 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_decap_4 FILLER_8_237 ();
 sg13g2_decap_4 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_fill_1 FILLER_8_286 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_decap_4 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_338 ();
 sg13g2_decap_4 FILLER_8_344 ();
 sg13g2_fill_2 FILLER_8_348 ();
 sg13g2_decap_4 FILLER_8_359 ();
 sg13g2_fill_1 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_fill_2 FILLER_8_393 ();
 sg13g2_fill_1 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_4 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_54 ();
 sg13g2_fill_1 FILLER_9_61 ();
 sg13g2_decap_8 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_decap_4 FILLER_9_85 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_4 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_decap_4 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_4 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_4 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_344 ();
 sg13g2_decap_4 FILLER_9_358 ();
 sg13g2_fill_1 FILLER_9_362 ();
 sg13g2_fill_1 FILLER_9_393 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_fill_2 FILLER_10_51 ();
 sg13g2_fill_2 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_266 ();
 sg13g2_decap_4 FILLER_10_272 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_decap_4 FILLER_10_338 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_364 ();
 sg13g2_decap_4 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_44 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_73 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_decap_4 FILLER_11_85 ();
 sg13g2_decap_8 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_100 ();
 sg13g2_fill_2 FILLER_11_107 ();
 sg13g2_decap_4 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_decap_8 FILLER_11_176 ();
 sg13g2_decap_8 FILLER_11_183 ();
 sg13g2_decap_8 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_decap_4 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_282 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_fill_2 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_25 ();
 sg13g2_decap_4 FILLER_12_32 ();
 sg13g2_decap_4 FILLER_12_40 ();
 sg13g2_fill_2 FILLER_12_44 ();
 sg13g2_fill_2 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_4 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_150 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_4 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_fill_2 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_4 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_312 ();
 sg13g2_fill_2 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_334 ();
 sg13g2_fill_1 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_decap_4 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_4 FILLER_12_393 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_1 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_4 FILLER_12_416 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_decap_4 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_4 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_decap_8 FILLER_13_145 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_177 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_decap_4 FILLER_13_363 ();
 sg13g2_decap_4 FILLER_13_387 ();
 sg13g2_fill_2 FILLER_13_391 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_2 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_51 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_decap_4 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_322 ();
 sg13g2_decap_4 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_102 ();
 sg13g2_fill_1 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_4 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_4 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_384 ();
 sg13g2_fill_1 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_decap_4 FILLER_16_37 ();
 sg13g2_fill_1 FILLER_16_41 ();
 sg13g2_decap_4 FILLER_16_46 ();
 sg13g2_decap_4 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_decap_4 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_fill_2 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_decap_4 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_111 ();
 sg13g2_fill_1 FILLER_16_121 ();
 sg13g2_decap_4 FILLER_16_127 ();
 sg13g2_decap_4 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_4 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_decap_4 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_decap_4 FILLER_17_62 ();
 sg13g2_decap_4 FILLER_17_80 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_decap_8 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_decap_4 FILLER_17_166 ();
 sg13g2_decap_4 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_decap_4 FILLER_17_270 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_4 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_393 ();
 sg13g2_decap_4 FILLER_17_418 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_27 ();
 sg13g2_fill_2 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_4 FILLER_18_95 ();
 sg13g2_fill_2 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_118 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_decap_4 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_4 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_4 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_decap_4 FILLER_18_362 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_55 ();
 sg13g2_decap_4 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_79 ();
 sg13g2_decap_8 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_decap_4 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_120 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_decap_4 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_fill_2 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_4 FILLER_20_29 ();
 sg13g2_fill_2 FILLER_20_33 ();
 sg13g2_decap_4 FILLER_20_40 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_decap_4 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_4 FILLER_20_179 ();
 sg13g2_fill_1 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_262 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_decap_4 FILLER_20_393 ();
 sg13g2_decap_4 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_4 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_decap_4 FILLER_21_142 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_decap_4 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_254 ();
 sg13g2_decap_4 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_296 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_4 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_decap_4 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_4 FILLER_22_306 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_decap_4 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_decap_8 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_decap_8 FILLER_23_43 ();
 sg13g2_decap_8 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_57 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_8 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_135 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_fill_2 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_4 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_85 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_decap_4 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_206 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_fill_2 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_386 ();
 sg13g2_decap_4 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_401 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_decap_4 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_4 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_243 ();
 sg13g2_decap_4 FILLER_25_255 ();
 sg13g2_decap_4 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_391 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_44 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_86 ();
 sg13g2_decap_4 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_decap_4 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_decap_4 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_410 ();
 sg13g2_fill_2 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_decap_4 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_decap_4 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_decap_4 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_4 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_374 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_384 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_decap_4 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_43 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_120 ();
 sg13g2_decap_4 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_144 ();
 sg13g2_decap_4 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_4 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_decap_4 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_4 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_4 FILLER_28_374 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_28_388 ();
 sg13g2_fill_1 FILLER_28_397 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_4 FILLER_29_26 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_4 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_decap_4 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_decap_4 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_decap_4 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_decap_8 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_29_415 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_85 ();
 sg13g2_decap_8 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_decap_4 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_decap_4 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_decap_4 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_405 ();
 sg13g2_fill_2 FILLER_30_411 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_decap_8 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_4 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_149 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_decap_4 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_decap_4 FILLER_31_424 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_30 ();
 sg13g2_decap_8 FILLER_32_38 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_61 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_411 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_decap_8 FILLER_33_36 ();
 sg13g2_decap_4 FILLER_33_43 ();
 sg13g2_decap_8 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_decap_4 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_decap_4 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_190 ();
 sg13g2_decap_4 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_258 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_33_404 ();
 sg13g2_decap_8 FILLER_33_411 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_decap_4 FILLER_34_65 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_decap_4 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_4 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_4 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_decap_4 FILLER_34_394 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_426 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_31 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_decap_4 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_128 ();
 sg13g2_decap_4 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_150 ();
 sg13g2_decap_8 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_fill_1 FILLER_36_140 ();
 sg13g2_decap_4 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_173 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_2 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_decap_4 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_decap_4 FILLER_37_394 ();
 sg13g2_fill_2 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_411 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_decap_8 FILLER_38_64 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_127 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_fill_1 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
