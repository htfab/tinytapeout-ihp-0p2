module tt_um_rebeccargb_hardware_utf8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire clknet_0_clk;
 wire retry;
 wire \u8.empty ;
 wire \u8.hs[0] ;
 wire \u8.hs[1] ;
 wire \u8.hs[2] ;
 wire \u8.hs[3] ;
 wire \u8.hs[4] ;
 wire \u8.hs[5] ;
 wire \u8.ls[0] ;
 wire \u8.ls[1] ;
 wire \u8.ls[2] ;
 wire \u8.ls[3] ;
 wire \u8.ls[4] ;
 wire \u8.ls[5] ;
 wire \u8.ls[6] ;
 wire \u8.ls[7] ;
 wire \u8.ls[8] ;
 wire \u8.ls[9] ;
 wire \u8.rbop[0] ;
 wire \u8.rbop[1] ;
 wire \u8.rbop[2] ;
 wire \u8.rc[16] ;
 wire \u8.rc[17] ;
 wire \u8.rc[18] ;
 wire \u8.rc[19] ;
 wire \u8.rc[20] ;
 wire \u8.rc[21] ;
 wire \u8.rc[22] ;
 wire \u8.rc[23] ;
 wire \u8.rc[24] ;
 wire \u8.rc[25] ;
 wire \u8.rc[26] ;
 wire \u8.rc[27] ;
 wire \u8.rc[28] ;
 wire \u8.rc[29] ;
 wire \u8.rc[30] ;
 wire \u8.rc[31] ;
 wire \u8.rcip[0] ;
 wire \u8.rcip[1] ;
 wire \u8.rcip[2] ;
 wire \u8.rcop[0] ;
 wire \u8.rcop[1] ;
 wire \u8.rcop[2] ;
 wire \u8.ruop[0] ;
 wire \u8.ruop[1] ;
 wire \u8.ruop[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_inv_1 _1491_ (.Y(_0654_),
    .A(net21));
 sg13g2_buf_2 _1492_ (.A(ui_in[6]),
    .X(_0655_));
 sg13g2_buf_8 _1493_ (.A(\u8.rc[30] ),
    .X(_0656_));
 sg13g2_buf_1 _1494_ (.A(\u8.rc[31] ),
    .X(_0657_));
 sg13g2_and2_1 _1495_ (.A(_0656_),
    .B(net140),
    .X(_0658_));
 sg13g2_buf_2 _1496_ (.A(_0658_),
    .X(_0659_));
 sg13g2_buf_2 _1497_ (.A(\u8.rc[27] ),
    .X(_0660_));
 sg13g2_buf_2 _1498_ (.A(\u8.rc[26] ),
    .X(_0661_));
 sg13g2_and2_1 _1499_ (.A(_0660_),
    .B(_0661_),
    .X(_0662_));
 sg13g2_buf_1 _1500_ (.A(_0662_),
    .X(_0663_));
 sg13g2_buf_8 _1501_ (.A(\u8.rc[23] ),
    .X(_0664_));
 sg13g2_buf_1 _1502_ (.A(\u8.rc[22] ),
    .X(_0665_));
 sg13g2_and2_1 _1503_ (.A(_0664_),
    .B(net139),
    .X(_0666_));
 sg13g2_buf_1 _1504_ (.A(\u8.rc[29] ),
    .X(_0667_));
 sg13g2_buf_8 _1505_ (.A(\u8.rc[28] ),
    .X(_0668_));
 sg13g2_nor2b_1 _1506_ (.A(net138),
    .B_N(net137),
    .Y(_0669_));
 sg13g2_buf_8 _1507_ (.A(\u8.rc[25] ),
    .X(_0670_));
 sg13g2_buf_8 _1508_ (.A(\u8.rc[24] ),
    .X(_0671_));
 sg13g2_nor2b_1 _1509_ (.A(net136),
    .B_N(_0671_),
    .Y(_0672_));
 sg13g2_and4_1 _1510_ (.A(_0663_),
    .B(_0666_),
    .C(_0669_),
    .D(_0672_),
    .X(_0673_));
 sg13g2_buf_1 _1511_ (.A(\u8.rc[21] ),
    .X(_0674_));
 sg13g2_buf_1 _1512_ (.A(\u8.rc[20] ),
    .X(_0675_));
 sg13g2_nand2b_1 _1513_ (.Y(_0676_),
    .B(net134),
    .A_N(net135));
 sg13g2_buf_1 _1514_ (.A(\u8.rc[19] ),
    .X(_0677_));
 sg13g2_buf_1 _1515_ (.A(\u8.rc[18] ),
    .X(_0678_));
 sg13g2_nand2_1 _1516_ (.Y(_0679_),
    .A(net133),
    .B(net132));
 sg13g2_buf_1 _1517_ (.A(_0020_),
    .X(_0680_));
 sg13g2_o21ai_1 _1518_ (.B1(net131),
    .Y(_0681_),
    .A1(_0676_),
    .A2(_0679_));
 sg13g2_buf_2 _1519_ (.A(_0019_),
    .X(_0682_));
 sg13g2_nor2b_1 _1520_ (.A(_0682_),
    .B_N(net137),
    .Y(_0683_));
 sg13g2_a21o_1 _1521_ (.A2(_0683_),
    .A1(_0663_),
    .B1(net138),
    .X(_0684_));
 sg13g2_a21o_1 _1522_ (.A2(_0681_),
    .A1(_0673_),
    .B1(_0684_),
    .X(_0685_));
 sg13g2_nand2_1 _1523_ (.Y(_0686_),
    .A(_0659_),
    .B(_0685_));
 sg13g2_and2_1 _1524_ (.A(_0659_),
    .B(_0685_),
    .X(_0687_));
 sg13g2_nor2b_1 _1525_ (.A(net135),
    .B_N(net134),
    .Y(_0688_));
 sg13g2_nor2b_1 _1526_ (.A(net138),
    .B_N(_0682_),
    .Y(_0689_));
 sg13g2_nand3_1 _1527_ (.B(_0689_),
    .C(_0659_),
    .A(_0688_),
    .Y(_0690_));
 sg13g2_nand4_1 _1528_ (.B(_0666_),
    .C(_0669_),
    .A(_0663_),
    .Y(_0691_),
    .D(_0672_));
 sg13g2_nor2_1 _1529_ (.A(_0690_),
    .B(_0691_),
    .Y(_0692_));
 sg13g2_buf_1 _1530_ (.A(\u8.hs[0] ),
    .X(_0693_));
 sg13g2_nand3_1 _1531_ (.B(\u8.hs[1] ),
    .C(net130),
    .A(\u8.hs[2] ),
    .Y(_0694_));
 sg13g2_buf_1 _1532_ (.A(_0694_),
    .X(_0695_));
 sg13g2_buf_2 _1533_ (.A(\u8.rc[16] ),
    .X(_0696_));
 sg13g2_buf_1 _1534_ (.A(\u8.hs[4] ),
    .X(_0697_));
 sg13g2_buf_2 _1535_ (.A(\u8.hs[5] ),
    .X(_0698_));
 sg13g2_nand3_1 _1536_ (.B(net129),
    .C(_0698_),
    .A(_0696_),
    .Y(_0699_));
 sg13g2_nor2_1 _1537_ (.A(_0695_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_nand2_1 _1538_ (.Y(_0701_),
    .A(_0664_),
    .B(net139));
 sg13g2_nor2_1 _1539_ (.A(net131),
    .B(_0701_),
    .Y(_0702_));
 sg13g2_buf_1 _1540_ (.A(\u8.ls[9] ),
    .X(_0703_));
 sg13g2_buf_1 _1541_ (.A(\u8.ls[8] ),
    .X(_0704_));
 sg13g2_nor2_1 _1542_ (.A(net128),
    .B(net127),
    .Y(_0705_));
 sg13g2_buf_1 _1543_ (.A(\u8.rc[17] ),
    .X(_0706_));
 sg13g2_inv_1 _1544_ (.Y(_0707_),
    .A(net126));
 sg13g2_buf_1 _1545_ (.A(\u8.hs[3] ),
    .X(_0708_));
 sg13g2_inv_1 _1546_ (.Y(_0709_),
    .A(net125));
 sg13g2_buf_2 _1547_ (.A(_0021_),
    .X(_0710_));
 sg13g2_nand4_1 _1548_ (.B(_0709_),
    .C(_0710_),
    .A(_0707_),
    .Y(_0711_),
    .D(_0022_));
 sg13g2_nor4_1 _1549_ (.A(_0679_),
    .B(_0702_),
    .C(_0705_),
    .D(_0711_),
    .Y(_0712_));
 sg13g2_nand3_1 _1550_ (.B(_0700_),
    .C(_0712_),
    .A(_0692_),
    .Y(_0713_));
 sg13g2_buf_1 _1551_ (.A(_0013_),
    .X(_0714_));
 sg13g2_inv_1 _1552_ (.Y(_0715_),
    .A(_0680_));
 sg13g2_a21oi_1 _1553_ (.A1(net133),
    .A2(_0688_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_a21oi_1 _1554_ (.A1(_0663_),
    .A2(_0683_),
    .Y(_0717_),
    .B1(net138));
 sg13g2_o21ai_1 _1555_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_0691_),
    .A2(_0716_));
 sg13g2_nand3_1 _1556_ (.B(_0659_),
    .C(_0718_),
    .A(net124),
    .Y(_0719_));
 sg13g2_a21o_1 _1557_ (.A2(_0713_),
    .A1(_0687_),
    .B1(_0719_),
    .X(_0720_));
 sg13g2_buf_2 _1558_ (.A(_0720_),
    .X(_0721_));
 sg13g2_nor4_2 _1559_ (.A(net133),
    .B(net132),
    .C(net126),
    .Y(_0722_),
    .D(_0696_));
 sg13g2_buf_1 _1560_ (.A(_0722_),
    .X(_0723_));
 sg13g2_nor2_1 _1561_ (.A(_0656_),
    .B(\u8.rc[31] ),
    .Y(_0724_));
 sg13g2_nor4_2 _1562_ (.A(\u8.rc[29] ),
    .B(net137),
    .C(_0660_),
    .Y(_0725_),
    .D(_0661_));
 sg13g2_nor2_1 _1563_ (.A(net136),
    .B(_0671_),
    .Y(_0726_));
 sg13g2_nor4_1 _1564_ (.A(_0664_),
    .B(net139),
    .C(\u8.rc[21] ),
    .D(\u8.rc[20] ),
    .Y(_0727_));
 sg13g2_and4_1 _1565_ (.A(_0724_),
    .B(_0725_),
    .C(_0726_),
    .D(_0727_),
    .X(_0728_));
 sg13g2_buf_1 _1566_ (.A(_0728_),
    .X(_0729_));
 sg13g2_and3_1 _1567_ (.X(_0730_),
    .A(_0714_),
    .B(_0723_),
    .C(_0729_));
 sg13g2_inv_1 _1568_ (.Y(_0731_),
    .A(net132));
 sg13g2_nand4_1 _1569_ (.B(_0731_),
    .C(net124),
    .A(net133),
    .Y(_0732_),
    .D(net131));
 sg13g2_nor3_1 _1570_ (.A(_0690_),
    .B(_0691_),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_or2_1 _1571_ (.X(_0734_),
    .B(_0733_),
    .A(_0730_));
 sg13g2_buf_2 _1572_ (.A(\u8.ruop[2] ),
    .X(_0735_));
 sg13g2_inv_1 _1573_ (.Y(_0736_),
    .A(\u8.rc[21] ));
 sg13g2_nor4_1 _1574_ (.A(_0664_),
    .B(net139),
    .C(net136),
    .D(_0671_),
    .Y(_0737_));
 sg13g2_and4_1 _1575_ (.A(_0736_),
    .B(_0724_),
    .C(_0725_),
    .D(_0737_),
    .X(_0738_));
 sg13g2_buf_2 _1576_ (.A(_0738_),
    .X(_0739_));
 sg13g2_xnor2_1 _1577_ (.Y(_0740_),
    .A(net134),
    .B(net91));
 sg13g2_nand3_1 _1578_ (.B(_0739_),
    .C(_0740_),
    .A(_0714_),
    .Y(_0741_));
 sg13g2_buf_1 _1579_ (.A(ui_in[4]),
    .X(_0742_));
 sg13g2_o21ai_1 _1580_ (.B1(net144),
    .Y(_0743_),
    .A1(_0735_),
    .A2(_0741_));
 sg13g2_nor3_1 _1581_ (.A(_0655_),
    .B(_0734_),
    .C(_0743_),
    .Y(_0744_));
 sg13g2_o21ai_1 _1582_ (.B1(_0744_),
    .Y(_0745_),
    .A1(_0686_),
    .A2(_0721_));
 sg13g2_buf_1 _1583_ (.A(net124),
    .X(_0746_));
 sg13g2_a21oi_1 _1584_ (.A1(_0673_),
    .A2(_0681_),
    .Y(_0747_),
    .B1(_0684_));
 sg13g2_nand4_1 _1585_ (.B(_0659_),
    .C(_0718_),
    .A(_0746_),
    .Y(_0748_),
    .D(_0747_));
 sg13g2_buf_1 _1586_ (.A(_0748_),
    .X(_0749_));
 sg13g2_inv_1 _1587_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_inv_1 _1588_ (.Y(_0751_),
    .A(net144));
 sg13g2_buf_1 _1589_ (.A(_0751_),
    .X(_0752_));
 sg13g2_buf_2 _1590_ (.A(_0032_),
    .X(_0753_));
 sg13g2_buf_1 _1591_ (.A(\u8.ruop[0] ),
    .X(_0754_));
 sg13g2_buf_2 _1592_ (.A(\u8.ruop[1] ),
    .X(_0755_));
 sg13g2_nor2b_1 _1593_ (.A(_0754_),
    .B_N(_0755_),
    .Y(_0756_));
 sg13g2_nor2b_1 _1594_ (.A(_0755_),
    .B_N(_0754_),
    .Y(_0757_));
 sg13g2_buf_2 _1595_ (.A(_0757_),
    .X(_0758_));
 sg13g2_or2_1 _1596_ (.X(_0759_),
    .B(_0758_),
    .A(_0756_));
 sg13g2_and2_1 _1597_ (.A(_0753_),
    .B(_0759_),
    .X(_0760_));
 sg13g2_buf_1 _1598_ (.A(_0754_),
    .X(_0761_));
 sg13g2_nor3_1 _1599_ (.A(net105),
    .B(_0755_),
    .C(_0735_),
    .Y(_0762_));
 sg13g2_nor3_1 _1600_ (.A(net106),
    .B(_0760_),
    .C(_0762_),
    .Y(_0763_));
 sg13g2_inv_1 _1601_ (.Y(_0764_),
    .A(_0755_));
 sg13g2_nand2_1 _1602_ (.Y(_0765_),
    .A(_0754_),
    .B(_0753_));
 sg13g2_o21ai_1 _1603_ (.B1(_0765_),
    .Y(_0766_),
    .A1(net105),
    .A2(_0735_));
 sg13g2_and2_1 _1604_ (.A(net91),
    .B(net84),
    .X(_0767_));
 sg13g2_buf_2 _1605_ (.A(_0767_),
    .X(_0768_));
 sg13g2_nand4_1 _1606_ (.B(_0663_),
    .C(_0688_),
    .A(net137),
    .Y(_0769_),
    .D(_0689_));
 sg13g2_nor2_1 _1607_ (.A(net138),
    .B(net136),
    .Y(_0770_));
 sg13g2_nand4_1 _1608_ (.B(_0666_),
    .C(_0659_),
    .A(_0671_),
    .Y(_0771_),
    .D(_0770_));
 sg13g2_nand3_1 _1609_ (.B(_0731_),
    .C(net131),
    .A(net133),
    .Y(_0772_));
 sg13g2_nor3_1 _1610_ (.A(_0769_),
    .B(_0771_),
    .C(_0772_),
    .Y(_0773_));
 sg13g2_o21ai_1 _1611_ (.B1(net124),
    .Y(_0774_),
    .A1(_0768_),
    .A2(_0773_));
 sg13g2_a21oi_1 _1612_ (.A1(_0764_),
    .A2(_0766_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_a22oi_1 _1613_ (.Y(_0776_),
    .B1(_0775_),
    .B2(_0721_),
    .A2(_0763_),
    .A1(_0750_));
 sg13g2_a21oi_2 _1614_ (.B1(_0719_),
    .Y(_0777_),
    .A2(_0713_),
    .A1(_0687_));
 sg13g2_xnor2_1 _1615_ (.Y(_0778_),
    .A(_0735_),
    .B(_0741_));
 sg13g2_inv_1 _1616_ (.Y(_0779_),
    .A(_0754_));
 sg13g2_nor2_1 _1617_ (.A(_0754_),
    .B(_0732_),
    .Y(_0780_));
 sg13g2_nor2_1 _1618_ (.A(_0754_),
    .B(_0755_),
    .Y(_0781_));
 sg13g2_a221oi_1 _1619_ (.B2(_0780_),
    .C1(_0781_),
    .B1(_0692_),
    .A1(_0779_),
    .Y(_0782_),
    .A2(_0730_));
 sg13g2_nor2_1 _1620_ (.A(_0778_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_buf_1 _1621_ (.A(_0755_),
    .X(_0784_));
 sg13g2_nand2_1 _1622_ (.Y(_0785_),
    .A(_0779_),
    .B(_0735_));
 sg13g2_a21o_1 _1623_ (.A2(_0774_),
    .A1(net104),
    .B1(_0785_),
    .X(_0786_));
 sg13g2_and3_1 _1624_ (.X(_0787_),
    .A(net107),
    .B(_0739_),
    .C(_0740_));
 sg13g2_and2_1 _1625_ (.A(_0753_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_nor3_1 _1626_ (.A(net104),
    .B(_0774_),
    .C(_0778_),
    .Y(_0789_));
 sg13g2_a221oi_1 _1627_ (.B2(_0788_),
    .C1(_0789_),
    .B1(_0786_),
    .A1(_0777_),
    .Y(_0790_),
    .A2(_0783_));
 sg13g2_a21oi_1 _1628_ (.A1(_0745_),
    .A2(_0776_),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_inv_1 _1629_ (.Y(_0792_),
    .A(net5));
 sg13g2_buf_1 _1630_ (.A(ui_in[5]),
    .X(_0793_));
 sg13g2_inv_2 _1631_ (.Y(_0794_),
    .A(net143));
 sg13g2_nor2_1 _1632_ (.A(_0792_),
    .B(_0794_),
    .Y(_0795_));
 sg13g2_o21ai_1 _1633_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0655_),
    .A2(_0791_));
 sg13g2_buf_1 _1634_ (.A(_0012_),
    .X(_0797_));
 sg13g2_nor2_2 _1635_ (.A(net106),
    .B(net143),
    .Y(_0798_));
 sg13g2_nand2_1 _1636_ (.Y(_0799_),
    .A(net123),
    .B(_0798_));
 sg13g2_buf_2 _1637_ (.A(\u8.rcop[1] ),
    .X(_0800_));
 sg13g2_buf_1 _1638_ (.A(\u8.rcop[0] ),
    .X(_0801_));
 sg13g2_nand2_1 _1639_ (.Y(_0802_),
    .A(_0800_),
    .B(net122));
 sg13g2_nor2_1 _1640_ (.A(_0799_),
    .B(_0802_),
    .Y(_0803_));
 sg13g2_a21oi_1 _1641_ (.A1(\u8.rcop[2] ),
    .A2(_0803_),
    .Y(_0804_),
    .B1(net106));
 sg13g2_nand4_1 _1642_ (.B(\u8.rc[31] ),
    .C(\u8.rc[29] ),
    .A(_0656_),
    .Y(_0805_),
    .D(_0668_));
 sg13g2_buf_2 _1643_ (.A(_0805_),
    .X(_0806_));
 sg13g2_nand4_1 _1644_ (.B(net139),
    .C(net136),
    .A(_0664_),
    .Y(_0807_),
    .D(_0671_));
 sg13g2_buf_2 _1645_ (.A(_0807_),
    .X(_0808_));
 sg13g2_nand4_1 _1646_ (.B(\u8.rc[20] ),
    .C(_0660_),
    .A(net135),
    .Y(_0809_),
    .D(_0661_));
 sg13g2_nand4_1 _1647_ (.B(net132),
    .C(\u8.rc[17] ),
    .A(\u8.rc[19] ),
    .Y(_0810_),
    .D(_0696_));
 sg13g2_buf_1 _1648_ (.A(_0810_),
    .X(_0811_));
 sg13g2_nor4_2 _1649_ (.A(_0806_),
    .B(_0808_),
    .C(_0809_),
    .Y(_0812_),
    .D(_0811_));
 sg13g2_inv_1 _1650_ (.Y(_0813_),
    .A(\u8.hs[2] ));
 sg13g2_nand3_1 _1651_ (.B(_0698_),
    .C(net125),
    .A(\u8.hs[4] ),
    .Y(_0814_));
 sg13g2_buf_1 _1652_ (.A(_0814_),
    .X(_0815_));
 sg13g2_nor2_1 _1653_ (.A(_0813_),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_and4_1 _1654_ (.A(_0656_),
    .B(net140),
    .C(net138),
    .D(net137),
    .X(_0817_));
 sg13g2_a22oi_1 _1655_ (.Y(_0818_),
    .B1(_0817_),
    .B2(_0660_),
    .A2(_0725_),
    .A1(_0724_));
 sg13g2_buf_1 _1656_ (.A(_0818_),
    .X(_0819_));
 sg13g2_nand2_1 _1657_ (.Y(_0820_),
    .A(_0660_),
    .B(_0661_));
 sg13g2_nor3_1 _1658_ (.A(_0820_),
    .B(_0806_),
    .C(_0808_),
    .Y(_0821_));
 sg13g2_or3_1 _1659_ (.A(_0739_),
    .B(_0819_),
    .C(_0821_),
    .X(_0822_));
 sg13g2_nand3_1 _1660_ (.B(net132),
    .C(\u8.rc[17] ),
    .A(\u8.rc[19] ),
    .Y(_0823_));
 sg13g2_nor4_2 _1661_ (.A(_0806_),
    .B(_0808_),
    .C(_0823_),
    .Y(_0824_),
    .D(_0809_));
 sg13g2_a21oi_1 _1662_ (.A1(_0722_),
    .A2(net84),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_or2_1 _1663_ (.X(_0826_),
    .B(\u8.hs[2] ),
    .A(\u8.hs[3] ));
 sg13g2_nor4_2 _1664_ (.A(\u8.hs[4] ),
    .B(_0698_),
    .C(\u8.hs[1] ),
    .Y(_0827_),
    .D(_0826_));
 sg13g2_and3_1 _1665_ (.X(_0828_),
    .A(_0722_),
    .B(_0728_),
    .C(_0827_));
 sg13g2_buf_1 _1666_ (.A(_0828_),
    .X(_0829_));
 sg13g2_a221oi_1 _1667_ (.B2(net76),
    .C1(_0829_),
    .B1(_0822_),
    .A1(_0812_),
    .Y(_0830_),
    .A2(_0816_));
 sg13g2_buf_2 _1668_ (.A(_0830_),
    .X(_0831_));
 sg13g2_nor3_2 _1669_ (.A(net130),
    .B(net128),
    .C(net127),
    .Y(_0832_));
 sg13g2_nand4_1 _1670_ (.B(net84),
    .C(_0827_),
    .A(net91),
    .Y(_0833_),
    .D(_0832_));
 sg13g2_nand2_1 _1671_ (.Y(_0834_),
    .A(net128),
    .B(net127));
 sg13g2_nor3_1 _1672_ (.A(_0695_),
    .B(_0834_),
    .C(_0815_),
    .Y(_0835_));
 sg13g2_nand2_1 _1673_ (.Y(_0836_),
    .A(_0812_),
    .B(_0835_));
 sg13g2_buf_2 _1674_ (.A(_0014_),
    .X(_0837_));
 sg13g2_buf_2 _1675_ (.A(\u8.ls[0] ),
    .X(_0838_));
 sg13g2_inv_1 _1676_ (.Y(_0839_),
    .A(_0838_));
 sg13g2_buf_2 _1677_ (.A(\u8.ls[7] ),
    .X(_0840_));
 sg13g2_buf_1 _1678_ (.A(\u8.ls[3] ),
    .X(_0841_));
 sg13g2_buf_1 _1679_ (.A(\u8.ls[2] ),
    .X(_0842_));
 sg13g2_buf_1 _1680_ (.A(\u8.ls[1] ),
    .X(_0843_));
 sg13g2_buf_1 _1681_ (.A(\u8.ls[4] ),
    .X(_0844_));
 sg13g2_nor4_2 _1682_ (.A(net121),
    .B(net120),
    .C(net119),
    .Y(_0845_),
    .D(_0844_));
 sg13g2_buf_2 _1683_ (.A(\u8.ls[5] ),
    .X(_0846_));
 sg13g2_nor2_1 _1684_ (.A(_0846_),
    .B(\u8.ls[6] ),
    .Y(_0847_));
 sg13g2_nand4_1 _1685_ (.B(_0840_),
    .C(_0845_),
    .A(_0839_),
    .Y(_0848_),
    .D(_0847_));
 sg13g2_nand2_1 _1686_ (.Y(_0849_),
    .A(_0837_),
    .B(_0848_));
 sg13g2_mux2_1 _1687_ (.A0(_0833_),
    .A1(_0836_),
    .S(_0849_),
    .X(_0850_));
 sg13g2_buf_1 _1688_ (.A(_0850_),
    .X(_0851_));
 sg13g2_buf_1 _1689_ (.A(\u8.rbop[0] ),
    .X(_0852_));
 sg13g2_nand3b_1 _1690_ (.B(net57),
    .C(net118),
    .Y(_0853_),
    .A_N(_0831_));
 sg13g2_and4_1 _1691_ (.A(_0722_),
    .B(net84),
    .C(_0827_),
    .D(_0832_),
    .X(_0854_));
 sg13g2_and2_1 _1692_ (.A(_0812_),
    .B(_0835_),
    .X(_0855_));
 sg13g2_mux2_1 _1693_ (.A0(_0854_),
    .A1(_0855_),
    .S(_0849_),
    .X(_0856_));
 sg13g2_buf_1 _1694_ (.A(_0856_),
    .X(_0857_));
 sg13g2_nand3_1 _1695_ (.B(net138),
    .C(net137),
    .A(_0656_),
    .Y(_0858_));
 sg13g2_nand2_1 _1696_ (.Y(_0859_),
    .A(net140),
    .B(_0858_));
 sg13g2_a221oi_1 _1697_ (.B2(_0819_),
    .C1(_0824_),
    .B1(_0859_),
    .A1(net91),
    .Y(_0860_),
    .A2(net84));
 sg13g2_buf_1 _1698_ (.A(_0860_),
    .X(_0861_));
 sg13g2_nand2b_2 _1699_ (.Y(_0862_),
    .B(net124),
    .A_N(\u8.rbop[1] ));
 sg13g2_buf_1 _1700_ (.A(\u8.rbop[2] ),
    .X(_0863_));
 sg13g2_inv_1 _1701_ (.Y(_0864_),
    .A(net117));
 sg13g2_a221oi_1 _1702_ (.B2(net140),
    .C1(_0824_),
    .B1(_0858_),
    .A1(net91),
    .Y(_0865_),
    .A2(net84));
 sg13g2_xnor2_1 _1703_ (.Y(_0866_),
    .A(_0864_),
    .B(_0865_));
 sg13g2_nor4_2 _1704_ (.A(net56),
    .B(net65),
    .C(_0862_),
    .Y(_0867_),
    .D(_0866_));
 sg13g2_buf_1 _1705_ (.A(_0018_),
    .X(_0868_));
 sg13g2_inv_1 _1706_ (.Y(_0869_),
    .A(_0013_));
 sg13g2_a21oi_1 _1707_ (.A1(net140),
    .A2(_0858_),
    .Y(_0870_),
    .B1(net116));
 sg13g2_nand3_1 _1708_ (.B(net76),
    .C(_0870_),
    .A(_0868_),
    .Y(_0871_));
 sg13g2_buf_1 _1709_ (.A(_0871_),
    .X(_0872_));
 sg13g2_buf_1 _1710_ (.A(_0822_),
    .X(_0873_));
 sg13g2_a21oi_1 _1711_ (.A1(net65),
    .A2(net64),
    .Y(_0874_),
    .B1(net116));
 sg13g2_and2_1 _1712_ (.A(net118),
    .B(\u8.rbop[1] ),
    .X(_0875_));
 sg13g2_nand2_1 _1713_ (.Y(_0876_),
    .A(net117),
    .B(_0875_));
 sg13g2_nor3_1 _1714_ (.A(net55),
    .B(_0874_),
    .C(_0876_),
    .Y(_0877_));
 sg13g2_a21o_1 _1715_ (.A2(_0867_),
    .A1(_0853_),
    .B1(_0877_),
    .X(_0878_));
 sg13g2_nand2b_1 _1716_ (.Y(_0879_),
    .B(net57),
    .A_N(_0831_));
 sg13g2_or4_1 _1717_ (.A(net56),
    .B(net65),
    .C(_0862_),
    .D(_0866_),
    .X(_0880_));
 sg13g2_nor2_1 _1718_ (.A(net116),
    .B(_0861_),
    .Y(_0881_));
 sg13g2_buf_1 _1719_ (.A(_0870_),
    .X(_0882_));
 sg13g2_buf_1 _1720_ (.A(\u8.rbop[1] ),
    .X(_0883_));
 sg13g2_nor2b_1 _1721_ (.A(_0863_),
    .B_N(net115),
    .Y(_0884_));
 sg13g2_nand4_1 _1722_ (.B(net76),
    .C(net83),
    .A(_0868_),
    .Y(_0885_),
    .D(_0884_));
 sg13g2_a21o_1 _1723_ (.A2(_0881_),
    .A1(net57),
    .B1(_0885_),
    .X(_0886_));
 sg13g2_inv_1 _1724_ (.Y(_0887_),
    .A(net118));
 sg13g2_a221oi_1 _1725_ (.B2(_0886_),
    .C1(_0887_),
    .B1(_0880_),
    .A1(net107),
    .Y(_0888_),
    .A2(_0879_));
 sg13g2_and3_1 _1726_ (.X(_0889_),
    .A(_0861_),
    .B(net64),
    .C(_0875_));
 sg13g2_nor3_1 _1727_ (.A(net117),
    .B(net55),
    .C(_0889_),
    .Y(_0890_));
 sg13g2_nand2_1 _1728_ (.Y(_0891_),
    .A(net135),
    .B(\u8.rc[20] ));
 sg13g2_or4_1 _1729_ (.A(_0820_),
    .B(_0806_),
    .C(_0891_),
    .D(_0808_),
    .X(_0892_));
 sg13g2_nor4_2 _1730_ (.A(_0813_),
    .B(_0892_),
    .C(_0811_),
    .Y(_0893_),
    .D(_0815_));
 sg13g2_o21ai_1 _1731_ (.B1(net118),
    .Y(_0894_),
    .A1(_0829_),
    .A2(_0893_));
 sg13g2_nand3_1 _1732_ (.B(net76),
    .C(net64),
    .A(net118),
    .Y(_0895_));
 sg13g2_nor2_1 _1733_ (.A(net65),
    .B(_0862_),
    .Y(_0896_));
 sg13g2_nand4_1 _1734_ (.B(_0894_),
    .C(_0895_),
    .A(_0850_),
    .Y(_0897_),
    .D(_0896_));
 sg13g2_nor2_2 _1735_ (.A(net118),
    .B(\u8.rbop[1] ),
    .Y(_0898_));
 sg13g2_and2_1 _1736_ (.A(_0868_),
    .B(_0898_),
    .X(_0899_));
 sg13g2_buf_1 _1737_ (.A(_0899_),
    .X(_0900_));
 sg13g2_a21o_1 _1738_ (.A2(_0897_),
    .A1(_0890_),
    .B1(_0900_),
    .X(_0901_));
 sg13g2_nor2_1 _1739_ (.A(net116),
    .B(\u8.rbop[0] ),
    .Y(_0902_));
 sg13g2_nand2b_1 _1740_ (.Y(_0903_),
    .B(_0902_),
    .A_N(_0883_));
 sg13g2_a21o_1 _1741_ (.A2(_0873_),
    .A1(net57),
    .B1(_0903_),
    .X(_0904_));
 sg13g2_a21o_1 _1742_ (.A2(net84),
    .A1(net91),
    .B1(_0824_),
    .X(_0905_));
 sg13g2_buf_1 _1743_ (.A(_0905_),
    .X(_0906_));
 sg13g2_nor2_1 _1744_ (.A(_0829_),
    .B(_0893_),
    .Y(_0907_));
 sg13g2_nand4_1 _1745_ (.B(_0906_),
    .C(_0907_),
    .A(net115),
    .Y(_0908_),
    .D(_0902_));
 sg13g2_a21oi_1 _1746_ (.A1(net76),
    .A2(net83),
    .Y(_0909_),
    .B1(_0864_));
 sg13g2_nand2_1 _1747_ (.Y(_0910_),
    .A(net124),
    .B(_0859_));
 sg13g2_buf_1 _1748_ (.A(_0910_),
    .X(_0911_));
 sg13g2_nor3_1 _1749_ (.A(net117),
    .B(_0906_),
    .C(net75),
    .Y(_0912_));
 sg13g2_or2_1 _1750_ (.X(_0913_),
    .B(_0912_),
    .A(_0909_));
 sg13g2_a21oi_1 _1751_ (.A1(_0904_),
    .A2(_0908_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_nor4_1 _1752_ (.A(_0878_),
    .B(_0888_),
    .C(_0901_),
    .D(_0914_),
    .Y(_0915_));
 sg13g2_nor2_2 _1753_ (.A(net116),
    .B(_0819_),
    .Y(_0916_));
 sg13g2_nand3_1 _1754_ (.B(net83),
    .C(_0819_),
    .A(_0825_),
    .Y(_0917_));
 sg13g2_and2_1 _1755_ (.A(_0900_),
    .B(_0917_),
    .X(_0918_));
 sg13g2_nor2b_1 _1756_ (.A(_0916_),
    .B_N(_0918_),
    .Y(_0919_));
 sg13g2_nor2_2 _1757_ (.A(net5),
    .B(_0751_),
    .Y(_0920_));
 sg13g2_inv_1 _1758_ (.Y(_0921_),
    .A(_0920_));
 sg13g2_nor4_1 _1759_ (.A(net116),
    .B(net76),
    .C(_0829_),
    .D(_0893_),
    .Y(_0922_));
 sg13g2_a21oi_1 _1760_ (.A1(net65),
    .A2(net64),
    .Y(_0923_),
    .B1(_0862_));
 sg13g2_or3_1 _1761_ (.A(_0922_),
    .B(_0923_),
    .C(_0898_),
    .X(_0924_));
 sg13g2_nand2b_1 _1762_ (.Y(_0925_),
    .B(_0902_),
    .A_N(net65));
 sg13g2_o21ai_1 _1763_ (.B1(net55),
    .Y(_0926_),
    .A1(net56),
    .A2(_0925_));
 sg13g2_o21ai_1 _1764_ (.B1(net55),
    .Y(_0927_),
    .A1(_0909_),
    .A2(_0912_));
 sg13g2_o21ai_1 _1765_ (.B1(_0927_),
    .Y(_0928_),
    .A1(_0924_),
    .A2(_0926_));
 sg13g2_nand2_1 _1766_ (.Y(_0929_),
    .A(net124),
    .B(net115));
 sg13g2_or4_1 _1767_ (.A(_0856_),
    .B(net65),
    .C(_0831_),
    .D(_0929_),
    .X(_0930_));
 sg13g2_nand2_1 _1768_ (.Y(_0931_),
    .A(net124),
    .B(_0887_));
 sg13g2_and2_1 _1769_ (.A(_0860_),
    .B(net64),
    .X(_0932_));
 sg13g2_nand2_1 _1770_ (.Y(_0933_),
    .A(_0887_),
    .B(net115));
 sg13g2_o21ai_1 _1771_ (.B1(_0933_),
    .Y(_0934_),
    .A1(_0931_),
    .A2(_0932_));
 sg13g2_a21o_1 _1772_ (.A2(net64),
    .A1(_0850_),
    .B1(_0862_),
    .X(_0935_));
 sg13g2_a21oi_1 _1773_ (.A1(net115),
    .A2(_0922_),
    .Y(_0936_),
    .B1(_0887_));
 sg13g2_a221oi_1 _1774_ (.B2(_0936_),
    .C1(_0913_),
    .B1(_0935_),
    .A1(_0930_),
    .Y(_0937_),
    .A2(_0934_));
 sg13g2_nor4_1 _1775_ (.A(_0798_),
    .B(_0921_),
    .C(_0928_),
    .D(_0937_),
    .Y(_0938_));
 sg13g2_buf_1 _1776_ (.A(_0938_),
    .X(_0939_));
 sg13g2_o21ai_1 _1777_ (.B1(net42),
    .Y(_0940_),
    .A1(_0915_),
    .A2(_0919_));
 sg13g2_nand3_1 _1778_ (.B(_0804_),
    .C(_0940_),
    .A(_0796_),
    .Y(_0941_));
 sg13g2_buf_8 _1779_ (.A(_0941_),
    .X(_0942_));
 sg13g2_buf_8 _1780_ (.A(_0942_),
    .X(_0943_));
 sg13g2_o21ai_1 _1781_ (.B1(net107),
    .Y(_0944_),
    .A1(net56),
    .A2(_0831_));
 sg13g2_nand2_1 _1782_ (.Y(_0945_),
    .A(_0852_),
    .B(_0944_));
 sg13g2_nand2_1 _1783_ (.Y(_0946_),
    .A(net83),
    .B(net57));
 sg13g2_nand2_1 _1784_ (.Y(_0947_),
    .A(_0859_),
    .B(_0819_));
 sg13g2_mux2_1 _1785_ (.A0(net76),
    .A1(_0947_),
    .S(_0864_),
    .X(_0948_));
 sg13g2_nand3_1 _1786_ (.B(_0863_),
    .C(_0859_),
    .A(net115),
    .Y(_0949_));
 sg13g2_or3_1 _1787_ (.A(_0906_),
    .B(_0819_),
    .C(_0949_),
    .X(_0950_));
 sg13g2_o21ai_1 _1788_ (.B1(_0950_),
    .Y(_0951_),
    .A1(_0883_),
    .A2(_0948_));
 sg13g2_nor2_1 _1789_ (.A(net116),
    .B(net56),
    .Y(_0952_));
 sg13g2_a22oi_1 _1790_ (.Y(_0953_),
    .B1(_0951_),
    .B2(_0952_),
    .A2(_0884_),
    .A1(_0946_));
 sg13g2_nor2_1 _1791_ (.A(_0909_),
    .B(_0912_),
    .Y(_0954_));
 sg13g2_a21o_1 _1792_ (.A2(_0908_),
    .A1(_0904_),
    .B1(_0954_),
    .X(_0955_));
 sg13g2_o21ai_1 _1793_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0945_),
    .A2(_0953_));
 sg13g2_buf_2 _1794_ (.A(_0956_),
    .X(_0957_));
 sg13g2_nor2_1 _1795_ (.A(_0015_),
    .B(net55),
    .Y(_0958_));
 sg13g2_xnor2_1 _1796_ (.Y(_0959_),
    .A(_0852_),
    .B(_0944_));
 sg13g2_a21oi_2 _1797_ (.B1(_0959_),
    .Y(_0960_),
    .A2(_0886_),
    .A1(_0880_));
 sg13g2_buf_1 _1798_ (.A(\u8.ls[6] ),
    .X(_0961_));
 sg13g2_a221oi_1 _1799_ (.B2(net114),
    .C1(_0900_),
    .B1(_0960_),
    .A1(_0957_),
    .Y(_0962_),
    .A2(_0958_));
 sg13g2_nor2_2 _1800_ (.A(_0906_),
    .B(net75),
    .Y(_0963_));
 sg13g2_and2_1 _1801_ (.A(_0868_),
    .B(_0963_),
    .X(_0964_));
 sg13g2_a22oi_1 _1802_ (.Y(_0965_),
    .B1(_0935_),
    .B2(_0936_),
    .A2(_0934_),
    .A1(_0930_));
 sg13g2_nor2_1 _1803_ (.A(net56),
    .B(_0925_),
    .Y(_0966_));
 sg13g2_or3_1 _1804_ (.A(net117),
    .B(_0966_),
    .C(_0924_),
    .X(_0967_));
 sg13g2_o21ai_1 _1805_ (.B1(net117),
    .Y(_0968_),
    .A1(_0966_),
    .A2(_0924_));
 sg13g2_and4_1 _1806_ (.A(_0964_),
    .B(_0965_),
    .C(_0967_),
    .D(_0968_),
    .X(_0969_));
 sg13g2_buf_1 _1807_ (.A(_0969_),
    .X(_0970_));
 sg13g2_a21oi_1 _1808_ (.A1(net57),
    .A2(net64),
    .Y(_0971_),
    .B1(_0933_));
 sg13g2_nor3_1 _1809_ (.A(_0887_),
    .B(net115),
    .C(_0874_),
    .Y(_0972_));
 sg13g2_nor2_1 _1810_ (.A(net117),
    .B(net55),
    .Y(_0973_));
 sg13g2_o21ai_1 _1811_ (.B1(_0973_),
    .Y(_0974_),
    .A1(_0971_),
    .A2(_0972_));
 sg13g2_nor3_1 _1812_ (.A(_0887_),
    .B(net55),
    .C(_0831_),
    .Y(_0975_));
 sg13g2_nand3b_1 _1813_ (.B(_0884_),
    .C(_0975_),
    .Y(_0976_),
    .A_N(net65));
 sg13g2_nand3_1 _1814_ (.B(_0879_),
    .C(_0867_),
    .A(_0902_),
    .Y(_0977_));
 sg13g2_nand3_1 _1815_ (.B(_0976_),
    .C(_0977_),
    .A(_0974_),
    .Y(_0978_));
 sg13g2_buf_1 _1816_ (.A(_0978_),
    .X(_0979_));
 sg13g2_buf_1 _1817_ (.A(\u8.hs[2] ),
    .X(_0980_));
 sg13g2_buf_2 _1818_ (.A(_0000_),
    .X(_0981_));
 sg13g2_a221oi_1 _1819_ (.B2(_0897_),
    .C1(_0877_),
    .B1(_0890_),
    .A1(_0853_),
    .Y(_0982_),
    .A2(_0867_));
 sg13g2_buf_2 _1820_ (.A(_0982_),
    .X(_0983_));
 sg13g2_nor2b_1 _1821_ (.A(_0981_),
    .B_N(_0983_),
    .Y(_0984_));
 sg13g2_a221oi_1 _1822_ (.B2(net113),
    .C1(_0984_),
    .B1(_0979_),
    .A1(net132),
    .Y(_0985_),
    .A2(_0970_));
 sg13g2_nor2_1 _1823_ (.A(net116),
    .B(net76),
    .Y(_0986_));
 sg13g2_nand2_1 _1824_ (.Y(_0987_),
    .A(net57),
    .B(_0986_));
 sg13g2_buf_1 _1825_ (.A(_0987_),
    .X(_0988_));
 sg13g2_inv_2 _1826_ (.Y(_0989_),
    .A(_0003_));
 sg13g2_buf_1 _1827_ (.A(_0831_),
    .X(_0990_));
 sg13g2_nor2_1 _1828_ (.A(_0027_),
    .B(net52),
    .Y(_0991_));
 sg13g2_a21oi_1 _1829_ (.A1(_0989_),
    .A2(net52),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_nor2_1 _1830_ (.A(net46),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_nor2_1 _1831_ (.A(net75),
    .B(net56),
    .Y(_0994_));
 sg13g2_inv_1 _1832_ (.Y(_0995_),
    .A(_0671_));
 sg13g2_inv_1 _1833_ (.Y(_0996_),
    .A(net140));
 sg13g2_nand2_1 _1834_ (.Y(_0997_),
    .A(_0656_),
    .B(_0996_));
 sg13g2_o21ai_1 _1835_ (.B1(_0997_),
    .Y(_0998_),
    .A1(_0995_),
    .A2(net64));
 sg13g2_and2_1 _1836_ (.A(_0963_),
    .B(_0932_),
    .X(_0999_));
 sg13g2_buf_1 _1837_ (.A(_0999_),
    .X(_1000_));
 sg13g2_nand2_2 _1838_ (.Y(_1001_),
    .A(_0868_),
    .B(_0898_));
 sg13g2_a221oi_1 _1839_ (.B2(net132),
    .C1(_1001_),
    .B1(_1000_),
    .A1(_0963_),
    .Y(_1002_),
    .A2(_0998_));
 sg13g2_o21ai_1 _1840_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0981_),
    .A2(_0994_));
 sg13g2_o21ai_1 _1841_ (.B1(net42),
    .Y(_1004_),
    .A1(_0993_),
    .A2(_1003_));
 sg13g2_a21oi_1 _1842_ (.A1(_0962_),
    .A2(_0985_),
    .Y(_1005_),
    .B1(_1004_));
 sg13g2_nor2_1 _1843_ (.A(_1005_),
    .B(_0943_),
    .Y(_1006_));
 sg13g2_buf_1 _1844_ (.A(_0741_),
    .X(_1007_));
 sg13g2_buf_1 _1845_ (.A(_0774_),
    .X(_1008_));
 sg13g2_buf_1 _1846_ (.A(net51),
    .X(_1009_));
 sg13g2_nand2_1 _1847_ (.Y(_1010_),
    .A(_1007_),
    .B(net45));
 sg13g2_buf_1 _1848_ (.A(ui_in[3]),
    .X(_1011_));
 sg13g2_buf_1 _1849_ (.A(net142),
    .X(_1012_));
 sg13g2_inv_1 _1850_ (.Y(_1013_),
    .A(net112));
 sg13g2_buf_1 _1851_ (.A(_1013_),
    .X(_1014_));
 sg13g2_buf_2 _1852_ (.A(net90),
    .X(_1015_));
 sg13g2_buf_1 _1853_ (.A(net82),
    .X(_1016_));
 sg13g2_buf_1 _1854_ (.A(_0001_),
    .X(_1017_));
 sg13g2_buf_1 _1855_ (.A(net112),
    .X(_1018_));
 sg13g2_buf_1 _1856_ (.A(net103),
    .X(_1019_));
 sg13g2_and2_1 _1857_ (.A(net89),
    .B(_0006_),
    .X(_1020_));
 sg13g2_a21oi_1 _1858_ (.A1(net74),
    .A2(net111),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_buf_1 _1859_ (.A(_0753_),
    .X(_1022_));
 sg13g2_nand2_1 _1860_ (.Y(_1023_),
    .A(net102),
    .B(_0759_));
 sg13g2_nand2_1 _1861_ (.Y(_1024_),
    .A(_1021_),
    .B(_1023_));
 sg13g2_nand2_1 _1862_ (.Y(_1025_),
    .A(_0755_),
    .B(_0753_));
 sg13g2_nor2_2 _1863_ (.A(net105),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_and2_1 _1864_ (.A(_0753_),
    .B(_0758_),
    .X(_1027_));
 sg13g2_buf_1 _1865_ (.A(_1027_),
    .X(_1028_));
 sg13g2_and2_1 _1866_ (.A(net89),
    .B(net111),
    .X(_1029_));
 sg13g2_a21oi_1 _1867_ (.A1(net82),
    .A2(_0006_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_a22oi_1 _1868_ (.Y(_1031_),
    .B1(net73),
    .B2(_1030_),
    .A2(_1026_),
    .A1(_0838_));
 sg13g2_buf_1 _1869_ (.A(_0749_),
    .X(_1032_));
 sg13g2_a21oi_1 _1870_ (.A1(_1024_),
    .A2(_1031_),
    .Y(_1033_),
    .B1(net50));
 sg13g2_buf_1 _1871_ (.A(net103),
    .X(_1034_));
 sg13g2_buf_1 _1872_ (.A(_1034_),
    .X(_1035_));
 sg13g2_buf_2 _1873_ (.A(_0002_),
    .X(_1036_));
 sg13g2_nand2_2 _1874_ (.Y(_1037_),
    .A(_0753_),
    .B(_0758_));
 sg13g2_nor2b_2 _1875_ (.A(_0735_),
    .B_N(_0755_),
    .Y(_1038_));
 sg13g2_a21oi_1 _1876_ (.A1(_0753_),
    .A2(_0758_),
    .Y(_1039_),
    .B1(_1038_));
 sg13g2_buf_1 _1877_ (.A(_1039_),
    .X(_1040_));
 sg13g2_buf_1 _1878_ (.A(_0696_),
    .X(_1041_));
 sg13g2_nor2_1 _1879_ (.A(net126),
    .B(net101),
    .Y(_1042_));
 sg13g2_xnor2_1 _1880_ (.Y(_1043_),
    .A(_0008_),
    .B(_1042_));
 sg13g2_nand2_1 _1881_ (.Y(_1044_),
    .A(net72),
    .B(_1043_));
 sg13g2_o21ai_1 _1882_ (.B1(_1044_),
    .Y(_1045_),
    .A1(_1036_),
    .A2(_1037_));
 sg13g2_and2_1 _1883_ (.A(net102),
    .B(_1038_),
    .X(_1046_));
 sg13g2_nor2_1 _1884_ (.A(_1013_),
    .B(net105),
    .Y(_1047_));
 sg13g2_nor2_1 _1885_ (.A(net112),
    .B(_0779_),
    .Y(_1048_));
 sg13g2_nor2_2 _1886_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nand2b_1 _1887_ (.Y(_1050_),
    .B(_1049_),
    .A_N(_0981_));
 sg13g2_o21ai_1 _1888_ (.B1(_1050_),
    .Y(_1051_),
    .A1(net111),
    .A2(_1049_));
 sg13g2_buf_1 _1889_ (.A(net89),
    .X(_1052_));
 sg13g2_inv_1 _1890_ (.Y(_1053_),
    .A(_1036_));
 sg13g2_a22oi_1 _1891_ (.Y(_1054_),
    .B1(_1043_),
    .B2(net73),
    .A2(net72),
    .A1(_1053_));
 sg13g2_nor2_1 _1892_ (.A(net80),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_a221oi_1 _1893_ (.B2(_1051_),
    .C1(_1055_),
    .B1(_1046_),
    .A1(net81),
    .Y(_1056_),
    .A2(_1045_));
 sg13g2_nor2_1 _1894_ (.A(net63),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nand2_2 _1895_ (.Y(_1058_),
    .A(net107),
    .B(_0768_));
 sg13g2_xnor2_1 _1896_ (.Y(_1059_),
    .A(net103),
    .B(_1028_));
 sg13g2_mux2_1 _1897_ (.A0(net111),
    .A1(_0981_),
    .S(_1059_),
    .X(_1060_));
 sg13g2_nor2_1 _1898_ (.A(_1058_),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_nor3_1 _1899_ (.A(_1033_),
    .B(_1057_),
    .C(_1061_),
    .Y(_1062_));
 sg13g2_o21ai_1 _1900_ (.B1(_1062_),
    .Y(_1063_),
    .A1(_0981_),
    .A2(_1010_));
 sg13g2_nor3_2 _1901_ (.A(_0798_),
    .B(_0920_),
    .C(_0790_),
    .Y(_1064_));
 sg13g2_nor2b_2 _1902_ (.A(_0800_),
    .B_N(net122),
    .Y(_1065_));
 sg13g2_nor2b_1 _1903_ (.A(net122),
    .B_N(_0800_),
    .Y(_1066_));
 sg13g2_buf_2 _1904_ (.A(_1066_),
    .X(_1067_));
 sg13g2_a22oi_1 _1905_ (.Y(_1068_),
    .B1(_1030_),
    .B2(_1067_),
    .A2(_1021_),
    .A1(_1065_));
 sg13g2_nand2b_1 _1906_ (.Y(_1069_),
    .B(net123),
    .A_N(_1068_));
 sg13g2_or2_1 _1907_ (.X(_1070_),
    .B(_0802_),
    .A(\u8.rcop[2] ));
 sg13g2_inv_1 _1908_ (.Y(_1071_),
    .A(_1070_));
 sg13g2_buf_1 _1909_ (.A(_1052_),
    .X(_1072_));
 sg13g2_nand2_1 _1910_ (.Y(_1073_),
    .A(_0838_),
    .B(net81));
 sg13g2_o21ai_1 _1911_ (.B1(_1073_),
    .Y(_1074_),
    .A1(_0995_),
    .A2(net71));
 sg13g2_inv_1 _1912_ (.Y(_1075_),
    .A(net123));
 sg13g2_nand2b_1 _1913_ (.Y(_1076_),
    .B(net122),
    .A_N(_0800_));
 sg13g2_nor2b_1 _1914_ (.A(\u8.rcop[2] ),
    .B_N(net122),
    .Y(_1077_));
 sg13g2_nor2b_1 _1915_ (.A(net122),
    .B_N(net123),
    .Y(_1078_));
 sg13g2_o21ai_1 _1916_ (.B1(_0800_),
    .Y(_1079_),
    .A1(_1077_),
    .A2(_1078_));
 sg13g2_o21ai_1 _1917_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1075_),
    .A2(_1076_));
 sg13g2_inv_2 _1918_ (.Y(_1081_),
    .A(_1080_));
 sg13g2_buf_1 _1919_ (.A(net81),
    .X(_1082_));
 sg13g2_nor2b_1 _1920_ (.A(_1019_),
    .B_N(_0981_),
    .Y(_1083_));
 sg13g2_a21oi_1 _1921_ (.A1(net70),
    .A2(_0015_),
    .Y(_1084_),
    .B1(_1083_));
 sg13g2_a22oi_1 _1922_ (.Y(_1085_),
    .B1(_1081_),
    .B2(_1084_),
    .A2(_1074_),
    .A1(_1071_));
 sg13g2_nor2_1 _1923_ (.A(_0800_),
    .B(net122),
    .Y(_1086_));
 sg13g2_a21o_1 _1924_ (.A2(_1086_),
    .A1(\u8.rcop[2] ),
    .B1(_0799_),
    .X(_1087_));
 sg13g2_buf_2 _1925_ (.A(_1087_),
    .X(_1088_));
 sg13g2_a21oi_1 _1926_ (.A1(_1069_),
    .A2(_1085_),
    .Y(_1089_),
    .B1(_1088_));
 sg13g2_a21oi_1 _1927_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1090_),
    .B1(_1089_));
 sg13g2_nand2_1 _1928_ (.Y(_1091_),
    .A(net2),
    .B(net1));
 sg13g2_buf_1 _1929_ (.A(_1091_),
    .X(_1092_));
 sg13g2_a221oi_1 _1930_ (.B2(_1090_),
    .C1(net110),
    .B1(_1006_),
    .A1(_0654_),
    .Y(_0036_),
    .A2(net38));
 sg13g2_inv_1 _1931_ (.Y(_1093_),
    .A(net22));
 sg13g2_buf_2 _1932_ (.A(_0030_),
    .X(_1094_));
 sg13g2_buf_1 _1933_ (.A(_0730_),
    .X(_1095_));
 sg13g2_buf_1 _1934_ (.A(_0022_),
    .X(_1096_));
 sg13g2_nand2b_1 _1935_ (.Y(_1097_),
    .B(_1059_),
    .A_N(_1094_));
 sg13g2_o21ai_1 _1936_ (.B1(_1097_),
    .Y(_1098_),
    .A1(net109),
    .A2(_1059_));
 sg13g2_buf_2 _1937_ (.A(_0007_),
    .X(_1099_));
 sg13g2_nand2_1 _1938_ (.Y(_1100_),
    .A(_0764_),
    .B(net102));
 sg13g2_nand2_1 _1939_ (.Y(_1101_),
    .A(net89),
    .B(_0784_));
 sg13g2_o21ai_1 _1940_ (.B1(_1101_),
    .Y(_1102_),
    .A1(net88),
    .A2(_1100_));
 sg13g2_o21ai_1 _1941_ (.B1(net102),
    .Y(_1103_),
    .A1(net105),
    .A2(net104));
 sg13g2_a22oi_1 _1942_ (.Y(_1104_),
    .B1(_1103_),
    .B2(net80),
    .A2(_1102_),
    .A1(_0761_));
 sg13g2_nand2_1 _1943_ (.Y(_1105_),
    .A(net90),
    .B(_0784_));
 sg13g2_o21ai_1 _1944_ (.B1(_1105_),
    .Y(_1106_),
    .A1(net90),
    .A2(_1100_));
 sg13g2_a22oi_1 _1945_ (.Y(_1107_),
    .B1(_1106_),
    .B2(_0761_),
    .A2(_1103_),
    .A1(net82));
 sg13g2_nor2_1 _1946_ (.A(net109),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_a21oi_1 _1947_ (.A1(net119),
    .A2(_1026_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_o21ai_1 _1948_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_1099_),
    .A2(_1104_));
 sg13g2_buf_2 _1949_ (.A(_0029_),
    .X(_1111_));
 sg13g2_buf_2 _1950_ (.A(_0031_),
    .X(_1112_));
 sg13g2_nor3_1 _1951_ (.A(net132),
    .B(net126),
    .C(_0696_),
    .Y(_1113_));
 sg13g2_xnor2_1 _1952_ (.Y(_1114_),
    .A(_1112_),
    .B(_1113_));
 sg13g2_nand2_1 _1953_ (.Y(_1115_),
    .A(net72),
    .B(_1114_));
 sg13g2_o21ai_1 _1954_ (.B1(_1115_),
    .Y(_1116_),
    .A1(_1111_),
    .A2(_1037_));
 sg13g2_nand2b_1 _1955_ (.Y(_1117_),
    .B(_1049_),
    .A_N(_1094_));
 sg13g2_o21ai_1 _1956_ (.B1(_1117_),
    .Y(_1118_),
    .A1(net109),
    .A2(_1049_));
 sg13g2_inv_2 _1957_ (.Y(_1119_),
    .A(_1111_));
 sg13g2_a22oi_1 _1958_ (.Y(_1120_),
    .B1(_1114_),
    .B2(net73),
    .A2(net72),
    .A1(_1119_));
 sg13g2_nor2_1 _1959_ (.A(_1052_),
    .B(_1120_),
    .Y(_1121_));
 sg13g2_a221oi_1 _1960_ (.B2(_1046_),
    .C1(_1121_),
    .B1(_1118_),
    .A1(net81),
    .Y(_1122_),
    .A2(_1116_));
 sg13g2_nor2_1 _1961_ (.A(net63),
    .B(_1122_),
    .Y(_1123_));
 sg13g2_a221oi_1 _1962_ (.B2(_0750_),
    .C1(_1123_),
    .B1(_1110_),
    .A1(net62),
    .Y(_1124_),
    .A2(_1098_));
 sg13g2_o21ai_1 _1963_ (.B1(_1124_),
    .Y(_1125_),
    .A1(_1094_),
    .A2(_1010_));
 sg13g2_mux2_1 _1964_ (.A0(_0670_),
    .A1(net119),
    .S(net81),
    .X(_1126_));
 sg13g2_inv_1 _1965_ (.Y(_1127_),
    .A(_0682_));
 sg13g2_nor2_1 _1966_ (.A(net88),
    .B(_1094_),
    .Y(_1128_));
 sg13g2_a21o_1 _1967_ (.A2(net71),
    .A1(_1127_),
    .B1(_1128_),
    .X(_1129_));
 sg13g2_and2_1 _1968_ (.A(net88),
    .B(_1099_),
    .X(_1130_));
 sg13g2_a21oi_1 _1969_ (.A1(net109),
    .A2(net74),
    .Y(_1131_),
    .B1(_1130_));
 sg13g2_buf_1 _1970_ (.A(_1018_),
    .X(_1132_));
 sg13g2_and2_1 _1971_ (.A(net109),
    .B(net87),
    .X(_1133_));
 sg13g2_a21oi_1 _1972_ (.A1(net74),
    .A2(_1099_),
    .Y(_1134_),
    .B1(_1133_));
 sg13g2_a22oi_1 _1973_ (.Y(_1135_),
    .B1(_1134_),
    .B2(_1067_),
    .A2(_1131_),
    .A1(_1065_));
 sg13g2_nor2_1 _1974_ (.A(_1075_),
    .B(_1135_),
    .Y(_1136_));
 sg13g2_a221oi_1 _1975_ (.B2(_1081_),
    .C1(_1136_),
    .B1(_1129_),
    .A1(_1071_),
    .Y(_1137_),
    .A2(_1126_));
 sg13g2_nor2_1 _1976_ (.A(_1088_),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_a21oi_1 _1977_ (.A1(_1064_),
    .A2(_1125_),
    .Y(_1139_),
    .B1(_1138_));
 sg13g2_buf_1 _1978_ (.A(_0840_),
    .X(_1140_));
 sg13g2_nor2_1 _1979_ (.A(_0682_),
    .B(net55),
    .Y(_1141_));
 sg13g2_a22oi_1 _1980_ (.Y(_1142_),
    .B1(_1141_),
    .B2(_0957_),
    .A2(_0960_),
    .A1(net100));
 sg13g2_or2_1 _1981_ (.X(_1143_),
    .B(_0983_),
    .A(_0900_));
 sg13g2_buf_1 _1982_ (.A(_1143_),
    .X(_1144_));
 sg13g2_a221oi_1 _1983_ (.B2(net125),
    .C1(_1144_),
    .B1(_0979_),
    .A1(net133),
    .Y(_1145_),
    .A2(_0970_));
 sg13g2_inv_2 _1984_ (.Y(_1146_),
    .A(_0710_));
 sg13g2_nand2_1 _1985_ (.Y(_1147_),
    .A(_1146_),
    .B(net52));
 sg13g2_o21ai_1 _1986_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_0837_),
    .A2(_0990_));
 sg13g2_nand2_1 _1987_ (.Y(_1149_),
    .A(net107),
    .B(_0906_));
 sg13g2_nor2_1 _1988_ (.A(net56),
    .B(_1149_),
    .Y(_1150_));
 sg13g2_or2_1 _1989_ (.X(_1151_),
    .B(_0821_),
    .A(_0739_));
 sg13g2_nor2b_1 _1990_ (.A(_1151_),
    .B_N(_0916_),
    .Y(_1152_));
 sg13g2_a21o_1 _1991_ (.A2(_1152_),
    .A1(_0670_),
    .B1(_1001_),
    .X(_1153_));
 sg13g2_a221oi_1 _1992_ (.B2(_1150_),
    .C1(_1153_),
    .B1(_1148_),
    .A1(net133),
    .Y(_1154_),
    .A2(_1000_));
 sg13g2_a21o_1 _1993_ (.A2(_1154_),
    .A1(_0994_),
    .B1(_1094_),
    .X(_1155_));
 sg13g2_a21o_1 _1994_ (.A2(_0983_),
    .A1(_1001_),
    .B1(_1154_),
    .X(_1156_));
 sg13g2_nor2_1 _1995_ (.A(_0928_),
    .B(_0937_),
    .Y(_1157_));
 sg13g2_nand4_1 _1996_ (.B(net144),
    .C(_0793_),
    .A(_0792_),
    .Y(_1158_),
    .D(_1157_));
 sg13g2_a221oi_1 _1997_ (.B2(_1156_),
    .C1(_1158_),
    .B1(_1155_),
    .A1(_1142_),
    .Y(_1159_),
    .A2(_1145_));
 sg13g2_nor2_1 _1998_ (.A(_0942_),
    .B(_1159_),
    .Y(_1160_));
 sg13g2_a221oi_1 _1999_ (.B2(_1160_),
    .C1(net110),
    .B1(_1139_),
    .A1(_1093_),
    .Y(_0037_),
    .A2(net38));
 sg13g2_inv_1 _2000_ (.Y(_1161_),
    .A(net23));
 sg13g2_a21oi_1 _2001_ (.A1(_1059_),
    .A2(_0721_),
    .Y(_1162_),
    .B1(net51));
 sg13g2_or2_1 _2002_ (.X(_1163_),
    .B(_1162_),
    .A(_0787_));
 sg13g2_and2_1 _2003_ (.A(net89),
    .B(_0008_),
    .X(_1164_));
 sg13g2_a21oi_1 _2004_ (.A1(net82),
    .A2(_1036_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_nand2_1 _2005_ (.Y(_1166_),
    .A(_1023_),
    .B(_1165_));
 sg13g2_nor2_1 _2006_ (.A(net82),
    .B(_1053_),
    .Y(_1167_));
 sg13g2_a21oi_1 _2007_ (.A1(net82),
    .A2(_0008_),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_a22oi_1 _2008_ (.Y(_1169_),
    .B1(net73),
    .B2(_1168_),
    .A2(_1026_),
    .A1(net120));
 sg13g2_a21oi_1 _2009_ (.A1(_1166_),
    .A2(_1169_),
    .Y(_1170_),
    .B1(net50));
 sg13g2_nor3_1 _2010_ (.A(_1036_),
    .B(_1058_),
    .C(_1059_),
    .Y(_1171_));
 sg13g2_a21oi_1 _2011_ (.A1(net113),
    .A2(_0758_),
    .Y(_1172_),
    .B1(_0756_));
 sg13g2_o21ai_1 _2012_ (.B1(net104),
    .Y(_1173_),
    .A1(net120),
    .A2(_1048_));
 sg13g2_o21ai_1 _2013_ (.B1(_1173_),
    .Y(_1174_),
    .A1(net74),
    .A2(_1172_));
 sg13g2_nor2b_1 _2014_ (.A(net72),
    .B_N(net102),
    .Y(_1175_));
 sg13g2_nand2_1 _2015_ (.Y(_1176_),
    .A(_1174_),
    .B(_1175_));
 sg13g2_nand3_1 _2016_ (.B(net74),
    .C(net72),
    .A(net113),
    .Y(_1177_));
 sg13g2_a21oi_1 _2017_ (.A1(_1176_),
    .A2(_1177_),
    .Y(_1178_),
    .B1(net63));
 sg13g2_nor3_1 _2018_ (.A(_1170_),
    .B(_1171_),
    .C(_1178_),
    .Y(_1179_));
 sg13g2_o21ai_1 _2019_ (.B1(_1179_),
    .Y(_1180_),
    .A1(_0023_),
    .A2(_1163_));
 sg13g2_a22oi_1 _2020_ (.Y(_1181_),
    .B1(_1168_),
    .B2(_1067_),
    .A2(_1165_),
    .A1(_1065_));
 sg13g2_nand2b_1 _2021_ (.Y(_1182_),
    .B(net123),
    .A_N(_1181_));
 sg13g2_inv_1 _2022_ (.Y(_1183_),
    .A(_0661_));
 sg13g2_nand2_1 _2023_ (.Y(_1184_),
    .A(net120),
    .B(net81));
 sg13g2_o21ai_1 _2024_ (.B1(_1184_),
    .Y(_1185_),
    .A1(_1183_),
    .A2(net71));
 sg13g2_inv_1 _2025_ (.Y(_1186_),
    .A(_0023_));
 sg13g2_nor2_1 _2026_ (.A(_1186_),
    .B(net89),
    .Y(_1187_));
 sg13g2_a21oi_1 _2027_ (.A1(net70),
    .A2(_0016_),
    .Y(_1188_),
    .B1(_1187_));
 sg13g2_a22oi_1 _2028_ (.Y(_1189_),
    .B1(_1188_),
    .B2(_1081_),
    .A2(_1185_),
    .A1(_1071_));
 sg13g2_a21oi_1 _2029_ (.A1(_1182_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1088_));
 sg13g2_a21oi_1 _2030_ (.A1(_1064_),
    .A2(_1180_),
    .Y(_1191_),
    .B1(_1190_));
 sg13g2_nor2_1 _2031_ (.A(_0016_),
    .B(_0872_),
    .Y(_1192_));
 sg13g2_a22oi_1 _2032_ (.Y(_1193_),
    .B1(_1192_),
    .B2(_0957_),
    .A2(_0960_),
    .A1(net127));
 sg13g2_a221oi_1 _2033_ (.B2(net129),
    .C1(_1144_),
    .B1(_0979_),
    .A1(net134),
    .Y(_1194_),
    .A2(_0970_));
 sg13g2_a22oi_1 _2034_ (.Y(_1195_),
    .B1(_1152_),
    .B2(_0661_),
    .A2(_1000_),
    .A1(net134));
 sg13g2_nand2b_1 _2035_ (.Y(_1196_),
    .B(net111),
    .A_N(_0990_));
 sg13g2_buf_2 _2036_ (.A(_0004_),
    .X(_1197_));
 sg13g2_nand2_1 _2037_ (.Y(_1198_),
    .A(_1197_),
    .B(net52));
 sg13g2_nand3_1 _2038_ (.B(_1196_),
    .C(_1198_),
    .A(_1150_),
    .Y(_1199_));
 sg13g2_nand3_1 _2039_ (.B(_1195_),
    .C(_1199_),
    .A(_0918_),
    .Y(_1200_));
 sg13g2_o21ai_1 _2040_ (.B1(_1186_),
    .Y(_1201_),
    .A1(_0946_),
    .A2(_1200_));
 sg13g2_nand2_1 _2041_ (.Y(_1202_),
    .A(_1001_),
    .B(_0983_));
 sg13g2_nand2_1 _2042_ (.Y(_1203_),
    .A(_1202_),
    .B(_1200_));
 sg13g2_a221oi_1 _2043_ (.B2(_1203_),
    .C1(_1158_),
    .B1(_1201_),
    .A1(_1193_),
    .Y(_1204_),
    .A2(_1194_));
 sg13g2_nor2_1 _2044_ (.A(_0942_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_a221oi_1 _2045_ (.B2(_1205_),
    .C1(net110),
    .B1(_1191_),
    .A1(_1161_),
    .Y(_0038_),
    .A2(net38));
 sg13g2_inv_1 _2046_ (.Y(_1206_),
    .A(net24));
 sg13g2_inv_1 _2047_ (.Y(_1207_),
    .A(_1088_));
 sg13g2_and2_1 _2048_ (.A(net121),
    .B(net71),
    .X(_1208_));
 sg13g2_a21oi_1 _2049_ (.A1(_0660_),
    .A2(net74),
    .Y(_1209_),
    .B1(_1208_));
 sg13g2_nand2_1 _2050_ (.Y(_1210_),
    .A(net87),
    .B(_1112_));
 sg13g2_o21ai_1 _2051_ (.B1(_1210_),
    .Y(_1211_),
    .A1(net80),
    .A2(_1119_));
 sg13g2_inv_1 _2052_ (.Y(_1212_),
    .A(_1112_));
 sg13g2_mux2_1 _2053_ (.A0(_1119_),
    .A1(_1212_),
    .S(net82),
    .X(_1213_));
 sg13g2_nand2_1 _2054_ (.Y(_1214_),
    .A(_1067_),
    .B(_1213_));
 sg13g2_o21ai_1 _2055_ (.B1(_1214_),
    .Y(_1215_),
    .A1(_1076_),
    .A2(_1211_));
 sg13g2_nor2b_1 _2056_ (.A(_1019_),
    .B_N(_0024_),
    .Y(_1216_));
 sg13g2_a21oi_1 _2057_ (.A1(net71),
    .A2(_0017_),
    .Y(_1217_),
    .B1(_1216_));
 sg13g2_a22oi_1 _2058_ (.Y(_1218_),
    .B1(_1217_),
    .B2(_1081_),
    .A2(_1215_),
    .A1(net123));
 sg13g2_o21ai_1 _2059_ (.B1(_1218_),
    .Y(_1219_),
    .A1(_1070_),
    .A2(_1209_));
 sg13g2_and3_1 _2060_ (.X(_1220_),
    .A(net107),
    .B(_0739_),
    .C(_0740_));
 sg13g2_buf_1 _2061_ (.A(_1220_),
    .X(_1221_));
 sg13g2_or2_1 _2062_ (.X(_1222_),
    .B(_1048_),
    .A(_1047_));
 sg13g2_o21ai_1 _2063_ (.B1(_1022_),
    .Y(_1223_),
    .A1(net121),
    .A2(_1222_));
 sg13g2_and2_1 _2064_ (.A(net90),
    .B(_1040_),
    .X(_1224_));
 sg13g2_a21oi_1 _2065_ (.A1(net89),
    .A2(_1028_),
    .Y(_1225_),
    .B1(_1224_));
 sg13g2_nor2_1 _2066_ (.A(net125),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_a21oi_1 _2067_ (.A1(_1038_),
    .A2(_1223_),
    .Y(_1227_),
    .B1(_1226_));
 sg13g2_a22oi_1 _2068_ (.Y(_1228_),
    .B1(net73),
    .B2(_1213_),
    .A2(_1026_),
    .A1(net121));
 sg13g2_o21ai_1 _2069_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_0760_),
    .A2(_1211_));
 sg13g2_nor3_1 _2070_ (.A(_1111_),
    .B(_1058_),
    .C(_1059_),
    .Y(_1230_));
 sg13g2_a221oi_1 _2071_ (.B2(_0750_),
    .C1(_1230_),
    .B1(_1229_),
    .A1(net61),
    .Y(_1231_),
    .A2(_1227_));
 sg13g2_o21ai_1 _2072_ (.B1(_1231_),
    .Y(_1232_),
    .A1(_0024_),
    .A2(_1163_));
 sg13g2_a22oi_1 _2073_ (.Y(_1233_),
    .B1(_1232_),
    .B2(_1064_),
    .A2(_1219_),
    .A1(_1207_));
 sg13g2_nor2_1 _2074_ (.A(_0017_),
    .B(_0872_),
    .Y(_1234_));
 sg13g2_a22oi_1 _2075_ (.Y(_1235_),
    .B1(_1234_),
    .B2(_0957_),
    .A2(_0960_),
    .A1(net128));
 sg13g2_buf_1 _2076_ (.A(_0698_),
    .X(_1236_));
 sg13g2_a221oi_1 _2077_ (.B2(net99),
    .C1(_1144_),
    .B1(_0979_),
    .A1(net135),
    .Y(_1237_),
    .A2(_0970_));
 sg13g2_inv_1 _2078_ (.Y(_1238_),
    .A(_0005_));
 sg13g2_nand2_1 _2079_ (.Y(_1239_),
    .A(_1238_),
    .B(net52));
 sg13g2_o21ai_1 _2080_ (.B1(_1239_),
    .Y(_1240_),
    .A1(net109),
    .A2(net52));
 sg13g2_nand2b_1 _2081_ (.Y(_1241_),
    .B(_0916_),
    .A_N(_1151_));
 sg13g2_nand2_1 _2082_ (.Y(_1242_),
    .A(_0918_),
    .B(_1241_));
 sg13g2_a221oi_1 _2083_ (.B2(_1150_),
    .C1(_1242_),
    .B1(_1240_),
    .A1(net135),
    .Y(_1243_),
    .A2(_1000_));
 sg13g2_a21o_1 _2084_ (.A2(_1243_),
    .A1(_0994_),
    .B1(_0024_),
    .X(_1244_));
 sg13g2_a21o_1 _2085_ (.A2(_0983_),
    .A1(_1001_),
    .B1(_1243_),
    .X(_1245_));
 sg13g2_a221oi_1 _2086_ (.B2(_1245_),
    .C1(_1158_),
    .B1(_1244_),
    .A1(_1235_),
    .Y(_1246_),
    .A2(_1237_));
 sg13g2_nor2_1 _2087_ (.A(_0942_),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_a221oi_1 _2088_ (.B2(_1247_),
    .C1(_1092_),
    .B1(_1233_),
    .A1(_1206_),
    .Y(_0039_),
    .A2(net38));
 sg13g2_buf_1 _2089_ (.A(net1),
    .X(_1248_));
 sg13g2_nand3_1 _2090_ (.B(net141),
    .C(net25),
    .A(net2),
    .Y(_1249_));
 sg13g2_nand4_1 _2091_ (.B(net137),
    .C(_0964_),
    .A(_0996_),
    .Y(_1250_),
    .D(_0957_));
 sg13g2_inv_1 _2092_ (.Y(_1251_),
    .A(_0009_));
 sg13g2_mux2_1 _2093_ (.A0(_0989_),
    .A1(_1251_),
    .S(net112),
    .X(_1252_));
 sg13g2_nand2_1 _2094_ (.Y(_1253_),
    .A(_1023_),
    .B(_1252_));
 sg13g2_buf_1 _2095_ (.A(_0844_),
    .X(_1254_));
 sg13g2_mux2_1 _2096_ (.A0(_0989_),
    .A1(_1251_),
    .S(net90),
    .X(_1255_));
 sg13g2_a22oi_1 _2097_ (.Y(_1256_),
    .B1(net73),
    .B2(_1255_),
    .A2(_1026_),
    .A1(net98));
 sg13g2_nand2_1 _2098_ (.Y(_1257_),
    .A(_1253_),
    .B(_1256_));
 sg13g2_o21ai_1 _2099_ (.B1(_0756_),
    .Y(_1258_),
    .A1(_0844_),
    .A2(net112));
 sg13g2_o21ai_1 _2100_ (.B1(_0758_),
    .Y(_1259_),
    .A1(net129),
    .A2(_1014_));
 sg13g2_nand2_1 _2101_ (.Y(_1260_),
    .A(_1258_),
    .B(_1259_));
 sg13g2_nor2_1 _2102_ (.A(_0844_),
    .B(_1014_),
    .Y(_1261_));
 sg13g2_o21ai_1 _2103_ (.B1(_1038_),
    .Y(_1262_),
    .A1(_0765_),
    .A2(_1261_));
 sg13g2_a22oi_1 _2104_ (.Y(_1263_),
    .B1(_1262_),
    .B2(_1037_),
    .A2(_1260_),
    .A1(net102));
 sg13g2_nor2b_1 _2105_ (.A(net129),
    .B_N(_1224_),
    .Y(_1264_));
 sg13g2_o21ai_1 _2106_ (.B1(net61),
    .Y(_1265_),
    .A1(_1263_),
    .A2(_1264_));
 sg13g2_buf_1 _2107_ (.A(_0734_),
    .X(_1266_));
 sg13g2_o21ai_1 _2108_ (.B1(net63),
    .Y(_1267_),
    .A1(_0025_),
    .A2(_1266_));
 sg13g2_a22oi_1 _2109_ (.Y(_1268_),
    .B1(_1265_),
    .B2(_1267_),
    .A2(_1257_),
    .A1(_0750_));
 sg13g2_inv_1 _2110_ (.Y(_1269_),
    .A(_0025_));
 sg13g2_mux4_1 _2111_ (.S0(net103),
    .A0(net113),
    .A1(_1254_),
    .A2(_1269_),
    .A3(_0989_),
    .S1(_1037_),
    .X(_1270_));
 sg13g2_nand3_1 _2112_ (.B(_0721_),
    .C(_1270_),
    .A(_1266_),
    .Y(_1271_));
 sg13g2_nor2_1 _2113_ (.A(net62),
    .B(_0733_),
    .Y(_1272_));
 sg13g2_nor2_1 _2114_ (.A(net104),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_inv_1 _2115_ (.Y(_1274_),
    .A(_0778_));
 sg13g2_nand2b_1 _2116_ (.Y(_1275_),
    .B(net102),
    .A_N(_0735_));
 sg13g2_a21o_1 _2117_ (.A2(_0765_),
    .A1(_1275_),
    .B1(net63),
    .X(_1276_));
 sg13g2_o21ai_1 _2118_ (.B1(_1276_),
    .Y(_1277_),
    .A1(net63),
    .A2(_1025_));
 sg13g2_a221oi_1 _2119_ (.B2(_1274_),
    .C1(_1277_),
    .B1(_1273_),
    .A1(_0777_),
    .Y(_1278_),
    .A2(_0783_));
 sg13g2_a221oi_1 _2120_ (.B2(_1271_),
    .C1(_1278_),
    .B1(_1268_),
    .A1(_0792_),
    .Y(_1279_),
    .A2(net144));
 sg13g2_a221oi_1 _2121_ (.B2(net139),
    .C1(_1279_),
    .B1(_0970_),
    .A1(net130),
    .Y(_1280_),
    .A2(_0960_));
 sg13g2_a21oi_1 _2122_ (.A1(net101),
    .A2(_0979_),
    .Y(_1281_),
    .B1(_1144_));
 sg13g2_nand3_1 _2123_ (.B(_1280_),
    .C(_1281_),
    .A(_1250_),
    .Y(_1282_));
 sg13g2_nand2_1 _2124_ (.Y(_1283_),
    .A(_0006_),
    .B(net52));
 sg13g2_o21ai_1 _2125_ (.B1(_1283_),
    .Y(_1284_),
    .A1(_1053_),
    .A2(net52));
 sg13g2_nor2_1 _2126_ (.A(_0963_),
    .B(_1001_),
    .Y(_1285_));
 sg13g2_o21ai_1 _2127_ (.B1(_1285_),
    .Y(_1286_),
    .A1(net46),
    .A2(_1284_));
 sg13g2_nand3_1 _2128_ (.B(_1285_),
    .C(_1284_),
    .A(_0994_),
    .Y(_1287_));
 sg13g2_a221oi_1 _2129_ (.B2(_1269_),
    .C1(_1279_),
    .B1(_1287_),
    .A1(_1202_),
    .Y(_1288_),
    .A2(_1286_));
 sg13g2_a21oi_1 _2130_ (.A1(_0920_),
    .A2(_1157_),
    .Y(_1289_),
    .B1(_1279_));
 sg13g2_nor4_1 _2131_ (.A(_0798_),
    .B(net110),
    .C(_1288_),
    .D(_1289_),
    .Y(_1290_));
 sg13g2_nand2_1 _2132_ (.Y(_1291_),
    .A(_1282_),
    .B(_1290_));
 sg13g2_a22oi_1 _2133_ (.Y(_1292_),
    .B1(_1255_),
    .B2(_1067_),
    .A2(_1252_),
    .A1(_1065_));
 sg13g2_nand2_1 _2134_ (.Y(_1293_),
    .A(net80),
    .B(_1081_));
 sg13g2_o21ai_1 _2135_ (.B1(_1293_),
    .Y(_1294_),
    .A1(net80),
    .A2(_1070_));
 sg13g2_nand2_1 _2136_ (.Y(_1295_),
    .A(net87),
    .B(_1071_));
 sg13g2_o21ai_1 _2137_ (.B1(_1295_),
    .Y(_1296_),
    .A1(net87),
    .A2(_1080_));
 sg13g2_a22oi_1 _2138_ (.Y(_1297_),
    .B1(_1296_),
    .B2(net98),
    .A2(_1294_),
    .A1(net137));
 sg13g2_o21ai_1 _2139_ (.B1(_1297_),
    .Y(_1298_),
    .A1(_1075_),
    .A2(_1292_));
 sg13g2_nor2_1 _2140_ (.A(_1088_),
    .B(net110),
    .Y(_1299_));
 sg13g2_a21oi_1 _2141_ (.A1(_1298_),
    .A2(_1299_),
    .Y(_1300_),
    .B1(net38));
 sg13g2_a22oi_1 _2142_ (.Y(_0040_),
    .B1(_1291_),
    .B2(_1300_),
    .A2(_1249_),
    .A1(_0943_));
 sg13g2_mux2_1 _2143_ (.A0(_0715_),
    .A1(_1146_),
    .S(net74),
    .X(_1301_));
 sg13g2_mux2_1 _2144_ (.A0(_0715_),
    .A1(_1146_),
    .S(net80),
    .X(_1302_));
 sg13g2_a22oi_1 _2145_ (.Y(_1303_),
    .B1(_1302_),
    .B2(_1067_),
    .A2(_1301_),
    .A1(_1065_));
 sg13g2_nand2b_1 _2146_ (.Y(_1304_),
    .B(net123),
    .A_N(_1303_));
 sg13g2_buf_1 _2147_ (.A(_0846_),
    .X(_1305_));
 sg13g2_a22oi_1 _2148_ (.Y(_1306_),
    .B1(_1296_),
    .B2(net97),
    .A2(_1294_),
    .A1(_0667_));
 sg13g2_a21oi_1 _2149_ (.A1(_1304_),
    .A2(_1306_),
    .Y(_1307_),
    .B1(_1088_));
 sg13g2_nor2_1 _2150_ (.A(net45),
    .B(_0777_),
    .Y(_1308_));
 sg13g2_inv_1 _2151_ (.Y(_1309_),
    .A(_0026_));
 sg13g2_mux4_1 _2152_ (.S0(net74),
    .A0(net125),
    .A1(net97),
    .A2(_1309_),
    .A3(_1146_),
    .S1(net73),
    .X(_1310_));
 sg13g2_nor2_1 _2153_ (.A(_0710_),
    .B(_1107_),
    .Y(_1311_));
 sg13g2_a21oi_1 _2154_ (.A1(net97),
    .A2(_1026_),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_o21ai_1 _2155_ (.B1(_1312_),
    .Y(_1313_),
    .A1(net131),
    .A2(_1104_));
 sg13g2_nor2_1 _2156_ (.A(_0685_),
    .B(_0719_),
    .Y(_1314_));
 sg13g2_buf_1 _2157_ (.A(_1314_),
    .X(_1315_));
 sg13g2_nor2b_1 _2158_ (.A(net80),
    .B_N(net99),
    .Y(_1316_));
 sg13g2_nand2_1 _2159_ (.Y(_1317_),
    .A(_0846_),
    .B(net104));
 sg13g2_nand3_1 _2160_ (.B(net88),
    .C(_0758_),
    .A(net99),
    .Y(_1318_));
 sg13g2_o21ai_1 _2161_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_1222_),
    .A2(_1317_));
 sg13g2_a22oi_1 _2162_ (.Y(_1320_),
    .B1(_1319_),
    .B2(_1175_),
    .A2(_1316_),
    .A1(_1040_));
 sg13g2_a21oi_1 _2163_ (.A1(_1309_),
    .A2(net51),
    .Y(_1321_),
    .B1(net61));
 sg13g2_a21oi_1 _2164_ (.A1(net61),
    .A2(_1320_),
    .Y(_1322_),
    .B1(_1321_));
 sg13g2_a221oi_1 _2165_ (.B2(net49),
    .C1(_1322_),
    .B1(_1313_),
    .A1(_1308_),
    .Y(_1323_),
    .A2(_1310_));
 sg13g2_nor2b_1 _2166_ (.A(_1323_),
    .B_N(_1064_),
    .Y(_1324_));
 sg13g2_a22oi_1 _2167_ (.Y(_1325_),
    .B1(_0979_),
    .B2(net126),
    .A2(_0970_),
    .A1(_0664_));
 sg13g2_buf_1 _2168_ (.A(\u8.hs[1] ),
    .X(_1326_));
 sg13g2_and3_1 _2169_ (.X(_1327_),
    .A(_0996_),
    .B(_0667_),
    .C(_0964_));
 sg13g2_a221oi_1 _2170_ (.B2(_0957_),
    .C1(_1144_),
    .B1(_1327_),
    .A1(net108),
    .Y(_1328_),
    .A2(_0960_));
 sg13g2_or4_1 _2171_ (.A(_1119_),
    .B(_0857_),
    .C(_1149_),
    .D(_0907_),
    .X(_1329_));
 sg13g2_o21ai_1 _2172_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1309_),
    .A2(_1150_));
 sg13g2_a221oi_1 _2173_ (.B2(_0897_),
    .C1(_1309_),
    .B1(_0890_),
    .A1(_0868_),
    .Y(_1331_),
    .A2(_0898_));
 sg13g2_a21oi_1 _2174_ (.A1(_0853_),
    .A2(_0867_),
    .Y(_1332_),
    .B1(_0877_));
 sg13g2_a22oi_1 _2175_ (.Y(_1333_),
    .B1(_1331_),
    .B2(_1332_),
    .A2(_1330_),
    .A1(_1285_));
 sg13g2_nand2_1 _2176_ (.Y(_1334_),
    .A(_0939_),
    .B(_1333_));
 sg13g2_a21oi_1 _2177_ (.A1(_1325_),
    .A2(_1328_),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_nor4_1 _2178_ (.A(_0942_),
    .B(_1307_),
    .C(_1324_),
    .D(_1335_),
    .Y(_1336_));
 sg13g2_nor2b_1 _2179_ (.A(net26),
    .B_N(net38),
    .Y(_1337_));
 sg13g2_nor3_1 _2180_ (.A(net110),
    .B(_1336_),
    .C(_1337_),
    .Y(_0041_));
 sg13g2_inv_1 _2181_ (.Y(_1338_),
    .A(net114));
 sg13g2_a21oi_1 _2182_ (.A1(_1338_),
    .A2(_0946_),
    .Y(_1339_),
    .B1(_1001_));
 sg13g2_inv_1 _2183_ (.Y(_1340_),
    .A(_1197_));
 sg13g2_nand2_1 _2184_ (.Y(_1341_),
    .A(net103),
    .B(_0010_));
 sg13g2_o21ai_1 _2185_ (.B1(_1341_),
    .Y(_1342_),
    .A1(net89),
    .A2(_1340_));
 sg13g2_nor2_1 _2186_ (.A(net90),
    .B(_1340_),
    .Y(_1343_));
 sg13g2_a21oi_1 _2187_ (.A1(net90),
    .A2(_0010_),
    .Y(_1344_),
    .B1(_1343_));
 sg13g2_a22oi_1 _2188_ (.Y(_1345_),
    .B1(net73),
    .B2(_1344_),
    .A2(_1026_),
    .A1(net114));
 sg13g2_o21ai_1 _2189_ (.B1(_1345_),
    .Y(_1346_),
    .A1(_0760_),
    .A2(_1342_));
 sg13g2_inv_1 _2190_ (.Y(_1347_),
    .A(net101));
 sg13g2_nor2_1 _2191_ (.A(_1347_),
    .B(net87),
    .Y(_1348_));
 sg13g2_a21oi_1 _2192_ (.A1(_1347_),
    .A2(_0764_),
    .Y(_1349_),
    .B1(net90));
 sg13g2_o21ai_1 _2193_ (.B1(net104),
    .Y(_1350_),
    .A1(net114),
    .A2(_1047_));
 sg13g2_o21ai_1 _2194_ (.B1(_1350_),
    .Y(_1351_),
    .A1(_0779_),
    .A2(_1349_));
 sg13g2_a21oi_1 _2195_ (.A1(net102),
    .A2(_1351_),
    .Y(_1352_),
    .B1(net72));
 sg13g2_a21oi_1 _2196_ (.A1(net72),
    .A2(_1348_),
    .Y(_1353_),
    .B1(_1352_));
 sg13g2_nor3_1 _2197_ (.A(_1197_),
    .B(_1058_),
    .C(_1059_),
    .Y(_1354_));
 sg13g2_a221oi_1 _2198_ (.B2(net61),
    .C1(_1354_),
    .B1(_1353_),
    .A1(_0750_),
    .Y(_1355_),
    .A2(_1346_));
 sg13g2_o21ai_1 _2199_ (.B1(_1355_),
    .Y(_1356_),
    .A1(_0027_),
    .A2(_1163_));
 sg13g2_nand2_1 _2200_ (.Y(_1357_),
    .A(_0656_),
    .B(_1294_));
 sg13g2_nand2_1 _2201_ (.Y(_1358_),
    .A(_1067_),
    .B(_1344_));
 sg13g2_o21ai_1 _2202_ (.B1(_1358_),
    .Y(_1359_),
    .A1(_1076_),
    .A2(_1342_));
 sg13g2_a22oi_1 _2203_ (.Y(_1360_),
    .B1(_1359_),
    .B2(_0797_),
    .A2(_1296_),
    .A1(net114));
 sg13g2_a21oi_1 _2204_ (.A1(_1357_),
    .A2(_1360_),
    .Y(_1361_),
    .B1(_1088_));
 sg13g2_a221oi_1 _2205_ (.B2(_1064_),
    .C1(_1361_),
    .B1(_1356_),
    .A1(net42),
    .Y(_1362_),
    .A2(_1339_));
 sg13g2_or2_1 _2206_ (.X(_1363_),
    .B(_1362_),
    .A(_0942_));
 sg13g2_nand2_1 _2207_ (.Y(_1364_),
    .A(net27),
    .B(net38));
 sg13g2_buf_1 _2208_ (.A(net110),
    .X(_1365_));
 sg13g2_a21oi_1 _2209_ (.A1(_1363_),
    .A2(_1364_),
    .Y(_0042_),
    .B1(net96));
 sg13g2_nand2_1 _2210_ (.Y(_1366_),
    .A(net28),
    .B(net38));
 sg13g2_inv_1 _2211_ (.Y(_1367_),
    .A(_0011_));
 sg13g2_mux2_1 _2212_ (.A0(_1238_),
    .A1(_1367_),
    .S(net103),
    .X(_1368_));
 sg13g2_nand2_1 _2213_ (.Y(_1369_),
    .A(net103),
    .B(_0005_));
 sg13g2_o21ai_1 _2214_ (.B1(_1369_),
    .Y(_1370_),
    .A1(net103),
    .A2(_1367_));
 sg13g2_nor2_1 _2215_ (.A(_1037_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_a221oi_1 _2216_ (.B2(_1368_),
    .C1(_1371_),
    .B1(_1023_),
    .A1(net100),
    .Y(_1372_),
    .A2(_1026_));
 sg13g2_xnor2_1 _2217_ (.Y(_1373_),
    .A(net126),
    .B(net101));
 sg13g2_o21ai_1 _2218_ (.B1(_1022_),
    .Y(_1374_),
    .A1(_0840_),
    .A2(_1222_));
 sg13g2_nand2_1 _2219_ (.Y(_1375_),
    .A(_1038_),
    .B(_1374_));
 sg13g2_o21ai_1 _2220_ (.B1(_1375_),
    .Y(_1376_),
    .A1(_1225_),
    .A2(_1373_));
 sg13g2_inv_1 _2221_ (.Y(_1377_),
    .A(_0837_));
 sg13g2_mux4_1 _2222_ (.S0(net112),
    .A0(_0698_),
    .A1(_0840_),
    .A2(_1377_),
    .A3(_1238_),
    .S1(_1037_),
    .X(_1378_));
 sg13g2_and2_1 _2223_ (.A(net54),
    .B(_1378_),
    .X(_1379_));
 sg13g2_a221oi_1 _2224_ (.B2(_1379_),
    .C1(_1221_),
    .B1(_0721_),
    .A1(_1377_),
    .Y(_1380_),
    .A2(_1272_));
 sg13g2_a21o_1 _2225_ (.A2(_1376_),
    .A1(net61),
    .B1(_1380_),
    .X(_1381_));
 sg13g2_o21ai_1 _2226_ (.B1(_1381_),
    .Y(_1382_),
    .A1(net50),
    .A2(_1372_));
 sg13g2_nand3_1 _2227_ (.B(net46),
    .C(_1285_),
    .A(_0837_),
    .Y(_1383_));
 sg13g2_nand2_1 _2228_ (.Y(_1384_),
    .A(net100),
    .B(net87));
 sg13g2_o21ai_1 _2229_ (.B1(_1384_),
    .Y(_1385_),
    .A1(_0996_),
    .A2(net81));
 sg13g2_nor2_1 _2230_ (.A(net82),
    .B(_0028_),
    .Y(_1386_));
 sg13g2_nor2_1 _2231_ (.A(_0837_),
    .B(net88),
    .Y(_1387_));
 sg13g2_or2_1 _2232_ (.X(_1388_),
    .B(_1387_),
    .A(_1386_));
 sg13g2_nor2_1 _2233_ (.A(_0801_),
    .B(_1370_),
    .Y(_1389_));
 sg13g2_a22oi_1 _2234_ (.Y(_1390_),
    .B1(_1389_),
    .B2(_0800_),
    .A2(_1368_),
    .A1(_1065_));
 sg13g2_nor2_1 _2235_ (.A(_1075_),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_a221oi_1 _2236_ (.B2(_1081_),
    .C1(_1391_),
    .B1(_1388_),
    .A1(_1071_),
    .Y(_1392_),
    .A2(_1385_));
 sg13g2_nor2_1 _2237_ (.A(_1088_),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_a221oi_1 _2238_ (.B2(net42),
    .C1(_1393_),
    .B1(_1383_),
    .A1(_1064_),
    .Y(_1394_),
    .A2(_1382_));
 sg13g2_or2_1 _2239_ (.X(_1395_),
    .B(_1394_),
    .A(_0942_));
 sg13g2_a21oi_1 _2240_ (.A1(_1366_),
    .A2(_1395_),
    .Y(_0043_),
    .B1(net96));
 sg13g2_inv_1 _2241_ (.Y(_1396_),
    .A(\u8.empty ));
 sg13g2_inv_1 _2242_ (.Y(_1397_),
    .A(_0655_));
 sg13g2_nand3_1 _2243_ (.B(_0739_),
    .C(_0740_),
    .A(_0746_),
    .Y(_1398_));
 sg13g2_and3_1 _2244_ (.X(_1399_),
    .A(net51),
    .B(_1398_),
    .C(_0721_));
 sg13g2_nand2_1 _2245_ (.Y(_1400_),
    .A(net5),
    .B(net143));
 sg13g2_a21oi_1 _2246_ (.A1(_1397_),
    .A2(_1399_),
    .Y(_1401_),
    .B1(_1400_));
 sg13g2_nand2_2 _2247_ (.Y(_1402_),
    .A(_0792_),
    .B(_0751_));
 sg13g2_nor3_2 _2248_ (.A(_0794_),
    .B(net75),
    .C(_1402_),
    .Y(_1403_));
 sg13g2_nand2_2 _2249_ (.Y(_1404_),
    .A(net106),
    .B(_0794_));
 sg13g2_buf_1 _2250_ (.A(\u8.rcip[0] ),
    .X(_1405_));
 sg13g2_buf_2 _2251_ (.A(\u8.rcip[2] ),
    .X(_1406_));
 sg13g2_nor3_2 _2252_ (.A(_1405_),
    .B(\u8.rcip[1] ),
    .C(_1406_),
    .Y(_1407_));
 sg13g2_nor2_2 _2253_ (.A(_1404_),
    .B(_1407_),
    .Y(_1408_));
 sg13g2_nand2_1 _2254_ (.Y(_1409_),
    .A(net106),
    .B(net2));
 sg13g2_nor4_1 _2255_ (.A(_1401_),
    .B(_1403_),
    .C(_1408_),
    .D(_1409_),
    .Y(_1410_));
 sg13g2_o21ai_1 _2256_ (.B1(net141),
    .Y(_0044_),
    .A1(_1396_),
    .A2(_1410_));
 sg13g2_xnor2_1 _2257_ (.Y(_1411_),
    .A(net118),
    .B(net42));
 sg13g2_nor2_1 _2258_ (.A(net96),
    .B(_1411_),
    .Y(_0045_));
 sg13g2_nand2_1 _2259_ (.Y(_1412_),
    .A(net118),
    .B(net42));
 sg13g2_xor2_1 _2260_ (.B(_1412_),
    .A(net115),
    .X(_1413_));
 sg13g2_nor2_1 _2261_ (.A(net96),
    .B(_1413_),
    .Y(_0046_));
 sg13g2_o21ai_1 _2262_ (.B1(net42),
    .Y(_1414_),
    .A1(_0900_),
    .A2(_0875_));
 sg13g2_and2_1 _2263_ (.A(_0864_),
    .B(_0875_),
    .X(_1415_));
 sg13g2_a22oi_1 _2264_ (.Y(_1416_),
    .B1(_1415_),
    .B2(net42),
    .A2(_1414_),
    .A1(net117));
 sg13g2_nor2_1 _2265_ (.A(net96),
    .B(_1416_),
    .Y(_0047_));
 sg13g2_buf_1 _2266_ (.A(_1272_),
    .X(_1417_));
 sg13g2_inv_1 _2267_ (.Y(_1418_),
    .A(net6));
 sg13g2_a21oi_1 _2268_ (.A1(net87),
    .A2(_1418_),
    .Y(_1419_),
    .B1(_1083_));
 sg13g2_nor2_1 _2269_ (.A(net112),
    .B(net12),
    .Y(_1420_));
 sg13g2_a21oi_1 _2270_ (.A1(net112),
    .A2(_0027_),
    .Y(_1421_),
    .B1(_1420_));
 sg13g2_nor2_1 _2271_ (.A(net8),
    .B(net142),
    .Y(_1422_));
 sg13g2_a21oi_1 _2272_ (.A1(_0023_),
    .A2(_1012_),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_nor2b_1 _2273_ (.A(_0026_),
    .B_N(net142),
    .Y(_1424_));
 sg13g2_nor2b_1 _2274_ (.A(net142),
    .B_N(net11),
    .Y(_1425_));
 sg13g2_nor2_1 _2275_ (.A(_1011_),
    .B(net9),
    .Y(_1426_));
 sg13g2_and2_1 _2276_ (.A(net142),
    .B(_0024_),
    .X(_1427_));
 sg13g2_nor4_1 _2277_ (.A(_1424_),
    .B(_1425_),
    .C(_1426_),
    .D(_1427_),
    .Y(_1428_));
 sg13g2_buf_2 _2278_ (.A(uio_in[7]),
    .X(_1429_));
 sg13g2_nand2b_1 _2279_ (.Y(_1430_),
    .B(_1429_),
    .A_N(net142));
 sg13g2_nand2b_1 _2280_ (.Y(_1431_),
    .B(net142),
    .A_N(_0837_));
 sg13g2_nor2_1 _2281_ (.A(net142),
    .B(net10),
    .Y(_1432_));
 sg13g2_a221oi_1 _2282_ (.B2(_1431_),
    .C1(_1432_),
    .B1(_1430_),
    .A1(_1012_),
    .Y(_1433_),
    .A2(_0025_));
 sg13g2_and4_1 _2283_ (.A(_1421_),
    .B(_1423_),
    .C(_1428_),
    .D(_1433_),
    .X(_1434_));
 sg13g2_buf_1 _2284_ (.A(_1434_),
    .X(_1435_));
 sg13g2_buf_1 _2285_ (.A(_1435_),
    .X(_1436_));
 sg13g2_buf_1 _2286_ (.A(net60),
    .X(_1437_));
 sg13g2_buf_1 _2287_ (.A(_1435_),
    .X(_1438_));
 sg13g2_nand2_1 _2288_ (.Y(_1439_),
    .A(_1419_),
    .B(net59));
 sg13g2_o21ai_1 _2289_ (.B1(_1439_),
    .Y(_1440_),
    .A1(net111),
    .A2(net53));
 sg13g2_a22oi_1 _2290_ (.Y(_1441_),
    .B1(_1440_),
    .B2(net49),
    .A2(_1419_),
    .A1(net48));
 sg13g2_nor2_2 _2291_ (.A(net61),
    .B(_0777_),
    .Y(_1442_));
 sg13g2_nor2_1 _2292_ (.A(net5),
    .B(net144),
    .Y(_1443_));
 sg13g2_buf_1 _2293_ (.A(_1443_),
    .X(_1444_));
 sg13g2_a21oi_1 _2294_ (.A1(net51),
    .A2(_1442_),
    .Y(_1445_),
    .B1(net95));
 sg13g2_buf_1 _2295_ (.A(_1445_),
    .X(_1446_));
 sg13g2_nand2_1 _2296_ (.Y(_1447_),
    .A(_1404_),
    .B(net44));
 sg13g2_nor2_2 _2297_ (.A(net144),
    .B(net143),
    .Y(_1448_));
 sg13g2_nand2b_1 _2298_ (.Y(_1449_),
    .B(_1448_),
    .A_N(_1407_));
 sg13g2_buf_1 _2299_ (.A(_1449_),
    .X(_1450_));
 sg13g2_inv_1 _2300_ (.Y(_1451_),
    .A(\u8.rcip[1] ));
 sg13g2_nor2_2 _2301_ (.A(_1451_),
    .B(_1406_),
    .Y(_1452_));
 sg13g2_nor2_2 _2302_ (.A(net79),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_inv_1 _2303_ (.Y(_1454_),
    .A(_1405_));
 sg13g2_nand2b_1 _2304_ (.Y(_1455_),
    .B(\u8.rcip[1] ),
    .A_N(_1406_));
 sg13g2_buf_1 _2305_ (.A(_1455_),
    .X(_1456_));
 sg13g2_nor2_1 _2306_ (.A(_1454_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_inv_1 _2307_ (.Y(_1458_),
    .A(_0033_));
 sg13g2_nor3_1 _2308_ (.A(_1405_),
    .B(_1451_),
    .C(_1458_),
    .Y(_1459_));
 sg13g2_buf_1 _2309_ (.A(_1459_),
    .X(_1460_));
 sg13g2_o21ai_1 _2310_ (.B1(net87),
    .Y(_1461_),
    .A1(_1457_),
    .A2(_1460_));
 sg13g2_a21oi_1 _2311_ (.A1(net63),
    .A2(_0721_),
    .Y(_1462_),
    .B1(net95));
 sg13g2_a22oi_1 _2312_ (.Y(_1463_),
    .B1(_1462_),
    .B2(_1404_),
    .A2(_1461_),
    .A1(_1408_));
 sg13g2_a22oi_1 _2313_ (.Y(_1464_),
    .B1(_1463_),
    .B2(net6),
    .A2(_1453_),
    .A1(_1419_));
 sg13g2_o21ai_1 _2314_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1441_),
    .A2(_1447_));
 sg13g2_nor2_1 _2315_ (.A(_0820_),
    .B(_0806_),
    .Y(_1466_));
 sg13g2_inv_1 _2316_ (.Y(_1467_),
    .A(_1466_));
 sg13g2_nand2b_1 _2317_ (.Y(_1468_),
    .B(_1466_),
    .A_N(_0808_));
 sg13g2_inv_1 _2318_ (.Y(_1469_),
    .A(net134));
 sg13g2_and3_1 _2319_ (.X(_1470_),
    .A(_0736_),
    .B(_1469_),
    .C(net91));
 sg13g2_nor3_1 _2320_ (.A(net131),
    .B(_1468_),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_nand4_1 _2321_ (.B(net120),
    .C(_0844_),
    .A(net121),
    .Y(_0090_),
    .D(_0846_));
 sg13g2_and2_1 _2322_ (.A(net114),
    .B(_0840_),
    .X(_0091_));
 sg13g2_o21ai_1 _2323_ (.B1(_0091_),
    .Y(_0092_),
    .A1(_1094_),
    .A2(_0090_));
 sg13g2_nor4_1 _2324_ (.A(_0837_),
    .B(_0695_),
    .C(_0834_),
    .D(_0815_),
    .Y(_0093_));
 sg13g2_nor2_1 _2325_ (.A(net108),
    .B(_0840_),
    .Y(_0094_));
 sg13g2_a221oi_1 _2326_ (.B2(_0832_),
    .C1(_1111_),
    .B1(_0094_),
    .A1(_0092_),
    .Y(_0095_),
    .A2(_0093_));
 sg13g2_nand2_2 _2327_ (.Y(_0096_),
    .A(\u8.hs[4] ),
    .B(_0698_));
 sg13g2_nor2_1 _2328_ (.A(_0710_),
    .B(_0096_),
    .Y(_0097_));
 sg13g2_nor2_1 _2329_ (.A(_1112_),
    .B(_0891_),
    .Y(_0098_));
 sg13g2_o21ai_1 _2330_ (.B1(_0098_),
    .Y(_0099_),
    .A1(_0811_),
    .A2(_0097_));
 sg13g2_a21o_1 _2331_ (.A2(_0095_),
    .A1(_0893_),
    .B1(_0099_),
    .X(_0100_));
 sg13g2_a21oi_1 _2332_ (.A1(_1471_),
    .A2(_0100_),
    .Y(_0101_),
    .B1(_0682_));
 sg13g2_and2_1 _2333_ (.A(_0687_),
    .B(_0713_),
    .X(_0102_));
 sg13g2_o21ai_1 _2334_ (.B1(_0102_),
    .Y(_0103_),
    .A1(_1467_),
    .A2(_0101_));
 sg13g2_nand2_1 _2335_ (.Y(_0104_),
    .A(_0659_),
    .B(_0718_));
 sg13g2_nor2_1 _2336_ (.A(_0028_),
    .B(_0104_),
    .Y(_0105_));
 sg13g2_inv_1 _2337_ (.Y(_0106_),
    .A(_1429_));
 sg13g2_nor2_1 _2338_ (.A(net12),
    .B(_0106_),
    .Y(_0107_));
 sg13g2_nand4_1 _2339_ (.B(_0103_),
    .C(_0105_),
    .A(_0916_),
    .Y(_0108_),
    .D(_0107_));
 sg13g2_nand2_2 _2340_ (.Y(_0109_),
    .A(_0723_),
    .B(_0729_));
 sg13g2_a21oi_1 _2341_ (.A1(_0709_),
    .A2(_0695_),
    .Y(_0110_),
    .B1(_0096_));
 sg13g2_nor2_2 _2342_ (.A(_0109_),
    .B(_0110_),
    .Y(_0111_));
 sg13g2_a21oi_1 _2343_ (.A1(net113),
    .A2(net108),
    .Y(_0112_),
    .B1(net125));
 sg13g2_nor2_2 _2344_ (.A(_0096_),
    .B(_0112_),
    .Y(_0113_));
 sg13g2_a21oi_1 _2345_ (.A1(_0111_),
    .A2(_0113_),
    .Y(_0114_),
    .B1(_1058_));
 sg13g2_nor3_1 _2346_ (.A(_0655_),
    .B(_1220_),
    .C(_0114_),
    .Y(_0115_));
 sg13g2_a21oi_1 _2347_ (.A1(_0794_),
    .A2(_1458_),
    .Y(_0116_),
    .B1(_1409_));
 sg13g2_o21ai_1 _2348_ (.B1(_0116_),
    .Y(_0117_),
    .A1(_1400_),
    .A2(_0115_));
 sg13g2_a21oi_1 _2349_ (.A1(_1403_),
    .A2(_0108_),
    .Y(_0118_),
    .B1(_0117_));
 sg13g2_buf_2 _2350_ (.A(_0118_),
    .X(_0119_));
 sg13g2_nor3_1 _2351_ (.A(net88),
    .B(_1458_),
    .C(_1450_),
    .Y(_0120_));
 sg13g2_a21oi_1 _2352_ (.A1(_1405_),
    .A2(_1406_),
    .Y(_0121_),
    .B1(_1451_));
 sg13g2_nand2_1 _2353_ (.Y(_0122_),
    .A(_0120_),
    .B(_0121_));
 sg13g2_and2_1 _2354_ (.A(_0119_),
    .B(_0122_),
    .X(_0123_));
 sg13g2_buf_2 _2355_ (.A(_0123_),
    .X(_0124_));
 sg13g2_mux2_1 _2356_ (.A0(_0838_),
    .A1(_1465_),
    .S(_0124_),
    .X(_0125_));
 sg13g2_and2_1 _2357_ (.A(net141),
    .B(_0125_),
    .X(_0048_));
 sg13g2_inv_1 _2358_ (.Y(_0126_),
    .A(net141));
 sg13g2_buf_1 _2359_ (.A(_0126_),
    .X(_0127_));
 sg13g2_buf_1 _2360_ (.A(_1404_),
    .X(_0128_));
 sg13g2_buf_1 _2361_ (.A(net78),
    .X(_0129_));
 sg13g2_nand2b_1 _2362_ (.Y(_0130_),
    .B(_1436_),
    .A_N(net111));
 sg13g2_o21ai_1 _2363_ (.B1(_0130_),
    .Y(_0131_),
    .A1(_0008_),
    .A2(_1436_));
 sg13g2_a22oi_1 _2364_ (.Y(_0132_),
    .B1(_0131_),
    .B2(net49),
    .A2(_1442_),
    .A1(net120));
 sg13g2_o21ai_1 _2365_ (.B1(net51),
    .Y(_0133_),
    .A1(_1442_),
    .A2(_1423_));
 sg13g2_o21ai_1 _2366_ (.B1(_0133_),
    .Y(_0134_),
    .A1(net45),
    .A2(_0132_));
 sg13g2_buf_1 _2367_ (.A(net83),
    .X(_0135_));
 sg13g2_nand2_1 _2368_ (.Y(_0136_),
    .A(net98),
    .B(net83));
 sg13g2_o21ai_1 _2369_ (.B1(_0136_),
    .Y(_0137_),
    .A1(_0106_),
    .A2(net68));
 sg13g2_mux2_1 _2370_ (.A0(_0134_),
    .A1(_0137_),
    .S(net95),
    .X(_0138_));
 sg13g2_buf_1 _2371_ (.A(_1456_),
    .X(_0139_));
 sg13g2_nor2_1 _2372_ (.A(_1405_),
    .B(_1459_),
    .Y(_0140_));
 sg13g2_nor3_2 _2373_ (.A(_1016_),
    .B(_1456_),
    .C(_0140_),
    .Y(_0141_));
 sg13g2_a22oi_1 _2374_ (.Y(_0142_),
    .B1(_0141_),
    .B2(net120),
    .A2(_1423_),
    .A1(net77));
 sg13g2_inv_1 _2375_ (.Y(_0143_),
    .A(_0142_));
 sg13g2_nand2_2 _2376_ (.Y(_0144_),
    .A(_0119_),
    .B(_0122_));
 sg13g2_a221oi_1 _2377_ (.B2(_1408_),
    .C1(_0144_),
    .B1(_0143_),
    .A1(net69),
    .Y(_0145_),
    .A2(_0138_));
 sg13g2_buf_8 _2378_ (.A(_0124_),
    .X(_0146_));
 sg13g2_nor2_1 _2379_ (.A(net130),
    .B(net37),
    .Y(_0147_));
 sg13g2_nor3_1 _2380_ (.A(net94),
    .B(_0145_),
    .C(_0147_),
    .Y(_0049_));
 sg13g2_nor2_1 _2381_ (.A(net108),
    .B(net37),
    .Y(_0148_));
 sg13g2_buf_1 _2382_ (.A(_0144_),
    .X(_0149_));
 sg13g2_nor2_1 _2383_ (.A(_1426_),
    .B(_1427_),
    .Y(_0150_));
 sg13g2_a22oi_1 _2384_ (.Y(_0151_),
    .B1(_0141_),
    .B2(net121),
    .A2(_0150_),
    .A1(net77));
 sg13g2_nor2_1 _2385_ (.A(net79),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_nand2_1 _2386_ (.Y(_0153_),
    .A(net97),
    .B(net46));
 sg13g2_o21ai_1 _2387_ (.B1(_0153_),
    .Y(_0154_),
    .A1(_0026_),
    .A2(net46));
 sg13g2_o21ai_1 _2388_ (.B1(net95),
    .Y(_0155_),
    .A1(_0106_),
    .A2(net83));
 sg13g2_a21oi_1 _2389_ (.A1(net68),
    .A2(_0154_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_a21o_1 _2390_ (.A2(_1442_),
    .A1(net51),
    .B1(net95),
    .X(_0157_));
 sg13g2_nand2_1 _2391_ (.Y(_0158_),
    .A(net109),
    .B(net60));
 sg13g2_o21ai_1 _2392_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_1212_),
    .A2(net59));
 sg13g2_a22oi_1 _2393_ (.Y(_0160_),
    .B1(net48),
    .B2(_0150_),
    .A2(net62),
    .A1(net121));
 sg13g2_o21ai_1 _2394_ (.B1(_0160_),
    .Y(_0161_),
    .A1(net50),
    .A2(_0159_));
 sg13g2_o21ai_1 _2395_ (.B1(net78),
    .Y(_0162_),
    .A1(_0157_),
    .A2(_0161_));
 sg13g2_nor2_1 _2396_ (.A(_0156_),
    .B(_0162_),
    .Y(_0163_));
 sg13g2_nor3_1 _2397_ (.A(net39),
    .B(_0152_),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_nor3_1 _2398_ (.A(net94),
    .B(_0148_),
    .C(_0164_),
    .Y(_0050_));
 sg13g2_a21oi_1 _2399_ (.A1(net71),
    .A2(_0025_),
    .Y(_0165_),
    .B1(_1432_));
 sg13g2_nand2_1 _2400_ (.Y(_0166_),
    .A(_1053_),
    .B(net60));
 sg13g2_o21ai_1 _2401_ (.B1(_0166_),
    .Y(_0167_),
    .A1(_0009_),
    .A2(net60));
 sg13g2_a22oi_1 _2402_ (.Y(_0168_),
    .B1(net49),
    .B2(_0167_),
    .A2(net62),
    .A1(net98));
 sg13g2_nand2b_1 _2403_ (.Y(_0169_),
    .B(_0168_),
    .A_N(net45));
 sg13g2_o21ai_1 _2404_ (.B1(_0169_),
    .Y(_0170_),
    .A1(net54),
    .A2(_0165_));
 sg13g2_nor2_1 _2405_ (.A(_0709_),
    .B(_0846_),
    .Y(_0171_));
 sg13g2_or2_1 _2406_ (.X(_0172_),
    .B(_0699_),
    .A(_0695_));
 sg13g2_nand2b_1 _2407_ (.Y(_0173_),
    .B(_0091_),
    .A_N(_0834_));
 sg13g2_nor3_1 _2408_ (.A(_0172_),
    .B(_0845_),
    .C(_0173_),
    .Y(_0174_));
 sg13g2_nand3_1 _2409_ (.B(_0171_),
    .C(_0174_),
    .A(_0824_),
    .Y(_0175_));
 sg13g2_nand3_1 _2410_ (.B(_0987_),
    .C(_0175_),
    .A(net114),
    .Y(_0176_));
 sg13g2_o21ai_1 _2411_ (.B1(_0176_),
    .Y(_0177_),
    .A1(_0027_),
    .A2(net46));
 sg13g2_a21oi_1 _2412_ (.A1(net68),
    .A2(_0177_),
    .Y(_0178_),
    .B1(_0155_));
 sg13g2_a221oi_1 _2413_ (.B2(_0170_),
    .C1(_0178_),
    .B1(net44),
    .A1(net106),
    .Y(_0179_),
    .A2(_0794_));
 sg13g2_a22oi_1 _2414_ (.Y(_0180_),
    .B1(_0141_),
    .B2(net98),
    .A2(_0165_),
    .A1(net77));
 sg13g2_nor2_1 _2415_ (.A(net79),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_o21ai_1 _2416_ (.B1(net37),
    .Y(_0182_),
    .A1(_0179_),
    .A2(_0181_));
 sg13g2_nand2_1 _2417_ (.Y(_0183_),
    .A(net113),
    .B(_0149_));
 sg13g2_buf_1 _2418_ (.A(_0126_),
    .X(_0184_));
 sg13g2_a21oi_1 _2419_ (.A1(_0182_),
    .A2(_0183_),
    .Y(_0051_),
    .B1(net93));
 sg13g2_nor2_1 _2420_ (.A(_0708_),
    .B(net37),
    .Y(_0185_));
 sg13g2_or2_1 _2421_ (.X(_0186_),
    .B(_1425_),
    .A(_1424_));
 sg13g2_a22oi_1 _2422_ (.Y(_0187_),
    .B1(_0141_),
    .B2(net97),
    .A2(_0186_),
    .A1(net77));
 sg13g2_nor2_1 _2423_ (.A(net79),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_buf_1 _2424_ (.A(net75),
    .X(_0189_));
 sg13g2_nand3_1 _2425_ (.B(net46),
    .C(_0175_),
    .A(net100),
    .Y(_0190_));
 sg13g2_o21ai_1 _2426_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0837_),
    .A2(net46));
 sg13g2_a21oi_2 _2427_ (.B1(_1402_),
    .Y(_0192_),
    .A2(net75),
    .A1(_0106_));
 sg13g2_o21ai_1 _2428_ (.B1(_0192_),
    .Y(_0193_),
    .A1(net58),
    .A2(_0191_));
 sg13g2_nor2_1 _2429_ (.A(_0680_),
    .B(net59),
    .Y(_0194_));
 sg13g2_a21oi_1 _2430_ (.A1(_1119_),
    .A2(net59),
    .Y(_0195_),
    .B1(_0194_));
 sg13g2_a22oi_1 _2431_ (.Y(_0196_),
    .B1(net48),
    .B2(_0186_),
    .A2(net62),
    .A1(net97));
 sg13g2_o21ai_1 _2432_ (.B1(_0196_),
    .Y(_0197_),
    .A1(net50),
    .A2(_0195_));
 sg13g2_nand2_1 _2433_ (.Y(_0198_),
    .A(_1446_),
    .B(_0197_));
 sg13g2_buf_1 _2434_ (.A(_1448_),
    .X(_0199_));
 sg13g2_a21oi_1 _2435_ (.A1(_0193_),
    .A2(_0198_),
    .Y(_0200_),
    .B1(net92));
 sg13g2_nor3_1 _2436_ (.A(net39),
    .B(_0188_),
    .C(_0200_),
    .Y(_0201_));
 sg13g2_nor3_1 _2437_ (.A(net94),
    .B(_0185_),
    .C(_0201_),
    .Y(_0052_));
 sg13g2_nand2_1 _2438_ (.Y(_0202_),
    .A(net129),
    .B(net39));
 sg13g2_nand3_1 _2439_ (.B(_0987_),
    .C(_0175_),
    .A(net127),
    .Y(_0203_));
 sg13g2_o21ai_1 _2440_ (.B1(_0203_),
    .Y(_0204_),
    .A1(net111),
    .A2(_0988_));
 sg13g2_o21ai_1 _2441_ (.B1(_0192_),
    .Y(_0205_),
    .A1(net58),
    .A2(_0204_));
 sg13g2_nor3_2 _2442_ (.A(net61),
    .B(_0777_),
    .C(net95),
    .Y(_0206_));
 sg13g2_o21ai_1 _2443_ (.B1(_0206_),
    .Y(_0207_),
    .A1(net114),
    .A2(net45));
 sg13g2_a21oi_1 _2444_ (.A1(_0205_),
    .A2(_0207_),
    .Y(_0208_),
    .B1(net92));
 sg13g2_nor2_2 _2445_ (.A(_0742_),
    .B(_0795_),
    .Y(_0209_));
 sg13g2_nand2_1 _2446_ (.Y(_0210_),
    .A(_0989_),
    .B(net53));
 sg13g2_o21ai_1 _2447_ (.B1(_0210_),
    .Y(_0211_),
    .A1(_0010_),
    .A2(net53));
 sg13g2_a22oi_1 _2448_ (.Y(_0212_),
    .B1(_0211_),
    .B2(net49),
    .A2(_1421_),
    .A1(net48));
 sg13g2_a22oi_1 _2449_ (.Y(_0213_),
    .B1(_0141_),
    .B2(_0961_),
    .A2(_1421_),
    .A1(net77));
 sg13g2_nand2b_1 _2450_ (.Y(_0214_),
    .B(_1408_),
    .A_N(_0213_));
 sg13g2_o21ai_1 _2451_ (.B1(_0214_),
    .Y(_0215_),
    .A1(_0209_),
    .A2(_0212_));
 sg13g2_o21ai_1 _2452_ (.B1(_0124_),
    .Y(_0216_),
    .A1(_0208_),
    .A2(_0215_));
 sg13g2_a21oi_1 _2453_ (.A1(_0202_),
    .A2(_0216_),
    .Y(_0053_),
    .B1(net93));
 sg13g2_nand2_1 _2454_ (.Y(_0217_),
    .A(_1430_),
    .B(_1431_));
 sg13g2_nand2_1 _2455_ (.Y(_0218_),
    .A(_1146_),
    .B(net60));
 sg13g2_o21ai_1 _2456_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0011_),
    .A2(net60));
 sg13g2_a22oi_1 _2457_ (.Y(_0220_),
    .B1(net49),
    .B2(_0219_),
    .A2(net62),
    .A1(net100));
 sg13g2_nand2b_1 _2458_ (.Y(_0221_),
    .B(_0220_),
    .A_N(net45));
 sg13g2_o21ai_1 _2459_ (.B1(_0221_),
    .Y(_0222_),
    .A1(net54),
    .A2(_0217_));
 sg13g2_nand3_1 _2460_ (.B(_0987_),
    .C(_0175_),
    .A(_0703_),
    .Y(_0223_));
 sg13g2_o21ai_1 _2461_ (.B1(_0223_),
    .Y(_0224_),
    .A1(net109),
    .A2(_0988_));
 sg13g2_a21oi_1 _2462_ (.A1(net68),
    .A2(_0224_),
    .Y(_0225_),
    .B1(_0155_));
 sg13g2_a221oi_1 _2463_ (.B2(_0222_),
    .C1(_0225_),
    .B1(net44),
    .A1(_0752_),
    .Y(_0226_),
    .A2(_0794_));
 sg13g2_a22oi_1 _2464_ (.Y(_0227_),
    .B1(_0141_),
    .B2(net100),
    .A2(_0217_),
    .A1(net77));
 sg13g2_nor2_1 _2465_ (.A(net79),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_o21ai_1 _2466_ (.B1(net37),
    .Y(_0229_),
    .A1(_0226_),
    .A2(_0228_));
 sg13g2_nand2_1 _2467_ (.Y(_0230_),
    .A(net99),
    .B(net39));
 sg13g2_a21oi_1 _2468_ (.A1(_0229_),
    .A2(_0230_),
    .Y(_0054_),
    .B1(net93));
 sg13g2_buf_1 _2469_ (.A(_1457_),
    .X(_0231_));
 sg13g2_a221oi_1 _2470_ (.B2(_0231_),
    .C1(_0117_),
    .B1(_0120_),
    .A1(_1403_),
    .Y(_0232_),
    .A2(_0108_));
 sg13g2_buf_1 _2471_ (.A(_0232_),
    .X(_0233_));
 sg13g2_buf_1 _2472_ (.A(_0233_),
    .X(_0234_));
 sg13g2_nand2b_1 _2473_ (.Y(_0235_),
    .B(net101),
    .A_N(net41));
 sg13g2_inv_1 _2474_ (.Y(_0236_),
    .A(_1435_));
 sg13g2_nor2_2 _2475_ (.A(_0749_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_nand2b_1 _2476_ (.Y(_0238_),
    .B(_0237_),
    .A_N(net129));
 sg13g2_o21ai_1 _2477_ (.B1(_1442_),
    .Y(_0239_),
    .A1(net127),
    .A2(net45));
 sg13g2_a21oi_1 _2478_ (.A1(_0238_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(net95));
 sg13g2_and3_1 _2479_ (.X(_0241_),
    .A(_0824_),
    .B(_0171_),
    .C(_0174_));
 sg13g2_a21oi_1 _2480_ (.A1(net57),
    .A2(_0986_),
    .Y(_0242_),
    .B1(_0241_));
 sg13g2_nor2_1 _2481_ (.A(net127),
    .B(_0840_),
    .Y(_0243_));
 sg13g2_nand3_1 _2482_ (.B(_0847_),
    .C(_0243_),
    .A(_0022_),
    .Y(_0244_));
 sg13g2_nand3b_1 _2483_ (.B(_0244_),
    .C(net134),
    .Y(_0245_),
    .A_N(net130));
 sg13g2_nand2b_1 _2484_ (.Y(_0246_),
    .B(net135),
    .A_N(_0028_));
 sg13g2_or4_1 _2485_ (.A(_0820_),
    .B(_0808_),
    .C(_0858_),
    .D(_0246_),
    .X(_0247_));
 sg13g2_nand2_1 _2486_ (.Y(_0248_),
    .A(net108),
    .B(_0816_));
 sg13g2_nor4_1 _2487_ (.A(_0811_),
    .B(_0245_),
    .C(_0247_),
    .D(_0248_),
    .Y(_0249_));
 sg13g2_nor3_2 _2488_ (.A(_0857_),
    .B(_1149_),
    .C(_0249_),
    .Y(_0250_));
 sg13g2_a22oi_1 _2489_ (.Y(_0251_),
    .B1(_0250_),
    .B2(_1053_),
    .A2(net47),
    .A1(net130));
 sg13g2_o21ai_1 _2490_ (.B1(net95),
    .Y(_0252_),
    .A1(_1429_),
    .A2(_0882_));
 sg13g2_buf_1 _2491_ (.A(_0252_),
    .X(_0253_));
 sg13g2_a21oi_1 _2492_ (.A1(net68),
    .A2(_0251_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_nor3_1 _2493_ (.A(net92),
    .B(_0240_),
    .C(_0254_),
    .Y(_0255_));
 sg13g2_buf_1 _2494_ (.A(_1035_),
    .X(_0256_));
 sg13g2_nand3_1 _2495_ (.B(\u8.rcip[1] ),
    .C(_0033_),
    .A(_1454_),
    .Y(_0257_));
 sg13g2_buf_2 _2496_ (.A(_0257_),
    .X(_0258_));
 sg13g2_nand2_1 _2497_ (.Y(_0259_),
    .A(_0704_),
    .B(net67));
 sg13g2_o21ai_1 _2498_ (.B1(_0259_),
    .Y(_0260_),
    .A1(_1017_),
    .A2(_0258_));
 sg13g2_nor2_1 _2499_ (.A(net71),
    .B(_1418_),
    .Y(_0261_));
 sg13g2_a22oi_1 _2500_ (.Y(_0262_),
    .B1(_0261_),
    .B2(net86),
    .A2(_0260_),
    .A1(net66));
 sg13g2_o21ai_1 _2501_ (.B1(net92),
    .Y(_0263_),
    .A1(net77),
    .A2(_0262_));
 sg13g2_nand3b_1 _2502_ (.B(net41),
    .C(_0263_),
    .Y(_0264_),
    .A_N(_0255_));
 sg13g2_a21oi_1 _2503_ (.A1(_0235_),
    .A2(_0264_),
    .Y(_0055_),
    .B1(net93));
 sg13g2_nor2_1 _2504_ (.A(net126),
    .B(_0234_),
    .Y(_0265_));
 sg13g2_xor2_1 _2505_ (.B(net99),
    .A(_0697_),
    .X(_0266_));
 sg13g2_a22oi_1 _2506_ (.Y(_0267_),
    .B1(_0237_),
    .B2(_0266_),
    .A2(net62),
    .A1(net128));
 sg13g2_a22oi_1 _2507_ (.Y(_0268_),
    .B1(_0250_),
    .B2(_1119_),
    .A2(net47),
    .A1(net108));
 sg13g2_a21o_1 _2508_ (.A2(_0268_),
    .A1(_0882_),
    .B1(_0253_),
    .X(_0269_));
 sg13g2_o21ai_1 _2509_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_0157_),
    .A2(_0267_));
 sg13g2_nand2_2 _2510_ (.Y(_0271_),
    .A(_1448_),
    .B(_1452_));
 sg13g2_nand2_1 _2511_ (.Y(_0272_),
    .A(net128),
    .B(net67));
 sg13g2_o21ai_1 _2512_ (.B1(_0272_),
    .Y(_0273_),
    .A1(_1096_),
    .A2(_0258_));
 sg13g2_nor2b_1 _2513_ (.A(_1018_),
    .B_N(net7),
    .Y(_0274_));
 sg13g2_a22oi_1 _2514_ (.Y(_0275_),
    .B1(_0274_),
    .B2(net86),
    .A2(_0273_),
    .A1(net70));
 sg13g2_nor2_1 _2515_ (.A(_0271_),
    .B(_0275_),
    .Y(_0276_));
 sg13g2_a21oi_1 _2516_ (.A1(net78),
    .A2(_0270_),
    .Y(_0277_),
    .B1(_0276_));
 sg13g2_and2_1 _2517_ (.A(_0233_),
    .B(_0277_),
    .X(_0278_));
 sg13g2_nor3_1 _2518_ (.A(net94),
    .B(_0265_),
    .C(_0278_),
    .Y(_0056_));
 sg13g2_and2_1 _2519_ (.A(net129),
    .B(net99),
    .X(_0279_));
 sg13g2_xnor2_1 _2520_ (.Y(_0280_),
    .A(net101),
    .B(_0279_));
 sg13g2_nor2_1 _2521_ (.A(_0209_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_a221oi_1 _2522_ (.B2(_0989_),
    .C1(net75),
    .B1(_0250_),
    .A1(net113),
    .Y(_0282_),
    .A2(net47));
 sg13g2_o21ai_1 _2523_ (.B1(_0206_),
    .Y(_0283_),
    .A1(_0693_),
    .A2(net45));
 sg13g2_o21ai_1 _2524_ (.B1(_0283_),
    .Y(_0284_),
    .A1(_0253_),
    .A2(_0282_));
 sg13g2_inv_1 _2525_ (.Y(_0285_),
    .A(net8));
 sg13g2_nor2_1 _2526_ (.A(_0285_),
    .B(_1035_),
    .Y(_0286_));
 sg13g2_nand2_1 _2527_ (.Y(_0287_),
    .A(_0693_),
    .B(_0231_));
 sg13g2_o21ai_1 _2528_ (.B1(_0287_),
    .Y(_0288_),
    .A1(_1036_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2529_ (.Y(_0289_),
    .B1(_0288_),
    .B2(net66),
    .A2(_0286_),
    .A1(net86));
 sg13g2_nor2_1 _2530_ (.A(_0271_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_a221oi_1 _2531_ (.B2(net78),
    .C1(_0290_),
    .B1(_0284_),
    .A1(_0237_),
    .Y(_0291_),
    .A2(_0281_));
 sg13g2_mux2_1 _2532_ (.A0(_0731_),
    .A1(_0291_),
    .S(_0233_),
    .X(_0292_));
 sg13g2_nor2_1 _2533_ (.A(net93),
    .B(_0292_),
    .Y(_0057_));
 sg13g2_a22oi_1 _2534_ (.Y(_0293_),
    .B1(_0250_),
    .B2(_1146_),
    .A2(net47),
    .A1(net125));
 sg13g2_nand2_1 _2535_ (.Y(_0294_),
    .A(net68),
    .B(_0293_));
 sg13g2_nand2_1 _2536_ (.Y(_0295_),
    .A(net63),
    .B(_0721_));
 sg13g2_buf_1 _2537_ (.A(_0295_),
    .X(_0296_));
 sg13g2_nor2_1 _2538_ (.A(net108),
    .B(net51),
    .Y(_0297_));
 sg13g2_xor2_1 _2539_ (.B(_0699_),
    .A(_1099_),
    .X(_0298_));
 sg13g2_nand2_1 _2540_ (.Y(_0299_),
    .A(_0237_),
    .B(_0298_));
 sg13g2_o21ai_1 _2541_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net43),
    .A2(_0297_));
 sg13g2_a22oi_1 _2542_ (.Y(_0301_),
    .B1(_0300_),
    .B2(_1402_),
    .A2(_0294_),
    .A1(_0192_));
 sg13g2_nor2_1 _2543_ (.A(net92),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_inv_1 _2544_ (.Y(_0303_),
    .A(net9));
 sg13g2_nor2_1 _2545_ (.A(net71),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_nand2_1 _2546_ (.Y(_0305_),
    .A(_1326_),
    .B(net67));
 sg13g2_o21ai_1 _2547_ (.B1(_0305_),
    .Y(_0306_),
    .A1(_1111_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2548_ (.Y(_0307_),
    .B1(_0306_),
    .B2(net66),
    .A2(_0304_),
    .A1(net86));
 sg13g2_nor2_1 _2549_ (.A(_0271_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_o21ai_1 _2550_ (.B1(net41),
    .Y(_0309_),
    .A1(_0302_),
    .A2(_0308_));
 sg13g2_nand2b_1 _2551_ (.Y(_0310_),
    .B(_0677_),
    .A_N(net41));
 sg13g2_buf_1 _2552_ (.A(_0127_),
    .X(_0311_));
 sg13g2_a21oi_1 _2553_ (.A1(_0309_),
    .A2(_0310_),
    .Y(_0058_),
    .B1(net85));
 sg13g2_nor2_1 _2554_ (.A(net119),
    .B(net37),
    .Y(_0312_));
 sg13g2_a21oi_1 _2555_ (.A1(_1132_),
    .A2(net7),
    .Y(_0313_),
    .B1(_1128_));
 sg13g2_inv_1 _2556_ (.Y(_0314_),
    .A(_0313_));
 sg13g2_nor2_1 _2557_ (.A(_1096_),
    .B(net59),
    .Y(_0315_));
 sg13g2_a21oi_1 _2558_ (.A1(net53),
    .A2(_0314_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_nand2_1 _2559_ (.Y(_0317_),
    .A(net48),
    .B(_0314_));
 sg13g2_o21ai_1 _2560_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net50),
    .A2(_0316_));
 sg13g2_nand3_1 _2561_ (.B(net44),
    .C(_0318_),
    .A(net69),
    .Y(_0319_));
 sg13g2_a22oi_1 _2562_ (.Y(_0320_),
    .B1(_0314_),
    .B2(_1453_),
    .A2(_1463_),
    .A1(net7));
 sg13g2_and3_1 _2563_ (.X(_0321_),
    .A(_0124_),
    .B(_0319_),
    .C(_0320_));
 sg13g2_nor3_1 _2564_ (.A(net94),
    .B(_0312_),
    .C(_0321_),
    .Y(_0059_));
 sg13g2_a22oi_1 _2565_ (.Y(_0322_),
    .B1(_0250_),
    .B2(_1340_),
    .A2(net47),
    .A1(net129));
 sg13g2_nand2_1 _2566_ (.Y(_0323_),
    .A(net68),
    .B(_0322_));
 sg13g2_nor2_1 _2567_ (.A(_0980_),
    .B(_1008_),
    .Y(_0324_));
 sg13g2_nand4_1 _2568_ (.B(net101),
    .C(_0279_),
    .A(net126),
    .Y(_0325_),
    .D(_0237_));
 sg13g2_o21ai_1 _2569_ (.B1(_0325_),
    .Y(_0326_),
    .A1(net43),
    .A2(_0324_));
 sg13g2_a22oi_1 _2570_ (.Y(_0327_),
    .B1(_0326_),
    .B2(_1402_),
    .A2(_0323_),
    .A1(_0192_));
 sg13g2_nor2_1 _2571_ (.A(net92),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_nor2b_1 _2572_ (.A(net70),
    .B_N(net10),
    .Y(_0329_));
 sg13g2_nand2_1 _2573_ (.Y(_0330_),
    .A(_0980_),
    .B(net67));
 sg13g2_o21ai_1 _2574_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_0003_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2575_ (.Y(_0332_),
    .B1(_0331_),
    .B2(net66),
    .A2(_0329_),
    .A1(net86));
 sg13g2_nor2_1 _2576_ (.A(_0271_),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_o21ai_1 _2577_ (.B1(net41),
    .Y(_0334_),
    .A1(_0328_),
    .A2(_0333_));
 sg13g2_nand2b_1 _2578_ (.Y(_0335_),
    .B(_0675_),
    .A_N(net41));
 sg13g2_a21oi_1 _2579_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0060_),
    .B1(net85));
 sg13g2_nor2_1 _2580_ (.A(_0794_),
    .B(_0253_),
    .Y(_0336_));
 sg13g2_nor3_1 _2581_ (.A(net108),
    .B(net130),
    .C(_0826_),
    .Y(_0337_));
 sg13g2_a21oi_1 _2582_ (.A1(_1197_),
    .A2(_0337_),
    .Y(_0338_),
    .B1(net99));
 sg13g2_nand2_1 _2583_ (.Y(_0339_),
    .A(_0812_),
    .B(_0338_));
 sg13g2_nand2_2 _2584_ (.Y(_0340_),
    .A(_0250_),
    .B(_0339_));
 sg13g2_a21oi_1 _2585_ (.A1(_1236_),
    .A2(_0242_),
    .Y(_0341_),
    .B1(_0911_));
 sg13g2_o21ai_1 _2586_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0005_),
    .A2(_0340_));
 sg13g2_nor2_1 _2587_ (.A(_0710_),
    .B(_0209_),
    .Y(_0343_));
 sg13g2_nand2_1 _2588_ (.Y(_0344_),
    .A(_0708_),
    .B(net67));
 sg13g2_o21ai_1 _2589_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0710_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2590_ (.Y(_0346_),
    .B1(_0345_),
    .B2(net70),
    .A2(_1425_),
    .A1(net86));
 sg13g2_nor2_1 _2591_ (.A(_0271_),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_a221oi_1 _2592_ (.B2(_1095_),
    .C1(_0347_),
    .B1(_0343_),
    .A1(_0336_),
    .Y(_0348_),
    .A2(_0342_));
 sg13g2_nand2_1 _2593_ (.Y(_0349_),
    .A(_0233_),
    .B(_0348_));
 sg13g2_o21ai_1 _2594_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0674_),
    .A2(net41));
 sg13g2_nor2_1 _2595_ (.A(net93),
    .B(_0350_),
    .Y(_0061_));
 sg13g2_inv_1 _2596_ (.Y(_0351_),
    .A(net12));
 sg13g2_nor2_1 _2597_ (.A(_1072_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nand2_1 _2598_ (.Y(_0353_),
    .A(_0697_),
    .B(net67));
 sg13g2_o21ai_1 _2599_ (.B1(_0353_),
    .Y(_0354_),
    .A1(_1197_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2600_ (.Y(_0355_),
    .B1(_0354_),
    .B2(_0256_),
    .A2(_0352_),
    .A1(net86));
 sg13g2_nor2_1 _2601_ (.A(_0271_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_a21oi_1 _2602_ (.A1(_1041_),
    .A2(net47),
    .Y(_0357_),
    .B1(_0911_));
 sg13g2_o21ai_1 _2603_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0006_),
    .A2(_0340_));
 sg13g2_nand2_1 _2604_ (.Y(_0359_),
    .A(_1197_),
    .B(net54));
 sg13g2_a22oi_1 _2605_ (.Y(_0360_),
    .B1(_0359_),
    .B2(_0206_),
    .A2(_0358_),
    .A1(_0192_));
 sg13g2_nor2_1 _2606_ (.A(net92),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_o21ai_1 _2607_ (.B1(_0234_),
    .Y(_0362_),
    .A1(_0356_),
    .A2(_0361_));
 sg13g2_nand2b_1 _2608_ (.Y(_0363_),
    .B(net139),
    .A_N(_0233_));
 sg13g2_a21oi_1 _2609_ (.A1(_0362_),
    .A2(_0363_),
    .Y(_0062_),
    .B1(net85));
 sg13g2_nand2_1 _2610_ (.Y(_0364_),
    .A(_1238_),
    .B(net62));
 sg13g2_nand2_1 _2611_ (.Y(_0365_),
    .A(_0706_),
    .B(net47));
 sg13g2_o21ai_1 _2612_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_1099_),
    .A2(_0340_));
 sg13g2_a21oi_1 _2613_ (.A1(net68),
    .A2(_0366_),
    .Y(_0367_),
    .B1(_0155_));
 sg13g2_a221oi_1 _2614_ (.B2(_0364_),
    .C1(_0367_),
    .B1(net44),
    .A1(_0752_),
    .Y(_0368_),
    .A2(_0794_));
 sg13g2_nor2_1 _2615_ (.A(net70),
    .B(_0106_),
    .Y(_0369_));
 sg13g2_nand2_1 _2616_ (.Y(_0370_),
    .A(_1236_),
    .B(net67));
 sg13g2_o21ai_1 _2617_ (.B1(_0370_),
    .Y(_0371_),
    .A1(_0005_),
    .A2(_0258_));
 sg13g2_a22oi_1 _2618_ (.Y(_0372_),
    .B1(_0371_),
    .B2(_0256_),
    .A2(_0369_),
    .A1(net86));
 sg13g2_nor2_1 _2619_ (.A(_0271_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_o21ai_1 _2620_ (.B1(net41),
    .Y(_0374_),
    .A1(_0368_),
    .A2(_0373_));
 sg13g2_nand2b_1 _2621_ (.Y(_0375_),
    .B(_0664_),
    .A_N(_0233_));
 sg13g2_a21oi_1 _2622_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0063_),
    .B1(net85));
 sg13g2_nor2_2 _2623_ (.A(_1454_),
    .B(_0271_),
    .Y(_0376_));
 sg13g2_a21o_1 _2624_ (.A2(net66),
    .A1(net101),
    .B1(_0261_),
    .X(_0377_));
 sg13g2_a21oi_1 _2625_ (.A1(_0678_),
    .A2(net47),
    .Y(_0378_),
    .B1(net75));
 sg13g2_o21ai_1 _2626_ (.B1(_0378_),
    .Y(_0379_),
    .A1(_0008_),
    .A2(_0340_));
 sg13g2_a21o_1 _2627_ (.A2(_0379_),
    .A1(_0192_),
    .B1(_0206_),
    .X(_0380_));
 sg13g2_a22oi_1 _2628_ (.Y(_0381_),
    .B1(_0380_),
    .B2(net69),
    .A2(_0377_),
    .A1(_0376_));
 sg13g2_mux2_1 _2629_ (.A0(_0995_),
    .A1(_0381_),
    .S(_0119_),
    .X(_0382_));
 sg13g2_nor2_1 _2630_ (.A(net93),
    .B(_0382_),
    .Y(_0064_));
 sg13g2_buf_1 _2631_ (.A(_0119_),
    .X(_0383_));
 sg13g2_nand2_1 _2632_ (.Y(_0384_),
    .A(net143),
    .B(_0192_));
 sg13g2_a21oi_2 _2633_ (.B1(_0241_),
    .Y(_0385_),
    .A2(_0916_),
    .A1(_0851_));
 sg13g2_or2_1 _2634_ (.X(_0386_),
    .B(_0385_),
    .A(_1152_));
 sg13g2_nand2b_1 _2635_ (.Y(_0387_),
    .B(_0340_),
    .A_N(_0386_));
 sg13g2_a221oi_1 _2636_ (.B2(_1212_),
    .C1(net58),
    .B1(_0387_),
    .A1(_0677_),
    .Y(_0388_),
    .A2(_1000_));
 sg13g2_a21oi_1 _2637_ (.A1(_0706_),
    .A2(net70),
    .Y(_0389_),
    .B1(_0274_));
 sg13g2_nand2b_1 _2638_ (.Y(_0390_),
    .B(_0376_),
    .A_N(_0389_));
 sg13g2_o21ai_1 _2639_ (.B1(_0390_),
    .Y(_0391_),
    .A1(_0384_),
    .A2(_0388_));
 sg13g2_nand2_1 _2640_ (.Y(_0392_),
    .A(net40),
    .B(_0391_));
 sg13g2_nand2b_1 _2641_ (.Y(_0393_),
    .B(net136),
    .A_N(_0119_));
 sg13g2_a21oi_1 _2642_ (.A1(_0392_),
    .A2(_0393_),
    .Y(_0065_),
    .B1(net85));
 sg13g2_nand3b_1 _2643_ (.B(_1112_),
    .C(_1113_),
    .Y(_0394_),
    .A_N(net99));
 sg13g2_nand3b_1 _2644_ (.B(_0394_),
    .C(_1469_),
    .Y(_0395_),
    .A_N(_0247_));
 sg13g2_nand4_1 _2645_ (.B(_0947_),
    .C(_0873_),
    .A(_0963_),
    .Y(_0396_),
    .D(_0395_));
 sg13g2_nand2_1 _2646_ (.Y(_0397_),
    .A(_0340_),
    .B(_0396_));
 sg13g2_a221oi_1 _2647_ (.B2(_1251_),
    .C1(net58),
    .B1(_0397_),
    .A1(_0675_),
    .Y(_0398_),
    .A2(_0386_));
 sg13g2_a21o_1 _2648_ (.A2(net70),
    .A1(_0678_),
    .B1(_0286_),
    .X(_0399_));
 sg13g2_a22oi_1 _2649_ (.Y(_0400_),
    .B1(_0376_),
    .B2(_0399_),
    .A2(_0206_),
    .A1(net78));
 sg13g2_o21ai_1 _2650_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0384_),
    .A2(_0398_));
 sg13g2_nand2_1 _2651_ (.Y(_0402_),
    .A(net40),
    .B(_0401_));
 sg13g2_nand2b_1 _2652_ (.Y(_0403_),
    .B(_0661_),
    .A_N(_0119_));
 sg13g2_a21oi_1 _2653_ (.A1(_0402_),
    .A2(_0403_),
    .Y(_0066_),
    .B1(net85));
 sg13g2_a221oi_1 _2654_ (.B2(_0715_),
    .C1(net58),
    .B1(_0397_),
    .A1(net135),
    .Y(_0404_),
    .A2(_0386_));
 sg13g2_a21o_1 _2655_ (.A2(_1082_),
    .A1(net133),
    .B1(_0304_),
    .X(_0405_));
 sg13g2_a22oi_1 _2656_ (.Y(_0406_),
    .B1(_0376_),
    .B2(_0405_),
    .A2(_0206_),
    .A1(net78));
 sg13g2_o21ai_1 _2657_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_0384_),
    .A2(_0404_));
 sg13g2_nand2_1 _2658_ (.Y(_0408_),
    .A(net40),
    .B(_0407_));
 sg13g2_nand2b_1 _2659_ (.Y(_0409_),
    .B(_0660_),
    .A_N(_0119_));
 sg13g2_a21oi_1 _2660_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0067_),
    .B1(net85));
 sg13g2_nand3_1 _2661_ (.B(_0340_),
    .C(_0396_),
    .A(_1241_),
    .Y(_0410_));
 sg13g2_a21o_1 _2662_ (.A2(_0727_),
    .A1(_0015_),
    .B1(net136),
    .X(_0411_));
 sg13g2_o21ai_1 _2663_ (.B1(_1152_),
    .Y(_0412_),
    .A1(_1467_),
    .A2(_0411_));
 sg13g2_nand2_1 _2664_ (.Y(_0413_),
    .A(_0851_),
    .B(_0916_));
 sg13g2_a21oi_1 _2665_ (.A1(_0010_),
    .A2(_0412_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_a221oi_1 _2666_ (.B2(_0414_),
    .C1(net58),
    .B1(_0410_),
    .A1(net139),
    .Y(_0415_),
    .A2(_0385_));
 sg13g2_nand2_1 _2667_ (.Y(_0416_),
    .A(_1442_),
    .B(_1402_));
 sg13g2_o21ai_1 _2668_ (.B1(_0416_),
    .Y(_0417_),
    .A1(_0253_),
    .A2(_0415_));
 sg13g2_a21oi_1 _2669_ (.A1(net134),
    .A2(net66),
    .Y(_0418_),
    .B1(_0329_));
 sg13g2_nor2_1 _2670_ (.A(net69),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_a22oi_1 _2671_ (.Y(_0420_),
    .B1(_0419_),
    .B2(net67),
    .A2(_0417_),
    .A1(net69));
 sg13g2_o21ai_1 _2672_ (.B1(net141),
    .Y(_0421_),
    .A1(_0668_),
    .A2(net40));
 sg13g2_a21oi_1 _2673_ (.A1(_0383_),
    .A2(_0420_),
    .Y(_0068_),
    .B1(_0421_));
 sg13g2_nand2_1 _2674_ (.Y(_0422_),
    .A(net83),
    .B(_0412_));
 sg13g2_o21ai_1 _2675_ (.B1(_1367_),
    .Y(_0423_),
    .A1(_0385_),
    .A2(_0410_));
 sg13g2_nand2b_1 _2676_ (.Y(_0424_),
    .B(_0423_),
    .A_N(_0422_));
 sg13g2_a21o_1 _2677_ (.A2(net66),
    .A1(_0674_),
    .B1(_1425_),
    .X(_0425_));
 sg13g2_a22oi_1 _2678_ (.Y(_0426_),
    .B1(_0425_),
    .B2(_0376_),
    .A2(_0424_),
    .A1(_0336_));
 sg13g2_o21ai_1 _2679_ (.B1(net141),
    .Y(_0427_),
    .A1(net138),
    .A2(net40));
 sg13g2_a21oi_1 _2680_ (.A1(net40),
    .A2(_0426_),
    .Y(_0069_),
    .B1(_0427_));
 sg13g2_nand2_1 _2681_ (.Y(_0428_),
    .A(_0842_),
    .B(net39));
 sg13g2_nand2_1 _2682_ (.Y(_0429_),
    .A(net43),
    .B(_1402_));
 sg13g2_a21oi_2 _2683_ (.B1(_1187_),
    .Y(_0430_),
    .A2(net88),
    .A1(_0285_));
 sg13g2_nor2_1 _2684_ (.A(_1036_),
    .B(net59),
    .Y(_0431_));
 sg13g2_a21oi_1 _2685_ (.A1(_1437_),
    .A2(_0430_),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_nand2_1 _2686_ (.Y(_0433_),
    .A(net48),
    .B(_0430_));
 sg13g2_o21ai_1 _2687_ (.B1(_0433_),
    .Y(_0434_),
    .A1(net50),
    .A2(_0432_));
 sg13g2_a22oi_1 _2688_ (.Y(_0435_),
    .B1(net44),
    .B2(_0434_),
    .A2(_0429_),
    .A1(net8));
 sg13g2_nand2_1 _2689_ (.Y(_0436_),
    .A(_1448_),
    .B(_1407_));
 sg13g2_and2_1 _2690_ (.A(_1461_),
    .B(_0436_),
    .X(_0437_));
 sg13g2_nand2_1 _2691_ (.Y(_0438_),
    .A(_0139_),
    .B(_0430_));
 sg13g2_nand2_1 _2692_ (.Y(_0439_),
    .A(_0437_),
    .B(_0438_));
 sg13g2_a221oi_1 _2693_ (.B2(net8),
    .C1(_0128_),
    .B1(_0439_),
    .A1(_1453_),
    .Y(_0440_),
    .A2(_0430_));
 sg13g2_a21oi_1 _2694_ (.A1(net69),
    .A2(_0435_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nand2_1 _2695_ (.Y(_0442_),
    .A(net37),
    .B(_0441_));
 sg13g2_a21oi_1 _2696_ (.A1(_0428_),
    .A2(_0442_),
    .Y(_0070_),
    .B1(_0311_));
 sg13g2_nand2b_1 _2697_ (.Y(_0443_),
    .B(_0656_),
    .A_N(_0119_));
 sg13g2_nand2_1 _2698_ (.Y(_0444_),
    .A(_0015_),
    .B(_0412_));
 sg13g2_a221oi_1 _2699_ (.B2(_0444_),
    .C1(net58),
    .B1(_0410_),
    .A1(_0671_),
    .Y(_0445_),
    .A2(_0385_));
 sg13g2_a21o_1 _2700_ (.A2(_1082_),
    .A1(_0665_),
    .B1(_0352_),
    .X(_0446_));
 sg13g2_a22oi_1 _2701_ (.Y(_0447_),
    .B1(_0376_),
    .B2(_0446_),
    .A2(_0206_),
    .A1(net78));
 sg13g2_o21ai_1 _2702_ (.B1(_0447_),
    .Y(_0448_),
    .A1(_0384_),
    .A2(_0445_));
 sg13g2_nand2_1 _2703_ (.Y(_0449_),
    .A(_0383_),
    .B(_0448_));
 sg13g2_a21oi_1 _2704_ (.A1(_0443_),
    .A2(_0449_),
    .Y(_0071_),
    .B1(net85));
 sg13g2_a221oi_1 _2705_ (.B2(_1127_),
    .C1(_0422_),
    .B1(_0397_),
    .A1(net136),
    .Y(_0450_),
    .A2(_0385_));
 sg13g2_o21ai_1 _2706_ (.B1(_0416_),
    .Y(_0451_),
    .A1(_0253_),
    .A2(_0450_));
 sg13g2_a21o_1 _2707_ (.A2(net66),
    .A1(_0664_),
    .B1(_0369_),
    .X(_0452_));
 sg13g2_a22oi_1 _2708_ (.Y(_0453_),
    .B1(_0452_),
    .B2(_0376_),
    .A2(_0451_),
    .A1(net69));
 sg13g2_o21ai_1 _2709_ (.B1(net141),
    .Y(_0454_),
    .A1(net140),
    .A2(net40));
 sg13g2_a21oi_1 _2710_ (.A1(net40),
    .A2(_0453_),
    .Y(_0072_),
    .B1(_0454_));
 sg13g2_nand2_1 _2711_ (.Y(_0455_),
    .A(_0841_),
    .B(_0149_));
 sg13g2_a21oi_2 _2712_ (.B1(_1216_),
    .Y(_0456_),
    .A2(_0303_),
    .A1(_1132_));
 sg13g2_nor2_1 _2713_ (.A(_1111_),
    .B(net59),
    .Y(_0457_));
 sg13g2_a21oi_1 _2714_ (.A1(_1437_),
    .A2(_0456_),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_nand2_1 _2715_ (.Y(_0459_),
    .A(_1417_),
    .B(_0456_));
 sg13g2_o21ai_1 _2716_ (.B1(_0459_),
    .Y(_0460_),
    .A1(net50),
    .A2(_0458_));
 sg13g2_a22oi_1 _2717_ (.Y(_0461_),
    .B1(net44),
    .B2(_0460_),
    .A2(_0429_),
    .A1(net9));
 sg13g2_nand2_1 _2718_ (.Y(_0462_),
    .A(_1456_),
    .B(_0456_));
 sg13g2_nand2_1 _2719_ (.Y(_0463_),
    .A(_0437_),
    .B(_0462_));
 sg13g2_a221oi_1 _2720_ (.B2(net9),
    .C1(_0128_),
    .B1(_0463_),
    .A1(_1453_),
    .Y(_0464_),
    .A2(_0456_));
 sg13g2_a21oi_1 _2721_ (.A1(net69),
    .A2(_0461_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nand2_1 _2722_ (.Y(_0466_),
    .A(_0146_),
    .B(_0465_));
 sg13g2_a21oi_1 _2723_ (.A1(_0455_),
    .A2(_0466_),
    .Y(_0073_),
    .B1(_0311_));
 sg13g2_nand2_1 _2724_ (.Y(_0467_),
    .A(net98),
    .B(net39));
 sg13g2_mux2_1 _2725_ (.A0(net10),
    .A1(_1269_),
    .S(_1015_),
    .X(_0468_));
 sg13g2_nor2_1 _2726_ (.A(_0003_),
    .B(net60),
    .Y(_0469_));
 sg13g2_a21oi_1 _2727_ (.A1(_1438_),
    .A2(_0468_),
    .Y(_0470_),
    .B1(_0469_));
 sg13g2_nand2_1 _2728_ (.Y(_0471_),
    .A(_1417_),
    .B(_0468_));
 sg13g2_o21ai_1 _2729_ (.B1(_0471_),
    .Y(_0472_),
    .A1(_1032_),
    .A2(_0470_));
 sg13g2_a22oi_1 _2730_ (.Y(_0473_),
    .B1(net44),
    .B2(_0472_),
    .A2(_0429_),
    .A1(net10));
 sg13g2_nand2_1 _2731_ (.Y(_0474_),
    .A(_1456_),
    .B(_0468_));
 sg13g2_nand2_1 _2732_ (.Y(_0475_),
    .A(_0437_),
    .B(_0474_));
 sg13g2_a221oi_1 _2733_ (.B2(net10),
    .C1(net78),
    .B1(_0475_),
    .A1(_1453_),
    .Y(_0476_),
    .A2(_0468_));
 sg13g2_a21oi_1 _2734_ (.A1(_0129_),
    .A2(_0473_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nand2_1 _2735_ (.Y(_0478_),
    .A(_0146_),
    .B(_0477_));
 sg13g2_a21oi_1 _2736_ (.A1(_0467_),
    .A2(_0478_),
    .Y(_0074_),
    .B1(net94));
 sg13g2_mux2_1 _2737_ (.A0(_0846_),
    .A1(net11),
    .S(_1034_),
    .X(_0479_));
 sg13g2_nand2_1 _2738_ (.Y(_0480_),
    .A(_1438_),
    .B(_0479_));
 sg13g2_o21ai_1 _2739_ (.B1(_0480_),
    .Y(_0481_),
    .A1(_0710_),
    .A2(net53));
 sg13g2_a22oi_1 _2740_ (.Y(_0482_),
    .B1(_0481_),
    .B2(net49),
    .A2(_0479_),
    .A1(net48));
 sg13g2_nor2_1 _2741_ (.A(_1457_),
    .B(_1460_),
    .Y(_0483_));
 sg13g2_nor2_1 _2742_ (.A(_1016_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_a21oi_1 _2743_ (.A1(_0484_),
    .A2(_0479_),
    .Y(_0485_),
    .B1(net79));
 sg13g2_nor2b_1 _2744_ (.A(_0485_),
    .B_N(net11),
    .Y(_0486_));
 sg13g2_nand2_1 _2745_ (.Y(_0487_),
    .A(_1404_),
    .B(_1462_));
 sg13g2_a22oi_1 _2746_ (.Y(_0488_),
    .B1(_0486_),
    .B2(_0487_),
    .A2(_0479_),
    .A1(_1453_));
 sg13g2_o21ai_1 _2747_ (.B1(_0488_),
    .Y(_0489_),
    .A1(_1447_),
    .A2(_0482_));
 sg13g2_mux2_1 _2748_ (.A0(net97),
    .A1(_0489_),
    .S(_0124_),
    .X(_0490_));
 sg13g2_and2_1 _2749_ (.A(_1248_),
    .B(_0490_),
    .X(_0075_));
 sg13g2_mux2_1 _2750_ (.A0(_0351_),
    .A1(_0027_),
    .S(_1015_),
    .X(_0491_));
 sg13g2_nand2_1 _2751_ (.Y(_0492_),
    .A(net12),
    .B(_0484_));
 sg13g2_o21ai_1 _2752_ (.B1(_0492_),
    .Y(_0493_),
    .A1(_1452_),
    .A2(_0491_));
 sg13g2_nand3_1 _2753_ (.B(net58),
    .C(_1444_),
    .A(net143),
    .Y(_0494_));
 sg13g2_a21oi_1 _2754_ (.A1(_0436_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(_0351_));
 sg13g2_a221oi_1 _2755_ (.B2(_0493_),
    .C1(_0495_),
    .B1(_1408_),
    .A1(_0838_),
    .Y(_0496_),
    .A2(_1403_));
 sg13g2_o21ai_1 _2756_ (.B1(net43),
    .Y(_0497_),
    .A1(net54),
    .A2(_0491_));
 sg13g2_o21ai_1 _2757_ (.B1(_0497_),
    .Y(_0498_),
    .A1(net12),
    .A2(net43));
 sg13g2_nor3_1 _2758_ (.A(_1009_),
    .B(_0236_),
    .C(_0491_),
    .Y(_0499_));
 sg13g2_nor3_1 _2759_ (.A(_1197_),
    .B(_1399_),
    .C(net53),
    .Y(_0500_));
 sg13g2_o21ai_1 _2760_ (.B1(net49),
    .Y(_0501_),
    .A1(_0499_),
    .A2(_0500_));
 sg13g2_a21oi_1 _2761_ (.A1(_0498_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(_0209_));
 sg13g2_nor2_1 _2762_ (.A(_0144_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_a221oi_1 _2763_ (.B2(_0503_),
    .C1(_0127_),
    .B1(_0496_),
    .A1(_1338_),
    .Y(_0076_),
    .A2(net39));
 sg13g2_a21oi_2 _2764_ (.B1(_1387_),
    .Y(_0504_),
    .A2(_1429_),
    .A1(net80));
 sg13g2_o21ai_1 _2765_ (.B1(_0437_),
    .Y(_0505_),
    .A1(_1452_),
    .A2(_0504_));
 sg13g2_nor3_1 _2766_ (.A(_1407_),
    .B(_1452_),
    .C(_0504_),
    .Y(_0506_));
 sg13g2_a21oi_1 _2767_ (.A1(_1429_),
    .A2(_0505_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_o21ai_1 _2768_ (.B1(_0336_),
    .Y(_0508_),
    .A1(net119),
    .A2(_0189_));
 sg13g2_o21ai_1 _2769_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0129_),
    .A2(_0507_));
 sg13g2_o21ai_1 _2770_ (.B1(net43),
    .Y(_0510_),
    .A1(net54),
    .A2(_0504_));
 sg13g2_o21ai_1 _2771_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_1429_),
    .A2(net43));
 sg13g2_nor3_1 _2772_ (.A(_1009_),
    .B(_0236_),
    .C(_0504_),
    .Y(_0512_));
 sg13g2_nor3_1 _2773_ (.A(_0005_),
    .B(_1399_),
    .C(net53),
    .Y(_0513_));
 sg13g2_o21ai_1 _2774_ (.B1(_1315_),
    .Y(_0514_),
    .A1(_0512_),
    .A2(_0513_));
 sg13g2_a21oi_1 _2775_ (.A1(_0511_),
    .A2(_0514_),
    .Y(_0515_),
    .B1(_0209_));
 sg13g2_nor3_1 _2776_ (.A(net39),
    .B(_0509_),
    .C(_0515_),
    .Y(_0516_));
 sg13g2_o21ai_1 _2777_ (.B1(net141),
    .Y(_0517_),
    .A1(net100),
    .A2(net37));
 sg13g2_nor2_1 _2778_ (.A(_0516_),
    .B(_0517_),
    .Y(_0077_));
 sg13g2_nor2_1 _2779_ (.A(_0704_),
    .B(_0124_),
    .Y(_0518_));
 sg13g2_nor2_1 _2780_ (.A(net81),
    .B(net6),
    .Y(_0519_));
 sg13g2_a21oi_1 _2781_ (.A1(_1072_),
    .A2(_0981_),
    .Y(_0520_),
    .B1(_0519_));
 sg13g2_a22oi_1 _2782_ (.Y(_0521_),
    .B1(_0520_),
    .B2(_0139_),
    .A2(_0141_),
    .A1(_0838_));
 sg13g2_nor2_1 _2783_ (.A(net79),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_a21oi_1 _2784_ (.A1(_0842_),
    .A2(_0135_),
    .Y(_0523_),
    .B1(_0155_));
 sg13g2_or3_1 _2785_ (.A(_0006_),
    .B(_0749_),
    .C(net60),
    .X(_0524_));
 sg13g2_o21ai_1 _2786_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0839_),
    .A2(_0296_));
 sg13g2_or2_1 _2787_ (.X(_0526_),
    .B(_0237_),
    .A(_1008_));
 sg13g2_o21ai_1 _2788_ (.B1(_1402_),
    .Y(_0527_),
    .A1(net54),
    .A2(net43));
 sg13g2_a221oi_1 _2789_ (.B2(_0520_),
    .C1(_0527_),
    .B1(_0526_),
    .A1(net54),
    .Y(_0528_),
    .A2(_0525_));
 sg13g2_nor3_1 _2790_ (.A(_0199_),
    .B(_0523_),
    .C(_0528_),
    .Y(_0529_));
 sg13g2_nor3_1 _2791_ (.A(_0144_),
    .B(_0522_),
    .C(_0529_),
    .Y(_0530_));
 sg13g2_nor3_1 _2792_ (.A(net94),
    .B(_0518_),
    .C(_0530_),
    .Y(_0078_));
 sg13g2_nor2_1 _2793_ (.A(_0703_),
    .B(_0124_),
    .Y(_0531_));
 sg13g2_nand2b_1 _2794_ (.Y(_0532_),
    .B(net88),
    .A_N(_1094_));
 sg13g2_nand2b_1 _2795_ (.Y(_0533_),
    .B(_0532_),
    .A_N(_0274_));
 sg13g2_a22oi_1 _2796_ (.Y(_0534_),
    .B1(_0533_),
    .B2(net77),
    .A2(_0141_),
    .A1(net119));
 sg13g2_nor2_1 _2797_ (.A(net79),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_o21ai_1 _2798_ (.B1(_0192_),
    .Y(_0536_),
    .A1(_0841_),
    .A2(_0189_));
 sg13g2_nor2_1 _2799_ (.A(_1099_),
    .B(net59),
    .Y(_0537_));
 sg13g2_a21oi_1 _2800_ (.A1(net53),
    .A2(_0533_),
    .Y(_0538_),
    .B1(_0537_));
 sg13g2_a22oi_1 _2801_ (.Y(_0539_),
    .B1(net48),
    .B2(_0533_),
    .A2(_1095_),
    .A1(_0843_));
 sg13g2_o21ai_1 _2802_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_1032_),
    .A2(_0538_));
 sg13g2_nand2_1 _2803_ (.Y(_0541_),
    .A(_1446_),
    .B(_0540_));
 sg13g2_a21oi_1 _2804_ (.A1(_0536_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(net92));
 sg13g2_nor3_1 _2805_ (.A(_0144_),
    .B(_0535_),
    .C(_0542_),
    .Y(_0543_));
 sg13g2_nor3_1 _2806_ (.A(net94),
    .B(_0531_),
    .C(_0543_),
    .Y(_0079_));
 sg13g2_o21ai_1 _2807_ (.B1(_1458_),
    .Y(_0544_),
    .A1(\u8.rcip[1] ),
    .A2(_1406_));
 sg13g2_nand3_1 _2808_ (.B(_0199_),
    .C(_0544_),
    .A(net2),
    .Y(_0545_));
 sg13g2_nand4_1 _2809_ (.B(net2),
    .C(_0033_),
    .A(_1405_),
    .Y(_0546_),
    .D(_1448_));
 sg13g2_nand2_1 _2810_ (.Y(_0547_),
    .A(_1248_),
    .B(_0546_));
 sg13g2_a21oi_1 _2811_ (.A1(_1454_),
    .A2(_0545_),
    .Y(_0080_),
    .B1(_0547_));
 sg13g2_xnor2_1 _2812_ (.Y(_0548_),
    .A(_1451_),
    .B(_0546_));
 sg13g2_nor2_1 _2813_ (.A(_0184_),
    .B(_0548_),
    .Y(_0081_));
 sg13g2_nor2_1 _2814_ (.A(_1451_),
    .B(_0546_),
    .Y(_0549_));
 sg13g2_xnor2_1 _2815_ (.Y(_0550_),
    .A(_1406_),
    .B(_0549_));
 sg13g2_nor2_1 _2816_ (.A(_0184_),
    .B(_0550_),
    .Y(_0082_));
 sg13g2_a22oi_1 _2817_ (.Y(_0551_),
    .B1(_1207_),
    .B2(_0035_),
    .A2(_0799_),
    .A1(_0801_));
 sg13g2_nor2_1 _2818_ (.A(net96),
    .B(_0551_),
    .Y(_0083_));
 sg13g2_nand3_1 _2819_ (.B(net123),
    .C(_0798_),
    .A(net122),
    .Y(_0552_));
 sg13g2_xor2_1 _2820_ (.B(_0552_),
    .A(_0800_),
    .X(_0553_));
 sg13g2_nor2_1 _2821_ (.A(net96),
    .B(_0553_),
    .Y(_0084_));
 sg13g2_xnor2_1 _2822_ (.Y(_0554_),
    .A(\u8.rcop[2] ),
    .B(_0803_));
 sg13g2_nor2_1 _2823_ (.A(net96),
    .B(_0554_),
    .Y(_0085_));
 sg13g2_nor2_1 _2824_ (.A(_1221_),
    .B(_0209_),
    .Y(_0555_));
 sg13g2_a21o_1 _2825_ (.A2(_0113_),
    .A1(_0111_),
    .B1(_0526_),
    .X(_0556_));
 sg13g2_a21oi_1 _2826_ (.A1(_0655_),
    .A2(_0795_),
    .Y(_0557_),
    .B1(_1409_));
 sg13g2_o21ai_1 _2827_ (.B1(_0557_),
    .Y(_0558_),
    .A1(net143),
    .A2(_1406_));
 sg13g2_a21oi_1 _2828_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_nand3_1 _2829_ (.B(_0105_),
    .C(_0107_),
    .A(_0103_),
    .Y(_0560_));
 sg13g2_nand2_1 _2830_ (.Y(_0561_),
    .A(_0135_),
    .B(_0560_));
 sg13g2_nand3_1 _2831_ (.B(_1444_),
    .C(_0561_),
    .A(net143),
    .Y(_0562_));
 sg13g2_a21oi_1 _2832_ (.A1(_0559_),
    .A2(_0562_),
    .Y(_0563_),
    .B1(retry));
 sg13g2_nor2_1 _2833_ (.A(net93),
    .B(_0563_),
    .Y(_0086_));
 sg13g2_nor4_2 _2834_ (.A(net106),
    .B(_0655_),
    .C(_1278_),
    .Y(_0564_),
    .D(_1400_));
 sg13g2_nand2b_1 _2835_ (.Y(_0565_),
    .B(net105),
    .A_N(_0564_));
 sg13g2_nand2_1 _2836_ (.Y(_0566_),
    .A(_0034_),
    .B(_0564_));
 sg13g2_a21oi_1 _2837_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0087_),
    .B1(net110));
 sg13g2_nand2_1 _2838_ (.Y(_0567_),
    .A(net105),
    .B(_0564_));
 sg13g2_xnor2_1 _2839_ (.Y(_0568_),
    .A(_0764_),
    .B(_0567_));
 sg13g2_nor2_1 _2840_ (.A(_1365_),
    .B(_0568_),
    .Y(_0088_));
 sg13g2_nand3_1 _2841_ (.B(net104),
    .C(_0564_),
    .A(net105),
    .Y(_0569_));
 sg13g2_xor2_1 _2842_ (.B(_0569_),
    .A(_0735_),
    .X(_0570_));
 sg13g2_nor2_1 _2843_ (.A(_1365_),
    .B(_0570_),
    .Y(_0089_));
 sg13g2_and2_1 _2844_ (.A(net84),
    .B(_0811_),
    .X(_0571_));
 sg13g2_o21ai_1 _2845_ (.B1(_0739_),
    .Y(_0572_),
    .A1(_1469_),
    .A2(net91));
 sg13g2_a21oi_1 _2846_ (.A1(net4),
    .A2(_0572_),
    .Y(_0573_),
    .B1(_0768_));
 sg13g2_nor2_1 _2847_ (.A(_0695_),
    .B(_0815_),
    .Y(_0574_));
 sg13g2_and4_1 _2848_ (.A(net121),
    .B(net120),
    .C(_0844_),
    .D(_0846_),
    .X(_0575_));
 sg13g2_nand2_1 _2849_ (.Y(_0576_),
    .A(net119),
    .B(_0839_));
 sg13g2_a21oi_1 _2850_ (.A1(_1094_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0173_));
 sg13g2_nand3_1 _2851_ (.B(_0575_),
    .C(_0577_),
    .A(_0574_),
    .Y(_0578_));
 sg13g2_and2_1 _2852_ (.A(_0573_),
    .B(_0578_),
    .X(_0579_));
 sg13g2_inv_1 _2853_ (.Y(_0580_),
    .A(net128));
 sg13g2_xor2_1 _2854_ (.B(_0846_),
    .A(net98),
    .X(_0581_));
 sg13g2_nand2_1 _2855_ (.Y(_0582_),
    .A(net119),
    .B(_0575_));
 sg13g2_nor2_1 _2856_ (.A(_0580_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_a21oi_1 _2857_ (.A1(_0580_),
    .A2(_0581_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_nand2_1 _2858_ (.Y(_0585_),
    .A(net127),
    .B(_0091_));
 sg13g2_nor4_1 _2859_ (.A(_0695_),
    .B(_0815_),
    .C(_0584_),
    .D(_0585_),
    .Y(_0586_));
 sg13g2_and2_1 _2860_ (.A(_0839_),
    .B(_0845_),
    .X(_0587_));
 sg13g2_and2_1 _2861_ (.A(_0832_),
    .B(_0094_),
    .X(_0588_));
 sg13g2_nor2_1 _2862_ (.A(_0709_),
    .B(net113),
    .Y(_0589_));
 sg13g2_nand4_1 _2863_ (.B(_0847_),
    .C(_0588_),
    .A(_0587_),
    .Y(_0590_),
    .D(_0589_));
 sg13g2_a21oi_1 _2864_ (.A1(_0710_),
    .A2(_0590_),
    .Y(_0591_),
    .B1(_0096_));
 sg13g2_o21ai_1 _2865_ (.B1(_0768_),
    .Y(_0592_),
    .A1(_0832_),
    .A2(_0248_));
 sg13g2_o21ai_1 _2866_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_0109_),
    .A2(_0591_));
 sg13g2_o21ai_1 _2867_ (.B1(_0113_),
    .Y(_0594_),
    .A1(_0586_),
    .A2(_0593_));
 sg13g2_a22oi_1 _2868_ (.Y(_0595_),
    .B1(_0594_),
    .B2(_0768_),
    .A2(_0579_),
    .A1(_0571_));
 sg13g2_nor4_1 _2869_ (.A(_0839_),
    .B(_1338_),
    .C(_1140_),
    .D(_0582_),
    .Y(_0596_));
 sg13g2_nand2b_1 _2870_ (.Y(_0597_),
    .B(_1140_),
    .A_N(_0587_));
 sg13g2_a221oi_1 _2871_ (.B2(net97),
    .C1(_0961_),
    .B1(_0597_),
    .A1(net100),
    .Y(_0598_),
    .A2(_1309_));
 sg13g2_o21ai_1 _2872_ (.B1(_0854_),
    .Y(_0599_),
    .A1(_0596_),
    .A2(_0598_));
 sg13g2_nor3_1 _2873_ (.A(net140),
    .B(\u8.empty ),
    .C(net3),
    .Y(_0600_));
 sg13g2_nand2_1 _2874_ (.Y(_0601_),
    .A(_0599_),
    .B(_0600_));
 sg13g2_nand2_1 _2875_ (.Y(_0602_),
    .A(_0103_),
    .B(_0105_));
 sg13g2_nand3_1 _2876_ (.B(net3),
    .C(_0602_),
    .A(net107),
    .Y(_0603_));
 sg13g2_o21ai_1 _2877_ (.B1(_0603_),
    .Y(net29),
    .A1(_0595_),
    .A2(_0601_));
 sg13g2_nand2b_1 _2878_ (.Y(_0604_),
    .B(_0600_),
    .A_N(_0599_));
 sg13g2_nand2_1 _2879_ (.Y(_0605_),
    .A(retry),
    .B(net3));
 sg13g2_nand2_1 _2880_ (.Y(net30),
    .A(_0604_),
    .B(_0605_));
 sg13g2_o21ai_1 _2881_ (.B1(_0600_),
    .Y(_0606_),
    .A1(_0109_),
    .A2(_0113_));
 sg13g2_a21o_1 _2882_ (.A2(_0591_),
    .A1(_0110_),
    .B1(_0109_),
    .X(_0607_));
 sg13g2_nand2_1 _2883_ (.Y(_0608_),
    .A(_0736_),
    .B(_0737_));
 sg13g2_a21oi_1 _2884_ (.A1(_0660_),
    .A2(_0608_),
    .Y(_0609_),
    .B1(_0661_));
 sg13g2_a21o_1 _2885_ (.A2(_0663_),
    .A1(_0682_),
    .B1(_0609_),
    .X(_0610_));
 sg13g2_nand2_1 _2886_ (.Y(_0611_),
    .A(_0817_),
    .B(_0610_));
 sg13g2_o21ai_1 _2887_ (.B1(_0824_),
    .Y(_0612_),
    .A1(_1041_),
    .A2(_0827_));
 sg13g2_a21oi_1 _2888_ (.A1(_0092_),
    .A2(_0093_),
    .Y(_0613_),
    .B1(_1111_));
 sg13g2_o21ai_1 _2889_ (.B1(_0816_),
    .Y(_0614_),
    .A1(_0613_),
    .A2(_0588_));
 sg13g2_nand3_1 _2890_ (.B(_0097_),
    .C(_0614_),
    .A(_0812_),
    .Y(_0615_));
 sg13g2_nand2b_1 _2891_ (.Y(_0616_),
    .B(_0615_),
    .A_N(_0612_));
 sg13g2_a21oi_1 _2892_ (.A1(_0098_),
    .A2(_0616_),
    .Y(_0617_),
    .B1(net131));
 sg13g2_o21ai_1 _2893_ (.B1(_0821_),
    .Y(_0618_),
    .A1(_1470_),
    .A2(_0617_));
 sg13g2_and3_1 _2894_ (.X(_0619_),
    .A(_0102_),
    .B(_0611_),
    .C(_0618_));
 sg13g2_nand3_1 _2895_ (.B(net3),
    .C(_0572_),
    .A(net107),
    .Y(_0620_));
 sg13g2_nor2_1 _2896_ (.A(_0028_),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_o21ai_1 _2897_ (.B1(_0621_),
    .Y(_0622_),
    .A1(_0104_),
    .A2(_0619_));
 sg13g2_o21ai_1 _2898_ (.B1(_0622_),
    .Y(net31),
    .A1(_0606_),
    .A2(_0607_));
 sg13g2_nand3_1 _2899_ (.B(_0097_),
    .C(_0588_),
    .A(_0816_),
    .Y(_0623_));
 sg13g2_nand2_1 _2900_ (.Y(_0624_),
    .A(_0812_),
    .B(_0623_));
 sg13g2_nor4_1 _2901_ (.A(net131),
    .B(_1112_),
    .C(_1468_),
    .D(_0612_),
    .Y(_0625_));
 sg13g2_a21oi_1 _2902_ (.A1(_0624_),
    .A2(_0625_),
    .Y(_0626_),
    .B1(_1470_));
 sg13g2_nor4_1 _2903_ (.A(_1183_),
    .B(_0682_),
    .C(_1468_),
    .D(_0626_),
    .Y(_0627_));
 sg13g2_nor3_1 _2904_ (.A(_0028_),
    .B(_0806_),
    .C(_0620_),
    .Y(_0628_));
 sg13g2_o21ai_1 _2905_ (.B1(_0628_),
    .Y(_0629_),
    .A1(_0609_),
    .A2(_0627_));
 sg13g2_inv_1 _2906_ (.Y(_0630_),
    .A(_0606_));
 sg13g2_o21ai_1 _2907_ (.B1(_0630_),
    .Y(_0631_),
    .A1(_0111_),
    .A2(_0573_));
 sg13g2_nand2_1 _2908_ (.Y(net32),
    .A(_0629_),
    .B(_0631_));
 sg13g2_nor3_1 _2909_ (.A(net125),
    .B(net130),
    .C(_0848_),
    .Y(_0632_));
 sg13g2_a21oi_1 _2910_ (.A1(_1377_),
    .A2(_0848_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_nor2b_1 _2911_ (.A(_0834_),
    .B_N(_0826_),
    .Y(_0634_));
 sg13g2_nand4_1 _2912_ (.B(_0279_),
    .C(_0111_),
    .A(_1326_),
    .Y(_0635_),
    .D(_0634_));
 sg13g2_nand2_1 _2913_ (.Y(_0636_),
    .A(_0573_),
    .B(_0578_));
 sg13g2_o21ai_1 _2914_ (.B1(_0592_),
    .Y(_0637_),
    .A1(_0571_),
    .A2(_0636_));
 sg13g2_nand2_1 _2915_ (.Y(_0638_),
    .A(_0607_),
    .B(_0637_));
 sg13g2_o21ai_1 _2916_ (.B1(_0638_),
    .Y(_0639_),
    .A1(_0633_),
    .A2(_0635_));
 sg13g2_nand2_1 _2917_ (.Y(_0640_),
    .A(_0630_),
    .B(_0639_));
 sg13g2_o21ai_1 _2918_ (.B1(_0640_),
    .Y(net33),
    .A1(_0657_),
    .A2(_0620_));
 sg13g2_nand2_1 _2919_ (.Y(_0641_),
    .A(net4),
    .B(_0572_));
 sg13g2_nor3_1 _2920_ (.A(_0657_),
    .B(_0869_),
    .C(_0641_),
    .Y(_0642_));
 sg13g2_o21ai_1 _2921_ (.B1(net3),
    .Y(_0643_),
    .A1(retry),
    .A2(_0642_));
 sg13g2_nand2_1 _2922_ (.Y(_0644_),
    .A(_0109_),
    .B(_0641_));
 sg13g2_nor2_1 _2923_ (.A(net98),
    .B(_1305_),
    .Y(_0645_));
 sg13g2_o21ai_1 _2924_ (.B1(_0580_),
    .Y(_0646_),
    .A1(_0585_),
    .A2(_0645_));
 sg13g2_a21o_1 _2925_ (.A2(_1305_),
    .A1(_1254_),
    .B1(net128),
    .X(_0647_));
 sg13g2_o21ai_1 _2926_ (.B1(_0647_),
    .Y(_0648_),
    .A1(_0173_),
    .A2(_0582_));
 sg13g2_nand4_1 _2927_ (.B(_0574_),
    .C(_0646_),
    .A(_0768_),
    .Y(_0649_),
    .D(_0648_));
 sg13g2_o21ai_1 _2928_ (.B1(_0649_),
    .Y(_0650_),
    .A1(_0644_),
    .A2(_0578_));
 sg13g2_nand3b_1 _2929_ (.B(_0630_),
    .C(_0650_),
    .Y(_0651_),
    .A_N(_0593_));
 sg13g2_nand4_1 _2930_ (.B(_0629_),
    .C(_0643_),
    .A(_0622_),
    .Y(net34),
    .D(_0651_));
 sg13g2_nand2_1 _2931_ (.Y(_0652_),
    .A(net144),
    .B(_1278_));
 sg13g2_o21ai_1 _2932_ (.B1(_0652_),
    .Y(net35),
    .A1(net144),
    .A2(_1007_));
 sg13g2_mux2_1 _2933_ (.A0(_1157_),
    .A1(_0917_),
    .S(net106),
    .X(_0653_));
 sg13g2_inv_1 _2934_ (.Y(net36),
    .A(_0653_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2936_ (.A(ui_in[4]),
    .X(net13));
 sg13g2_buf_1 _2937_ (.A(ui_in[4]),
    .X(net14));
 sg13g2_buf_1 _2938_ (.A(ui_in[4]),
    .X(net15));
 sg13g2_buf_1 _2939_ (.A(ui_in[4]),
    .X(net16));
 sg13g2_buf_1 _2940_ (.A(ui_in[4]),
    .X(net17));
 sg13g2_buf_1 _2941_ (.A(ui_in[4]),
    .X(net18));
 sg13g2_buf_1 _2942_ (.A(ui_in[4]),
    .X(net19));
 sg13g2_buf_1 _2943_ (.A(ui_in[4]),
    .X(net20));
 sg13g2_dfrbp_1 \u8.dout[0]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net145),
    .D(_0036_),
    .Q_N(_1489_),
    .Q(net21));
 sg13g2_dfrbp_1 \u8.dout[1]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net146),
    .D(_0037_),
    .Q_N(_1488_),
    .Q(net22));
 sg13g2_dfrbp_1 \u8.dout[2]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net147),
    .D(_0038_),
    .Q_N(_1487_),
    .Q(net23));
 sg13g2_dfrbp_1 \u8.dout[3]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net148),
    .D(_0039_),
    .Q_N(_1486_),
    .Q(net24));
 sg13g2_dfrbp_1 \u8.dout[4]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net149),
    .D(_0040_),
    .Q_N(_1485_),
    .Q(net25));
 sg13g2_dfrbp_1 \u8.dout[5]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net150),
    .D(_0041_),
    .Q_N(_1484_),
    .Q(net26));
 sg13g2_dfrbp_1 \u8.dout[6]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net151),
    .D(_0042_),
    .Q_N(_1483_),
    .Q(net27));
 sg13g2_dfrbp_1 \u8.dout[7]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net152),
    .D(_0043_),
    .Q_N(_1482_),
    .Q(net28));
 sg13g2_dfrbp_1 \u8.empty$_SDFFE_PN1P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net153),
    .D(_0044_),
    .Q_N(_0013_),
    .Q(\u8.empty ));
 sg13g2_dfrbp_1 \u8.rbop[0]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net154),
    .D(_0045_),
    .Q_N(_1481_),
    .Q(\u8.rbop[0] ));
 sg13g2_dfrbp_1 \u8.rbop[1]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net155),
    .D(_0046_),
    .Q_N(_1480_),
    .Q(\u8.rbop[1] ));
 sg13g2_dfrbp_1 \u8.rbop[2]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net156),
    .D(_0047_),
    .Q_N(_0018_),
    .Q(\u8.rbop[2] ));
 sg13g2_dfrbp_1 \u8.rc[0]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net157),
    .D(_0048_),
    .Q_N(_0000_),
    .Q(\u8.ls[0] ));
 sg13g2_dfrbp_1 \u8.rc[10]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net158),
    .D(_0049_),
    .Q_N(_0002_),
    .Q(\u8.hs[0] ));
 sg13g2_dfrbp_1 \u8.rc[11]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net159),
    .D(_0050_),
    .Q_N(_0029_),
    .Q(\u8.hs[1] ));
 sg13g2_dfrbp_1 \u8.rc[12]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net160),
    .D(_0051_),
    .Q_N(_0003_),
    .Q(\u8.hs[2] ));
 sg13g2_dfrbp_1 \u8.rc[13]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net161),
    .D(_0052_),
    .Q_N(_0021_),
    .Q(\u8.hs[3] ));
 sg13g2_dfrbp_1 \u8.rc[14]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net162),
    .D(_0053_),
    .Q_N(_0004_),
    .Q(\u8.hs[4] ));
 sg13g2_dfrbp_1 \u8.rc[15]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net163),
    .D(_0054_),
    .Q_N(_0005_),
    .Q(\u8.hs[5] ));
 sg13g2_dfrbp_1 \u8.rc[16]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net164),
    .D(_0055_),
    .Q_N(_0006_),
    .Q(\u8.rc[16] ));
 sg13g2_dfrbp_1 \u8.rc[17]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net165),
    .D(_0056_),
    .Q_N(_0007_),
    .Q(\u8.rc[17] ));
 sg13g2_dfrbp_1 \u8.rc[18]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net166),
    .D(_0057_),
    .Q_N(_0008_),
    .Q(\u8.rc[18] ));
 sg13g2_dfrbp_1 \u8.rc[19]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net167),
    .D(_0058_),
    .Q_N(_0031_),
    .Q(\u8.rc[19] ));
 sg13g2_dfrbp_1 \u8.rc[1]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net168),
    .D(_0059_),
    .Q_N(_0030_),
    .Q(\u8.ls[1] ));
 sg13g2_dfrbp_1 \u8.rc[20]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net169),
    .D(_0060_),
    .Q_N(_0009_),
    .Q(\u8.rc[20] ));
 sg13g2_dfrbp_1 \u8.rc[21]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net170),
    .D(_0061_),
    .Q_N(_0020_),
    .Q(\u8.rc[21] ));
 sg13g2_dfrbp_1 \u8.rc[22]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net171),
    .D(_0062_),
    .Q_N(_0010_),
    .Q(\u8.rc[22] ));
 sg13g2_dfrbp_1 \u8.rc[23]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net172),
    .D(_0063_),
    .Q_N(_0011_),
    .Q(\u8.rc[23] ));
 sg13g2_dfrbp_1 \u8.rc[24]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net173),
    .D(_0064_),
    .Q_N(_0015_),
    .Q(\u8.rc[24] ));
 sg13g2_dfrbp_1 \u8.rc[25]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net174),
    .D(_0065_),
    .Q_N(_0019_),
    .Q(\u8.rc[25] ));
 sg13g2_dfrbp_1 \u8.rc[26]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net175),
    .D(_0066_),
    .Q_N(_0016_),
    .Q(\u8.rc[26] ));
 sg13g2_dfrbp_1 \u8.rc[27]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net176),
    .D(_0067_),
    .Q_N(_0017_),
    .Q(\u8.rc[27] ));
 sg13g2_dfrbp_1 \u8.rc[28]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net177),
    .D(_0068_),
    .Q_N(_1479_),
    .Q(\u8.rc[28] ));
 sg13g2_dfrbp_1 \u8.rc[29]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net178),
    .D(_0069_),
    .Q_N(_1478_),
    .Q(\u8.rc[29] ));
 sg13g2_dfrbp_1 \u8.rc[2]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net179),
    .D(_0070_),
    .Q_N(_0023_),
    .Q(\u8.ls[2] ));
 sg13g2_dfrbp_1 \u8.rc[30]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net180),
    .D(_0071_),
    .Q_N(_1477_),
    .Q(\u8.rc[30] ));
 sg13g2_dfrbp_1 \u8.rc[31]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net181),
    .D(_0072_),
    .Q_N(_0028_),
    .Q(\u8.rc[31] ));
 sg13g2_dfrbp_1 \u8.rc[3]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net182),
    .D(_0073_),
    .Q_N(_0024_),
    .Q(\u8.ls[3] ));
 sg13g2_dfrbp_1 \u8.rc[4]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net183),
    .D(_0074_),
    .Q_N(_0025_),
    .Q(\u8.ls[4] ));
 sg13g2_dfrbp_1 \u8.rc[5]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net184),
    .D(_0075_),
    .Q_N(_0026_),
    .Q(\u8.ls[5] ));
 sg13g2_dfrbp_1 \u8.rc[6]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net185),
    .D(_0076_),
    .Q_N(_0027_),
    .Q(\u8.ls[6] ));
 sg13g2_dfrbp_1 \u8.rc[7]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net186),
    .D(_0077_),
    .Q_N(_0014_),
    .Q(\u8.ls[7] ));
 sg13g2_dfrbp_1 \u8.rc[8]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net187),
    .D(_0078_),
    .Q_N(_0001_),
    .Q(\u8.ls[8] ));
 sg13g2_dfrbp_1 \u8.rc[9]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net188),
    .D(_0079_),
    .Q_N(_0022_),
    .Q(\u8.ls[9] ));
 sg13g2_dfrbp_1 \u8.rcip[0]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net189),
    .D(_0080_),
    .Q_N(_1476_),
    .Q(\u8.rcip[0] ));
 sg13g2_dfrbp_1 \u8.rcip[1]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net190),
    .D(_0081_),
    .Q_N(_1475_),
    .Q(\u8.rcip[1] ));
 sg13g2_dfrbp_1 \u8.rcip[2]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net191),
    .D(_0082_),
    .Q_N(_0033_),
    .Q(\u8.rcip[2] ));
 sg13g2_dfrbp_1 \u8.rcop[0]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net192),
    .D(_0083_),
    .Q_N(_0035_),
    .Q(\u8.rcop[0] ));
 sg13g2_dfrbp_1 \u8.rcop[1]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net193),
    .D(_0084_),
    .Q_N(_1474_),
    .Q(\u8.rcop[1] ));
 sg13g2_dfrbp_1 \u8.rcop[2]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net194),
    .D(_0085_),
    .Q_N(_0012_),
    .Q(\u8.rcop[2] ));
 sg13g2_dfrbp_1 \u8.retry$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net195),
    .D(_0086_),
    .Q_N(_1473_),
    .Q(retry));
 sg13g2_dfrbp_1 \u8.ruop[0]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net196),
    .D(_0087_),
    .Q_N(_0034_),
    .Q(\u8.ruop[0] ));
 sg13g2_dfrbp_1 \u8.ruop[1]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net197),
    .D(_0088_),
    .Q_N(_1472_),
    .Q(\u8.ruop[1] ));
 sg13g2_dfrbp_1 \u8.ruop[2]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net198),
    .D(_0089_),
    .Q_N(_0032_),
    .Q(\u8.ruop[2] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[7]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[0]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[1]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[3]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[4]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[5]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[6]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[7]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[0]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[1]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[2]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[3]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[4]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[5]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[6]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout37 (.A(_0146_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0943_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0149_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0383_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0234_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0939_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0296_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1446_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1009_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0988_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0242_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1417_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1315_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1032_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1008_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0990_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1437_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1266_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0872_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0857_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0851_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0189_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1438_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1436_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1221_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1095_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1007_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0873_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0861_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0256_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0231_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0135_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0129_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1082_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1072_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1040_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1028_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1016_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0911_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0825_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0139_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0128_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1450_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1052_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1035_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1015_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0882_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0729_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0311_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1460_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1132_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1034_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1019_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1014_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0723_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0199_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0184_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0127_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1444_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1365_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1305_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1254_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1236_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1140_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1041_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1022_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1018_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0784_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0761_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0752_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0746_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1326_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1096_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1092_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1017_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1012_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0980_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0961_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0883_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0869_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0863_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0852_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0843_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0842_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0841_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0801_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0797_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0714_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0708_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_0706_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_0704_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0703_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0697_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0693_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0680_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0678_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0677_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_0675_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0674_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_0670_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0668_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_0667_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0665_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0657_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1248_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1011_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0793_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0742_),
    .X(net144));
 sg13g2_tiehi \u8.dout[0]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \u8.dout[1]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \u8.dout[2]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \u8.dout[3]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \u8.dout[4]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \u8.dout[5]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \u8.dout[6]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \u8.dout[7]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \u8.empty$_SDFFE_PN1P__153  (.L_HI(net153));
 sg13g2_tiehi \u8.rbop[0]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \u8.rbop[1]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \u8.rbop[2]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \u8.rc[0]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \u8.rc[10]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \u8.rc[11]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \u8.rc[12]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \u8.rc[13]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \u8.rc[14]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \u8.rc[15]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \u8.rc[16]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \u8.rc[17]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \u8.rc[18]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \u8.rc[19]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \u8.rc[1]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \u8.rc[20]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \u8.rc[21]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \u8.rc[22]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \u8.rc[23]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \u8.rc[24]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \u8.rc[25]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \u8.rc[26]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \u8.rc[27]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \u8.rc[28]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \u8.rc[29]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \u8.rc[2]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \u8.rc[30]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \u8.rc[31]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \u8.rc[3]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \u8.rc[4]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \u8.rc[5]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \u8.rc[6]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \u8.rc[7]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \u8.rc[8]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \u8.rc[9]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \u8.rcip[0]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \u8.rcip[1]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \u8.rcip[2]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \u8.rcop[0]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \u8.rcop[1]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \u8.rcop[2]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \u8.retry$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \u8.ruop[0]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \u8.ruop[1]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \u8.ruop[2]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_227 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_fill_2 FILLER_3_239 ();
 sg13g2_decap_4 FILLER_3_285 ();
 sg13g2_decap_4 FILLER_3_332 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_411 ();
 sg13g2_decap_8 FILLER_3_418 ();
 sg13g2_decap_4 FILLER_3_425 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_119 ();
 sg13g2_fill_1 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_148 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_decap_4 FILLER_4_156 ();
 sg13g2_fill_1 FILLER_4_160 ();
 sg13g2_fill_2 FILLER_4_166 ();
 sg13g2_decap_8 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_180 ();
 sg13g2_decap_4 FILLER_4_186 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_2 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_fill_2 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_223 ();
 sg13g2_decap_4 FILLER_4_250 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_fill_2 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_fill_1 FILLER_4_273 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_decap_4 FILLER_4_287 ();
 sg13g2_fill_2 FILLER_4_291 ();
 sg13g2_fill_2 FILLER_4_321 ();
 sg13g2_fill_2 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_404 ();
 sg13g2_decap_8 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_12 ();
 sg13g2_decap_8 FILLER_5_19 ();
 sg13g2_fill_2 FILLER_5_26 ();
 sg13g2_fill_1 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_64 ();
 sg13g2_decap_8 FILLER_5_71 ();
 sg13g2_decap_8 FILLER_5_78 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_4 FILLER_5_99 ();
 sg13g2_fill_1 FILLER_5_103 ();
 sg13g2_decap_4 FILLER_5_130 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_decap_4 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_decap_4 FILLER_5_208 ();
 sg13g2_fill_1 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_2 FILLER_5_236 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_4 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_255 ();
 sg13g2_decap_4 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_decap_4 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_fill_2 FILLER_5_345 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_4 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_80 ();
 sg13g2_decap_8 FILLER_6_87 ();
 sg13g2_decap_8 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_108 ();
 sg13g2_fill_1 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_115 ();
 sg13g2_decap_8 FILLER_6_122 ();
 sg13g2_decap_8 FILLER_6_129 ();
 sg13g2_decap_8 FILLER_6_136 ();
 sg13g2_decap_4 FILLER_6_143 ();
 sg13g2_fill_2 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_179 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_8 FILLER_6_250 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_340 ();
 sg13g2_decap_4 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_8 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_6_412 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_4 FILLER_6_426 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_18 ();
 sg13g2_fill_1 FILLER_7_20 ();
 sg13g2_decap_8 FILLER_7_40 ();
 sg13g2_fill_1 FILLER_7_47 ();
 sg13g2_fill_2 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_61 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_decap_4 FILLER_7_90 ();
 sg13g2_decap_8 FILLER_7_99 ();
 sg13g2_decap_8 FILLER_7_106 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_decap_4 FILLER_7_120 ();
 sg13g2_fill_2 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_136 ();
 sg13g2_fill_2 FILLER_7_143 ();
 sg13g2_fill_2 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_158 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_fill_2 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_decap_4 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_decap_8 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_decap_4 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_259 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_decap_4 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_20 ();
 sg13g2_decap_4 FILLER_8_26 ();
 sg13g2_decap_8 FILLER_8_34 ();
 sg13g2_decap_4 FILLER_8_41 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_fill_2 FILLER_8_71 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_fill_2 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_159 ();
 sg13g2_fill_1 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_4 FILLER_8_186 ();
 sg13g2_fill_2 FILLER_8_190 ();
 sg13g2_decap_8 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_208 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_decap_4 FILLER_8_226 ();
 sg13g2_decap_4 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_238 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_4 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_fill_2 FILLER_8_308 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_fill_2 FILLER_8_320 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_fill_2 FILLER_8_340 ();
 sg13g2_decap_4 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_4 FILLER_8_386 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_404 ();
 sg13g2_decap_8 FILLER_8_411 ();
 sg13g2_decap_8 FILLER_8_418 ();
 sg13g2_decap_4 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_23 ();
 sg13g2_fill_1 FILLER_9_35 ();
 sg13g2_decap_4 FILLER_9_62 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_decap_4 FILLER_9_81 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_fill_2 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_103 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_decap_4 FILLER_9_232 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_decap_4 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_4 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_decap_4 FILLER_9_364 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_373 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_37 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_88 ();
 sg13g2_fill_1 FILLER_10_90 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_4 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_4 FILLER_10_144 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_186 ();
 sg13g2_fill_2 FILLER_10_214 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_decap_4 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_decap_4 FILLER_10_253 ();
 sg13g2_fill_2 FILLER_10_262 ();
 sg13g2_decap_4 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_decap_4 FILLER_10_298 ();
 sg13g2_decap_4 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_344 ();
 sg13g2_fill_2 FILLER_10_351 ();
 sg13g2_fill_1 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_fill_2 FILLER_10_399 ();
 sg13g2_fill_1 FILLER_10_401 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_26 ();
 sg13g2_fill_1 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_decap_4 FILLER_11_78 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_decap_4 FILLER_11_87 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_fill_2 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_4 FILLER_11_256 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_4 FILLER_11_294 ();
 sg13g2_decap_4 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_decap_4 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_fill_1 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_48 ();
 sg13g2_fill_1 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_79 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_decap_4 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_decap_4 FILLER_12_142 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_2 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_232 ();
 sg13g2_decap_4 FILLER_12_239 ();
 sg13g2_fill_2 FILLER_12_243 ();
 sg13g2_decap_4 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_2 FILLER_12_368 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_22 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_37 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_decap_4 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_74 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_114 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_decap_8 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_155 ();
 sg13g2_fill_2 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_212 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_4 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_fill_2 FILLER_13_359 ();
 sg13g2_decap_4 FILLER_13_365 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_29 ();
 sg13g2_decap_4 FILLER_14_36 ();
 sg13g2_decap_8 FILLER_14_51 ();
 sg13g2_fill_2 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_68 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_4 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_88 ();
 sg13g2_decap_4 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_4 FILLER_14_275 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_decap_4 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_370 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_fill_2 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_1 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_414 ();
 sg13g2_decap_8 FILLER_14_421 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_30 ();
 sg13g2_fill_2 FILLER_15_54 ();
 sg13g2_decap_8 FILLER_15_66 ();
 sg13g2_decap_4 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_decap_4 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_decap_4 FILLER_15_122 ();
 sg13g2_fill_2 FILLER_15_131 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_decap_4 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_173 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_2 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_4 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_2 FILLER_15_367 ();
 sg13g2_decap_4 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_decap_8 FILLER_16_47 ();
 sg13g2_decap_4 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_115 ();
 sg13g2_fill_1 FILLER_16_117 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_decap_4 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_decap_4 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_4 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_4 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_295 ();
 sg13g2_decap_4 FILLER_16_307 ();
 sg13g2_decap_4 FILLER_16_319 ();
 sg13g2_decap_4 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_decap_4 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_fill_2 FILLER_16_399 ();
 sg13g2_fill_1 FILLER_16_401 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_27 ();
 sg13g2_decap_8 FILLER_17_34 ();
 sg13g2_decap_4 FILLER_17_41 ();
 sg13g2_fill_2 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_4 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_decap_4 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_284 ();
 sg13g2_decap_4 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_decap_4 FILLER_17_336 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_fill_1 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_8 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_29 ();
 sg13g2_decap_8 FILLER_18_36 ();
 sg13g2_decap_8 FILLER_18_43 ();
 sg13g2_decap_8 FILLER_18_50 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_decap_4 FILLER_18_64 ();
 sg13g2_decap_4 FILLER_18_90 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_4 FILLER_18_193 ();
 sg13g2_decap_4 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_decap_4 FILLER_18_278 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_decap_4 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_8 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_decap_8 FILLER_19_50 ();
 sg13g2_decap_4 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_decap_8 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_decap_8 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_fill_2 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_222 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_decap_4 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_391 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_31 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_decap_8 FILLER_20_45 ();
 sg13g2_fill_2 FILLER_20_52 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_141 ();
 sg13g2_fill_1 FILLER_20_145 ();
 sg13g2_decap_4 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_167 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_decap_4 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_27 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_121 ();
 sg13g2_decap_4 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_185 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_412 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_18 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_41 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_decap_4 FILLER_22_113 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_decap_4 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_decap_4 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_decap_4 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_decap_4 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_4 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_4 FILLER_23_424 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_20 ();
 sg13g2_fill_1 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_33 ();
 sg13g2_fill_2 FILLER_24_45 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_76 ();
 sg13g2_decap_4 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_183 ();
 sg13g2_decap_4 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_decap_4 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_decap_4 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_324 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_393 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_decap_4 FILLER_25_19 ();
 sg13g2_decap_4 FILLER_25_31 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_136 ();
 sg13g2_decap_4 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_decap_4 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_4 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_decap_4 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_4 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_17 ();
 sg13g2_decap_8 FILLER_26_24 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_8 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_45 ();
 sg13g2_fill_2 FILLER_26_62 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_decap_4 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_decap_4 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_decap_4 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_30 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_decap_4 FILLER_27_79 ();
 sg13g2_decap_4 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_decap_4 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_decap_4 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_384 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_decap_4 FILLER_28_17 ();
 sg13g2_decap_8 FILLER_28_27 ();
 sg13g2_decap_8 FILLER_28_34 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_decap_4 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_2 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_decap_4 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_decap_4 FILLER_28_179 ();
 sg13g2_decap_4 FILLER_28_187 ();
 sg13g2_decap_4 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_decap_4 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_4 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_decap_4 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_decap_4 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_decap_8 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_12 ();
 sg13g2_fill_1 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_19 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_33 ();
 sg13g2_decap_8 FILLER_30_40 ();
 sg13g2_decap_4 FILLER_30_47 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_decap_4 FILLER_30_58 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_4 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_32 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_decap_8 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_decap_4 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_decap_4 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_decap_4 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_234 ();
 sg13g2_decap_4 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_decap_4 FILLER_31_400 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_fill_2 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_4 FILLER_31_422 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_12 ();
 sg13g2_decap_8 FILLER_32_19 ();
 sg13g2_decap_4 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_decap_4 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_decap_4 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_247 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_4 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_68 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_decap_4 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_decap_4 FILLER_34_32 ();
 sg13g2_fill_1 FILLER_34_41 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_4 FILLER_34_80 ();
 sg13g2_decap_8 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_118 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_decap_4 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_4 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_251 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_25 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_2 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_decap_4 FILLER_35_67 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_decap_4 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_decap_4 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_23 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_2 FILLER_36_43 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_decap_8 FILLER_36_51 ();
 sg13g2_decap_8 FILLER_36_58 ();
 sg13g2_decap_8 FILLER_36_65 ();
 sg13g2_decap_4 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_111 ();
 sg13g2_decap_8 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_4 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_293 ();
 sg13g2_decap_8 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_405 ();
 sg13g2_fill_1 FILLER_36_412 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_decap_4 FILLER_37_45 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_fill_1 FILLER_37_74 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_114 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_4 FILLER_37_190 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_11 ();
 sg13g2_fill_2 FILLER_38_18 ();
 sg13g2_fill_1 FILLER_38_20 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_decap_4 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_4 FILLER_38_349 ();
 sg13g2_decap_4 FILLER_38_361 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
