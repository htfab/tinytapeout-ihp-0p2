module tt_um_algofoogle_tinyvga_fun_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire clknet_0_clk;
 wire net83;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[2] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \depth[0] ;
 wire \depth[1] ;
 wire \depth[2] ;
 wire \dither_threshold[0] ;
 wire \dither_threshold[1] ;
 wire \dither_threshold[2] ;
 wire \dither_threshold[3] ;
 wire \dither_threshold[4] ;
 wire \dither_threshold[5] ;
 wire \dither_threshold[6] ;
 wire hsync;
 wire \i_project.controller_0.divider[0] ;
 wire \i_project.controller_0.divider[1] ;
 wire \i_project.controller_0.grey_pass[10] ;
 wire \i_project.controller_0.grey_pass[11] ;
 wire \i_project.controller_0.grey_pass[12] ;
 wire \i_project.controller_0.grey_pass[13] ;
 wire \i_project.controller_0.grey_pass[14] ;
 wire \i_project.controller_0.grey_pass[15] ;
 wire \i_project.controller_0.h[0] ;
 wire \i_project.controller_0.h[1] ;
 wire \i_project.controller_0.h[2] ;
 wire \i_project.controller_0.h[3] ;
 wire \i_project.controller_0.h[4] ;
 wire \i_project.controller_0.h[5] ;
 wire \i_project.controller_0.h[6] ;
 wire \i_project.controller_0.h[7] ;
 wire \i_project.controller_0.h[8] ;
 wire \i_project.controller_0.h[9] ;
 wire \i_project.controller_0.mode[0] ;
 wire \i_project.controller_0.mode[1] ;
 wire \i_project.controller_0.mode[2] ;
 wire \i_project.controller_0.mode_ramp_base[0] ;
 wire \i_project.controller_0.mode_ramp_base[1] ;
 wire \i_project.controller_0.mode_ramp_base[2] ;
 wire \i_project.controller_0.mode_ramp_base[3] ;
 wire \i_project.controller_0.mode_ramp_base[4] ;
 wire \i_project.controller_0.mode_ramp_base[5] ;
 wire \i_project.controller_0.mode_ramp_base[6] ;
 wire \i_project.controller_0.mode_ramp_base[7] ;
 wire \i_project.controller_0.rst_n ;
 wire \i_project.controller_0.t[10] ;
 wire \i_project.controller_0.t[11] ;
 wire \i_project.controller_0.t[8] ;
 wire \i_project.controller_0.t[9] ;
 wire \i_project.controller_0.v[0] ;
 wire \i_project.controller_0.v[1] ;
 wire \i_project.controller_0.v[2] ;
 wire \i_project.controller_0.v[3] ;
 wire \i_project.controller_0.v[4] ;
 wire \i_project.controller_0.v[5] ;
 wire \i_project.controller_0.v[6] ;
 wire \i_project.controller_0.v[7] ;
 wire \i_project.controller_0.v[8] ;
 wire \i_project.controller_0.v[9] ;
 wire \i_project.controller_0.vga_sync.hsync ;
 wire \i_project.controller_0.vga_sync.mode ;
 wire \i_project.controller_0.vga_sync.o_vsync ;
 wire \i_project.controller_0.vga_sync.vsync ;
 wire \i_project.controller_0.voffset[0] ;
 wire \i_project.controller_0.voffset[1] ;
 wire \i_project.controller_0.voffset[2] ;
 wire \i_project.controller_0.voffset[3] ;
 wire \i_project.controller_0.voffset[4] ;
 wire \i_project.controller_0.voffset[5] ;
 wire \i_project.controller_0.voffset[6] ;
 wire \i_project.controller_0.voffset[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_nor2b_1 _2265_ (.A(_0303_),
    .B_N(_0307_),
    .Y(_0308_));
 sg13g2_nand2_1 _2266_ (.Y(_0309_),
    .A(net18),
    .B(_0229_));
 sg13g2_nor2_1 _2267_ (.A(_0229_),
    .B(_0163_),
    .Y(_0310_));
 sg13g2_a21oi_1 _2268_ (.A1(_0309_),
    .A2(_0250_),
    .Y(_0311_),
    .B1(_0310_));
 sg13g2_nor2b_1 _2269_ (.A(_0308_),
    .B_N(_0311_),
    .Y(_0312_));
 sg13g2_nand2_1 _2270_ (.Y(_0313_),
    .A(_0305_),
    .B(_0312_));
 sg13g2_nand2_1 _2271_ (.Y(_0314_),
    .A(_0301_),
    .B(_0313_));
 sg13g2_nand3_1 _2272_ (.B(_0299_),
    .C(_0287_),
    .A(_0295_),
    .Y(_0315_));
 sg13g2_nand2_1 _2273_ (.Y(_0316_),
    .A(_0288_),
    .B(_0291_));
 sg13g2_nand2_1 _2274_ (.Y(_0317_),
    .A(_0316_),
    .B(_0294_));
 sg13g2_nand3_1 _2275_ (.B(_0291_),
    .C(_0298_),
    .A(_0288_),
    .Y(_0318_));
 sg13g2_inv_1 _2276_ (.Y(_0319_),
    .A(_0287_));
 sg13g2_nand3_1 _2277_ (.B(_0318_),
    .C(_0319_),
    .A(_0317_),
    .Y(_0320_));
 sg13g2_nand2_1 _2278_ (.Y(_0321_),
    .A(_0315_),
    .B(_0320_));
 sg13g2_xnor2_1 _2279_ (.Y(_0322_),
    .A(_0237_),
    .B(net19));
 sg13g2_xnor2_1 _2280_ (.Y(_0323_),
    .A(_0229_),
    .B(_0163_));
 sg13g2_nor2_1 _2281_ (.A(_0322_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_nand2_1 _2282_ (.Y(_0325_),
    .A(_0324_),
    .B(_0307_));
 sg13g2_nand2_1 _2283_ (.Y(_0326_),
    .A(_0325_),
    .B(_0311_));
 sg13g2_nor2_1 _2284_ (.A(_0304_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nand2_1 _2285_ (.Y(_0328_),
    .A(_0321_),
    .B(_0327_));
 sg13g2_nand2_1 _2286_ (.Y(_0329_),
    .A(_0314_),
    .B(_0328_));
 sg13g2_nand2_1 _2287_ (.Y(_0330_),
    .A(_0329_),
    .B(net48));
 sg13g2_xnor2_1 _2288_ (.Y(_0331_),
    .A(net60),
    .B(_0168_));
 sg13g2_a21o_1 _2289_ (.A2(net47),
    .A1(_0331_),
    .B1(_2026_),
    .X(_0332_));
 sg13g2_nand2_1 _2290_ (.Y(_0333_),
    .A(_0330_),
    .B(_0332_));
 sg13g2_a21oi_1 _2291_ (.A1(_0256_),
    .A2(net50),
    .Y(_0334_),
    .B1(_2111_));
 sg13g2_nand2_1 _2292_ (.Y(_0335_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_a21oi_1 _2293_ (.A1(_1852_),
    .A2(_1580_),
    .Y(_0336_),
    .B1(_1583_));
 sg13g2_nand2b_1 _2294_ (.Y(_0337_),
    .B(net57),
    .A_N(_0049_));
 sg13g2_nand2_1 _2295_ (.Y(_0338_),
    .A(_1750_),
    .B(_1579_));
 sg13g2_o21ai_1 _2296_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_1579_),
    .A2(_0048_));
 sg13g2_inv_1 _2297_ (.Y(_0340_),
    .A(_0339_));
 sg13g2_a22oi_1 _2298_ (.Y(_0341_),
    .B1(_1584_),
    .B2(_0340_),
    .A2(_0337_),
    .A1(_0336_));
 sg13g2_xnor2_1 _2299_ (.Y(_0342_),
    .A(_0341_),
    .B(_2129_));
 sg13g2_a21oi_1 _2300_ (.A1(_0342_),
    .A2(net40),
    .Y(_0343_),
    .B1(net45));
 sg13g2_nand2_1 _2301_ (.Y(_0344_),
    .A(_0335_),
    .B(_0343_));
 sg13g2_a21oi_1 _2302_ (.A1(_0341_),
    .A2(net45),
    .Y(_0345_),
    .B1(net28));
 sg13g2_nand2_1 _2303_ (.Y(_0346_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nand2_1 _2304_ (.Y(_0347_),
    .A(_0346_),
    .B(_0276_));
 sg13g2_nand2_1 _2305_ (.Y(_0348_),
    .A(_0347_),
    .B(_0197_));
 sg13g2_buf_8 _2306_ (.A(_0348_),
    .X(_0349_));
 sg13g2_nor3_1 _2307_ (.A(_0178_),
    .B(_0187_),
    .C(_0203_),
    .Y(_0350_));
 sg13g2_buf_2 _2308_ (.A(_0350_),
    .X(_0351_));
 sg13g2_nand2_1 _2309_ (.Y(_0352_),
    .A(_1764_),
    .B(_0047_));
 sg13g2_nand4_1 _2310_ (.B(_0199_),
    .C(_0351_),
    .A(_0349_),
    .Y(_0353_),
    .D(_0352_));
 sg13g2_nor2_1 _2311_ (.A(_0203_),
    .B(_0180_),
    .Y(_0354_));
 sg13g2_inv_1 _2312_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_inv_2 _2313_ (.Y(_0356_),
    .A(_0199_));
 sg13g2_nor2_1 _2314_ (.A(_0355_),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_buf_2 _2315_ (.A(_0357_),
    .X(_0358_));
 sg13g2_buf_1 _2316_ (.A(_0352_),
    .X(_0359_));
 sg13g2_nand3_1 _2317_ (.B(_0358_),
    .C(net44),
    .A(_0349_),
    .Y(_0360_));
 sg13g2_nand3_1 _2318_ (.B(_0353_),
    .C(_0360_),
    .A(_0284_),
    .Y(_0361_));
 sg13g2_xnor2_1 _2319_ (.Y(_0362_),
    .A(_1658_),
    .B(_2009_));
 sg13g2_a21oi_1 _2320_ (.A1(_0319_),
    .A2(_0293_),
    .Y(_0363_),
    .B1(_0292_));
 sg13g2_xor2_1 _2321_ (.B(_0363_),
    .A(_0362_),
    .X(_0364_));
 sg13g2_xor2_1 _2322_ (.B(_2191_),
    .A(_2009_),
    .X(_0365_));
 sg13g2_nor2_1 _2323_ (.A(_0323_),
    .B(_0316_),
    .Y(_0366_));
 sg13g2_inv_1 _2324_ (.Y(_0367_),
    .A(_0251_));
 sg13g2_nand2_1 _2325_ (.Y(_0368_),
    .A(_0288_),
    .B(_0310_));
 sg13g2_nand2_1 _2326_ (.Y(_0369_),
    .A(_0368_),
    .B(_0291_));
 sg13g2_a21oi_1 _2327_ (.A1(_0366_),
    .A2(_0367_),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_nor2b_1 _2328_ (.A(_0322_),
    .B_N(_0247_),
    .Y(_0371_));
 sg13g2_nand3_1 _2329_ (.B(_0371_),
    .C(_0236_),
    .A(_0366_),
    .Y(_0372_));
 sg13g2_nand2_1 _2330_ (.Y(_0373_),
    .A(_0370_),
    .B(_0372_));
 sg13g2_nand2b_1 _2331_ (.Y(_0374_),
    .B(_0373_),
    .A_N(_0365_));
 sg13g2_nand3_1 _2332_ (.B(_0372_),
    .C(_0365_),
    .A(_0370_),
    .Y(_0375_));
 sg13g2_nand2_1 _2333_ (.Y(_0376_),
    .A(_0374_),
    .B(_0375_));
 sg13g2_nand2b_1 _2334_ (.Y(_0377_),
    .B(_0376_),
    .A_N(_0364_));
 sg13g2_nand3_1 _2335_ (.B(_0375_),
    .C(_0364_),
    .A(_0374_),
    .Y(_0378_));
 sg13g2_nand3_1 _2336_ (.B(_0378_),
    .C(_2026_),
    .A(_0377_),
    .Y(_0379_));
 sg13g2_inv_2 _2337_ (.Y(_0380_),
    .A(net47));
 sg13g2_xnor2_1 _2338_ (.Y(_0381_),
    .A(_1659_),
    .B(_2191_));
 sg13g2_o21ai_1 _2339_ (.B1(net41),
    .Y(_0382_),
    .A1(_0380_),
    .A2(_0381_));
 sg13g2_nand2_1 _2340_ (.Y(_0383_),
    .A(_0379_),
    .B(_0382_));
 sg13g2_a21oi_1 _2341_ (.A1(_0331_),
    .A2(net50),
    .Y(_0384_),
    .B1(_2112_));
 sg13g2_nand2_1 _2342_ (.Y(_0385_),
    .A(_0383_),
    .B(_0384_));
 sg13g2_inv_1 _2343_ (.Y(_0386_),
    .A(_0267_));
 sg13g2_o21ai_1 _2344_ (.B1(_1582_),
    .Y(_0387_),
    .A1(net57),
    .A2(_1679_));
 sg13g2_o21ai_1 _2345_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_1582_),
    .A2(_0386_));
 sg13g2_inv_1 _2346_ (.Y(_0389_),
    .A(_0388_));
 sg13g2_xnor2_1 _2347_ (.Y(_0390_),
    .A(_0389_),
    .B(net29));
 sg13g2_a21oi_1 _2348_ (.A1(_0390_),
    .A2(net40),
    .Y(_0391_),
    .B1(net45));
 sg13g2_nand2_1 _2349_ (.Y(_0392_),
    .A(_0385_),
    .B(_0391_));
 sg13g2_a21oi_1 _2350_ (.A1(_0389_),
    .A2(net45),
    .Y(_0393_),
    .B1(net28));
 sg13g2_nand2_1 _2351_ (.Y(_0394_),
    .A(_0392_),
    .B(_0393_));
 sg13g2_nand2_1 _2352_ (.Y(_0395_),
    .A(_0394_),
    .B(_0276_));
 sg13g2_nand2_1 _2353_ (.Y(_0396_),
    .A(_0395_),
    .B(net38));
 sg13g2_a21oi_1 _2354_ (.A1(_0036_),
    .A2(_1764_),
    .Y(_0397_),
    .B1(_0356_));
 sg13g2_buf_8 _2355_ (.A(_0397_),
    .X(_0398_));
 sg13g2_nor3_1 _2356_ (.A(_0178_),
    .B(_0179_),
    .C(_0183_),
    .Y(_0399_));
 sg13g2_buf_1 _2357_ (.A(_0399_),
    .X(_0400_));
 sg13g2_nand3_1 _2358_ (.B(_0398_),
    .C(_0400_),
    .A(_0396_),
    .Y(_0401_));
 sg13g2_nor2b_1 _2359_ (.A(_0361_),
    .B_N(_0401_),
    .Y(_0402_));
 sg13g2_nand2_1 _2360_ (.Y(_0403_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_buf_8 _2361_ (.A(_0403_),
    .X(_0404_));
 sg13g2_buf_8 _2362_ (.A(_0209_),
    .X(_0405_));
 sg13g2_nand2_1 _2363_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_nor2b_2 _2364_ (.A(_0402_),
    .B_N(_0406_),
    .Y(_0407_));
 sg13g2_buf_1 _2365_ (.A(_0199_),
    .X(_0408_));
 sg13g2_nand4_1 _2366_ (.B(_0408_),
    .C(net56),
    .A(_0349_),
    .Y(_0409_),
    .D(net44));
 sg13g2_buf_1 _2367_ (.A(net48),
    .X(_0410_));
 sg13g2_a21oi_1 _2368_ (.A1(_2106_),
    .A2(net47),
    .Y(_0411_),
    .B1(net43));
 sg13g2_xnor2_1 _2369_ (.Y(_0412_),
    .A(_2070_),
    .B(_2086_));
 sg13g2_xor2_1 _2370_ (.B(_2034_),
    .A(_2029_),
    .X(_0413_));
 sg13g2_o21ai_1 _2371_ (.B1(net43),
    .Y(_0414_),
    .A1(_0413_),
    .A2(_0412_));
 sg13g2_a21oi_1 _2372_ (.A1(_0412_),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_xnor2_1 _2373_ (.Y(_0416_),
    .A(_1669_),
    .B(_2068_));
 sg13g2_inv_1 _2374_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_buf_1 _2375_ (.A(net35),
    .X(_0418_));
 sg13g2_a21oi_1 _2376_ (.A1(_0417_),
    .A2(net46),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_o21ai_1 _2377_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0411_),
    .A2(_0415_));
 sg13g2_inv_1 _2378_ (.Y(_0421_),
    .A(_2129_));
 sg13g2_buf_1 _2379_ (.A(_0421_),
    .X(_0422_));
 sg13g2_nand2_1 _2380_ (.Y(_0423_),
    .A(_1580_),
    .B(_0038_));
 sg13g2_a21oi_1 _2381_ (.A1(net57),
    .A2(_0037_),
    .Y(_0424_),
    .B1(_1582_));
 sg13g2_nand2_1 _2382_ (.Y(_0425_),
    .A(net57),
    .B(_0053_));
 sg13g2_o21ai_1 _2383_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net57),
    .A2(_1741_));
 sg13g2_inv_1 _2384_ (.Y(_0427_),
    .A(_0426_));
 sg13g2_a22oi_1 _2385_ (.Y(_0428_),
    .B1(_1582_),
    .B2(_0427_),
    .A2(_0424_),
    .A1(_0423_));
 sg13g2_inv_1 _2386_ (.Y(_0429_),
    .A(_0428_));
 sg13g2_buf_1 _2387_ (.A(_2140_),
    .X(_0430_));
 sg13g2_a21oi_1 _2388_ (.A1(_0422_),
    .A2(_0429_),
    .Y(_0431_),
    .B1(net31));
 sg13g2_o21ai_1 _2389_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0422_),
    .A2(_0429_));
 sg13g2_nand3_1 _2390_ (.B(_2119_),
    .C(_0432_),
    .A(_0420_),
    .Y(_0433_));
 sg13g2_buf_1 _2391_ (.A(net33),
    .X(_0434_));
 sg13g2_a21oi_1 _2392_ (.A1(_0429_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(_2148_));
 sg13g2_nand2_1 _2393_ (.Y(_0436_),
    .A(_0433_),
    .B(_0435_));
 sg13g2_nor2_1 _2394_ (.A(_1764_),
    .B(_0196_),
    .Y(_0437_));
 sg13g2_inv_1 _2395_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nor3_1 _2396_ (.A(_0438_),
    .B(_0185_),
    .C(_0176_),
    .Y(_0439_));
 sg13g2_inv_1 _2397_ (.Y(_0440_),
    .A(_0358_));
 sg13g2_nand2_1 _2398_ (.Y(_0441_),
    .A(_0279_),
    .B(net37));
 sg13g2_nor2_1 _2399_ (.A(_0440_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_a21oi_1 _2400_ (.A1(_0436_),
    .A2(_0439_),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_nand2_1 _2401_ (.Y(_0444_),
    .A(_0409_),
    .B(_0443_));
 sg13g2_nor2b_1 _2402_ (.A(_0205_),
    .B_N(_0204_),
    .Y(_0445_));
 sg13g2_nor2_1 _2403_ (.A(_0188_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_inv_1 _2404_ (.Y(_0447_),
    .A(_0446_));
 sg13g2_nor2_1 _2405_ (.A(_0206_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_nor2_1 _2406_ (.A(_0448_),
    .B(_0404_),
    .Y(_0449_));
 sg13g2_nor2_2 _2407_ (.A(_0444_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_inv_2 _2408_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_nand2_1 _2409_ (.Y(_0452_),
    .A(_0407_),
    .B(_0451_));
 sg13g2_nand4_1 _2410_ (.B(_0199_),
    .C(_0213_),
    .A(_0349_),
    .Y(_0453_),
    .D(net44));
 sg13g2_a21oi_1 _2411_ (.A1(_2034_),
    .A2(_0225_),
    .Y(_0454_),
    .B1(_0217_));
 sg13g2_xor2_1 _2412_ (.B(_0454_),
    .A(_0219_),
    .X(_0455_));
 sg13g2_xnor2_1 _2413_ (.Y(_0456_),
    .A(_0247_),
    .B(_0236_));
 sg13g2_xnor2_1 _2414_ (.Y(_0457_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_xnor2_1 _2415_ (.Y(_0458_),
    .A(net66),
    .B(net20));
 sg13g2_a21o_1 _2416_ (.A2(net47),
    .A1(_0458_),
    .B1(net48),
    .X(_0459_));
 sg13g2_o21ai_1 _2417_ (.B1(_0459_),
    .Y(_0460_),
    .A1(_2027_),
    .A2(_0457_));
 sg13g2_a21oi_1 _2418_ (.A1(_2099_),
    .A2(net46),
    .Y(_0461_),
    .B1(net35));
 sg13g2_nand2_1 _2419_ (.Y(_0462_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_nor2_1 _2420_ (.A(net55),
    .B(_0265_),
    .Y(_0463_));
 sg13g2_a21oi_2 _2421_ (.B1(_0463_),
    .Y(_0464_),
    .A2(_0426_),
    .A1(net55));
 sg13g2_a21oi_1 _2422_ (.A1(_0421_),
    .A2(_0464_),
    .Y(_0465_),
    .B1(_2140_));
 sg13g2_o21ai_1 _2423_ (.B1(_0465_),
    .Y(_0466_),
    .A1(net26),
    .A2(_0464_));
 sg13g2_nand3_1 _2424_ (.B(net34),
    .C(_0466_),
    .A(_0462_),
    .Y(_0467_));
 sg13g2_a21oi_1 _2425_ (.A1(_0464_),
    .A2(net33),
    .Y(_0468_),
    .B1(net24));
 sg13g2_nand2_1 _2426_ (.Y(_0469_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_buf_1 _2427_ (.A(_0276_),
    .X(_0470_));
 sg13g2_nand2_1 _2428_ (.Y(_0471_),
    .A(_0469_),
    .B(net16));
 sg13g2_nor2_1 _2429_ (.A(_0206_),
    .B(_0356_),
    .Y(_0472_));
 sg13g2_a21oi_1 _2430_ (.A1(_1765_),
    .A2(_0017_),
    .Y(_0473_),
    .B1(_0354_));
 sg13g2_nand2_1 _2431_ (.Y(_0474_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_a21oi_1 _2432_ (.A1(_0471_),
    .A2(_0278_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_nor2_1 _2433_ (.A(_0209_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nand2_1 _2434_ (.Y(_0477_),
    .A(_0453_),
    .B(_0476_));
 sg13g2_nand2_1 _2435_ (.Y(_0478_),
    .A(_0406_),
    .B(_0477_));
 sg13g2_nor2_1 _2436_ (.A(_0354_),
    .B(_0351_),
    .Y(_0479_));
 sg13g2_nor2_1 _2437_ (.A(_0479_),
    .B(_0404_),
    .Y(_0480_));
 sg13g2_inv_1 _2438_ (.Y(_0481_),
    .A(_0480_));
 sg13g2_nand2_2 _2439_ (.Y(_0482_),
    .A(_0478_),
    .B(_0481_));
 sg13g2_inv_2 _2440_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_inv_1 _2441_ (.Y(_0484_),
    .A(_0472_));
 sg13g2_nand2_1 _2442_ (.Y(_0485_),
    .A(net49),
    .B(_0052_));
 sg13g2_inv_1 _2443_ (.Y(_0486_),
    .A(_0485_));
 sg13g2_o21ai_1 _2444_ (.B1(_0221_),
    .Y(_0487_),
    .A1(_0219_),
    .A2(_0454_));
 sg13g2_xnor2_1 _2445_ (.Y(_0488_),
    .A(_0218_),
    .B(_0487_));
 sg13g2_nor2b_1 _2446_ (.A(_0250_),
    .B_N(_0249_),
    .Y(_0489_));
 sg13g2_xnor2_1 _2447_ (.Y(_0490_),
    .A(_0488_),
    .B(_0489_));
 sg13g2_inv_1 _2448_ (.Y(_0491_),
    .A(_0246_));
 sg13g2_a21oi_1 _2449_ (.A1(_0236_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(_0243_));
 sg13g2_xnor2_1 _2450_ (.Y(_0493_),
    .A(_0490_),
    .B(_0492_));
 sg13g2_nand2_1 _2451_ (.Y(_0494_),
    .A(_0493_),
    .B(net43));
 sg13g2_a21oi_1 _2452_ (.A1(_0261_),
    .A2(net47),
    .Y(_0495_),
    .B1(_2025_));
 sg13g2_inv_1 _2453_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_nand2_1 _2454_ (.Y(_0497_),
    .A(_0494_),
    .B(_0496_));
 sg13g2_a21oi_1 _2455_ (.A1(_0458_),
    .A2(net50),
    .Y(_0498_),
    .B1(net35));
 sg13g2_nand2_1 _2456_ (.Y(_0499_),
    .A(_0497_),
    .B(_0498_));
 sg13g2_nor2_1 _2457_ (.A(net55),
    .B(_0339_),
    .Y(_0500_));
 sg13g2_a21oi_2 _2458_ (.B1(_0500_),
    .Y(_0501_),
    .A2(_2136_),
    .A1(net55));
 sg13g2_nor2b_1 _2459_ (.A(_2130_),
    .B_N(_0501_),
    .Y(_0502_));
 sg13g2_nor2_1 _2460_ (.A(_0501_),
    .B(_0421_),
    .Y(_0503_));
 sg13g2_nor3_1 _2461_ (.A(_2140_),
    .B(_0502_),
    .C(_0503_),
    .Y(_0504_));
 sg13g2_nor2_1 _2462_ (.A(net39),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_nand2_1 _2463_ (.Y(_0506_),
    .A(_0499_),
    .B(_0505_));
 sg13g2_a21oi_1 _2464_ (.A1(_0501_),
    .A2(net39),
    .Y(_0507_),
    .B1(net28));
 sg13g2_nand2_1 _2465_ (.Y(_0508_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_a21oi_1 _2466_ (.A1(_0508_),
    .A2(net16),
    .Y(_0509_),
    .B1(net49));
 sg13g2_nor3_1 _2467_ (.A(_0484_),
    .B(_0486_),
    .C(_0509_),
    .Y(_0510_));
 sg13g2_nor2_1 _2468_ (.A(_0209_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_nand2_1 _2469_ (.Y(_0512_),
    .A(_0353_),
    .B(_0511_));
 sg13g2_nand3_1 _2470_ (.B(_0404_),
    .C(_0210_),
    .A(_0512_),
    .Y(_0513_));
 sg13g2_a21oi_1 _2471_ (.A1(_0452_),
    .A2(_0483_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nor2_1 _2472_ (.A(_0214_),
    .B(_0404_),
    .Y(_0515_));
 sg13g2_a21oi_1 _2473_ (.A1(_0406_),
    .A2(_0512_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_buf_2 _2474_ (.A(_0516_),
    .X(_0517_));
 sg13g2_nor2_1 _2475_ (.A(_0402_),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_inv_1 _2476_ (.Y(_0519_),
    .A(net56));
 sg13g2_nor2_1 _2477_ (.A(_0519_),
    .B(_0282_),
    .Y(_0520_));
 sg13g2_nor2b_1 _2478_ (.A(_0356_),
    .B_N(_0188_),
    .Y(_0521_));
 sg13g2_nand3_1 _2479_ (.B(net44),
    .C(_0521_),
    .A(_0349_),
    .Y(_0522_));
 sg13g2_nor3_1 _2480_ (.A(_0440_),
    .B(_0486_),
    .C(_0509_),
    .Y(_0523_));
 sg13g2_nor2b_1 _2481_ (.A(_0438_),
    .B_N(_0181_),
    .Y(_0524_));
 sg13g2_nand2_1 _2482_ (.Y(_0525_),
    .A(_0276_),
    .B(_0524_));
 sg13g2_inv_1 _2483_ (.Y(_0526_),
    .A(_0525_));
 sg13g2_inv_1 _2484_ (.Y(_0527_),
    .A(_2126_));
 sg13g2_xnor2_1 _2485_ (.Y(_0528_),
    .A(_0527_),
    .B(net29));
 sg13g2_xnor2_1 _2486_ (.Y(_0529_),
    .A(net64),
    .B(_2066_));
 sg13g2_a21oi_1 _2487_ (.A1(_0529_),
    .A2(_2109_),
    .Y(_0530_),
    .B1(net35));
 sg13g2_xor2_1 _2488_ (.B(_2031_),
    .A(_2030_),
    .X(_0531_));
 sg13g2_nand2b_1 _2489_ (.Y(_0532_),
    .B(_2063_),
    .A_N(_2069_));
 sg13g2_xnor2_1 _2490_ (.Y(_0533_),
    .A(_2067_),
    .B(_0532_));
 sg13g2_xor2_1 _2491_ (.B(_0533_),
    .A(_0531_),
    .X(_0534_));
 sg13g2_a21oi_1 _2492_ (.A1(_0417_),
    .A2(net47),
    .Y(_0535_),
    .B1(net43));
 sg13g2_inv_1 _2493_ (.Y(_0536_),
    .A(_0535_));
 sg13g2_o21ai_1 _2494_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net41),
    .A2(_0534_));
 sg13g2_a22oi_1 _2495_ (.Y(_0538_),
    .B1(_0530_),
    .B2(_0537_),
    .A2(_0528_),
    .A1(net32));
 sg13g2_nand2_1 _2496_ (.Y(_0539_),
    .A(_2126_),
    .B(net33));
 sg13g2_o21ai_1 _2497_ (.B1(_0539_),
    .Y(_0540_),
    .A1(net33),
    .A2(_0538_));
 sg13g2_nand2_1 _2498_ (.Y(_0541_),
    .A(_0540_),
    .B(_2146_));
 sg13g2_a21oi_1 _2499_ (.A1(_0526_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(_0209_));
 sg13g2_nor2b_1 _2500_ (.A(_0523_),
    .B_N(_0542_),
    .Y(_0543_));
 sg13g2_nand2_1 _2501_ (.Y(_0544_),
    .A(_0522_),
    .B(_0543_));
 sg13g2_nor2_1 _2502_ (.A(_0520_),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_nand4_1 _2503_ (.B(_0408_),
    .C(_0359_),
    .A(_0349_),
    .Y(_0546_),
    .D(_0445_));
 sg13g2_nand2_1 _2504_ (.Y(_0547_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_nand2_1 _2505_ (.Y(_0548_),
    .A(_0547_),
    .B(_0406_));
 sg13g2_inv_4 _2506_ (.A(_0404_),
    .Y(_0549_));
 sg13g2_nand2_1 _2507_ (.Y(_0550_),
    .A(_0549_),
    .B(_0184_));
 sg13g2_nand2_1 _2508_ (.Y(_0551_),
    .A(_0548_),
    .B(_0550_));
 sg13g2_nand2_1 _2509_ (.Y(_0552_),
    .A(_0518_),
    .B(_0551_));
 sg13g2_nand2_1 _2510_ (.Y(_0553_),
    .A(_0349_),
    .B(_0359_));
 sg13g2_nor2_1 _2511_ (.A(_0200_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_nand2_1 _2512_ (.Y(_0555_),
    .A(_0360_),
    .B(net23));
 sg13g2_nand2_1 _2513_ (.Y(_0556_),
    .A(_0409_),
    .B(_0546_));
 sg13g2_nor3_1 _2514_ (.A(_0554_),
    .B(_0555_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_nor2b_1 _2515_ (.A(_0557_),
    .B_N(_0406_),
    .Y(_0558_));
 sg13g2_nor2_1 _2516_ (.A(_0477_),
    .B(_0480_),
    .Y(_0559_));
 sg13g2_nor2_1 _2517_ (.A(_0559_),
    .B(_0450_),
    .Y(_0560_));
 sg13g2_o21ai_1 _2518_ (.B1(net23),
    .Y(_0561_),
    .A1(_0484_),
    .A2(_0441_));
 sg13g2_nor2_1 _2519_ (.A(_0283_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_nand3_1 _2520_ (.B(_0398_),
    .C(_0351_),
    .A(_0396_),
    .Y(_0563_));
 sg13g2_a22oi_1 _2521_ (.Y(_0564_),
    .B1(_0562_),
    .B2(_0563_),
    .A2(net27),
    .A1(_0404_));
 sg13g2_buf_8 _2522_ (.A(_0564_),
    .X(_0565_));
 sg13g2_a21oi_1 _2523_ (.A1(_0560_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(_0404_));
 sg13g2_a21oi_1 _2524_ (.A1(_0552_),
    .A2(_0558_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_nor2_1 _2525_ (.A(_0514_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_nand4_1 _2526_ (.B(net17),
    .C(_0213_),
    .A(_0279_),
    .Y(_0569_),
    .D(_0281_));
 sg13g2_nand2_1 _2527_ (.Y(_0570_),
    .A(_0569_),
    .B(_0202_));
 sg13g2_nor2_1 _2528_ (.A(_0570_),
    .B(_0555_),
    .Y(_0571_));
 sg13g2_nand3_1 _2529_ (.B(_0401_),
    .C(_0353_),
    .A(_0571_),
    .Y(_0572_));
 sg13g2_nand2_1 _2530_ (.Y(_0573_),
    .A(_0482_),
    .B(_0572_));
 sg13g2_nand2_1 _2531_ (.Y(_0574_),
    .A(_0573_),
    .B(_0517_));
 sg13g2_nand2_1 _2532_ (.Y(_0575_),
    .A(_0574_),
    .B(_0557_));
 sg13g2_nand2_1 _2533_ (.Y(_0576_),
    .A(_0575_),
    .B(_0549_));
 sg13g2_nand2_1 _2534_ (.Y(_0577_),
    .A(_0576_),
    .B(_0565_));
 sg13g2_nand2_1 _2535_ (.Y(_0578_),
    .A(_0568_),
    .B(_0577_));
 sg13g2_inv_1 _2536_ (.Y(_0579_),
    .A(_0558_));
 sg13g2_nand2_1 _2537_ (.Y(_0580_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_nand3_1 _2538_ (.B(_0577_),
    .C(_0558_),
    .A(_0568_),
    .Y(_0581_));
 sg13g2_nand2_1 _2539_ (.Y(_0582_),
    .A(_0580_),
    .B(_0581_));
 sg13g2_nand2_1 _2540_ (.Y(_0583_),
    .A(_0582_),
    .B(_0407_));
 sg13g2_inv_1 _2541_ (.Y(_0584_),
    .A(_0583_));
 sg13g2_nand3_1 _2542_ (.B(_0577_),
    .C(_0579_),
    .A(_0568_),
    .Y(_0585_));
 sg13g2_buf_2 _2543_ (.A(_0585_),
    .X(_0586_));
 sg13g2_nand3_1 _2544_ (.B(_0549_),
    .C(_0483_),
    .A(_0586_),
    .Y(_0587_));
 sg13g2_nand2_1 _2545_ (.Y(_0588_),
    .A(_0586_),
    .B(_0549_));
 sg13g2_buf_8 _2546_ (.A(_0588_),
    .X(_0589_));
 sg13g2_nand2_1 _2547_ (.Y(_0590_),
    .A(_0589_),
    .B(_0482_));
 sg13g2_inv_1 _2548_ (.Y(_0591_),
    .A(_0590_));
 sg13g2_a21oi_1 _2549_ (.A1(_0584_),
    .A2(_0587_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_xnor2_1 _2550_ (.Y(_0593_),
    .A(_0565_),
    .B(_0589_));
 sg13g2_inv_2 _2551_ (.Y(_0594_),
    .A(_0593_));
 sg13g2_nand2_1 _2552_ (.Y(_0595_),
    .A(_0578_),
    .B(_0558_));
 sg13g2_nand2_1 _2553_ (.Y(_0596_),
    .A(_0595_),
    .B(_0586_));
 sg13g2_buf_8 _2554_ (.A(_0596_),
    .X(_0597_));
 sg13g2_nand2b_1 _2555_ (.Y(_0598_),
    .B(_0597_),
    .A_N(_0517_));
 sg13g2_nand3_1 _2556_ (.B(_0586_),
    .C(_0517_),
    .A(_0595_),
    .Y(_0599_));
 sg13g2_nand2_1 _2557_ (.Y(_0600_),
    .A(_0598_),
    .B(_0599_));
 sg13g2_nand2_1 _2558_ (.Y(_0601_),
    .A(_0594_),
    .B(_0600_));
 sg13g2_nor2_1 _2559_ (.A(_0592_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_inv_1 _2560_ (.Y(_0603_),
    .A(_0589_));
 sg13g2_inv_1 _2561_ (.Y(_0604_),
    .A(_0565_));
 sg13g2_nand2_1 _2562_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_nor2_1 _2563_ (.A(_0517_),
    .B(_0597_),
    .Y(_0606_));
 sg13g2_nor2_1 _2564_ (.A(_0604_),
    .B(_0603_),
    .Y(_0607_));
 sg13g2_a21oi_1 _2565_ (.A1(_0605_),
    .A2(_0606_),
    .Y(_0608_),
    .B1(_0607_));
 sg13g2_nor2b_1 _2566_ (.A(_0602_),
    .B_N(_0608_),
    .Y(_0609_));
 sg13g2_inv_1 _2567_ (.Y(_0610_),
    .A(_0551_));
 sg13g2_nand3_1 _2568_ (.B(_0581_),
    .C(_0610_),
    .A(_0580_),
    .Y(_0611_));
 sg13g2_buf_2 _2569_ (.A(_0611_),
    .X(_0612_));
 sg13g2_nand3_1 _2570_ (.B(_0549_),
    .C(_0450_),
    .A(_0586_),
    .Y(_0613_));
 sg13g2_a21oi_1 _2571_ (.A1(_0586_),
    .A2(_0549_),
    .Y(_0614_),
    .B1(_0450_));
 sg13g2_a21oi_1 _2572_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_inv_1 _2573_ (.Y(_0616_),
    .A(_0615_));
 sg13g2_xnor2_1 _2574_ (.Y(_0617_),
    .A(_0517_),
    .B(_0597_));
 sg13g2_nor2_1 _2575_ (.A(_0593_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_nand2_1 _2576_ (.Y(_0619_),
    .A(_0590_),
    .B(_0587_));
 sg13g2_inv_1 _2577_ (.Y(_0620_),
    .A(_0407_));
 sg13g2_nand3_1 _2578_ (.B(_0581_),
    .C(_0620_),
    .A(_0580_),
    .Y(_0621_));
 sg13g2_nand2_1 _2579_ (.Y(_0622_),
    .A(_0583_),
    .B(_0621_));
 sg13g2_nor2_1 _2580_ (.A(_0619_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_nand3_1 _2581_ (.B(_0618_),
    .C(_0623_),
    .A(_0616_),
    .Y(_0624_));
 sg13g2_nand2_1 _2582_ (.Y(_0625_),
    .A(_0609_),
    .B(_0624_));
 sg13g2_inv_1 _2583_ (.Y(_0626_),
    .A(_0578_));
 sg13g2_nand2_1 _2584_ (.Y(_0627_),
    .A(_0625_),
    .B(_0626_));
 sg13g2_inv_1 _2585_ (.Y(_0628_),
    .A(\dither_threshold[6] ));
 sg13g2_nand2_1 _2586_ (.Y(_0629_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_nand3_1 _2587_ (.B(\dither_threshold[6] ),
    .C(_0626_),
    .A(_0625_),
    .Y(_0630_));
 sg13g2_nand2_1 _2588_ (.Y(_0631_),
    .A(_0629_),
    .B(_0630_));
 sg13g2_inv_1 _2589_ (.Y(_0632_),
    .A(_0631_));
 sg13g2_nand2_1 _2590_ (.Y(_0633_),
    .A(_0589_),
    .B(_0483_));
 sg13g2_nand3_1 _2591_ (.B(_0549_),
    .C(_0482_),
    .A(_0586_),
    .Y(_0634_));
 sg13g2_nand2_1 _2592_ (.Y(_0635_),
    .A(_0633_),
    .B(_0634_));
 sg13g2_nand2_1 _2593_ (.Y(_0636_),
    .A(_0600_),
    .B(_0635_));
 sg13g2_a21oi_1 _2594_ (.A1(_0614_),
    .A2(_0621_),
    .Y(_0637_),
    .B1(_0584_));
 sg13g2_nor2_1 _2595_ (.A(_0636_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nand2_1 _2596_ (.Y(_0639_),
    .A(_0597_),
    .B(_0517_));
 sg13g2_a21oi_1 _2597_ (.A1(_0591_),
    .A2(_0639_),
    .Y(_0640_),
    .B1(_0606_));
 sg13g2_nor2b_1 _2598_ (.A(_0638_),
    .B_N(_0640_),
    .Y(_0641_));
 sg13g2_nor2_1 _2599_ (.A(_0619_),
    .B(_0617_),
    .Y(_0642_));
 sg13g2_nand2_1 _2600_ (.Y(_0643_),
    .A(_0589_),
    .B(_0451_));
 sg13g2_nand2_1 _2601_ (.Y(_0644_),
    .A(_0643_),
    .B(_0613_));
 sg13g2_nor2_1 _2602_ (.A(_0644_),
    .B(_0622_),
    .Y(_0645_));
 sg13g2_nand3_1 _2603_ (.B(_0645_),
    .C(_0612_),
    .A(_0642_),
    .Y(_0646_));
 sg13g2_nand2_1 _2604_ (.Y(_0647_),
    .A(_0641_),
    .B(_0646_));
 sg13g2_nand2_1 _2605_ (.Y(_0648_),
    .A(_0647_),
    .B(_0594_));
 sg13g2_nand3_1 _2606_ (.B(_0646_),
    .C(_0593_),
    .A(_0641_),
    .Y(_0649_));
 sg13g2_nand2_1 _2607_ (.Y(_0650_),
    .A(_0648_),
    .B(_0649_));
 sg13g2_inv_1 _2608_ (.Y(_0651_),
    .A(_1840_));
 sg13g2_nand2_1 _2609_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_));
 sg13g2_nand3_1 _2610_ (.B(_0649_),
    .C(_1840_),
    .A(_0648_),
    .Y(_0653_));
 sg13g2_nand2_1 _2611_ (.Y(_0654_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_nor2_1 _2612_ (.A(_0632_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_nand2_1 _2613_ (.Y(_0656_),
    .A(_0616_),
    .B(_0623_));
 sg13g2_nand2_1 _2614_ (.Y(_0657_),
    .A(_0656_),
    .B(_0592_));
 sg13g2_nand2_1 _2615_ (.Y(_0658_),
    .A(_0657_),
    .B(_0617_));
 sg13g2_nand3_1 _2616_ (.B(_0600_),
    .C(_0592_),
    .A(_0656_),
    .Y(_0659_));
 sg13g2_nand2_1 _2617_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_nand2_1 _2618_ (.Y(_0661_),
    .A(_0660_),
    .B(_1835_));
 sg13g2_nand3_1 _2619_ (.B(_0659_),
    .C(_1841_),
    .A(_0658_),
    .Y(_0662_));
 sg13g2_xnor2_1 _2620_ (.Y(_0663_),
    .A(_0407_),
    .B(_0597_));
 sg13g2_nand2_1 _2621_ (.Y(_0664_),
    .A(_0589_),
    .B(_0450_));
 sg13g2_nand3_1 _2622_ (.B(_0549_),
    .C(_0451_),
    .A(_0586_),
    .Y(_0665_));
 sg13g2_nand2_1 _2623_ (.Y(_0666_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_nand3_1 _2624_ (.B(_0612_),
    .C(_0666_),
    .A(_0663_),
    .Y(_0667_));
 sg13g2_nand2_1 _2625_ (.Y(_0668_),
    .A(_0667_),
    .B(_0637_));
 sg13g2_nand2_1 _2626_ (.Y(_0669_),
    .A(_0668_),
    .B(_0635_));
 sg13g2_nand3_1 _2627_ (.B(_0619_),
    .C(_0637_),
    .A(_0667_),
    .Y(_0670_));
 sg13g2_nand2_1 _2628_ (.Y(_0671_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_nor2b_1 _2629_ (.A(_0671_),
    .B_N(_1805_),
    .Y(_0672_));
 sg13g2_nand3_1 _2630_ (.B(_0662_),
    .C(_0672_),
    .A(_0661_),
    .Y(_0673_));
 sg13g2_nand2_1 _2631_ (.Y(_0674_),
    .A(_0660_),
    .B(_1807_));
 sg13g2_nand2_1 _2632_ (.Y(_0675_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_nor2_1 _2633_ (.A(\dither_threshold[5] ),
    .B(_0650_),
    .Y(_0676_));
 sg13g2_nand2_1 _2634_ (.Y(_0677_),
    .A(_0631_),
    .B(_0676_));
 sg13g2_nand3_1 _2635_ (.B(_0628_),
    .C(_0626_),
    .A(_0625_),
    .Y(_0678_));
 sg13g2_nand2_1 _2636_ (.Y(_0679_),
    .A(_0677_),
    .B(_0678_));
 sg13g2_a21oi_1 _2637_ (.A1(_0655_),
    .A2(_0675_),
    .Y(_0680_),
    .B1(_0679_));
 sg13g2_nand2_1 _2638_ (.Y(_0681_),
    .A(_0582_),
    .B(_0551_));
 sg13g2_nand2_1 _2639_ (.Y(_0682_),
    .A(_0681_),
    .B(_0612_));
 sg13g2_nor2_1 _2640_ (.A(_1799_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_xnor2_1 _2641_ (.Y(_0684_),
    .A(_0663_),
    .B(_0615_));
 sg13g2_inv_1 _2642_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_nand2_1 _2643_ (.Y(_0686_),
    .A(_0685_),
    .B(_1808_));
 sg13g2_xnor2_1 _2644_ (.Y(_0687_),
    .A(_0612_),
    .B(_0666_));
 sg13g2_xnor2_1 _2645_ (.Y(_0688_),
    .A(_0031_),
    .B(_0687_));
 sg13g2_nand2_1 _2646_ (.Y(_0689_),
    .A(_0684_),
    .B(_1809_));
 sg13g2_nand3_1 _2647_ (.B(_0688_),
    .C(_0689_),
    .A(_0686_),
    .Y(_0690_));
 sg13g2_o21ai_1 _2648_ (.B1(_0689_),
    .Y(_0691_),
    .A1(_1801_),
    .A2(_0687_));
 sg13g2_nand2_1 _2649_ (.Y(_0692_),
    .A(_0691_),
    .B(_0686_));
 sg13g2_o21ai_1 _2650_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0683_),
    .A2(_0690_));
 sg13g2_xnor2_1 _2651_ (.Y(_0694_),
    .A(_1827_),
    .B(_0671_));
 sg13g2_nand2_1 _2652_ (.Y(_0695_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_nor2_1 _2653_ (.A(_0694_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_nand3_1 _2654_ (.B(_0693_),
    .C(_0696_),
    .A(_0655_),
    .Y(_0697_));
 sg13g2_nand2_1 _2655_ (.Y(_0698_),
    .A(_0680_),
    .B(_0697_));
 sg13g2_nor2_1 _2656_ (.A(_0695_),
    .B(_0654_),
    .Y(_0699_));
 sg13g2_xnor2_1 _2657_ (.Y(_0700_),
    .A(_1800_),
    .B(_0682_));
 sg13g2_nor3_1 _2658_ (.A(_0690_),
    .B(_0700_),
    .C(_0694_),
    .Y(_0701_));
 sg13g2_nand3_1 _2659_ (.B(_0701_),
    .C(_0631_),
    .A(_0699_),
    .Y(_0702_));
 sg13g2_nand3_1 _2660_ (.B(_0597_),
    .C(_0702_),
    .A(_0698_),
    .Y(_0703_));
 sg13g2_nand2_1 _2661_ (.Y(_0704_),
    .A(_0703_),
    .B(_0603_));
 sg13g2_nand4_1 _2662_ (.B(_0589_),
    .C(_0597_),
    .A(_0698_),
    .Y(_0705_),
    .D(_0702_));
 sg13g2_nand2_1 _2663_ (.Y(net8),
    .A(_0704_),
    .B(_0705_));
 sg13g2_nor2_1 _2664_ (.A(_0044_),
    .B(_2083_),
    .Y(_0706_));
 sg13g2_inv_1 _2665_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_xnor2_1 _2666_ (.Y(_0708_),
    .A(_1986_),
    .B(net22));
 sg13g2_nor2_1 _2667_ (.A(_0043_),
    .B(net22),
    .Y(_0709_));
 sg13g2_inv_1 _2668_ (.Y(_0710_),
    .A(_0709_));
 sg13g2_o21ai_1 _2669_ (.B1(_0710_),
    .Y(_0711_),
    .A1(_0707_),
    .A2(_0708_));
 sg13g2_xnor2_1 _2670_ (.Y(_0712_),
    .A(_1983_),
    .B(net20));
 sg13g2_nand2_1 _2671_ (.Y(_0713_),
    .A(_0240_),
    .B(_0234_));
 sg13g2_nand2_1 _2672_ (.Y(_0714_),
    .A(net19),
    .B(_0041_));
 sg13g2_nand2_1 _2673_ (.Y(_0715_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_nor2_1 _2674_ (.A(_0712_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_nor2_1 _2675_ (.A(_0042_),
    .B(net20),
    .Y(_0717_));
 sg13g2_inv_1 _2676_ (.Y(_0718_),
    .A(_0713_));
 sg13g2_a21oi_1 _2677_ (.A1(_0714_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(_0718_));
 sg13g2_inv_1 _2678_ (.Y(_0720_),
    .A(_0719_));
 sg13g2_a21oi_1 _2679_ (.A1(_0711_),
    .A2(_0716_),
    .Y(_0721_),
    .B1(_0720_));
 sg13g2_nor2_1 _2680_ (.A(_0045_),
    .B(net36),
    .Y(_0722_));
 sg13g2_xnor2_1 _2681_ (.Y(_0723_),
    .A(_1993_),
    .B(net36));
 sg13g2_nor2_1 _2682_ (.A(_1990_),
    .B(_2066_),
    .Y(_0724_));
 sg13g2_nand2_1 _2683_ (.Y(_0725_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_nand2b_1 _2684_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0722_));
 sg13g2_inv_1 _2685_ (.Y(_0727_),
    .A(_0044_));
 sg13g2_xnor2_1 _2686_ (.Y(_0728_),
    .A(_0727_),
    .B(_2083_));
 sg13g2_nor2b_1 _2687_ (.A(_0708_),
    .B_N(_0728_),
    .Y(_0729_));
 sg13g2_nand3_1 _2688_ (.B(_0726_),
    .C(_0729_),
    .A(_0716_),
    .Y(_0730_));
 sg13g2_xnor2_1 _2689_ (.Y(_0731_),
    .A(_0244_),
    .B(net18));
 sg13g2_nor2_1 _2690_ (.A(net61),
    .B(_2002_),
    .Y(_0732_));
 sg13g2_nand2_1 _2691_ (.Y(_0733_),
    .A(net61),
    .B(_2002_));
 sg13g2_inv_1 _2692_ (.Y(_0734_),
    .A(_0733_));
 sg13g2_nor2_1 _2693_ (.A(_0732_),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_nand2_1 _2694_ (.Y(_0736_),
    .A(net63),
    .B(net59));
 sg13g2_xnor2_1 _2695_ (.Y(_0737_),
    .A(net62),
    .B(net58));
 sg13g2_nand2_1 _2696_ (.Y(_0738_),
    .A(net62),
    .B(net58));
 sg13g2_o21ai_1 _2697_ (.B1(_0738_),
    .Y(_0739_),
    .A1(_0736_),
    .A2(_0737_));
 sg13g2_xor2_1 _2698_ (.B(_1978_),
    .A(_1654_),
    .X(_0740_));
 sg13g2_inv_1 _2699_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_xor2_1 _2700_ (.B(net70),
    .A(_1651_),
    .X(_0742_));
 sg13g2_inv_1 _2701_ (.Y(_0743_),
    .A(_0742_));
 sg13g2_nor2_1 _2702_ (.A(_0741_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand2_1 _2703_ (.Y(_0745_),
    .A(net66),
    .B(net70));
 sg13g2_nor2_1 _2704_ (.A(_0745_),
    .B(_0741_),
    .Y(_0746_));
 sg13g2_a221oi_1 _2705_ (.B2(_0744_),
    .C1(_0746_),
    .B1(_0739_),
    .A1(net65),
    .Y(_0747_),
    .A2(_1978_));
 sg13g2_nand2_1 _2706_ (.Y(_0748_),
    .A(net64),
    .B(_1993_));
 sg13g2_xnor2_1 _2707_ (.Y(_0749_),
    .A(net73),
    .B(net69));
 sg13g2_nand2_1 _2708_ (.Y(_0750_),
    .A(net73),
    .B(net69));
 sg13g2_o21ai_1 _2709_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0748_),
    .A2(_0749_));
 sg13g2_buf_1 _2710_ (.A(_0751_),
    .X(_0752_));
 sg13g2_xor2_1 _2711_ (.B(net59),
    .A(net63),
    .X(_0753_));
 sg13g2_inv_1 _2712_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_nor2_1 _2713_ (.A(_0737_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_nand3_1 _2714_ (.B(_0755_),
    .C(_0744_),
    .A(_0752_),
    .Y(_0756_));
 sg13g2_nand2_1 _2715_ (.Y(_0757_),
    .A(_0747_),
    .B(_0756_));
 sg13g2_xnor2_1 _2716_ (.Y(_0758_),
    .A(_0735_),
    .B(_0757_));
 sg13g2_xnor2_1 _2717_ (.Y(_0759_),
    .A(_0731_),
    .B(_0758_));
 sg13g2_a21oi_1 _2718_ (.A1(_0721_),
    .A2(_0730_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_nand3_1 _2719_ (.B(_0721_),
    .C(_0730_),
    .A(_0759_),
    .Y(_0761_));
 sg13g2_nand2_1 _2720_ (.Y(_0762_),
    .A(_0761_),
    .B(net48));
 sg13g2_inv_1 _2721_ (.Y(_0763_),
    .A(_0341_));
 sg13g2_inv_1 _2722_ (.Y(_0764_),
    .A(net50));
 sg13g2_nand2_1 _2723_ (.Y(_0765_),
    .A(_0380_),
    .B(_0764_));
 sg13g2_o21ai_1 _2724_ (.B1(_0257_),
    .Y(_0766_),
    .A1(_0763_),
    .A2(_0765_));
 sg13g2_o21ai_1 _2725_ (.B1(_0766_),
    .Y(_0767_),
    .A1(_0760_),
    .A2(_0762_));
 sg13g2_inv_1 _2726_ (.Y(_0768_),
    .A(net18));
 sg13g2_nor2_1 _2727_ (.A(_0048_),
    .B(_0764_),
    .Y(_0769_));
 sg13g2_a21oi_1 _2728_ (.A1(_0768_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(_2111_));
 sg13g2_nand2_1 _2729_ (.Y(_0771_),
    .A(_0767_),
    .B(_0770_));
 sg13g2_xnor2_1 _2730_ (.Y(_0772_),
    .A(_0421_),
    .B(_0164_));
 sg13g2_a21oi_1 _2731_ (.A1(_0772_),
    .A2(net40),
    .Y(_0773_),
    .B1(net45));
 sg13g2_nand2_1 _2732_ (.Y(_0774_),
    .A(_0771_),
    .B(_0773_));
 sg13g2_a21oi_1 _2733_ (.A1(_0768_),
    .A2(net45),
    .Y(_0775_),
    .B1(net28));
 sg13g2_nand2_1 _2734_ (.Y(_0776_),
    .A(_0774_),
    .B(_0775_));
 sg13g2_nand2_1 _2735_ (.Y(_0777_),
    .A(_0776_),
    .B(_0276_));
 sg13g2_nand2_1 _2736_ (.Y(_0778_),
    .A(_0777_),
    .B(_0197_));
 sg13g2_nand3_1 _2737_ (.B(_0358_),
    .C(net44),
    .A(_0778_),
    .Y(_0779_));
 sg13g2_nand2_1 _2738_ (.Y(_0780_),
    .A(_0779_),
    .B(net23));
 sg13g2_xnor2_1 _2739_ (.Y(_0781_),
    .A(_0754_),
    .B(_0752_));
 sg13g2_xnor2_1 _2740_ (.Y(_0782_),
    .A(_0728_),
    .B(_0726_));
 sg13g2_xnor2_1 _2741_ (.Y(_0783_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_o21ai_1 _2742_ (.B1(_0411_),
    .Y(_0784_),
    .A1(_2139_),
    .A2(_0765_));
 sg13g2_o21ai_1 _2743_ (.B1(_0784_),
    .Y(_0785_),
    .A1(net41),
    .A2(_0783_));
 sg13g2_buf_1 _2744_ (.A(_0764_),
    .X(_0786_));
 sg13g2_nor2_1 _2745_ (.A(_0037_),
    .B(net42),
    .Y(_0787_));
 sg13g2_a21oi_1 _2746_ (.A1(_2089_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(net32));
 sg13g2_nand2_1 _2747_ (.Y(_0789_),
    .A(_0785_),
    .B(_0788_));
 sg13g2_a21oi_1 _2748_ (.A1(net26),
    .A2(_2089_),
    .Y(_0790_),
    .B1(_2140_));
 sg13g2_o21ai_1 _2749_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_2089_),
    .A2(net26));
 sg13g2_nor2b_1 _2750_ (.A(net30),
    .B_N(_0791_),
    .Y(_0792_));
 sg13g2_a221oi_1 _2751_ (.B2(_0792_),
    .C1(net24),
    .B1(_0789_),
    .A1(_2089_),
    .Y(_0793_),
    .A2(net30));
 sg13g2_o21ai_1 _2752_ (.B1(net38),
    .Y(_0794_),
    .A1(_0176_),
    .A2(_0793_));
 sg13g2_nand2_1 _2753_ (.Y(_0795_),
    .A(_0794_),
    .B(_0201_));
 sg13g2_nor2b_1 _2754_ (.A(_0780_),
    .B_N(_0795_),
    .Y(_0796_));
 sg13g2_a21o_1 _2755_ (.A2(_0755_),
    .A1(_0752_),
    .B1(_0739_),
    .X(_0797_));
 sg13g2_nand2_1 _2756_ (.Y(_0798_),
    .A(_0797_),
    .B(_0742_));
 sg13g2_nand2_1 _2757_ (.Y(_0799_),
    .A(_0798_),
    .B(_0745_));
 sg13g2_xnor2_1 _2758_ (.Y(_0800_),
    .A(_0741_),
    .B(_0799_));
 sg13g2_nor2_1 _2759_ (.A(_0708_),
    .B(_0712_),
    .Y(_0801_));
 sg13g2_nand4_1 _2760_ (.B(_0728_),
    .C(_0724_),
    .A(_0801_),
    .Y(_0802_),
    .D(_0723_));
 sg13g2_a21oi_1 _2761_ (.A1(_0728_),
    .A2(_0722_),
    .Y(_0803_),
    .B1(_0706_));
 sg13g2_inv_1 _2762_ (.Y(_0804_),
    .A(_0803_));
 sg13g2_xnor2_1 _2763_ (.Y(_0805_),
    .A(net58),
    .B(net20));
 sg13g2_nand2_1 _2764_ (.Y(_0806_),
    .A(_0805_),
    .B(_0709_));
 sg13g2_inv_1 _2765_ (.Y(_0807_),
    .A(_0717_));
 sg13g2_nand2_1 _2766_ (.Y(_0808_),
    .A(_0806_),
    .B(_0807_));
 sg13g2_a21oi_1 _2767_ (.A1(_0804_),
    .A2(_0801_),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_nand2_1 _2768_ (.Y(_0810_),
    .A(_0802_),
    .B(_0809_));
 sg13g2_nand2b_1 _2769_ (.Y(_0811_),
    .B(_0810_),
    .A_N(_0715_));
 sg13g2_nand3_1 _2770_ (.B(_0809_),
    .C(_0715_),
    .A(_0802_),
    .Y(_0812_));
 sg13g2_nand2_1 _2771_ (.Y(_0813_),
    .A(_0811_),
    .B(_0812_));
 sg13g2_nor2_1 _2772_ (.A(_0800_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_a21oi_1 _2773_ (.A1(_0813_),
    .A2(_0800_),
    .Y(_0815_),
    .B1(net41));
 sg13g2_nand2b_1 _2774_ (.Y(_0816_),
    .B(_0815_),
    .A_N(_0814_));
 sg13g2_inv_1 _2775_ (.Y(_0817_),
    .A(_0270_));
 sg13g2_o21ai_1 _2776_ (.B1(_0495_),
    .Y(_0818_),
    .A1(_0817_),
    .A2(_0765_));
 sg13g2_nand2_1 _2777_ (.Y(_0819_),
    .A(_0816_),
    .B(_0818_));
 sg13g2_nor2_1 _2778_ (.A(_0051_),
    .B(net42),
    .Y(_0820_));
 sg13g2_a21oi_1 _2779_ (.A1(_0240_),
    .A2(_0820_),
    .Y(_0821_),
    .B1(net32));
 sg13g2_nand2_1 _2780_ (.Y(_0822_),
    .A(_0819_),
    .B(_0821_));
 sg13g2_xnor2_1 _2781_ (.Y(_0823_),
    .A(net26),
    .B(_0154_));
 sg13g2_a21oi_1 _2782_ (.A1(_0823_),
    .A2(net32),
    .Y(_0824_),
    .B1(net33));
 sg13g2_nand2_1 _2783_ (.Y(_0825_),
    .A(_0822_),
    .B(_0824_));
 sg13g2_a21oi_1 _2784_ (.A1(_0240_),
    .A2(net30),
    .Y(_0826_),
    .B1(net24));
 sg13g2_nand2_1 _2785_ (.Y(_0827_),
    .A(_0825_),
    .B(_0826_));
 sg13g2_nand2_1 _2786_ (.Y(_0828_),
    .A(_0827_),
    .B(net16));
 sg13g2_nand2_1 _2787_ (.Y(_0829_),
    .A(_0828_),
    .B(net38));
 sg13g2_nand4_1 _2788_ (.B(net17),
    .C(_0213_),
    .A(_0829_),
    .Y(_0830_),
    .D(net37));
 sg13g2_nand2_1 _2789_ (.Y(_0831_),
    .A(_0778_),
    .B(_0352_));
 sg13g2_nor2_2 _2790_ (.A(_0356_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_nand2_1 _2791_ (.Y(_0833_),
    .A(_0832_),
    .B(_0351_));
 sg13g2_inv_1 _2792_ (.Y(_0834_),
    .A(_0732_));
 sg13g2_o21ai_1 _2793_ (.B1(_0834_),
    .Y(_0835_),
    .A1(_0734_),
    .A2(_0757_));
 sg13g2_xnor2_1 _2794_ (.Y(_0836_),
    .A(net60),
    .B(_2004_));
 sg13g2_inv_1 _2795_ (.Y(_0837_),
    .A(_0039_));
 sg13g2_xnor2_1 _2796_ (.Y(_0838_),
    .A(_0837_),
    .B(_0168_));
 sg13g2_xnor2_1 _2797_ (.Y(_0839_),
    .A(_0836_),
    .B(_0838_));
 sg13g2_xnor2_1 _2798_ (.Y(_0840_),
    .A(_0835_),
    .B(_0839_));
 sg13g2_inv_2 _2799_ (.Y(_0841_),
    .A(_0731_));
 sg13g2_nor2_1 _2800_ (.A(_0715_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_nand2_1 _2801_ (.Y(_0843_),
    .A(_0842_),
    .B(_0808_));
 sg13g2_nor2_1 _2802_ (.A(_0242_),
    .B(net18),
    .Y(_0844_));
 sg13g2_a21oi_1 _2803_ (.A1(_0731_),
    .A2(_0718_),
    .Y(_0845_),
    .B1(_0844_));
 sg13g2_nand2_1 _2804_ (.Y(_0846_),
    .A(_0843_),
    .B(_0845_));
 sg13g2_nand2_1 _2805_ (.Y(_0847_),
    .A(_0726_),
    .B(_0728_));
 sg13g2_nand2_1 _2806_ (.Y(_0848_),
    .A(_0847_),
    .B(_0707_));
 sg13g2_nand3_1 _2807_ (.B(_0848_),
    .C(_0801_),
    .A(_0842_),
    .Y(_0849_));
 sg13g2_nor2b_1 _2808_ (.A(_0846_),
    .B_N(_0849_),
    .Y(_0850_));
 sg13g2_nor2_1 _2809_ (.A(_0840_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_nand2_1 _2810_ (.Y(_0852_),
    .A(_0850_),
    .B(_0840_));
 sg13g2_nand2_1 _2811_ (.Y(_0853_),
    .A(_0852_),
    .B(net43));
 sg13g2_a21oi_1 _2812_ (.A1(_0380_),
    .A2(_0389_),
    .Y(_0854_),
    .B1(_0332_));
 sg13g2_nor2_1 _2813_ (.A(net50),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_o21ai_1 _2814_ (.B1(_0855_),
    .Y(_0856_),
    .A1(_0851_),
    .A2(_0853_));
 sg13g2_inv_1 _2815_ (.Y(_0857_),
    .A(_0168_));
 sg13g2_nor2_1 _2816_ (.A(_0026_),
    .B(_0786_),
    .Y(_0858_));
 sg13g2_a21oi_1 _2817_ (.A1(_0857_),
    .A2(_0858_),
    .Y(_0859_),
    .B1(net35));
 sg13g2_nand2_1 _2818_ (.Y(_0860_),
    .A(_0856_),
    .B(_0859_));
 sg13g2_xnor2_1 _2819_ (.Y(_0861_),
    .A(_0421_),
    .B(_0168_));
 sg13g2_a21oi_1 _2820_ (.A1(_0861_),
    .A2(_2113_),
    .Y(_0862_),
    .B1(net39));
 sg13g2_nand2_1 _2821_ (.Y(_0863_),
    .A(_0860_),
    .B(_0862_));
 sg13g2_a21oi_1 _2822_ (.A1(_0857_),
    .A2(_2118_),
    .Y(_0864_),
    .B1(net28));
 sg13g2_nand2_1 _2823_ (.Y(_0865_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_nand2_1 _2824_ (.Y(_0866_),
    .A(_0865_),
    .B(_0470_));
 sg13g2_nand2_1 _2825_ (.Y(_0867_),
    .A(_0866_),
    .B(_0278_));
 sg13g2_nand2_1 _2826_ (.Y(_0868_),
    .A(_0867_),
    .B(_0398_));
 sg13g2_buf_8 _2827_ (.A(_0868_),
    .X(_0869_));
 sg13g2_inv_8 _2828_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_nand2_1 _2829_ (.Y(_0871_),
    .A(_0870_),
    .B(net56));
 sg13g2_nand4_1 _2830_ (.B(_0830_),
    .C(_0833_),
    .A(_0796_),
    .Y(_0872_),
    .D(_0871_));
 sg13g2_nand2_1 _2831_ (.Y(_0873_),
    .A(_0869_),
    .B(net27));
 sg13g2_nand2_1 _2832_ (.Y(_0874_),
    .A(_0832_),
    .B(net56));
 sg13g2_inv_1 _2833_ (.Y(_0875_),
    .A(_0874_));
 sg13g2_nor2_1 _2834_ (.A(_0446_),
    .B(_0869_),
    .Y(_0876_));
 sg13g2_nand3_1 _2835_ (.B(net37),
    .C(_0358_),
    .A(_0829_),
    .Y(_0877_));
 sg13g2_xor2_1 _2836_ (.B(_0749_),
    .A(_0748_),
    .X(_0878_));
 sg13g2_xor2_1 _2837_ (.B(_0723_),
    .A(_0724_),
    .X(_0879_));
 sg13g2_xor2_1 _2838_ (.B(_0879_),
    .A(_0878_),
    .X(_0880_));
 sg13g2_o21ai_1 _2839_ (.B1(_0535_),
    .Y(_0881_),
    .A1(_0428_),
    .A2(_0765_));
 sg13g2_o21ai_1 _2840_ (.B1(_0881_),
    .Y(_0882_),
    .A1(net41),
    .A2(_0880_));
 sg13g2_inv_1 _2841_ (.Y(_0883_),
    .A(net36));
 sg13g2_nor2_1 _2842_ (.A(_0038_),
    .B(net42),
    .Y(_0884_));
 sg13g2_a21oi_1 _2843_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(net32));
 sg13g2_nand2_1 _2844_ (.Y(_0886_),
    .A(_0882_),
    .B(_0885_));
 sg13g2_a21oi_1 _2845_ (.A1(net25),
    .A2(net36),
    .Y(_0887_),
    .B1(net31));
 sg13g2_o21ai_1 _2846_ (.B1(_0887_),
    .Y(_0888_),
    .A1(net36),
    .A2(net25));
 sg13g2_nand3_1 _2847_ (.B(net34),
    .C(_0888_),
    .A(_0886_),
    .Y(_0889_));
 sg13g2_a21oi_1 _2848_ (.A1(_0883_),
    .A2(net30),
    .Y(_0890_),
    .B1(net24));
 sg13g2_nand2_1 _2849_ (.Y(_0891_),
    .A(_0889_),
    .B(_0890_));
 sg13g2_a21oi_1 _2850_ (.A1(_0439_),
    .A2(_0891_),
    .Y(_0892_),
    .B1(_0405_));
 sg13g2_nand2_1 _2851_ (.Y(_0893_),
    .A(_0877_),
    .B(_0892_));
 sg13g2_nor3_1 _2852_ (.A(_0875_),
    .B(_0876_),
    .C(_0893_),
    .Y(_0894_));
 sg13g2_inv_1 _2853_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_nand3_1 _2854_ (.B(_0873_),
    .C(_0895_),
    .A(_0872_),
    .Y(_0896_));
 sg13g2_nand2_1 _2855_ (.Y(_0897_),
    .A(net23),
    .B(_0479_));
 sg13g2_nand2_1 _2856_ (.Y(_0898_),
    .A(_0832_),
    .B(_0213_));
 sg13g2_nand2_1 _2857_ (.Y(_0899_),
    .A(_0464_),
    .B(_0380_));
 sg13g2_nand2_1 _2858_ (.Y(_0900_),
    .A(_0752_),
    .B(_0753_));
 sg13g2_nand2_1 _2859_ (.Y(_0901_),
    .A(_0900_),
    .B(_0736_));
 sg13g2_xnor2_1 _2860_ (.Y(_0902_),
    .A(_0737_),
    .B(_0901_));
 sg13g2_xnor2_1 _2861_ (.Y(_0903_),
    .A(_0708_),
    .B(_0848_));
 sg13g2_xnor2_1 _2862_ (.Y(_0904_),
    .A(_0902_),
    .B(_0903_));
 sg13g2_a22oi_1 _2863_ (.Y(_0905_),
    .B1(_0410_),
    .B2(_0904_),
    .A2(_0899_),
    .A1(_2102_));
 sg13g2_o21ai_1 _2864_ (.B1(net46),
    .Y(_0906_),
    .A1(_0023_),
    .A2(net22));
 sg13g2_o21ai_1 _2865_ (.B1(_0906_),
    .Y(_0907_),
    .A1(net46),
    .A2(_0905_));
 sg13g2_nand2_1 _2866_ (.Y(_0908_),
    .A(_0907_),
    .B(_0430_));
 sg13g2_a21oi_1 _2867_ (.A1(_2131_),
    .A2(net22),
    .Y(_0909_),
    .B1(net31));
 sg13g2_o21ai_1 _2868_ (.B1(_0909_),
    .Y(_0910_),
    .A1(net22),
    .A2(_2131_));
 sg13g2_nand3_1 _2869_ (.B(net34),
    .C(_0910_),
    .A(_0908_),
    .Y(_0911_));
 sg13g2_a21oi_1 _2870_ (.A1(_0233_),
    .A2(_0434_),
    .Y(_0912_),
    .B1(net24));
 sg13g2_a21oi_1 _2871_ (.A1(_0911_),
    .A2(_0912_),
    .Y(_0913_),
    .B1(_0176_));
 sg13g2_inv_1 _2872_ (.Y(_0914_),
    .A(_0474_));
 sg13g2_o21ai_1 _2873_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net49),
    .A2(_0913_));
 sg13g2_nand2_1 _2874_ (.Y(_0916_),
    .A(_0898_),
    .B(_0915_));
 sg13g2_a21oi_2 _2875_ (.B1(_0916_),
    .Y(_0917_),
    .A2(_0897_),
    .A1(_0870_));
 sg13g2_xnor2_1 _2876_ (.Y(_0918_),
    .A(_0743_),
    .B(_0797_));
 sg13g2_inv_1 _2877_ (.Y(_0919_),
    .A(_0708_));
 sg13g2_a21oi_1 _2878_ (.A1(_0848_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(_0709_));
 sg13g2_xnor2_1 _2879_ (.Y(_0921_),
    .A(_0712_),
    .B(_0920_));
 sg13g2_xnor2_1 _2880_ (.Y(_0922_),
    .A(_0918_),
    .B(_0921_));
 sg13g2_a21oi_1 _2881_ (.A1(_0380_),
    .A2(_0501_),
    .Y(_0923_),
    .B1(_0459_));
 sg13g2_nor2_1 _2882_ (.A(net50),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_o21ai_1 _2883_ (.B1(_0924_),
    .Y(_0925_),
    .A1(_2027_),
    .A2(_0922_));
 sg13g2_nor2_1 _2884_ (.A(_0053_),
    .B(net42),
    .Y(_0926_));
 sg13g2_a21oi_1 _2885_ (.A1(_0245_),
    .A2(_0926_),
    .Y(_0927_),
    .B1(_2113_));
 sg13g2_nand2_1 _2886_ (.Y(_0928_),
    .A(_0925_),
    .B(_0927_));
 sg13g2_xor2_1 _2887_ (.B(net29),
    .A(_0145_),
    .X(_0929_));
 sg13g2_a21oi_1 _2888_ (.A1(_0929_),
    .A2(_0418_),
    .Y(_0930_),
    .B1(_2118_));
 sg13g2_nand2_1 _2889_ (.Y(_0931_),
    .A(_0928_),
    .B(_0930_));
 sg13g2_a21oi_1 _2890_ (.A1(_0245_),
    .A2(_2144_),
    .Y(_0932_),
    .B1(net24));
 sg13g2_nand2_1 _2891_ (.Y(_0933_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_a21oi_1 _2892_ (.A1(_0933_),
    .A2(_0470_),
    .Y(_0934_),
    .B1(net49));
 sg13g2_nor3_1 _2893_ (.A(_0484_),
    .B(_0486_),
    .C(_0934_),
    .Y(_0935_));
 sg13g2_nor2_1 _2894_ (.A(net27),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_nand2_1 _2895_ (.Y(_0937_),
    .A(_0833_),
    .B(_0936_));
 sg13g2_nand3_1 _2896_ (.B(net23),
    .C(_0869_),
    .A(_0937_),
    .Y(_0938_));
 sg13g2_a21oi_1 _2897_ (.A1(_0896_),
    .A2(_0917_),
    .Y(_0939_),
    .B1(_0938_));
 sg13g2_nor2_1 _2898_ (.A(_0214_),
    .B(_0869_),
    .Y(_0940_));
 sg13g2_nand2_1 _2899_ (.Y(_0941_),
    .A(_0937_),
    .B(_0873_));
 sg13g2_nand2b_1 _2900_ (.Y(_0942_),
    .B(_0941_),
    .A_N(_0940_));
 sg13g2_inv_2 _2901_ (.Y(_0943_),
    .A(_0942_));
 sg13g2_inv_1 _2902_ (.Y(_0944_),
    .A(_0871_));
 sg13g2_inv_1 _2903_ (.Y(_0945_),
    .A(_0796_));
 sg13g2_nand2_1 _2904_ (.Y(_0946_),
    .A(_0830_),
    .B(_0833_));
 sg13g2_nor3_1 _2905_ (.A(_0944_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0947_));
 sg13g2_nor2_1 _2906_ (.A(_0943_),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_inv_1 _2907_ (.Y(_0949_),
    .A(_0184_));
 sg13g2_inv_1 _2908_ (.Y(_0950_),
    .A(_2066_));
 sg13g2_inv_1 _2909_ (.Y(_0951_),
    .A(_1993_));
 sg13g2_xnor2_1 _2910_ (.Y(_0952_),
    .A(net64),
    .B(_1989_));
 sg13g2_xnor2_1 _2911_ (.Y(_0953_),
    .A(_0951_),
    .B(_0952_));
 sg13g2_a21oi_1 _2912_ (.A1(_0953_),
    .A2(_0950_),
    .Y(_0954_),
    .B1(net41));
 sg13g2_o21ai_1 _2913_ (.B1(_0954_),
    .Y(_0955_),
    .A1(_0950_),
    .A2(_0953_));
 sg13g2_nand4_1 _2914_ (.B(net42),
    .C(_0380_),
    .A(_0955_),
    .Y(_0956_),
    .D(_0527_));
 sg13g2_a21oi_1 _2915_ (.A1(_0529_),
    .A2(net47),
    .Y(_0957_),
    .B1(_0410_));
 sg13g2_inv_1 _2916_ (.Y(_0958_),
    .A(_0957_));
 sg13g2_a21oi_1 _2917_ (.A1(_0955_),
    .A2(_0958_),
    .Y(_0959_),
    .B1(net32));
 sg13g2_nand3_1 _2918_ (.B(_1850_),
    .C(net46),
    .A(_0950_),
    .Y(_0960_));
 sg13g2_nand3_1 _2919_ (.B(_0959_),
    .C(_0960_),
    .A(_0956_),
    .Y(_0961_));
 sg13g2_a21oi_1 _2920_ (.A1(net26),
    .A2(_0950_),
    .Y(_0962_),
    .B1(_0430_));
 sg13g2_o21ai_1 _2921_ (.B1(_0962_),
    .Y(_0963_),
    .A1(_0950_),
    .A2(net26));
 sg13g2_nand3_1 _2922_ (.B(net34),
    .C(_0963_),
    .A(_0961_),
    .Y(_0964_));
 sg13g2_nand2_1 _2923_ (.Y(_0965_),
    .A(_0950_),
    .B(net30));
 sg13g2_nand3_1 _2924_ (.B(_2146_),
    .C(_0965_),
    .A(_0964_),
    .Y(_0966_));
 sg13g2_nand2_1 _2925_ (.Y(_0967_),
    .A(_0526_),
    .B(_0966_));
 sg13g2_o21ai_1 _2926_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_0949_),
    .A2(_0869_));
 sg13g2_nand4_1 _2927_ (.B(net17),
    .C(net56),
    .A(_0829_),
    .Y(_0969_),
    .D(net37));
 sg13g2_nand2_1 _2928_ (.Y(_0970_),
    .A(_0832_),
    .B(_0188_));
 sg13g2_nand2_1 _2929_ (.Y(_0971_),
    .A(_0969_),
    .B(_0970_));
 sg13g2_nor2_1 _2930_ (.A(_0968_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_nor3_1 _2931_ (.A(_0440_),
    .B(_0486_),
    .C(_0934_),
    .Y(_0973_));
 sg13g2_nand2b_1 _2932_ (.Y(_0974_),
    .B(_0898_),
    .A_N(_0973_));
 sg13g2_nor2b_1 _2933_ (.A(_0974_),
    .B_N(_0833_),
    .Y(_0975_));
 sg13g2_nand2_1 _2934_ (.Y(_0976_),
    .A(_0870_),
    .B(net27));
 sg13g2_nand3_1 _2935_ (.B(_0975_),
    .C(_0976_),
    .A(_0972_),
    .Y(_0977_));
 sg13g2_nand2_1 _2936_ (.Y(_0978_),
    .A(_0948_),
    .B(_0977_));
 sg13g2_inv_1 _2937_ (.Y(_0979_),
    .A(_0873_));
 sg13g2_inv_1 _2938_ (.Y(_0980_),
    .A(_0780_));
 sg13g2_nand2_1 _2939_ (.Y(_0981_),
    .A(_0446_),
    .B(_0185_));
 sg13g2_nand2_1 _2940_ (.Y(_0982_),
    .A(_0832_),
    .B(_0981_));
 sg13g2_nand3_1 _2941_ (.B(_0982_),
    .C(_0874_),
    .A(_0980_),
    .Y(_0983_));
 sg13g2_inv_1 _2942_ (.Y(_0984_),
    .A(_0983_));
 sg13g2_nor2_2 _2943_ (.A(_0979_),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_nor2_1 _2944_ (.A(_0917_),
    .B(_0894_),
    .Y(_0986_));
 sg13g2_nor2_1 _2945_ (.A(_0213_),
    .B(_0188_),
    .Y(_0987_));
 sg13g2_nand3_1 _2946_ (.B(_0180_),
    .C(_0949_),
    .A(_0987_),
    .Y(_0988_));
 sg13g2_nand4_1 _2947_ (.B(net17),
    .C(net37),
    .A(_0829_),
    .Y(_0989_),
    .D(_0988_));
 sg13g2_nand2_1 _2948_ (.Y(_0990_),
    .A(_0870_),
    .B(_0351_));
 sg13g2_nand4_1 _2949_ (.B(_0989_),
    .C(_0990_),
    .A(_0969_),
    .Y(_0991_),
    .D(net23));
 sg13g2_a21oi_1 _2950_ (.A1(_0986_),
    .A2(_0991_),
    .Y(_0992_),
    .B1(_0869_));
 sg13g2_a21oi_1 _2951_ (.A1(_0978_),
    .A2(_0985_),
    .Y(_0993_),
    .B1(_0992_));
 sg13g2_nor2_1 _2952_ (.A(_0939_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_inv_1 _2953_ (.Y(_0995_),
    .A(_0917_));
 sg13g2_nand2_1 _2954_ (.Y(_0996_),
    .A(_0872_),
    .B(_0995_));
 sg13g2_nand2_1 _2955_ (.Y(_0997_),
    .A(_0996_),
    .B(_0943_));
 sg13g2_nand2_1 _2956_ (.Y(_0998_),
    .A(_0997_),
    .B(_0984_));
 sg13g2_nand2_1 _2957_ (.Y(_0999_),
    .A(_0998_),
    .B(_0870_));
 sg13g2_nand2_1 _2958_ (.Y(_1000_),
    .A(_0991_),
    .B(_0873_));
 sg13g2_inv_1 _2959_ (.Y(_1001_),
    .A(_1000_));
 sg13g2_nand2_1 _2960_ (.Y(_1002_),
    .A(_0999_),
    .B(_1001_));
 sg13g2_inv_1 _2961_ (.Y(_1003_),
    .A(_0985_));
 sg13g2_nand3_1 _2962_ (.B(_1002_),
    .C(_1003_),
    .A(_0994_),
    .Y(_1004_));
 sg13g2_buf_2 _2963_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nand2_2 _2964_ (.Y(_1006_),
    .A(_1005_),
    .B(_0870_));
 sg13g2_nor2_1 _2965_ (.A(_0979_),
    .B(_0894_),
    .Y(_1007_));
 sg13g2_nand2_1 _2966_ (.Y(_1008_),
    .A(_1006_),
    .B(_1007_));
 sg13g2_inv_1 _2967_ (.Y(_1009_),
    .A(_1007_));
 sg13g2_nand3_1 _2968_ (.B(_0870_),
    .C(_1009_),
    .A(_1005_),
    .Y(_1010_));
 sg13g2_nand2_1 _2969_ (.Y(_1011_),
    .A(_1008_),
    .B(_1010_));
 sg13g2_nand2_1 _2970_ (.Y(_1012_),
    .A(_0994_),
    .B(_1002_));
 sg13g2_nand2_1 _2971_ (.Y(_1013_),
    .A(_1012_),
    .B(_1003_));
 sg13g2_nand3_1 _2972_ (.B(_1002_),
    .C(_0985_),
    .A(_0994_),
    .Y(_1014_));
 sg13g2_nand2_1 _2973_ (.Y(_1015_),
    .A(_1013_),
    .B(_1014_));
 sg13g2_nor2_1 _2974_ (.A(_0979_),
    .B(_0947_),
    .Y(_1016_));
 sg13g2_nand2_1 _2975_ (.Y(_1017_),
    .A(_1015_),
    .B(_1016_));
 sg13g2_inv_1 _2976_ (.Y(_1018_),
    .A(_1016_));
 sg13g2_nand3_1 _2977_ (.B(_1014_),
    .C(_1018_),
    .A(_1013_),
    .Y(_1019_));
 sg13g2_nand2_1 _2978_ (.Y(_1020_),
    .A(_1017_),
    .B(_1019_));
 sg13g2_nor2_1 _2979_ (.A(_1011_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_inv_1 _2980_ (.Y(_1022_),
    .A(_0977_));
 sg13g2_nand3_1 _2981_ (.B(_1014_),
    .C(_1022_),
    .A(_1013_),
    .Y(_1023_));
 sg13g2_buf_2 _2982_ (.A(_1023_),
    .X(_1024_));
 sg13g2_nand2_1 _2983_ (.Y(_1025_),
    .A(_1021_),
    .B(_1024_));
 sg13g2_inv_1 _2984_ (.Y(_1026_),
    .A(_1008_));
 sg13g2_nand2_1 _2985_ (.Y(_1027_),
    .A(_1012_),
    .B(_0985_));
 sg13g2_nand2_1 _2986_ (.Y(_1028_),
    .A(_1027_),
    .B(_1005_));
 sg13g2_buf_2 _2987_ (.A(_1028_),
    .X(_1029_));
 sg13g2_nor2_1 _2988_ (.A(_1018_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_a21oi_1 _2989_ (.A1(_1026_),
    .A2(_1019_),
    .Y(_1031_),
    .B1(_1030_));
 sg13g2_nand2_1 _2990_ (.Y(_1032_),
    .A(_1025_),
    .B(_1031_));
 sg13g2_nand2_1 _2991_ (.Y(_1033_),
    .A(_1006_),
    .B(_0995_));
 sg13g2_nand3_1 _2992_ (.B(_0870_),
    .C(_0917_),
    .A(_1005_),
    .Y(_1034_));
 sg13g2_nand2_1 _2993_ (.Y(_1035_),
    .A(_1033_),
    .B(_1034_));
 sg13g2_inv_1 _2994_ (.Y(_1036_),
    .A(_1035_));
 sg13g2_nand2_1 _2995_ (.Y(_1037_),
    .A(_1032_),
    .B(_1036_));
 sg13g2_nand3_1 _2996_ (.B(_1031_),
    .C(_1035_),
    .A(_1025_),
    .Y(_1038_));
 sg13g2_nand2_1 _2997_ (.Y(_1039_),
    .A(_1037_),
    .B(_1038_));
 sg13g2_xnor2_1 _2998_ (.Y(_1040_),
    .A(_1827_),
    .B(_1039_));
 sg13g2_a21oi_1 _2999_ (.A1(_1024_),
    .A2(_1010_),
    .Y(_1041_),
    .B1(_1026_));
 sg13g2_inv_1 _3000_ (.Y(_1042_),
    .A(_1041_));
 sg13g2_nor2_1 _3001_ (.A(_1035_),
    .B(_1020_),
    .Y(_1043_));
 sg13g2_nand2_1 _3002_ (.Y(_1044_),
    .A(_1042_),
    .B(_1043_));
 sg13g2_inv_1 _3003_ (.Y(_1045_),
    .A(_1033_));
 sg13g2_a21oi_1 _3004_ (.A1(_1030_),
    .A2(_1034_),
    .Y(_1046_),
    .B1(_1045_));
 sg13g2_nand2_1 _3005_ (.Y(_1047_),
    .A(_1044_),
    .B(_1046_));
 sg13g2_nor2_1 _3006_ (.A(_0943_),
    .B(_1029_),
    .Y(_1048_));
 sg13g2_nand2_1 _3007_ (.Y(_1049_),
    .A(_1029_),
    .B(_0943_));
 sg13g2_nor2b_1 _3008_ (.A(_1048_),
    .B_N(_1049_),
    .Y(_1050_));
 sg13g2_nand2_1 _3009_ (.Y(_1051_),
    .A(_1047_),
    .B(_1050_));
 sg13g2_nand2b_1 _3010_ (.Y(_1052_),
    .B(_1049_),
    .A_N(_1048_));
 sg13g2_nand3_1 _3011_ (.B(_1052_),
    .C(_1046_),
    .A(_1044_),
    .Y(_1053_));
 sg13g2_buf_1 _3012_ (.A(_1053_),
    .X(_1054_));
 sg13g2_nand2_1 _3013_ (.Y(_1055_),
    .A(_1051_),
    .B(_1054_));
 sg13g2_nand2_1 _3014_ (.Y(_1056_),
    .A(_1055_),
    .B(_1841_));
 sg13g2_nand3_1 _3015_ (.B(_1054_),
    .C(_1835_),
    .A(_1051_),
    .Y(_1057_));
 sg13g2_nand2_1 _3016_ (.Y(_1058_),
    .A(_1056_),
    .B(_1057_));
 sg13g2_nor2_1 _3017_ (.A(_1040_),
    .B(_1058_),
    .Y(_1059_));
 sg13g2_xor2_1 _3018_ (.B(_1011_),
    .A(_1024_),
    .X(_1060_));
 sg13g2_nand2_1 _3019_ (.Y(_1061_),
    .A(_1029_),
    .B(_0977_));
 sg13g2_nand2_1 _3020_ (.Y(_1062_),
    .A(_1015_),
    .B(_1022_));
 sg13g2_nand3_1 _3021_ (.B(_1062_),
    .C(_1800_),
    .A(_1061_),
    .Y(_1063_));
 sg13g2_nand2_1 _3022_ (.Y(_1064_),
    .A(_1063_),
    .B(_0031_));
 sg13g2_nand3_1 _3023_ (.B(_1064_),
    .C(_1802_),
    .A(_1060_),
    .Y(_1065_));
 sg13g2_nand2_1 _3024_ (.Y(_1066_),
    .A(_1063_),
    .B(_1821_));
 sg13g2_nand2b_1 _3025_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1060_));
 sg13g2_nand2_1 _3026_ (.Y(_1068_),
    .A(_1065_),
    .B(_1067_));
 sg13g2_nand2_1 _3027_ (.Y(_1069_),
    .A(_1068_),
    .B(_1809_));
 sg13g2_xnor2_1 _3028_ (.Y(_1070_),
    .A(_1020_),
    .B(_1041_));
 sg13g2_nand2_1 _3029_ (.Y(_1071_),
    .A(_1069_),
    .B(_1070_));
 sg13g2_nand3_1 _3030_ (.B(_1067_),
    .C(_1808_),
    .A(_1065_),
    .Y(_1072_));
 sg13g2_nand2_1 _3031_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_nand2_1 _3032_ (.Y(_1074_),
    .A(_1059_),
    .B(_1073_));
 sg13g2_nand2_1 _3033_ (.Y(_1075_),
    .A(_1055_),
    .B(_1835_));
 sg13g2_nand3_1 _3034_ (.B(_1054_),
    .C(_1841_),
    .A(_1051_),
    .Y(_1076_));
 sg13g2_nand2_1 _3035_ (.Y(_1077_),
    .A(_1075_),
    .B(_1076_));
 sg13g2_a21oi_1 _3036_ (.A1(_1037_),
    .A2(_1038_),
    .Y(_1078_),
    .B1(_0032_));
 sg13g2_a21oi_1 _3037_ (.A1(_1051_),
    .A2(_1054_),
    .Y(_1079_),
    .B1(_1807_));
 sg13g2_a21oi_1 _3038_ (.A1(_1077_),
    .A2(_1078_),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_nand2_1 _3039_ (.Y(_1081_),
    .A(_1074_),
    .B(_1080_));
 sg13g2_nor3_1 _3040_ (.A(_1052_),
    .B(_1035_),
    .C(_1031_),
    .Y(_1082_));
 sg13g2_a21oi_1 _3041_ (.A1(_1045_),
    .A2(_1049_),
    .Y(_1083_),
    .B1(_1048_));
 sg13g2_nor2b_1 _3042_ (.A(_1082_),
    .B_N(_1083_),
    .Y(_1084_));
 sg13g2_nand4_1 _3043_ (.B(_1050_),
    .C(_1024_),
    .A(_1021_),
    .Y(_1085_),
    .D(_1036_));
 sg13g2_nand2_1 _3044_ (.Y(_1086_),
    .A(_1084_),
    .B(_1085_));
 sg13g2_xnor2_1 _3045_ (.Y(_1087_),
    .A(_1000_),
    .B(_1006_));
 sg13g2_nand2_1 _3046_ (.Y(_1088_),
    .A(_1086_),
    .B(_1087_));
 sg13g2_inv_2 _3047_ (.Y(_1089_),
    .A(_1087_));
 sg13g2_nand3_1 _3048_ (.B(_1089_),
    .C(_1085_),
    .A(_1084_),
    .Y(_1090_));
 sg13g2_nand2_1 _3049_ (.Y(_1091_),
    .A(_1088_),
    .B(_1090_));
 sg13g2_nand2_1 _3050_ (.Y(_1092_),
    .A(_1091_),
    .B(_0651_));
 sg13g2_nand3_1 _3051_ (.B(_1090_),
    .C(_1840_),
    .A(_1088_),
    .Y(_1093_));
 sg13g2_nand2_1 _3052_ (.Y(_1094_),
    .A(_1092_),
    .B(_1093_));
 sg13g2_nor3_1 _3053_ (.A(_1089_),
    .B(_1052_),
    .C(_1046_),
    .Y(_1095_));
 sg13g2_nand2_1 _3054_ (.Y(_1096_),
    .A(_1006_),
    .B(_1001_));
 sg13g2_inv_1 _3055_ (.Y(_1097_),
    .A(_1096_));
 sg13g2_a21oi_1 _3056_ (.A1(_1087_),
    .A2(_1048_),
    .Y(_1098_),
    .B1(_1097_));
 sg13g2_nor2b_1 _3057_ (.A(_1095_),
    .B_N(_1098_),
    .Y(_1099_));
 sg13g2_nand4_1 _3058_ (.B(_1043_),
    .C(_1050_),
    .A(_1042_),
    .Y(_1100_),
    .D(_1087_));
 sg13g2_nand2_1 _3059_ (.Y(_1101_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_inv_1 _3060_ (.Y(_1102_),
    .A(_1012_));
 sg13g2_nand2_1 _3061_ (.Y(_1103_),
    .A(_1101_),
    .B(_1102_));
 sg13g2_xnor2_1 _3062_ (.Y(_1104_),
    .A(_1846_),
    .B(_1103_));
 sg13g2_nor2b_1 _3063_ (.A(_1094_),
    .B_N(_1104_),
    .Y(_1105_));
 sg13g2_nand2_1 _3064_ (.Y(_1106_),
    .A(_1081_),
    .B(_1105_));
 sg13g2_a21oi_1 _3065_ (.A1(_1088_),
    .A2(_1090_),
    .Y(_1107_),
    .B1(_1804_));
 sg13g2_a21oi_1 _3066_ (.A1(_1101_),
    .A2(_1102_),
    .Y(_1108_),
    .B1(_1846_));
 sg13g2_a21oi_1 _3067_ (.A1(_1104_),
    .A2(_1107_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_nand3_1 _3068_ (.B(_1029_),
    .C(_1109_),
    .A(_1106_),
    .Y(_1110_));
 sg13g2_nor2_1 _3069_ (.A(_0985_),
    .B(_1012_),
    .Y(_1111_));
 sg13g2_nor2_1 _3070_ (.A(_0869_),
    .B(_1111_),
    .Y(_1112_));
 sg13g2_nand2_1 _3071_ (.Y(_1113_),
    .A(_1110_),
    .B(_1112_));
 sg13g2_nand4_1 _3072_ (.B(_1006_),
    .C(_1029_),
    .A(_1106_),
    .Y(_1114_),
    .D(_1109_));
 sg13g2_nand2_1 _3073_ (.Y(net9),
    .A(_1113_),
    .B(_1114_));
 sg13g2_nand2_1 _3074_ (.Y(_1115_),
    .A(_1745_),
    .B(_1988_));
 sg13g2_nand2_1 _3075_ (.Y(_1116_),
    .A(net62),
    .B(net69));
 sg13g2_inv_1 _3076_ (.Y(_1117_),
    .A(_1116_));
 sg13g2_a21oi_2 _3077_ (.B1(_1117_),
    .Y(_1118_),
    .A2(_1115_),
    .A1(net22));
 sg13g2_xnor2_1 _3078_ (.Y(_1119_),
    .A(_1651_),
    .B(_1985_));
 sg13g2_nand2_1 _3079_ (.Y(_1120_),
    .A(_0245_),
    .B(_1119_));
 sg13g2_nand2b_1 _3080_ (.Y(_1121_),
    .B(net20),
    .A_N(_1119_));
 sg13g2_nand2_1 _3081_ (.Y(_1122_),
    .A(_1120_),
    .B(_1121_));
 sg13g2_xor2_1 _3082_ (.B(_1122_),
    .A(_1118_),
    .X(_1123_));
 sg13g2_inv_1 _3083_ (.Y(_1124_),
    .A(_1123_));
 sg13g2_xor2_1 _3084_ (.B(_1993_),
    .A(net63),
    .X(_1125_));
 sg13g2_nand2_1 _3085_ (.Y(_1126_),
    .A(_2083_),
    .B(_1125_));
 sg13g2_o21ai_1 _3086_ (.B1(_1126_),
    .Y(_1127_),
    .A1(_1859_),
    .A2(_0951_));
 sg13g2_nand2_1 _3087_ (.Y(_1128_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_inv_1 _3088_ (.Y(_1129_),
    .A(_1128_));
 sg13g2_xnor2_1 _3089_ (.Y(_1130_),
    .A(_1129_),
    .B(_2057_));
 sg13g2_nand2b_1 _3090_ (.Y(_1131_),
    .B(_1130_),
    .A_N(_1127_));
 sg13g2_xnor2_1 _3091_ (.Y(_1132_),
    .A(_1125_),
    .B(_2083_));
 sg13g2_xor2_1 _3092_ (.B(_1989_),
    .A(net73),
    .X(_1133_));
 sg13g2_nand2_1 _3093_ (.Y(_1134_),
    .A(net36),
    .B(_1133_));
 sg13g2_o21ai_1 _3094_ (.B1(_1134_),
    .Y(_1135_),
    .A1(_1669_),
    .A2(_1990_));
 sg13g2_nor2b_1 _3095_ (.A(_1132_),
    .B_N(_1135_),
    .Y(_1136_));
 sg13g2_xnor2_1 _3096_ (.Y(_1137_),
    .A(_1128_),
    .B(net22));
 sg13g2_nand2_1 _3097_ (.Y(_1138_),
    .A(_1137_),
    .B(_1127_));
 sg13g2_inv_1 _3098_ (.Y(_1139_),
    .A(_1138_));
 sg13g2_a21oi_1 _3099_ (.A1(_1131_),
    .A2(_1136_),
    .Y(_1140_),
    .B1(_1139_));
 sg13g2_xor2_1 _3100_ (.B(net58),
    .A(_1654_),
    .X(_1141_));
 sg13g2_nand2_1 _3101_ (.Y(_1142_),
    .A(net19),
    .B(_1141_));
 sg13g2_inv_1 _3102_ (.Y(_1143_),
    .A(_1141_));
 sg13g2_nand2_1 _3103_ (.Y(_1144_),
    .A(_0240_),
    .B(_1143_));
 sg13g2_nand2_1 _3104_ (.Y(_1145_),
    .A(_1142_),
    .B(_1144_));
 sg13g2_nand2_1 _3105_ (.Y(_1146_),
    .A(net66),
    .B(net59));
 sg13g2_nand2_1 _3106_ (.Y(_1147_),
    .A(_1121_),
    .B(_1146_));
 sg13g2_inv_1 _3107_ (.Y(_1148_),
    .A(_1147_));
 sg13g2_nand2_1 _3108_ (.Y(_1149_),
    .A(_1145_),
    .B(_1148_));
 sg13g2_nand3_1 _3109_ (.B(_1144_),
    .C(_1147_),
    .A(_1142_),
    .Y(_1150_));
 sg13g2_nand2_1 _3110_ (.Y(_1151_),
    .A(_1149_),
    .B(_1150_));
 sg13g2_nor3_1 _3111_ (.A(_1124_),
    .B(_1140_),
    .C(_1151_),
    .Y(_1152_));
 sg13g2_nor2_1 _3112_ (.A(_1118_),
    .B(_1122_),
    .Y(_1153_));
 sg13g2_inv_1 _3113_ (.Y(_1154_),
    .A(_1150_));
 sg13g2_a21oi_1 _3114_ (.A1(_1149_),
    .A2(_1153_),
    .Y(_1155_),
    .B1(_1154_));
 sg13g2_nor2b_1 _3115_ (.A(_1152_),
    .B_N(_1155_),
    .Y(_1156_));
 sg13g2_xnor2_1 _3116_ (.Y(_1157_),
    .A(_1147_),
    .B(_1145_));
 sg13g2_xnor2_1 _3117_ (.Y(_1158_),
    .A(_1135_),
    .B(_1132_));
 sg13g2_inv_1 _3118_ (.Y(_1159_),
    .A(_1158_));
 sg13g2_nand2_1 _3119_ (.Y(_1160_),
    .A(_1131_),
    .B(_1138_));
 sg13g2_nor2_1 _3120_ (.A(_1159_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_xnor2_1 _3121_ (.Y(_1162_),
    .A(_1133_),
    .B(net36));
 sg13g2_nor2_1 _3122_ (.A(_1975_),
    .B(_2066_),
    .Y(_1163_));
 sg13g2_nand2_1 _3123_ (.Y(_1164_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_xnor2_1 _3124_ (.Y(_1165_),
    .A(_1991_),
    .B(_2066_));
 sg13g2_nor2_1 _3125_ (.A(_2174_),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_nor2_1 _3126_ (.A(_1163_),
    .B(_1162_),
    .Y(_1167_));
 sg13g2_a21oi_1 _3127_ (.A1(_1164_),
    .A2(_1166_),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_inv_1 _3128_ (.Y(_1169_),
    .A(_1168_));
 sg13g2_nand4_1 _3129_ (.B(_1161_),
    .C(_1169_),
    .A(_1157_),
    .Y(_1170_),
    .D(_1123_));
 sg13g2_nand2_1 _3130_ (.Y(_1171_),
    .A(_1156_),
    .B(_1170_));
 sg13g2_nand2_1 _3131_ (.Y(_1172_),
    .A(net65),
    .B(_2016_));
 sg13g2_nand2_1 _3132_ (.Y(_1173_),
    .A(_1142_),
    .B(_1172_));
 sg13g2_xor2_1 _3133_ (.B(_1980_),
    .A(_1662_),
    .X(_1174_));
 sg13g2_xnor2_1 _3134_ (.Y(_1175_),
    .A(_1174_),
    .B(net18));
 sg13g2_xnor2_1 _3135_ (.Y(_1176_),
    .A(_1173_),
    .B(_1175_));
 sg13g2_nand2_1 _3136_ (.Y(_1177_),
    .A(_1171_),
    .B(_1176_));
 sg13g2_inv_1 _3137_ (.Y(_1178_),
    .A(_1176_));
 sg13g2_nand3_1 _3138_ (.B(_1170_),
    .C(_1178_),
    .A(_1156_),
    .Y(_1179_));
 sg13g2_nand3_1 _3139_ (.B(_1179_),
    .C(net50),
    .A(_1177_),
    .Y(_1180_));
 sg13g2_xnor2_1 _3140_ (.Y(_1181_),
    .A(net65),
    .B(net70));
 sg13g2_xnor2_1 _3141_ (.Y(_1182_),
    .A(net66),
    .B(net58));
 sg13g2_xor2_1 _3142_ (.B(_1993_),
    .A(net73),
    .X(_1183_));
 sg13g2_nand2_1 _3143_ (.Y(_1184_),
    .A(_1666_),
    .B(_1989_));
 sg13g2_inv_1 _3144_ (.Y(_1185_),
    .A(_1184_));
 sg13g2_nand2_1 _3145_ (.Y(_1186_),
    .A(net73),
    .B(_1993_));
 sg13g2_inv_1 _3146_ (.Y(_1187_),
    .A(_1186_));
 sg13g2_a21oi_2 _3147_ (.B1(_1187_),
    .Y(_1188_),
    .A2(_1185_),
    .A1(_1183_));
 sg13g2_inv_1 _3148_ (.Y(_1189_),
    .A(_1188_));
 sg13g2_xor2_1 _3149_ (.B(net59),
    .A(net62),
    .X(_1190_));
 sg13g2_inv_1 _3150_ (.Y(_1191_),
    .A(_1190_));
 sg13g2_nor2_1 _3151_ (.A(net63),
    .B(net69),
    .Y(_1192_));
 sg13g2_nand2_1 _3152_ (.Y(_1193_),
    .A(_1671_),
    .B(net69));
 sg13g2_nand2b_1 _3153_ (.Y(_1194_),
    .B(_1193_),
    .A_N(_1192_));
 sg13g2_nor2_1 _3154_ (.A(_1191_),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_nand2_1 _3155_ (.Y(_1196_),
    .A(net62),
    .B(net59));
 sg13g2_o21ai_1 _3156_ (.B1(_1196_),
    .Y(_1197_),
    .A1(_1193_),
    .A2(_1191_));
 sg13g2_a21oi_1 _3157_ (.A1(_1189_),
    .A2(_1195_),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_nand2_1 _3158_ (.Y(_1199_),
    .A(net66),
    .B(net58));
 sg13g2_o21ai_1 _3159_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_1182_),
    .A2(_1198_));
 sg13g2_xnor2_1 _3160_ (.Y(_1201_),
    .A(_1181_),
    .B(_1200_));
 sg13g2_nor2_1 _3161_ (.A(_0242_),
    .B(net19),
    .Y(_1202_));
 sg13g2_nand2_1 _3162_ (.Y(_1203_),
    .A(net19),
    .B(_0242_));
 sg13g2_nand2b_1 _3163_ (.Y(_1204_),
    .B(_1203_),
    .A_N(_1202_));
 sg13g2_xnor2_1 _3164_ (.Y(_1205_),
    .A(_1201_),
    .B(_1204_));
 sg13g2_xnor2_1 _3165_ (.Y(_1206_),
    .A(net69),
    .B(_2062_));
 sg13g2_nor2_1 _3166_ (.A(_0951_),
    .B(_2066_),
    .Y(_1207_));
 sg13g2_nand2_1 _3167_ (.Y(_1208_),
    .A(_1206_),
    .B(_1207_));
 sg13g2_nand2_1 _3168_ (.Y(_1209_),
    .A(_0883_),
    .B(_0727_));
 sg13g2_nand2_1 _3169_ (.Y(_1210_),
    .A(_1208_),
    .B(_1209_));
 sg13g2_xnor2_1 _3170_ (.Y(_1211_),
    .A(_1985_),
    .B(_2083_));
 sg13g2_nand2_1 _3171_ (.Y(_1212_),
    .A(_1210_),
    .B(_1211_));
 sg13g2_inv_1 _3172_ (.Y(_1213_),
    .A(_0043_));
 sg13g2_nand2_1 _3173_ (.Y(_1214_),
    .A(_2089_),
    .B(_1213_));
 sg13g2_nand2_1 _3174_ (.Y(_1215_),
    .A(_1212_),
    .B(_1214_));
 sg13g2_xnor2_1 _3175_ (.Y(_1216_),
    .A(net58),
    .B(_2057_));
 sg13g2_nand2_1 _3176_ (.Y(_1217_),
    .A(_1215_),
    .B(_1216_));
 sg13g2_nand2_1 _3177_ (.Y(_1218_),
    .A(_0233_),
    .B(_2090_));
 sg13g2_nand2_1 _3178_ (.Y(_1219_),
    .A(_1217_),
    .B(_1218_));
 sg13g2_xnor2_1 _3179_ (.Y(_1220_),
    .A(_1981_),
    .B(net20));
 sg13g2_inv_1 _3180_ (.Y(_1221_),
    .A(_1220_));
 sg13g2_nand2_1 _3181_ (.Y(_1222_),
    .A(_1219_),
    .B(_1221_));
 sg13g2_nor2_1 _3182_ (.A(_0041_),
    .B(_0145_),
    .Y(_1223_));
 sg13g2_inv_1 _3183_ (.Y(_1224_),
    .A(_1223_));
 sg13g2_nand2_1 _3184_ (.Y(_1225_),
    .A(_1222_),
    .B(_1224_));
 sg13g2_xnor2_1 _3185_ (.Y(_1226_),
    .A(_1205_),
    .B(_1225_));
 sg13g2_nand2_1 _3186_ (.Y(_1227_),
    .A(_1226_),
    .B(_2025_));
 sg13g2_a21oi_1 _3187_ (.A1(_1227_),
    .A2(_0496_),
    .Y(_1228_),
    .B1(_2111_));
 sg13g2_nand2_1 _3188_ (.Y(_1229_),
    .A(_1180_),
    .B(_1228_));
 sg13g2_xnor2_1 _3189_ (.Y(_1230_),
    .A(net70),
    .B(_2129_));
 sg13g2_a21oi_1 _3190_ (.A1(_1230_),
    .A2(_2111_),
    .Y(_1231_),
    .B1(_2116_));
 sg13g2_nand2_1 _3191_ (.Y(_1232_),
    .A(_1229_),
    .B(_1231_));
 sg13g2_a21oi_1 _3192_ (.A1(_0234_),
    .A2(_2116_),
    .Y(_1233_),
    .B1(net28));
 sg13g2_nand2_1 _3193_ (.Y(_1234_),
    .A(_1232_),
    .B(_1233_));
 sg13g2_nand2_1 _3194_ (.Y(_1235_),
    .A(_1234_),
    .B(_0276_));
 sg13g2_nand2_1 _3195_ (.Y(_1236_),
    .A(_1235_),
    .B(_0197_));
 sg13g2_nand4_1 _3196_ (.B(net17),
    .C(_0213_),
    .A(_1236_),
    .Y(_1237_),
    .D(net44));
 sg13g2_inv_1 _3197_ (.Y(_1238_),
    .A(_1160_));
 sg13g2_nand2_1 _3198_ (.Y(_1239_),
    .A(_1158_),
    .B(_1169_));
 sg13g2_nand2b_1 _3199_ (.Y(_1240_),
    .B(_1239_),
    .A_N(_1136_));
 sg13g2_xnor2_1 _3200_ (.Y(_1241_),
    .A(_1238_),
    .B(_1240_));
 sg13g2_xnor2_1 _3201_ (.Y(_1242_),
    .A(_1194_),
    .B(_1188_));
 sg13g2_xnor2_1 _3202_ (.Y(_1243_),
    .A(_1211_),
    .B(_1210_));
 sg13g2_xnor2_1 _3203_ (.Y(_1244_),
    .A(_1242_),
    .B(_1243_));
 sg13g2_a21oi_1 _3204_ (.A1(_1244_),
    .A2(net43),
    .Y(_1245_),
    .B1(_0411_));
 sg13g2_nor2_1 _3205_ (.A(net32),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_o21ai_1 _3206_ (.B1(_1246_),
    .Y(_1247_),
    .A1(net42),
    .A2(_1241_));
 sg13g2_a21oi_1 _3207_ (.A1(net25),
    .A2(_1988_),
    .Y(_1248_),
    .B1(_2140_));
 sg13g2_o21ai_1 _3208_ (.B1(_1248_),
    .Y(_1249_),
    .A1(_1988_),
    .A2(net25));
 sg13g2_nand3_1 _3209_ (.B(net34),
    .C(_1249_),
    .A(_1247_),
    .Y(_1250_));
 sg13g2_nand2_1 _3210_ (.Y(_1251_),
    .A(net33),
    .B(_0727_));
 sg13g2_nand3_1 _3211_ (.B(_2146_),
    .C(_1251_),
    .A(_1250_),
    .Y(_1252_));
 sg13g2_nand2_1 _3212_ (.Y(_1253_),
    .A(_1252_),
    .B(net16));
 sg13g2_nand2_1 _3213_ (.Y(_1254_),
    .A(_1253_),
    .B(net38));
 sg13g2_a21oi_1 _3214_ (.A1(_1254_),
    .A2(_0914_),
    .Y(_1255_),
    .B1(net27));
 sg13g2_nand2_1 _3215_ (.Y(_1256_),
    .A(_1237_),
    .B(_1255_));
 sg13g2_nand3_1 _3216_ (.B(_1240_),
    .C(_1238_),
    .A(_1123_),
    .Y(_1257_));
 sg13g2_nand2_1 _3217_ (.Y(_1258_),
    .A(_1176_),
    .B(_1157_));
 sg13g2_nor2_1 _3218_ (.A(_1257_),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_nand2_1 _3219_ (.Y(_1260_),
    .A(net18),
    .B(_1174_));
 sg13g2_o21ai_1 _3220_ (.B1(_1260_),
    .Y(_1261_),
    .A1(_1695_),
    .A2(_1981_));
 sg13g2_xnor2_1 _3221_ (.Y(_1262_),
    .A(_1979_),
    .B(_0331_));
 sg13g2_xnor2_1 _3222_ (.Y(_1263_),
    .A(_1261_),
    .B(_1262_));
 sg13g2_nor2_1 _3223_ (.A(_1153_),
    .B(_1139_),
    .Y(_1264_));
 sg13g2_nand2_1 _3224_ (.Y(_1265_),
    .A(_1122_),
    .B(_1118_));
 sg13g2_nor2b_1 _3225_ (.A(_1264_),
    .B_N(_1265_),
    .Y(_1266_));
 sg13g2_nand3_1 _3226_ (.B(_1266_),
    .C(_1157_),
    .A(_1176_),
    .Y(_1267_));
 sg13g2_inv_1 _3227_ (.Y(_1268_),
    .A(_1175_));
 sg13g2_inv_1 _3228_ (.Y(_1269_),
    .A(_1173_));
 sg13g2_a21oi_1 _3229_ (.A1(_1269_),
    .A2(_1175_),
    .Y(_1270_),
    .B1(_1150_));
 sg13g2_a21oi_1 _3230_ (.A1(_1173_),
    .A2(_1268_),
    .Y(_1271_),
    .B1(_1270_));
 sg13g2_nand2_1 _3231_ (.Y(_1272_),
    .A(_1267_),
    .B(_1271_));
 sg13g2_nor3_1 _3232_ (.A(_1259_),
    .B(_1263_),
    .C(_1272_),
    .Y(_1273_));
 sg13g2_nor2_1 _3233_ (.A(_0786_),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_o21ai_1 _3234_ (.B1(_1263_),
    .Y(_1275_),
    .A1(_1259_),
    .A2(_1272_));
 sg13g2_nand2_1 _3235_ (.Y(_1276_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_nor2_1 _3236_ (.A(_1220_),
    .B(_1204_),
    .Y(_1277_));
 sg13g2_nand2_1 _3237_ (.Y(_1278_),
    .A(_1277_),
    .B(_1219_));
 sg13g2_o21ai_1 _3238_ (.B1(_1203_),
    .Y(_1279_),
    .A1(_1223_),
    .A2(_1202_));
 sg13g2_xor2_1 _3239_ (.B(_1978_),
    .A(net61),
    .X(_1280_));
 sg13g2_nor2_1 _3240_ (.A(_1182_),
    .B(_1181_),
    .Y(_1281_));
 sg13g2_nand2_1 _3241_ (.Y(_1282_),
    .A(net65),
    .B(net70));
 sg13g2_o21ai_1 _3242_ (.B1(_1282_),
    .Y(_1283_),
    .A1(_1199_),
    .A2(_1181_));
 sg13g2_a21oi_1 _3243_ (.A1(_1197_),
    .A2(_1281_),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_nand3_1 _3244_ (.B(_1195_),
    .C(_1281_),
    .A(_1189_),
    .Y(_1285_));
 sg13g2_nand2_1 _3245_ (.Y(_1286_),
    .A(_1284_),
    .B(_1285_));
 sg13g2_xnor2_1 _3246_ (.Y(_1287_),
    .A(_1280_),
    .B(_1286_));
 sg13g2_xnor2_1 _3247_ (.Y(_1288_),
    .A(_0837_),
    .B(net18));
 sg13g2_xnor2_1 _3248_ (.Y(_1289_),
    .A(_1287_),
    .B(_1288_));
 sg13g2_a21oi_1 _3249_ (.A1(_1278_),
    .A2(_1279_),
    .Y(_1290_),
    .B1(_1289_));
 sg13g2_nand3_1 _3250_ (.B(_1289_),
    .C(_1279_),
    .A(_1278_),
    .Y(_1291_));
 sg13g2_nand3b_1 _3251_ (.B(net48),
    .C(_1291_),
    .Y(_1292_),
    .A_N(_1290_));
 sg13g2_a21oi_1 _3252_ (.A1(_1292_),
    .A2(_0258_),
    .Y(_1293_),
    .B1(net40));
 sg13g2_nand2_1 _3253_ (.Y(_1294_),
    .A(_1276_),
    .B(_1293_));
 sg13g2_xnor2_1 _3254_ (.Y(_1295_),
    .A(_1978_),
    .B(net29));
 sg13g2_a21oi_1 _3255_ (.A1(_1295_),
    .A2(net40),
    .Y(_1296_),
    .B1(net45));
 sg13g2_nand2_1 _3256_ (.Y(_1297_),
    .A(_1294_),
    .B(_1296_));
 sg13g2_a21oi_1 _3257_ (.A1(_0244_),
    .A2(net45),
    .Y(_1298_),
    .B1(net28));
 sg13g2_nand2_1 _3258_ (.Y(_1299_),
    .A(_1297_),
    .B(_1298_));
 sg13g2_nand2_1 _3259_ (.Y(_1300_),
    .A(_1299_),
    .B(_0276_));
 sg13g2_nand2_1 _3260_ (.Y(_1301_),
    .A(_1300_),
    .B(net38));
 sg13g2_nand3b_1 _3261_ (.B(_1301_),
    .C(_0398_),
    .Y(_1302_),
    .A_N(_0479_));
 sg13g2_nor2b_1 _3262_ (.A(_1256_),
    .B_N(_1302_),
    .Y(_1303_));
 sg13g2_nand2_1 _3263_ (.Y(_1304_),
    .A(_1301_),
    .B(_0398_));
 sg13g2_buf_8 _3264_ (.A(_1304_),
    .X(_1305_));
 sg13g2_nand2_1 _3265_ (.Y(_1306_),
    .A(_1305_),
    .B(net27));
 sg13g2_nor2b_1 _3266_ (.A(_1303_),
    .B_N(_1306_),
    .Y(_1307_));
 sg13g2_nand3_1 _3267_ (.B(_1220_),
    .C(_1218_),
    .A(_1217_),
    .Y(_1308_));
 sg13g2_nand2_1 _3268_ (.Y(_1309_),
    .A(_1222_),
    .B(_1308_));
 sg13g2_xor2_1 _3269_ (.B(_1198_),
    .A(_1182_),
    .X(_1310_));
 sg13g2_nand2_1 _3270_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_inv_1 _3271_ (.Y(_1312_),
    .A(_1310_));
 sg13g2_nand3_1 _3272_ (.B(_1308_),
    .C(_1312_),
    .A(_1222_),
    .Y(_1313_));
 sg13g2_nand3_1 _3273_ (.B(_1313_),
    .C(net43),
    .A(_1311_),
    .Y(_1314_));
 sg13g2_nand2_1 _3274_ (.Y(_1315_),
    .A(_1314_),
    .B(_0459_));
 sg13g2_inv_1 _3275_ (.Y(_1316_),
    .A(_1266_));
 sg13g2_nand2_1 _3276_ (.Y(_1317_),
    .A(_1257_),
    .B(_1316_));
 sg13g2_nand2_1 _3277_ (.Y(_1318_),
    .A(_1317_),
    .B(_1157_));
 sg13g2_nand3_1 _3278_ (.B(_1316_),
    .C(_1151_),
    .A(_1257_),
    .Y(_1319_));
 sg13g2_nand3_1 _3279_ (.B(_1319_),
    .C(net46),
    .A(_1318_),
    .Y(_1320_));
 sg13g2_nand3_1 _3280_ (.B(_1320_),
    .C(_2140_),
    .A(_1315_),
    .Y(_1321_));
 sg13g2_xnor2_1 _3281_ (.Y(_1322_),
    .A(_2016_),
    .B(net29));
 sg13g2_a21oi_1 _3282_ (.A1(_1322_),
    .A2(net32),
    .Y(_1323_),
    .B1(net39));
 sg13g2_nand2_1 _3283_ (.Y(_1324_),
    .A(_1321_),
    .B(_1323_));
 sg13g2_a21oi_1 _3284_ (.A1(_2090_),
    .A2(net33),
    .Y(_1325_),
    .B1(net24));
 sg13g2_nand2_1 _3285_ (.Y(_1326_),
    .A(_1324_),
    .B(_1325_));
 sg13g2_nand2_1 _3286_ (.Y(_1327_),
    .A(_1326_),
    .B(net16));
 sg13g2_nand2_1 _3287_ (.Y(_1328_),
    .A(_1327_),
    .B(net38));
 sg13g2_nand4_1 _3288_ (.B(net17),
    .C(_0213_),
    .A(_1328_),
    .Y(_1329_),
    .D(net37));
 sg13g2_xnor2_1 _3289_ (.Y(_1330_),
    .A(_1184_),
    .B(_1183_));
 sg13g2_xor2_1 _3290_ (.B(_1206_),
    .A(_1207_),
    .X(_1331_));
 sg13g2_xor2_1 _3291_ (.B(_1331_),
    .A(_1330_),
    .X(_1332_));
 sg13g2_o21ai_1 _3292_ (.B1(_0536_),
    .Y(_1333_),
    .A1(net41),
    .A2(_1332_));
 sg13g2_nand2_1 _3293_ (.Y(_1334_),
    .A(_1159_),
    .B(_1168_));
 sg13g2_nand3_1 _3294_ (.B(net46),
    .C(_1239_),
    .A(_1334_),
    .Y(_1335_));
 sg13g2_nand3_1 _3295_ (.B(net31),
    .C(_1335_),
    .A(_1333_),
    .Y(_1336_));
 sg13g2_a21oi_1 _3296_ (.A1(net25),
    .A2(_0951_),
    .Y(_1337_),
    .B1(net31));
 sg13g2_o21ai_1 _3297_ (.B1(_1337_),
    .Y(_1338_),
    .A1(_0951_),
    .A2(net25));
 sg13g2_nand3_1 _3298_ (.B(net34),
    .C(_1338_),
    .A(_1336_),
    .Y(_1339_));
 sg13g2_nand2b_1 _3299_ (.Y(_1340_),
    .B(net30),
    .A_N(_0045_));
 sg13g2_nand3_1 _3300_ (.B(_2146_),
    .C(_1340_),
    .A(_1339_),
    .Y(_1341_));
 sg13g2_a21o_1 _3301_ (.A2(_1341_),
    .A1(net16),
    .B1(net49),
    .X(_1342_));
 sg13g2_a21oi_1 _3302_ (.A1(_1342_),
    .A2(_0201_),
    .Y(_1343_),
    .B1(net27));
 sg13g2_nand2_1 _3303_ (.Y(_1344_),
    .A(_1329_),
    .B(_1343_));
 sg13g2_nand3_1 _3304_ (.B(_0398_),
    .C(net56),
    .A(_1301_),
    .Y(_1345_));
 sg13g2_nand3_1 _3305_ (.B(_0358_),
    .C(net44),
    .A(_1236_),
    .Y(_1346_));
 sg13g2_nand2_1 _3306_ (.Y(_1347_),
    .A(_1345_),
    .B(_1346_));
 sg13g2_nor2_1 _3307_ (.A(_1344_),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_nand2_1 _3308_ (.Y(_1349_),
    .A(_1236_),
    .B(_0352_));
 sg13g2_nor2_1 _3309_ (.A(_0356_),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_nand2_1 _3310_ (.Y(_1351_),
    .A(_1350_),
    .B(_0351_));
 sg13g2_nand2_1 _3311_ (.Y(_1352_),
    .A(_1348_),
    .B(_1351_));
 sg13g2_nand2_1 _3312_ (.Y(_1353_),
    .A(_1307_),
    .B(_1352_));
 sg13g2_inv_2 _3313_ (.Y(_1354_),
    .A(_1306_));
 sg13g2_o21ai_1 _3314_ (.B1(_1193_),
    .Y(_1355_),
    .A1(_1192_),
    .A2(_1188_));
 sg13g2_xnor2_1 _3315_ (.Y(_1356_),
    .A(_1191_),
    .B(_1355_));
 sg13g2_xnor2_1 _3316_ (.Y(_1357_),
    .A(_1216_),
    .B(_1215_));
 sg13g2_xor2_1 _3317_ (.B(_1357_),
    .A(_1356_),
    .X(_1358_));
 sg13g2_nand2_1 _3318_ (.Y(_1359_),
    .A(_1358_),
    .B(net43));
 sg13g2_a21oi_1 _3319_ (.A1(_1359_),
    .A2(_2103_),
    .Y(_1360_),
    .B1(net35));
 sg13g2_a21oi_1 _3320_ (.A1(_1240_),
    .A2(_1131_),
    .Y(_1361_),
    .B1(_1139_));
 sg13g2_xnor2_1 _3321_ (.Y(_1362_),
    .A(_1123_),
    .B(_1361_));
 sg13g2_nand2_1 _3322_ (.Y(_1363_),
    .A(_1362_),
    .B(net46));
 sg13g2_nand2_1 _3323_ (.Y(_1364_),
    .A(_1360_),
    .B(_1363_));
 sg13g2_xnor2_1 _3324_ (.Y(_1365_),
    .A(net59),
    .B(net29));
 sg13g2_a21oi_1 _3325_ (.A1(_1365_),
    .A2(net35),
    .Y(_1366_),
    .B1(net39));
 sg13g2_nand2_1 _3326_ (.Y(_1367_),
    .A(_1364_),
    .B(_1366_));
 sg13g2_a21oi_1 _3327_ (.A1(_1213_),
    .A2(net33),
    .Y(_1368_),
    .B1(net24));
 sg13g2_nand2_1 _3328_ (.Y(_1369_),
    .A(_1367_),
    .B(_1368_));
 sg13g2_nand2_1 _3329_ (.Y(_1370_),
    .A(_1369_),
    .B(net16));
 sg13g2_a21oi_1 _3330_ (.A1(_1370_),
    .A2(net38),
    .Y(_1371_),
    .B1(_0486_));
 sg13g2_nand2_1 _3331_ (.Y(_1372_),
    .A(_1371_),
    .B(_0472_));
 sg13g2_o21ai_1 _3332_ (.B1(_1372_),
    .Y(_1373_),
    .A1(_0214_),
    .A2(_1305_));
 sg13g2_nand2_1 _3333_ (.Y(_1374_),
    .A(_1351_),
    .B(net23));
 sg13g2_nor2_1 _3334_ (.A(_1373_),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_nor2_2 _3335_ (.A(_1354_),
    .B(_1375_),
    .Y(_1376_));
 sg13g2_inv_4 _3336_ (.A(_1376_),
    .Y(_1377_));
 sg13g2_nand2_1 _3337_ (.Y(_1378_),
    .A(_1353_),
    .B(_1377_));
 sg13g2_nand2_1 _3338_ (.Y(_1379_),
    .A(_1346_),
    .B(net23));
 sg13g2_inv_1 _3339_ (.Y(_1380_),
    .A(_1379_));
 sg13g2_nand2_1 _3340_ (.Y(_1381_),
    .A(_1350_),
    .B(_0981_));
 sg13g2_nand2_1 _3341_ (.Y(_1382_),
    .A(_1350_),
    .B(net56));
 sg13g2_nand3_1 _3342_ (.B(_1381_),
    .C(_1382_),
    .A(_1380_),
    .Y(_1383_));
 sg13g2_inv_1 _3343_ (.Y(_1384_),
    .A(_1383_));
 sg13g2_nand2_1 _3344_ (.Y(_1385_),
    .A(_1378_),
    .B(_1384_));
 sg13g2_inv_8 _3345_ (.Y(_1386_),
    .A(_1305_));
 sg13g2_nand2_1 _3346_ (.Y(_1387_),
    .A(_1385_),
    .B(_1386_));
 sg13g2_inv_1 _3347_ (.Y(_1388_),
    .A(net37));
 sg13g2_a21oi_1 _3348_ (.A1(_1326_),
    .A2(net16),
    .Y(_1389_),
    .B1(net49));
 sg13g2_nor3_1 _3349_ (.A(_1388_),
    .B(_0484_),
    .C(_1389_),
    .Y(_1390_));
 sg13g2_nor2_1 _3350_ (.A(net27),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_nand3_1 _3351_ (.B(_0398_),
    .C(_0351_),
    .A(_1301_),
    .Y(_1392_));
 sg13g2_nand3_1 _3352_ (.B(_1392_),
    .C(_1329_),
    .A(_1391_),
    .Y(_1393_));
 sg13g2_nor2b_1 _3353_ (.A(_1354_),
    .B_N(_1393_),
    .Y(_1394_));
 sg13g2_nand2_1 _3354_ (.Y(_1395_),
    .A(_1387_),
    .B(_1394_));
 sg13g2_nand2b_1 _3355_ (.Y(_1396_),
    .B(_1386_),
    .A_N(_0448_));
 sg13g2_nor2b_1 _3356_ (.A(_1167_),
    .B_N(_1164_),
    .Y(_1397_));
 sg13g2_xnor2_1 _3357_ (.Y(_1398_),
    .A(_1166_),
    .B(_1397_));
 sg13g2_o21ai_1 _3358_ (.B1(_0959_),
    .Y(_1399_),
    .A1(net42),
    .A2(_1398_));
 sg13g2_a21oi_1 _3359_ (.A1(net26),
    .A2(_1989_),
    .Y(_1400_),
    .B1(net31));
 sg13g2_o21ai_1 _3360_ (.B1(_1400_),
    .Y(_1401_),
    .A1(_1989_),
    .A2(net26));
 sg13g2_nand3_1 _3361_ (.B(net34),
    .C(_1401_),
    .A(_1399_),
    .Y(_1402_));
 sg13g2_nand2b_1 _3362_ (.Y(_1403_),
    .B(net30),
    .A_N(_0021_));
 sg13g2_nand3_1 _3363_ (.B(_2146_),
    .C(_1403_),
    .A(_1402_),
    .Y(_1404_));
 sg13g2_nor2_1 _3364_ (.A(_1388_),
    .B(_1389_),
    .Y(_1405_));
 sg13g2_a22oi_1 _3365_ (.Y(_1406_),
    .B1(_0358_),
    .B2(_1405_),
    .A2(_1404_),
    .A1(_0439_));
 sg13g2_nand3_1 _3366_ (.B(_1396_),
    .C(_1406_),
    .A(_1382_),
    .Y(_1407_));
 sg13g2_nand3_1 _3367_ (.B(_1407_),
    .C(_1306_),
    .A(_1352_),
    .Y(_1408_));
 sg13g2_inv_1 _3368_ (.Y(_1409_),
    .A(_1307_));
 sg13g2_nand2_1 _3369_ (.Y(_1410_),
    .A(_1376_),
    .B(_1305_));
 sg13g2_a21oi_1 _3370_ (.A1(_1408_),
    .A2(_1409_),
    .Y(_1411_),
    .B1(_1410_));
 sg13g2_nand3_1 _3371_ (.B(net17),
    .C(net44),
    .A(_1236_),
    .Y(_1412_));
 sg13g2_nor2b_1 _3372_ (.A(_1412_),
    .B_N(_0351_),
    .Y(_1413_));
 sg13g2_nor3_1 _3373_ (.A(_1413_),
    .B(_1344_),
    .C(_1347_),
    .Y(_1414_));
 sg13g2_nor2_1 _3374_ (.A(_1375_),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_nor2_1 _3375_ (.A(_0949_),
    .B(_1305_),
    .Y(_1416_));
 sg13g2_nor2_1 _3376_ (.A(_0987_),
    .B(_1412_),
    .Y(_1417_));
 sg13g2_nand4_1 _3377_ (.B(net17),
    .C(net56),
    .A(_1328_),
    .Y(_1418_),
    .D(net37));
 sg13g2_xnor2_1 _3378_ (.Y(_1419_),
    .A(_1991_),
    .B(net25));
 sg13g2_xnor2_1 _3379_ (.Y(_1420_),
    .A(_0054_),
    .B(_1165_));
 sg13g2_o21ai_1 _3380_ (.B1(net31),
    .Y(_1421_),
    .A1(net42),
    .A2(_1420_));
 sg13g2_o21ai_1 _3381_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net31),
    .A2(_1419_));
 sg13g2_nand2_1 _3382_ (.Y(_1423_),
    .A(net30),
    .B(_1975_));
 sg13g2_nand3_1 _3383_ (.B(_2146_),
    .C(_1423_),
    .A(_1422_),
    .Y(_1424_));
 sg13g2_a22oi_1 _3384_ (.Y(_1425_),
    .B1(_0358_),
    .B2(_1371_),
    .A2(_1424_),
    .A1(_0526_));
 sg13g2_nand2_1 _3385_ (.Y(_1426_),
    .A(_1418_),
    .B(_1425_));
 sg13g2_nor3_1 _3386_ (.A(_1416_),
    .B(_1417_),
    .C(_1426_),
    .Y(_1427_));
 sg13g2_nand2b_1 _3387_ (.Y(_1428_),
    .B(_1427_),
    .A_N(_1374_));
 sg13g2_nand2_1 _3388_ (.Y(_1429_),
    .A(_1415_),
    .B(_1428_));
 sg13g2_nor2_1 _3389_ (.A(_1354_),
    .B(_1384_),
    .Y(_1430_));
 sg13g2_inv_4 _3390_ (.A(_1407_),
    .Y(_1431_));
 sg13g2_nand3_1 _3391_ (.B(_1302_),
    .C(_1255_),
    .A(_1237_),
    .Y(_1432_));
 sg13g2_nand2_1 _3392_ (.Y(_1433_),
    .A(_1432_),
    .B(_1393_));
 sg13g2_nor2_1 _3393_ (.A(_1431_),
    .B(_1433_),
    .Y(_1434_));
 sg13g2_nor2_1 _3394_ (.A(_1305_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_a21oi_1 _3395_ (.A1(_1429_),
    .A2(_1430_),
    .Y(_1436_),
    .B1(_1435_));
 sg13g2_nor2_1 _3396_ (.A(_1411_),
    .B(_1436_),
    .Y(_1437_));
 sg13g2_nand2_1 _3397_ (.Y(_1438_),
    .A(_1395_),
    .B(_1437_));
 sg13g2_inv_1 _3398_ (.Y(_1439_),
    .A(_1430_));
 sg13g2_nand2_1 _3399_ (.Y(_1440_),
    .A(_1438_),
    .B(_1439_));
 sg13g2_nand3_1 _3400_ (.B(_1430_),
    .C(_1437_),
    .A(_1395_),
    .Y(_1441_));
 sg13g2_nand2_1 _3401_ (.Y(_1442_),
    .A(_1440_),
    .B(_1441_));
 sg13g2_nand2_1 _3402_ (.Y(_1443_),
    .A(_1442_),
    .B(_1376_));
 sg13g2_nand3_1 _3403_ (.B(_1439_),
    .C(_1437_),
    .A(_1395_),
    .Y(_1444_));
 sg13g2_buf_8 _3404_ (.A(_1444_),
    .X(_1445_));
 sg13g2_nand2_1 _3405_ (.Y(_1446_),
    .A(_1445_),
    .B(_1386_));
 sg13g2_buf_8 _3406_ (.A(_1446_),
    .X(_1447_));
 sg13g2_xnor2_1 _3407_ (.Y(_1448_),
    .A(_1394_),
    .B(_1447_));
 sg13g2_nand2_1 _3408_ (.Y(_1449_),
    .A(_1447_),
    .B(_1394_));
 sg13g2_o21ai_1 _3409_ (.B1(_1449_),
    .Y(_1450_),
    .A1(_1443_),
    .A2(_1448_));
 sg13g2_nor2_1 _3410_ (.A(_1354_),
    .B(_1414_),
    .Y(_1451_));
 sg13g2_nand2_1 _3411_ (.Y(_1452_),
    .A(_1442_),
    .B(_1451_));
 sg13g2_inv_1 _3412_ (.Y(_1453_),
    .A(_1452_));
 sg13g2_nand3_1 _3413_ (.B(_1386_),
    .C(_1409_),
    .A(_1445_),
    .Y(_1454_));
 sg13g2_nand2_1 _3414_ (.Y(_1455_),
    .A(_1447_),
    .B(_1307_));
 sg13g2_inv_1 _3415_ (.Y(_1456_),
    .A(_1455_));
 sg13g2_a21oi_1 _3416_ (.A1(_1453_),
    .A2(_1454_),
    .Y(_1457_),
    .B1(_1456_));
 sg13g2_inv_2 _3417_ (.Y(_1458_),
    .A(_1448_));
 sg13g2_nand2_1 _3418_ (.Y(_1459_),
    .A(_1438_),
    .B(_1430_));
 sg13g2_nand2_2 _3419_ (.Y(_1460_),
    .A(_1459_),
    .B(_1445_));
 sg13g2_nand2_1 _3420_ (.Y(_1461_),
    .A(_1460_),
    .B(_1376_));
 sg13g2_nand3_1 _3421_ (.B(_1445_),
    .C(_1377_),
    .A(_1459_),
    .Y(_1462_));
 sg13g2_nand2_1 _3422_ (.Y(_1463_),
    .A(_1461_),
    .B(_1462_));
 sg13g2_nand2_1 _3423_ (.Y(_1464_),
    .A(_1458_),
    .B(_1463_));
 sg13g2_nor2_1 _3424_ (.A(_1457_),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_nor2_1 _3425_ (.A(_1450_),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_nand2_1 _3426_ (.Y(_1467_),
    .A(_1428_),
    .B(_1306_));
 sg13g2_nand3_1 _3427_ (.B(_1441_),
    .C(_1467_),
    .A(_1440_),
    .Y(_1468_));
 sg13g2_buf_2 _3428_ (.A(_1468_),
    .X(_1469_));
 sg13g2_nand3_1 _3429_ (.B(_1386_),
    .C(_1431_),
    .A(_1445_),
    .Y(_1470_));
 sg13g2_a21oi_1 _3430_ (.A1(_1445_),
    .A2(_1386_),
    .Y(_1471_),
    .B1(_1431_));
 sg13g2_a21oi_2 _3431_ (.B1(_1471_),
    .Y(_1472_),
    .A2(_1470_),
    .A1(_1469_));
 sg13g2_inv_1 _3432_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_nand2_1 _3433_ (.Y(_1474_),
    .A(_1460_),
    .B(_1377_));
 sg13g2_nand2_1 _3434_ (.Y(_1475_),
    .A(_1443_),
    .B(_1474_));
 sg13g2_nor2_1 _3435_ (.A(_1448_),
    .B(_1475_),
    .Y(_1476_));
 sg13g2_nand2_1 _3436_ (.Y(_1477_),
    .A(_1455_),
    .B(_1454_));
 sg13g2_inv_1 _3437_ (.Y(_1478_),
    .A(_1451_));
 sg13g2_nand3_1 _3438_ (.B(_1441_),
    .C(_1478_),
    .A(_1440_),
    .Y(_1479_));
 sg13g2_buf_8 _3439_ (.A(_1479_),
    .X(_1480_));
 sg13g2_nand2_2 _3440_ (.Y(_1481_),
    .A(_1452_),
    .B(_1480_));
 sg13g2_nor2_1 _3441_ (.A(_1477_),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_nand3_1 _3442_ (.B(_1476_),
    .C(_1482_),
    .A(_1473_),
    .Y(_1483_));
 sg13g2_nand2_1 _3443_ (.Y(_1484_),
    .A(_1466_),
    .B(_1483_));
 sg13g2_inv_1 _3444_ (.Y(_1485_),
    .A(_1438_));
 sg13g2_nand2_1 _3445_ (.Y(_1486_),
    .A(_1484_),
    .B(_1485_));
 sg13g2_nand2_1 _3446_ (.Y(_1487_),
    .A(_1486_),
    .B(\dither_threshold[6] ));
 sg13g2_nand3_1 _3447_ (.B(_0628_),
    .C(_1485_),
    .A(_1484_),
    .Y(_1488_));
 sg13g2_nand2_1 _3448_ (.Y(_1489_),
    .A(_1487_),
    .B(_1488_));
 sg13g2_nand2_1 _3449_ (.Y(_1490_),
    .A(_1447_),
    .B(_1409_));
 sg13g2_nand3_1 _3450_ (.B(_1386_),
    .C(_1307_),
    .A(_1445_),
    .Y(_1491_));
 sg13g2_nand2_1 _3451_ (.Y(_1492_),
    .A(_1490_),
    .B(_1491_));
 sg13g2_nand2_1 _3452_ (.Y(_1493_),
    .A(_1463_),
    .B(_1492_));
 sg13g2_a21oi_1 _3453_ (.A1(_1471_),
    .A2(_1480_),
    .Y(_1494_),
    .B1(_1453_));
 sg13g2_nor2_1 _3454_ (.A(_1493_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_inv_1 _3455_ (.Y(_1496_),
    .A(_1443_));
 sg13g2_a21oi_1 _3456_ (.A1(_1456_),
    .A2(_1474_),
    .Y(_1497_),
    .B1(_1496_));
 sg13g2_nor2b_1 _3457_ (.A(_1495_),
    .B_N(_1497_),
    .Y(_1498_));
 sg13g2_nor2_1 _3458_ (.A(_1477_),
    .B(_1475_),
    .Y(_1499_));
 sg13g2_nand2_1 _3459_ (.Y(_1500_),
    .A(_1447_),
    .B(_1407_));
 sg13g2_nand2_1 _3460_ (.Y(_1501_),
    .A(_1500_),
    .B(_1470_));
 sg13g2_nor2_1 _3461_ (.A(_1501_),
    .B(_1481_),
    .Y(_1502_));
 sg13g2_nand3_1 _3462_ (.B(_1502_),
    .C(_1469_),
    .A(_1499_),
    .Y(_1503_));
 sg13g2_nand2_1 _3463_ (.Y(_1504_),
    .A(_1498_),
    .B(_1503_));
 sg13g2_nand2_1 _3464_ (.Y(_1505_),
    .A(_1504_),
    .B(_1448_));
 sg13g2_nand3_1 _3465_ (.B(_1503_),
    .C(_1458_),
    .A(_1498_),
    .Y(_1506_));
 sg13g2_nand2_1 _3466_ (.Y(_1507_),
    .A(_1505_),
    .B(_1506_));
 sg13g2_nand2_1 _3467_ (.Y(_1508_),
    .A(_1507_),
    .B(_1840_));
 sg13g2_nand3_1 _3468_ (.B(_1506_),
    .C(_0651_),
    .A(_1505_),
    .Y(_1509_));
 sg13g2_nand2_1 _3469_ (.Y(_1510_),
    .A(_1508_),
    .B(_1509_));
 sg13g2_nor2_1 _3470_ (.A(_1489_),
    .B(_1510_),
    .Y(_1511_));
 sg13g2_nand2_1 _3471_ (.Y(_1512_),
    .A(_1473_),
    .B(_1482_));
 sg13g2_nand2_1 _3472_ (.Y(_1513_),
    .A(_1512_),
    .B(_1457_));
 sg13g2_nand2_1 _3473_ (.Y(_1514_),
    .A(_1513_),
    .B(_1475_));
 sg13g2_nand3_1 _3474_ (.B(_1463_),
    .C(_1457_),
    .A(_1512_),
    .Y(_1515_));
 sg13g2_nand2_1 _3475_ (.Y(_1516_),
    .A(_1514_),
    .B(_1515_));
 sg13g2_nand2_1 _3476_ (.Y(_1517_),
    .A(_1516_),
    .B(_1835_));
 sg13g2_nand3_1 _3477_ (.B(_1515_),
    .C(_1841_),
    .A(_1514_),
    .Y(_1518_));
 sg13g2_nand2_1 _3478_ (.Y(_1519_),
    .A(_1472_),
    .B(_1452_));
 sg13g2_nand2_1 _3479_ (.Y(_1520_),
    .A(_1519_),
    .B(_1480_));
 sg13g2_nand2_1 _3480_ (.Y(_1521_),
    .A(_1520_),
    .B(_1477_));
 sg13g2_nand3_1 _3481_ (.B(_1480_),
    .C(_1492_),
    .A(_1519_),
    .Y(_1522_));
 sg13g2_nand2_1 _3482_ (.Y(_1523_),
    .A(_1521_),
    .B(_1522_));
 sg13g2_nor2_1 _3483_ (.A(\dither_threshold[3] ),
    .B(_1523_),
    .Y(_1524_));
 sg13g2_nand3_1 _3484_ (.B(_1518_),
    .C(_1524_),
    .A(_1517_),
    .Y(_1525_));
 sg13g2_nand2_1 _3485_ (.Y(_1526_),
    .A(_1516_),
    .B(_1807_));
 sg13g2_nand2_1 _3486_ (.Y(_1527_),
    .A(_1525_),
    .B(_1526_));
 sg13g2_nand3_1 _3487_ (.B(_1507_),
    .C(_1804_),
    .A(_1487_),
    .Y(_1528_));
 sg13g2_nand2_1 _3488_ (.Y(_1529_),
    .A(_1528_),
    .B(_1488_));
 sg13g2_a21oi_1 _3489_ (.A1(_1511_),
    .A2(_1527_),
    .Y(_1530_),
    .B1(_1529_));
 sg13g2_xnor2_1 _3490_ (.Y(_1531_),
    .A(_1467_),
    .B(_1460_));
 sg13g2_xor2_1 _3491_ (.B(_1501_),
    .A(_1469_),
    .X(_1532_));
 sg13g2_xnor2_1 _3492_ (.Y(_1533_),
    .A(_1821_),
    .B(_1532_));
 sg13g2_xor2_1 _3493_ (.B(_1472_),
    .A(_1481_),
    .X(_1534_));
 sg13g2_nand2_1 _3494_ (.Y(_1535_),
    .A(_1534_),
    .B(_1809_));
 sg13g2_xnor2_1 _3495_ (.Y(_1536_),
    .A(_1481_),
    .B(_1472_));
 sg13g2_nand2_1 _3496_ (.Y(_1537_),
    .A(_1536_),
    .B(_1808_));
 sg13g2_nand2_1 _3497_ (.Y(_1538_),
    .A(_1535_),
    .B(_1537_));
 sg13g2_nor2_1 _3498_ (.A(_1533_),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_o21ai_1 _3499_ (.B1(_1539_),
    .Y(_1540_),
    .A1(_1799_),
    .A2(_1531_));
 sg13g2_nor2_1 _3500_ (.A(_1801_),
    .B(_1532_),
    .Y(_1541_));
 sg13g2_inv_1 _3501_ (.Y(_1542_),
    .A(_1535_));
 sg13g2_a21oi_1 _3502_ (.A1(_1537_),
    .A2(_1541_),
    .Y(_1543_),
    .B1(_1542_));
 sg13g2_nand2_1 _3503_ (.Y(_1544_),
    .A(_1540_),
    .B(_1543_));
 sg13g2_xnor2_1 _3504_ (.Y(_1545_),
    .A(_1827_),
    .B(_1523_));
 sg13g2_nand2_1 _3505_ (.Y(_1546_),
    .A(_1517_),
    .B(_1518_));
 sg13g2_nor2_1 _3506_ (.A(_1545_),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_nand3_1 _3507_ (.B(_1544_),
    .C(_1547_),
    .A(_1511_),
    .Y(_1548_));
 sg13g2_nand2_1 _3508_ (.Y(_1549_),
    .A(_1530_),
    .B(_1548_));
 sg13g2_xnor2_1 _3509_ (.Y(_1550_),
    .A(_1800_),
    .B(_1531_));
 sg13g2_nor3_1 _3510_ (.A(_1533_),
    .B(_1550_),
    .C(_1538_),
    .Y(_1551_));
 sg13g2_nand3_1 _3511_ (.B(_1547_),
    .C(_1551_),
    .A(_1511_),
    .Y(_1552_));
 sg13g2_nand3_1 _3512_ (.B(_1460_),
    .C(_1552_),
    .A(_1549_),
    .Y(_1553_));
 sg13g2_inv_1 _3513_ (.Y(_1554_),
    .A(_1447_));
 sg13g2_nand2_1 _3514_ (.Y(_1555_),
    .A(_1553_),
    .B(_1554_));
 sg13g2_nand4_1 _3515_ (.B(_1447_),
    .C(_1460_),
    .A(_1549_),
    .Y(_1556_),
    .D(_1552_));
 sg13g2_nand2_1 _3516_ (.Y(net10),
    .A(_1555_),
    .B(_1556_));
 sg13g2_a21oi_1 _3517_ (.A1(_0698_),
    .A2(_0702_),
    .Y(_1557_),
    .B1(_0597_));
 sg13g2_nor2b_1 _3518_ (.A(_1557_),
    .B_N(_0703_),
    .Y(net12));
 sg13g2_a21oi_1 _3519_ (.A1(_1106_),
    .A2(_1109_),
    .Y(_1558_),
    .B1(_1029_));
 sg13g2_nor2b_1 _3520_ (.A(_1558_),
    .B_N(_1110_),
    .Y(net13));
 sg13g2_a21oi_1 _3521_ (.A1(_1549_),
    .A2(_1552_),
    .Y(_1559_),
    .B1(_1460_));
 sg13g2_nor2b_1 _3522_ (.A(_1559_),
    .B_N(_1553_),
    .Y(net14));
 sg13g2_nor4_1 _3523_ (.A(\counter[21] ),
    .B(\counter[20] ),
    .C(\counter[23] ),
    .D(\counter[22] ),
    .Y(_1560_));
 sg13g2_nor4_1 _3524_ (.A(\counter[17] ),
    .B(\counter[16] ),
    .C(\counter[19] ),
    .D(\counter[18] ),
    .Y(_1561_));
 sg13g2_buf_1 _3525_ (.A(\counter[26] ),
    .X(_1562_));
 sg13g2_nor3_1 _3526_ (.A(\counter[25] ),
    .B(\counter[24] ),
    .C(_1562_),
    .Y(_1563_));
 sg13g2_and3_1 _3527_ (.X(_1564_),
    .A(_1560_),
    .B(_1561_),
    .C(_1563_));
 sg13g2_inv_1 _3528_ (.Y(_1565_),
    .A(\counter[4] ));
 sg13g2_inv_1 _3529_ (.Y(_1566_),
    .A(\counter[7] ));
 sg13g2_nand2_1 _3530_ (.Y(_1567_),
    .A(_1565_),
    .B(_1566_));
 sg13g2_nor2_1 _3531_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1568_));
 sg13g2_inv_1 _3532_ (.Y(_1569_),
    .A(\counter[2] ));
 sg13g2_nand3b_1 _3533_ (.B(_1568_),
    .C(_1569_),
    .Y(_1570_),
    .A_N(\counter[3] ));
 sg13g2_nor4_1 _3534_ (.A(\counter[5] ),
    .B(\counter[6] ),
    .C(_1567_),
    .D(_1570_),
    .Y(_1571_));
 sg13g2_buf_1 _3535_ (.A(\counter[13] ),
    .X(_1572_));
 sg13g2_buf_1 _3536_ (.A(\counter[12] ),
    .X(_1573_));
 sg13g2_buf_1 _3537_ (.A(\counter[14] ),
    .X(_1574_));
 sg13g2_nor4_1 _3538_ (.A(_1572_),
    .B(_1573_),
    .C(\counter[15] ),
    .D(_1574_),
    .Y(_1575_));
 sg13g2_nor4_1 _3539_ (.A(\counter[9] ),
    .B(\counter[8] ),
    .C(\counter[11] ),
    .D(\counter[10] ),
    .Y(_1576_));
 sg13g2_nand4_1 _3540_ (.B(_1571_),
    .C(_1575_),
    .A(_1564_),
    .Y(_0008_),
    .D(_1576_));
 sg13g2_buf_1 _3541_ (.A(\i_project.controller_0.rst_n ),
    .X(_1577_));
 sg13g2_buf_1 _3542_ (.A(_1577_),
    .X(_1578_));
 sg13g2_buf_2 _3543_ (.A(\i_project.controller_0.divider[0] ),
    .X(_1579_));
 sg13g2_inv_1 _3544_ (.Y(_1580_),
    .A(_1579_));
 sg13g2_nor2_1 _3545_ (.A(net68),
    .B(\i_project.controller_0.grey_pass[10] ),
    .Y(_1581_));
 sg13g2_a21oi_1 _3546_ (.A1(net68),
    .A2(_1580_),
    .Y(_0003_),
    .B1(_1581_));
 sg13g2_buf_2 _3547_ (.A(\i_project.controller_0.divider[1] ),
    .X(_1582_));
 sg13g2_inv_1 _3548_ (.Y(_1583_),
    .A(_1582_));
 sg13g2_buf_1 _3549_ (.A(_1583_),
    .X(_1584_));
 sg13g2_nor2_1 _3550_ (.A(net68),
    .B(\i_project.controller_0.grey_pass[11] ),
    .Y(_1585_));
 sg13g2_a21oi_1 _3551_ (.A1(net68),
    .A2(_1584_),
    .Y(_0004_),
    .B1(_1585_));
 sg13g2_buf_1 _3552_ (.A(rst_n),
    .X(_1586_));
 sg13g2_inv_1 _3553_ (.Y(_1587_),
    .A(_1586_));
 sg13g2_buf_1 _3554_ (.A(_1587_),
    .X(_1588_));
 sg13g2_inv_1 _3555_ (.Y(_1589_),
    .A(\counter[25] ));
 sg13g2_inv_1 _3556_ (.Y(_1590_),
    .A(\counter[24] ));
 sg13g2_nand2_1 _3557_ (.Y(_1591_),
    .A(\counter[23] ),
    .B(\counter[22] ));
 sg13g2_nor3_1 _3558_ (.A(_1589_),
    .B(_1590_),
    .C(_1591_),
    .Y(_1592_));
 sg13g2_inv_1 _3559_ (.Y(_1593_),
    .A(_1592_));
 sg13g2_inv_1 _3560_ (.Y(_1594_),
    .A(\counter[21] ));
 sg13g2_inv_1 _3561_ (.Y(_1595_),
    .A(\counter[20] ));
 sg13g2_inv_1 _3562_ (.Y(_1596_),
    .A(_1572_));
 sg13g2_inv_1 _3563_ (.Y(_1597_),
    .A(\counter[11] ));
 sg13g2_inv_1 _3564_ (.Y(_1598_),
    .A(\counter[10] ));
 sg13g2_inv_1 _3565_ (.Y(_1599_),
    .A(\counter[9] ));
 sg13g2_inv_1 _3566_ (.Y(_1600_),
    .A(\counter[8] ));
 sg13g2_inv_1 _3567_ (.Y(_1601_),
    .A(\counter[6] ));
 sg13g2_nand2_1 _3568_ (.Y(_1602_),
    .A(\counter[5] ),
    .B(\counter[4] ));
 sg13g2_nand2_1 _3569_ (.Y(_1603_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_nor2_1 _3570_ (.A(_1569_),
    .B(_1603_),
    .Y(_1604_));
 sg13g2_nand2_1 _3571_ (.Y(_1605_),
    .A(_1604_),
    .B(\counter[3] ));
 sg13g2_nor2_1 _3572_ (.A(_1602_),
    .B(_1605_),
    .Y(_1606_));
 sg13g2_inv_1 _3573_ (.Y(_1607_),
    .A(_1606_));
 sg13g2_nor2_1 _3574_ (.A(_1601_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_nand2_1 _3575_ (.Y(_1609_),
    .A(_1608_),
    .B(\counter[7] ));
 sg13g2_nor2_1 _3576_ (.A(_1600_),
    .B(_1609_),
    .Y(_1610_));
 sg13g2_inv_1 _3577_ (.Y(_1611_),
    .A(_1610_));
 sg13g2_nor2_1 _3578_ (.A(_1599_),
    .B(_1611_),
    .Y(_1612_));
 sg13g2_inv_1 _3579_ (.Y(_1613_),
    .A(_1612_));
 sg13g2_nor3_1 _3580_ (.A(_1597_),
    .B(_1598_),
    .C(_1613_),
    .Y(_1614_));
 sg13g2_nand2_1 _3581_ (.Y(_1615_),
    .A(_1614_),
    .B(_1573_));
 sg13g2_nor2_1 _3582_ (.A(_1596_),
    .B(_1615_),
    .Y(_1616_));
 sg13g2_nand3_1 _3583_ (.B(\counter[15] ),
    .C(_1574_),
    .A(_1616_),
    .Y(_1617_));
 sg13g2_nor2b_1 _3584_ (.A(_1617_),
    .B_N(\counter[16] ),
    .Y(_1618_));
 sg13g2_nand2_1 _3585_ (.Y(_1619_),
    .A(_1618_),
    .B(\counter[17] ));
 sg13g2_nor2b_1 _3586_ (.A(_1619_),
    .B_N(\counter[18] ),
    .Y(_1620_));
 sg13g2_nand2_1 _3587_ (.Y(_1621_),
    .A(_1620_),
    .B(\counter[19] ));
 sg13g2_nor2_1 _3588_ (.A(_1595_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_inv_1 _3589_ (.Y(_1623_),
    .A(_1622_));
 sg13g2_nor2_2 _3590_ (.A(_1594_),
    .B(_1623_),
    .Y(_1624_));
 sg13g2_inv_2 _3591_ (.Y(_1625_),
    .A(_1624_));
 sg13g2_nor2_1 _3592_ (.A(_1593_),
    .B(_1625_),
    .Y(_1626_));
 sg13g2_nand2_1 _3593_ (.Y(_1627_),
    .A(_1626_),
    .B(_1562_));
 sg13g2_nor2b_1 _3594_ (.A(_1627_),
    .B_N(\counter[27] ),
    .Y(_1628_));
 sg13g2_a21oi_1 _3595_ (.A1(_1628_),
    .A2(\counter[28] ),
    .Y(_1629_),
    .B1(\counter[29] ));
 sg13g2_nand3_1 _3596_ (.B(\counter[28] ),
    .C(\counter[29] ),
    .A(_1628_),
    .Y(_1630_));
 sg13g2_inv_1 _3597_ (.Y(_1631_),
    .A(_1630_));
 sg13g2_nor3_2 _3598_ (.A(net67),
    .B(_1629_),
    .C(_1631_),
    .Y(_0079_));
 sg13g2_inv_1 _3599_ (.Y(_1632_),
    .A(_1627_));
 sg13g2_nor2_1 _3600_ (.A(\counter[27] ),
    .B(_1632_),
    .Y(_1633_));
 sg13g2_nor3_1 _3601_ (.A(_1587_),
    .B(_1628_),
    .C(_1633_),
    .Y(_0077_));
 sg13g2_inv_1 _3602_ (.Y(_1634_),
    .A(_0077_));
 sg13g2_nand4_1 _3603_ (.B(\counter[20] ),
    .C(_1562_),
    .A(\counter[21] ),
    .Y(_1635_),
    .D(\counter[27] ));
 sg13g2_nand4_1 _3604_ (.B(\counter[16] ),
    .C(\counter[19] ),
    .A(\counter[17] ),
    .Y(_1636_),
    .D(\counter[18] ));
 sg13g2_nand4_1 _3605_ (.B(_1573_),
    .C(\counter[15] ),
    .A(_1572_),
    .Y(_1637_),
    .D(_1574_));
 sg13g2_nor4_1 _3606_ (.A(_1635_),
    .B(_1636_),
    .C(_1593_),
    .D(_1637_),
    .Y(_1638_));
 sg13g2_inv_1 _3607_ (.Y(_1639_),
    .A(_1605_));
 sg13g2_nor3_1 _3608_ (.A(_1566_),
    .B(_1601_),
    .C(_1602_),
    .Y(_1640_));
 sg13g2_nor4_1 _3609_ (.A(_1599_),
    .B(_1600_),
    .C(_1597_),
    .D(_1598_),
    .Y(_1641_));
 sg13g2_nand4_1 _3610_ (.B(_1639_),
    .C(_1640_),
    .A(_1638_),
    .Y(_1642_),
    .D(_1641_));
 sg13g2_xor2_1 _3611_ (.B(_1642_),
    .A(\counter[28] ),
    .X(_1643_));
 sg13g2_nor2_1 _3612_ (.A(_1587_),
    .B(_1643_),
    .Y(_0078_));
 sg13g2_nand2_1 _3613_ (.Y(_1644_),
    .A(_1634_),
    .B(_0078_));
 sg13g2_nor2_1 _3614_ (.A(_0078_),
    .B(_1634_),
    .Y(_1645_));
 sg13g2_a21oi_1 _3615_ (.A1(_0079_),
    .A2(_1644_),
    .Y(_0000_),
    .B1(_1645_));
 sg13g2_inv_1 _3616_ (.Y(_1646_),
    .A(_0079_));
 sg13g2_o21ai_1 _3617_ (.B1(_1644_),
    .Y(_0001_),
    .A1(_1645_),
    .A2(_1646_));
 sg13g2_a21o_1 _3618_ (.A2(_0078_),
    .A1(_0079_),
    .B1(_0077_),
    .X(_0002_));
 sg13g2_buf_1 _3619_ (.A(ui_in[7]),
    .X(_1647_));
 sg13g2_mux2_1 _3620_ (.A0(_0012_),
    .A1(net1),
    .S(net74),
    .X(_0009_));
 sg13g2_mux2_1 _3621_ (.A0(_0013_),
    .A1(net2),
    .S(net74),
    .X(_0010_));
 sg13g2_mux2_1 _3622_ (.A0(_0014_),
    .A1(net3),
    .S(net74),
    .X(_0011_));
 sg13g2_nand2_1 _3623_ (.Y(_1648_),
    .A(net74),
    .B(net5));
 sg13g2_o21ai_1 _3624_ (.B1(_1648_),
    .Y(_0005_),
    .A1(net74),
    .A2(_1590_));
 sg13g2_nand2_1 _3625_ (.Y(_1649_),
    .A(net74),
    .B(net6));
 sg13g2_o21ai_1 _3626_ (.B1(_1649_),
    .Y(_0006_),
    .A1(_1647_),
    .A2(_1589_));
 sg13g2_mux2_1 _3627_ (.A0(_1562_),
    .A1(net7),
    .S(net74),
    .X(_0007_));
 sg13g2_nor2_2 _3628_ (.A(_1577_),
    .B(_1586_),
    .Y(_1650_));
 sg13g2_buf_2 _3629_ (.A(\i_project.controller_0.h[4] ),
    .X(_1651_));
 sg13g2_buf_1 _3630_ (.A(_1651_),
    .X(_1652_));
 sg13g2_inv_1 _3631_ (.Y(_1653_),
    .A(net66));
 sg13g2_buf_2 _3632_ (.A(\i_project.controller_0.h[5] ),
    .X(_1654_));
 sg13g2_buf_1 _3633_ (.A(_1654_),
    .X(_1655_));
 sg13g2_nand2_1 _3634_ (.Y(_1656_),
    .A(_1653_),
    .B(net65));
 sg13g2_buf_1 _3635_ (.A(\i_project.controller_0.h[9] ),
    .X(_1657_));
 sg13g2_buf_2 _3636_ (.A(\i_project.controller_0.h[8] ),
    .X(_1658_));
 sg13g2_inv_1 _3637_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_nor2_1 _3638_ (.A(_1657_),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_inv_1 _3639_ (.Y(_1661_),
    .A(_1660_));
 sg13g2_buf_2 _3640_ (.A(\i_project.controller_0.h[6] ),
    .X(_1662_));
 sg13g2_buf_1 _3641_ (.A(\i_project.controller_0.h[7] ),
    .X(_1663_));
 sg13g2_inv_1 _3642_ (.Y(_1664_),
    .A(_1663_));
 sg13g2_nor2_1 _3643_ (.A(_1662_),
    .B(_1664_),
    .Y(_1665_));
 sg13g2_buf_1 _3644_ (.A(\i_project.controller_0.h[0] ),
    .X(_1666_));
 sg13g2_buf_1 _3645_ (.A(_1666_),
    .X(_1667_));
 sg13g2_buf_1 _3646_ (.A(\i_project.controller_0.h[1] ),
    .X(_1668_));
 sg13g2_inv_1 _3647_ (.Y(_1669_),
    .A(net73));
 sg13g2_nor2_1 _3648_ (.A(_1667_),
    .B(_1669_),
    .Y(_1670_));
 sg13g2_buf_1 _3649_ (.A(\i_project.controller_0.h[2] ),
    .X(_1671_));
 sg13g2_buf_1 _3650_ (.A(_1671_),
    .X(_1672_));
 sg13g2_buf_1 _3651_ (.A(\i_project.controller_0.h[3] ),
    .X(_1673_));
 sg13g2_buf_1 _3652_ (.A(_1673_),
    .X(_1674_));
 sg13g2_nor2_1 _3653_ (.A(net63),
    .B(net62),
    .Y(_1675_));
 sg13g2_inv_1 _3654_ (.Y(_1676_),
    .A(_0025_));
 sg13g2_nand4_1 _3655_ (.B(_1670_),
    .C(_1675_),
    .A(_1665_),
    .Y(_1677_),
    .D(_1676_));
 sg13g2_nor3_1 _3656_ (.A(_1656_),
    .B(_1661_),
    .C(_1677_),
    .Y(_1678_));
 sg13g2_inv_1 _3657_ (.Y(_1679_),
    .A(_1657_));
 sg13g2_nor2_1 _3658_ (.A(_1658_),
    .B(_1679_),
    .Y(_1680_));
 sg13g2_inv_1 _3659_ (.Y(_1681_),
    .A(_1680_));
 sg13g2_nor2_1 _3660_ (.A(_1668_),
    .B(net64),
    .Y(_1682_));
 sg13g2_nand2_1 _3661_ (.Y(_1683_),
    .A(_1675_),
    .B(_1682_));
 sg13g2_buf_1 _3662_ (.A(_1662_),
    .X(_1684_));
 sg13g2_buf_1 _3663_ (.A(_1663_),
    .X(_1685_));
 sg13g2_nand4_1 _3664_ (.B(net66),
    .C(net61),
    .A(net65),
    .Y(_1686_),
    .D(net60));
 sg13g2_nor4_1 _3665_ (.A(_1676_),
    .B(_1681_),
    .C(_1683_),
    .D(_1686_),
    .Y(_1687_));
 sg13g2_nor2_1 _3666_ (.A(net65),
    .B(_1653_),
    .Y(_1688_));
 sg13g2_nand2_1 _3667_ (.Y(_1689_),
    .A(_1665_),
    .B(_1688_));
 sg13g2_nor3_1 _3668_ (.A(_1681_),
    .B(_1683_),
    .C(_1689_),
    .Y(_1690_));
 sg13g2_nand2_1 _3669_ (.Y(_1691_),
    .A(net63),
    .B(net62));
 sg13g2_inv_1 _3670_ (.Y(_1692_),
    .A(_1682_));
 sg13g2_nor4_1 _3671_ (.A(_0025_),
    .B(_1691_),
    .C(_1692_),
    .D(_1661_),
    .Y(_1693_));
 sg13g2_inv_1 _3672_ (.Y(_1694_),
    .A(net65));
 sg13g2_inv_1 _3673_ (.Y(_1695_),
    .A(_1662_));
 sg13g2_nor4_1 _3674_ (.A(_1685_),
    .B(_1694_),
    .C(_1653_),
    .D(_1695_),
    .Y(_1696_));
 sg13g2_a221oi_1 _3675_ (.B2(_1696_),
    .C1(\i_project.controller_0.vga_sync.hsync ),
    .B1(_1693_),
    .A1(_1690_),
    .Y(_1697_),
    .A2(_0025_));
 sg13g2_nor4_1 _3676_ (.A(_1650_),
    .B(_1678_),
    .C(_1687_),
    .D(_1697_),
    .Y(_0123_));
 sg13g2_buf_2 _3677_ (.A(\i_project.controller_0.v[8] ),
    .X(_1698_));
 sg13g2_inv_1 _3678_ (.Y(_1699_),
    .A(_1698_));
 sg13g2_buf_1 _3679_ (.A(\i_project.controller_0.v[9] ),
    .X(_1700_));
 sg13g2_buf_1 _3680_ (.A(\i_project.controller_0.v[7] ),
    .X(_1701_));
 sg13g2_buf_1 _3681_ (.A(\i_project.controller_0.v[6] ),
    .X(_1702_));
 sg13g2_nand2_1 _3682_ (.Y(_1703_),
    .A(_1701_),
    .B(net72));
 sg13g2_inv_1 _3683_ (.Y(_1704_),
    .A(_1703_));
 sg13g2_buf_8 _3684_ (.A(\i_project.controller_0.v[4] ),
    .X(_1705_));
 sg13g2_buf_8 _3685_ (.A(\i_project.controller_0.v[5] ),
    .X(_1706_));
 sg13g2_inv_1 _3686_ (.Y(_1707_),
    .A(_1706_));
 sg13g2_nor2_1 _3687_ (.A(_1705_),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_nand2_1 _3688_ (.Y(_1709_),
    .A(_1704_),
    .B(_1708_));
 sg13g2_nor3_1 _3689_ (.A(_1699_),
    .B(_1700_),
    .C(_1709_),
    .Y(_1710_));
 sg13g2_buf_1 _3690_ (.A(\i_project.controller_0.vga_sync.mode ),
    .X(_1711_));
 sg13g2_buf_8 _3691_ (.A(\i_project.controller_0.v[2] ),
    .X(_1712_));
 sg13g2_buf_8 _3692_ (.A(\i_project.controller_0.v[3] ),
    .X(_1713_));
 sg13g2_nand2_1 _3693_ (.Y(_1714_),
    .A(_1712_),
    .B(_1713_));
 sg13g2_buf_8 _3694_ (.A(\i_project.controller_0.v[0] ),
    .X(_1715_));
 sg13g2_buf_8 _3695_ (.A(\i_project.controller_0.v[1] ),
    .X(_1716_));
 sg13g2_nor2_1 _3696_ (.A(_1715_),
    .B(_1716_),
    .Y(_1717_));
 sg13g2_inv_1 _3697_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_nor3_1 _3698_ (.A(net71),
    .B(_1714_),
    .C(_1718_),
    .Y(_1719_));
 sg13g2_nand2_1 _3699_ (.Y(_1720_),
    .A(_1710_),
    .B(_1719_));
 sg13g2_inv_2 _3700_ (.Y(_1721_),
    .A(_1712_));
 sg13g2_nand2_1 _3701_ (.Y(_1722_),
    .A(_1721_),
    .B(_1713_));
 sg13g2_inv_1 _3702_ (.Y(_1723_),
    .A(_1701_));
 sg13g2_nor2_1 _3703_ (.A(net72),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_nor2_1 _3704_ (.A(_1705_),
    .B(_1706_),
    .Y(_1725_));
 sg13g2_nand2_1 _3705_ (.Y(_1726_),
    .A(_1724_),
    .B(_1725_));
 sg13g2_nor3_1 _3706_ (.A(_1718_),
    .B(_1722_),
    .C(_1726_),
    .Y(_1727_));
 sg13g2_inv_1 _3707_ (.Y(_1728_),
    .A(net71));
 sg13g2_inv_1 _3708_ (.Y(_1729_),
    .A(_1700_));
 sg13g2_nor3_1 _3709_ (.A(_1728_),
    .B(_1699_),
    .C(_1729_),
    .Y(_1730_));
 sg13g2_nand2_1 _3710_ (.Y(_1731_),
    .A(_1727_),
    .B(_1730_));
 sg13g2_inv_1 _3711_ (.Y(_1732_),
    .A(_1650_));
 sg13g2_nand3_1 _3712_ (.B(_1731_),
    .C(_1732_),
    .A(_1720_),
    .Y(_1733_));
 sg13g2_inv_1 _3713_ (.Y(_1734_),
    .A(_1716_));
 sg13g2_nor4_1 _3714_ (.A(net71),
    .B(_1715_),
    .C(_1734_),
    .D(_1722_),
    .Y(_1735_));
 sg13g2_and3_1 _3715_ (.X(_1736_),
    .A(_1730_),
    .B(_1715_),
    .C(_1734_));
 sg13g2_nor3_1 _3716_ (.A(_1721_),
    .B(_1713_),
    .C(_1726_),
    .Y(_1737_));
 sg13g2_a221oi_1 _3717_ (.B2(_1737_),
    .C1(\i_project.controller_0.vga_sync.vsync ),
    .B1(_1736_),
    .A1(_1710_),
    .Y(_1738_),
    .A2(_1735_));
 sg13g2_nor2_1 _3718_ (.A(_1733_),
    .B(_1738_),
    .Y(_0134_));
 sg13g2_inv_1 _3719_ (.Y(_1739_),
    .A(\i_project.controller_0.voffset[0] ));
 sg13g2_o21ai_1 _3720_ (.B1(_1658_),
    .Y(_1740_),
    .A1(net61),
    .A2(net60));
 sg13g2_inv_1 _3721_ (.Y(_1741_),
    .A(_0023_));
 sg13g2_o21ai_1 _3722_ (.B1(_1655_),
    .Y(_1742_),
    .A1(net66),
    .A2(_1741_));
 sg13g2_nor3_1 _3723_ (.A(_1695_),
    .B(net60),
    .C(_1661_),
    .Y(_1743_));
 sg13g2_a22oi_1 _3724_ (.Y(_1744_),
    .B1(_1742_),
    .B2(_1743_),
    .A2(_1740_),
    .A1(_1679_));
 sg13g2_inv_1 _3725_ (.Y(_1745_),
    .A(_1673_));
 sg13g2_nor2_1 _3726_ (.A(_1672_),
    .B(_1745_),
    .Y(_1746_));
 sg13g2_nor2_1 _3727_ (.A(_1656_),
    .B(_1692_),
    .Y(_1747_));
 sg13g2_nand3_1 _3728_ (.B(_1746_),
    .C(_1747_),
    .A(_1743_),
    .Y(_1748_));
 sg13g2_nand2_1 _3729_ (.Y(_1749_),
    .A(_1748_),
    .B(net71));
 sg13g2_inv_1 _3730_ (.Y(_1750_),
    .A(_0026_));
 sg13g2_nand3_1 _3731_ (.B(_1694_),
    .C(_1653_),
    .A(_1665_),
    .Y(_1751_));
 sg13g2_nor2_1 _3732_ (.A(_1683_),
    .B(_1751_),
    .Y(_1752_));
 sg13g2_nor3_1 _3733_ (.A(_1658_),
    .B(_1750_),
    .C(_1752_),
    .Y(_1753_));
 sg13g2_o21ai_1 _3734_ (.B1(_1728_),
    .Y(_1754_),
    .A1(_1679_),
    .A2(_1753_));
 sg13g2_o21ai_1 _3735_ (.B1(_1754_),
    .Y(_1755_),
    .A1(_1744_),
    .A2(_1749_));
 sg13g2_xor2_1 _3736_ (.B(\i_project.controller_0.grey_pass[14] ),
    .A(\i_project.controller_0.mode[2] ),
    .X(_1756_));
 sg13g2_buf_2 _3737_ (.A(\i_project.controller_0.mode[1] ),
    .X(_1757_));
 sg13g2_xor2_1 _3738_ (.B(\i_project.controller_0.grey_pass[13] ),
    .A(_1757_),
    .X(_1758_));
 sg13g2_nor2_1 _3739_ (.A(_1756_),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_buf_1 _3740_ (.A(\i_project.controller_0.mode[0] ),
    .X(_1760_));
 sg13g2_xnor2_1 _3741_ (.Y(_1761_),
    .A(_1760_),
    .B(\i_project.controller_0.grey_pass[12] ));
 sg13g2_inv_1 _3742_ (.Y(_1762_),
    .A(_0027_));
 sg13g2_nor3_1 _3743_ (.A(_1757_),
    .B(_1760_),
    .C(_1762_),
    .Y(_1763_));
 sg13g2_buf_2 _3744_ (.A(_1763_),
    .X(_1764_));
 sg13g2_buf_1 _3745_ (.A(_1764_),
    .X(_1765_));
 sg13g2_a21oi_1 _3746_ (.A1(_1759_),
    .A2(_1761_),
    .Y(_1766_),
    .B1(net49));
 sg13g2_nand2b_1 _3747_ (.Y(_1767_),
    .B(_1766_),
    .A_N(_1755_));
 sg13g2_nand2_2 _3748_ (.Y(_1768_),
    .A(_1767_),
    .B(_1577_));
 sg13g2_inv_2 _3749_ (.Y(_1769_),
    .A(_1768_));
 sg13g2_nand2b_1 _3750_ (.Y(_1770_),
    .B(net68),
    .A_N(_1761_));
 sg13g2_inv_1 _3751_ (.Y(_1771_),
    .A(\i_project.controller_0.mode[2] ));
 sg13g2_nor3_1 _3752_ (.A(_1757_),
    .B(_1577_),
    .C(_1771_),
    .Y(_1772_));
 sg13g2_nand2_1 _3753_ (.Y(_1773_),
    .A(_1772_),
    .B(_0016_));
 sg13g2_nor2b_2 _3754_ (.A(_1769_),
    .B_N(_1773_),
    .Y(_1774_));
 sg13g2_a22oi_1 _3755_ (.Y(_0135_),
    .B1(_1770_),
    .B2(_1774_),
    .A2(_1769_),
    .A1(_1739_));
 sg13g2_a22oi_1 _3756_ (.Y(_1775_),
    .B1(net68),
    .B2(_1758_),
    .A2(_0015_),
    .A1(_1772_));
 sg13g2_buf_8 _3757_ (.A(\i_project.controller_0.voffset[1] ),
    .X(_1776_));
 sg13g2_nor2_1 _3758_ (.A(_1776_),
    .B(_1768_),
    .Y(_1777_));
 sg13g2_a21oi_1 _3759_ (.A1(_1768_),
    .A2(_1775_),
    .Y(_0136_),
    .B1(_1777_));
 sg13g2_inv_1 _3760_ (.Y(_1778_),
    .A(\i_project.controller_0.voffset[2] ));
 sg13g2_nand2_1 _3761_ (.Y(_1779_),
    .A(_1756_),
    .B(net68));
 sg13g2_a22oi_1 _3762_ (.Y(_0137_),
    .B1(_1779_),
    .B2(_1774_),
    .A2(_1769_),
    .A1(_1778_));
 sg13g2_inv_1 _3763_ (.Y(_1780_),
    .A(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _3764_ (.Y(_1781_),
    .A(_1772_),
    .B(_0144_));
 sg13g2_o21ai_1 _3765_ (.B1(_1781_),
    .Y(_0138_),
    .A1(_1780_),
    .A2(_1768_));
 sg13g2_inv_1 _3766_ (.Y(_1782_),
    .A(\i_project.controller_0.voffset[4] ));
 sg13g2_o21ai_1 _3767_ (.B1(_1773_),
    .Y(_0139_),
    .A1(_1782_),
    .A2(_1768_));
 sg13g2_buf_8 _3768_ (.A(\i_project.controller_0.voffset[5] ),
    .X(_1783_));
 sg13g2_inv_1 _3769_ (.Y(_1784_),
    .A(_1783_));
 sg13g2_buf_1 _3770_ (.A(_1578_),
    .X(_1785_));
 sg13g2_nand2_1 _3771_ (.Y(_1786_),
    .A(net54),
    .B(\i_project.controller_0.grey_pass[10] ));
 sg13g2_a22oi_1 _3772_ (.Y(_0140_),
    .B1(_1786_),
    .B2(_1774_),
    .A2(_1769_),
    .A1(_1784_));
 sg13g2_inv_1 _3773_ (.Y(_1787_),
    .A(\i_project.controller_0.voffset[6] ));
 sg13g2_nand2_1 _3774_ (.Y(_1788_),
    .A(net54),
    .B(\i_project.controller_0.grey_pass[11] ));
 sg13g2_a22oi_1 _3775_ (.Y(_0141_),
    .B1(_1788_),
    .B2(_1774_),
    .A2(_1769_),
    .A1(_1787_));
 sg13g2_inv_1 _3776_ (.Y(_1789_),
    .A(_1577_));
 sg13g2_inv_1 _3777_ (.Y(_1790_),
    .A(\i_project.controller_0.grey_pass[15] ));
 sg13g2_nor3_1 _3778_ (.A(_1789_),
    .B(_1790_),
    .C(_1767_),
    .Y(_1791_));
 sg13g2_a21o_1 _3779_ (.A2(_1769_),
    .A1(\i_project.controller_0.voffset[7] ),
    .B1(_1791_),
    .X(_0142_));
 sg13g2_inv_1 _3780_ (.Y(_1792_),
    .A(_1760_));
 sg13g2_nor2_1 _3781_ (.A(net54),
    .B(\i_project.controller_0.grey_pass[12] ),
    .Y(_1793_));
 sg13g2_a21oi_1 _3782_ (.A1(_1792_),
    .A2(net54),
    .Y(_0097_),
    .B1(_1793_));
 sg13g2_inv_1 _3783_ (.Y(_1794_),
    .A(_1757_));
 sg13g2_nor2_1 _3784_ (.A(_1785_),
    .B(\i_project.controller_0.grey_pass[13] ),
    .Y(_1795_));
 sg13g2_a21oi_1 _3785_ (.A1(_1794_),
    .A2(_1785_),
    .Y(_0098_),
    .B1(_1795_));
 sg13g2_nor2_1 _3786_ (.A(net54),
    .B(\i_project.controller_0.grey_pass[14] ),
    .Y(_1796_));
 sg13g2_a21oi_1 _3787_ (.A1(_1771_),
    .A2(net54),
    .Y(_0099_),
    .B1(_1796_));
 sg13g2_nand2_1 _3788_ (.Y(_1797_),
    .A(net71),
    .B(net54));
 sg13g2_o21ai_1 _3789_ (.B1(_1797_),
    .Y(_0100_),
    .A1(net54),
    .A2(_1790_));
 sg13g2_buf_1 _3790_ (.A(\dither_threshold[0] ),
    .X(_1798_));
 sg13g2_inv_1 _3791_ (.Y(_1799_),
    .A(_1798_));
 sg13g2_buf_2 _3792_ (.A(_0022_),
    .X(_1800_));
 sg13g2_buf_2 _3793_ (.A(\dither_threshold[1] ),
    .X(_1801_));
 sg13g2_inv_1 _3794_ (.Y(_1802_),
    .A(_1801_));
 sg13g2_a21oi_1 _3795_ (.A1(_1800_),
    .A2(_1798_),
    .Y(_1803_),
    .B1(_1802_));
 sg13g2_inv_1 _3796_ (.Y(_1804_),
    .A(\dither_threshold[5] ));
 sg13g2_inv_1 _3797_ (.Y(_1805_),
    .A(\dither_threshold[3] ));
 sg13g2_buf_1 _3798_ (.A(\dither_threshold[4] ),
    .X(_1806_));
 sg13g2_inv_1 _3799_ (.Y(_1807_),
    .A(_1806_));
 sg13g2_buf_2 _3800_ (.A(\dither_threshold[2] ),
    .X(_1808_));
 sg13g2_inv_2 _3801_ (.Y(_1809_),
    .A(_1808_));
 sg13g2_nand4_1 _3802_ (.B(_1805_),
    .C(_1807_),
    .A(_1804_),
    .Y(_1810_),
    .D(_1809_));
 sg13g2_o21ai_1 _3803_ (.B1(\dither_threshold[6] ),
    .Y(_1811_),
    .A1(_1803_),
    .A2(_1810_));
 sg13g2_buf_2 _3804_ (.A(_1811_),
    .X(_1812_));
 sg13g2_inv_2 _3805_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_xor2_1 _3806_ (.B(\i_project.controller_0.vga_sync.vsync ),
    .A(net71),
    .X(_1814_));
 sg13g2_inv_1 _3807_ (.Y(\i_project.controller_0.vga_sync.o_vsync ),
    .A(_1814_));
 sg13g2_nand2_1 _3808_ (.Y(_1815_),
    .A(\i_project.controller_0.vga_sync.o_vsync ),
    .B(\i_project.controller_0.grey_pass[15] ));
 sg13g2_nand2_1 _3809_ (.Y(_1816_),
    .A(_1814_),
    .B(_1790_));
 sg13g2_nand3_1 _3810_ (.B(_1586_),
    .C(_1816_),
    .A(_1815_),
    .Y(_1817_));
 sg13g2_buf_1 _3811_ (.A(_1817_),
    .X(_1818_));
 sg13g2_inv_1 _3812_ (.Y(_1819_),
    .A(_1818_));
 sg13g2_o21ai_1 _3813_ (.B1(_1819_),
    .Y(_1820_),
    .A1(_1799_),
    .A2(_1813_));
 sg13g2_a21oi_1 _3814_ (.A1(_1799_),
    .A2(_1813_),
    .Y(_0090_),
    .B1(_1820_));
 sg13g2_inv_1 _3815_ (.Y(_1821_),
    .A(_0031_));
 sg13g2_nor2_1 _3816_ (.A(_1801_),
    .B(_1798_),
    .Y(_1822_));
 sg13g2_nor2_1 _3817_ (.A(_1822_),
    .B(_1813_),
    .Y(_1823_));
 sg13g2_nand2_1 _3818_ (.Y(_1824_),
    .A(_1801_),
    .B(_1798_));
 sg13g2_a221oi_1 _3819_ (.B2(_1824_),
    .C1(_1818_),
    .B1(_1823_),
    .A1(_1821_),
    .Y(_0091_),
    .A2(_1813_));
 sg13g2_a21oi_1 _3820_ (.A1(_1802_),
    .A2(_1813_),
    .Y(_1825_),
    .B1(_1823_));
 sg13g2_xnor2_1 _3821_ (.Y(_1826_),
    .A(_1809_),
    .B(_1825_));
 sg13g2_nor2_1 _3822_ (.A(_1818_),
    .B(_1826_),
    .Y(_0092_));
 sg13g2_inv_2 _3823_ (.Y(_1827_),
    .A(_0032_));
 sg13g2_a21oi_1 _3824_ (.A1(_1802_),
    .A2(_1800_),
    .Y(_1828_),
    .B1(_1809_));
 sg13g2_xnor2_1 _3825_ (.Y(_1829_),
    .A(_1827_),
    .B(_1828_));
 sg13g2_o21ai_1 _3826_ (.B1(\dither_threshold[3] ),
    .Y(_1830_),
    .A1(_1808_),
    .A2(_1801_));
 sg13g2_nor2_1 _3827_ (.A(_1808_),
    .B(_1801_),
    .Y(_1831_));
 sg13g2_nand2_1 _3828_ (.Y(_1832_),
    .A(_1831_),
    .B(_1805_));
 sg13g2_nand2_1 _3829_ (.Y(_1833_),
    .A(_1830_),
    .B(_1832_));
 sg13g2_o21ai_1 _3830_ (.B1(_1819_),
    .Y(_1834_),
    .A1(_1812_),
    .A2(_1833_));
 sg13g2_a21oi_1 _3831_ (.A1(_1812_),
    .A2(_1829_),
    .Y(_0093_),
    .B1(_1834_));
 sg13g2_buf_2 _3832_ (.A(_0033_),
    .X(_1835_));
 sg13g2_nor3_2 _3833_ (.A(_1805_),
    .B(_1809_),
    .C(_1822_),
    .Y(_1836_));
 sg13g2_xnor2_1 _3834_ (.Y(_1837_),
    .A(_1835_),
    .B(_1836_));
 sg13g2_xnor2_1 _3835_ (.Y(_1838_),
    .A(_1806_),
    .B(_1832_));
 sg13g2_o21ai_1 _3836_ (.B1(_1819_),
    .Y(_1839_),
    .A1(_1838_),
    .A2(_1812_));
 sg13g2_a21oi_1 _3837_ (.A1(_1812_),
    .A2(_1837_),
    .Y(_0094_),
    .B1(_1839_));
 sg13g2_buf_2 _3838_ (.A(_0034_),
    .X(_1840_));
 sg13g2_inv_1 _3839_ (.Y(_1841_),
    .A(_1835_));
 sg13g2_a21oi_1 _3840_ (.A1(_1836_),
    .A2(_1807_),
    .Y(_1842_),
    .B1(_1841_));
 sg13g2_xnor2_1 _3841_ (.Y(_1843_),
    .A(_1840_),
    .B(_1842_));
 sg13g2_o21ai_1 _3842_ (.B1(\dither_threshold[5] ),
    .Y(_1844_),
    .A1(_1806_),
    .A2(_1832_));
 sg13g2_a21o_1 _3843_ (.A2(_1844_),
    .A1(_1813_),
    .B1(_1818_),
    .X(_1845_));
 sg13g2_a21oi_1 _3844_ (.A1(_1843_),
    .A2(_1812_),
    .Y(_0095_),
    .B1(_1845_));
 sg13g2_buf_1 _3845_ (.A(_0035_),
    .X(_1846_));
 sg13g2_o21ai_1 _3846_ (.B1(\dither_threshold[5] ),
    .Y(_1847_),
    .A1(_1806_),
    .A2(_1836_));
 sg13g2_nor2b_1 _3847_ (.A(_1813_),
    .B_N(_1847_),
    .Y(_1848_));
 sg13g2_o21ai_1 _3848_ (.B1(_1819_),
    .Y(_1849_),
    .A1(_1846_),
    .A2(_1848_));
 sg13g2_a21oi_1 _3849_ (.A1(_1846_),
    .A2(_1848_),
    .Y(_0096_),
    .B1(_1849_));
 sg13g2_inv_1 _3850_ (.Y(_1850_),
    .A(_0054_));
 sg13g2_nand2_1 _3851_ (.Y(_1851_),
    .A(net73),
    .B(_1667_));
 sg13g2_inv_1 _3852_ (.Y(_1852_),
    .A(_0024_));
 sg13g2_nand3_1 _3853_ (.B(_1741_),
    .C(_1852_),
    .A(_1688_),
    .Y(_1853_));
 sg13g2_nand2_1 _3854_ (.Y(_1854_),
    .A(_1672_),
    .B(_1657_));
 sg13g2_inv_1 _3855_ (.Y(_1855_),
    .A(_1854_));
 sg13g2_nor2_1 _3856_ (.A(net61),
    .B(net60),
    .Y(_1856_));
 sg13g2_a21oi_1 _3857_ (.A1(_1855_),
    .A2(_1856_),
    .Y(_1857_),
    .B1(net71));
 sg13g2_nor3_1 _3858_ (.A(_1851_),
    .B(_1853_),
    .C(_1857_),
    .Y(_1858_));
 sg13g2_inv_1 _3859_ (.Y(_1859_),
    .A(net63));
 sg13g2_nand4_1 _3860_ (.B(_1679_),
    .C(net61),
    .A(_1859_),
    .Y(_1860_),
    .D(net60));
 sg13g2_nand2_1 _3861_ (.Y(_1861_),
    .A(_1860_),
    .B(net71));
 sg13g2_nand2_1 _3862_ (.Y(_1862_),
    .A(_1858_),
    .B(_1861_));
 sg13g2_buf_2 _3863_ (.A(_1862_),
    .X(_1863_));
 sg13g2_nand2_1 _3864_ (.Y(_1864_),
    .A(_1863_),
    .B(_1732_));
 sg13g2_buf_1 _3865_ (.A(_1864_),
    .X(_1865_));
 sg13g2_nor2_1 _3866_ (.A(_1850_),
    .B(net21),
    .Y(_0113_));
 sg13g2_inv_1 _3867_ (.Y(_1866_),
    .A(_1851_));
 sg13g2_nor3_1 _3868_ (.A(_1682_),
    .B(_1866_),
    .C(net21),
    .Y(_0114_));
 sg13g2_nor2_1 _3869_ (.A(net63),
    .B(_1866_),
    .Y(_1867_));
 sg13g2_nor2_1 _3870_ (.A(_1859_),
    .B(_1851_),
    .Y(_1868_));
 sg13g2_nor3_1 _3871_ (.A(_1867_),
    .B(_1868_),
    .C(net21),
    .Y(_0115_));
 sg13g2_nor2_1 _3872_ (.A(_1674_),
    .B(_1868_),
    .Y(_1869_));
 sg13g2_nor2_1 _3873_ (.A(_1691_),
    .B(_1851_),
    .Y(_1870_));
 sg13g2_nor3_1 _3874_ (.A(_1869_),
    .B(_1870_),
    .C(net21),
    .Y(_0116_));
 sg13g2_nor2_1 _3875_ (.A(_1652_),
    .B(_1870_),
    .Y(_1871_));
 sg13g2_nand2_1 _3876_ (.Y(_1872_),
    .A(_1870_),
    .B(_1652_));
 sg13g2_inv_1 _3877_ (.Y(_1873_),
    .A(_1872_));
 sg13g2_nor3_1 _3878_ (.A(_1871_),
    .B(_1873_),
    .C(net21),
    .Y(_0117_));
 sg13g2_nor2_1 _3879_ (.A(_1655_),
    .B(_1873_),
    .Y(_1874_));
 sg13g2_nor2_1 _3880_ (.A(_1694_),
    .B(_1872_),
    .Y(_1875_));
 sg13g2_nor3_1 _3881_ (.A(_1874_),
    .B(_1875_),
    .C(net21),
    .Y(_0118_));
 sg13g2_nor2_1 _3882_ (.A(net61),
    .B(_1875_),
    .Y(_1876_));
 sg13g2_nand2_1 _3883_ (.Y(_1877_),
    .A(_1875_),
    .B(_1684_));
 sg13g2_inv_1 _3884_ (.Y(_1878_),
    .A(_1877_));
 sg13g2_nor3_1 _3885_ (.A(_1876_),
    .B(_1878_),
    .C(net21),
    .Y(_0119_));
 sg13g2_nor2_1 _3886_ (.A(_1685_),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_nor2_1 _3887_ (.A(_1664_),
    .B(_1877_),
    .Y(_1880_));
 sg13g2_nor3_1 _3888_ (.A(_1879_),
    .B(_1880_),
    .C(net21),
    .Y(_0120_));
 sg13g2_nor2_1 _3889_ (.A(_1658_),
    .B(_1880_),
    .Y(_1881_));
 sg13g2_nand2_1 _3890_ (.Y(_1882_),
    .A(_1880_),
    .B(_1658_));
 sg13g2_inv_1 _3891_ (.Y(_1883_),
    .A(_1882_));
 sg13g2_nor3_1 _3892_ (.A(_1864_),
    .B(_1881_),
    .C(_1883_),
    .Y(_0121_));
 sg13g2_nor2_1 _3893_ (.A(_1679_),
    .B(_1882_),
    .Y(_1884_));
 sg13g2_nor2_1 _3894_ (.A(_1657_),
    .B(_1883_),
    .Y(_1885_));
 sg13g2_nor3_1 _3895_ (.A(_1864_),
    .B(_1884_),
    .C(_1885_),
    .Y(_0122_));
 sg13g2_inv_1 _3896_ (.Y(_1886_),
    .A(_1715_));
 sg13g2_nor2_1 _3897_ (.A(_1886_),
    .B(_1863_),
    .Y(_1887_));
 sg13g2_nand3_1 _3898_ (.B(_1711_),
    .C(_1698_),
    .A(_1708_),
    .Y(_1888_));
 sg13g2_nor2_1 _3899_ (.A(_1712_),
    .B(_1713_),
    .Y(_1889_));
 sg13g2_nand4_1 _3900_ (.B(_1889_),
    .C(_1715_),
    .A(_1724_),
    .Y(_1890_),
    .D(_1716_));
 sg13g2_nor3_1 _3901_ (.A(_1701_),
    .B(net72),
    .C(_1698_),
    .Y(_1891_));
 sg13g2_nand3_1 _3902_ (.B(_1725_),
    .C(_1891_),
    .A(_1719_),
    .Y(_1892_));
 sg13g2_o21ai_1 _3903_ (.B1(_1892_),
    .Y(_1893_),
    .A1(_1888_),
    .A2(_1890_));
 sg13g2_inv_1 _3904_ (.Y(_1894_),
    .A(_0028_));
 sg13g2_nand2_1 _3905_ (.Y(_1895_),
    .A(_1893_),
    .B(_1894_));
 sg13g2_inv_1 _3906_ (.Y(_1896_),
    .A(_1863_));
 sg13g2_a21oi_1 _3907_ (.A1(_1895_),
    .A2(_1896_),
    .Y(_1897_),
    .B1(_1715_));
 sg13g2_nor3_1 _3908_ (.A(_1650_),
    .B(_1887_),
    .C(_1897_),
    .Y(_0124_));
 sg13g2_nor2_1 _3909_ (.A(_1716_),
    .B(_1887_),
    .Y(_1898_));
 sg13g2_inv_1 _3910_ (.Y(_1899_),
    .A(_1887_));
 sg13g2_nor2_1 _3911_ (.A(_1734_),
    .B(_1899_),
    .Y(_1900_));
 sg13g2_nor3_1 _3912_ (.A(_1650_),
    .B(_1898_),
    .C(_1900_),
    .Y(_0125_));
 sg13g2_nor3_1 _3913_ (.A(_1734_),
    .B(_1721_),
    .C(_1899_),
    .Y(_1901_));
 sg13g2_nor2_1 _3914_ (.A(_1712_),
    .B(_1900_),
    .Y(_1902_));
 sg13g2_nor2_2 _3915_ (.A(_1863_),
    .B(_1895_),
    .Y(_1903_));
 sg13g2_inv_1 _3916_ (.Y(_1904_),
    .A(_1903_));
 sg13g2_nand2_1 _3917_ (.Y(_1905_),
    .A(_1904_),
    .B(_1732_));
 sg13g2_nor3_1 _3918_ (.A(_1901_),
    .B(_1902_),
    .C(_1905_),
    .Y(_0126_));
 sg13g2_nor3_1 _3919_ (.A(_1886_),
    .B(_1734_),
    .C(_1714_),
    .Y(_1906_));
 sg13g2_inv_1 _3920_ (.Y(_1907_),
    .A(_1906_));
 sg13g2_nor2_1 _3921_ (.A(_1907_),
    .B(_1863_),
    .Y(_1908_));
 sg13g2_nor2_1 _3922_ (.A(_1713_),
    .B(_1901_),
    .Y(_1909_));
 sg13g2_nor3_1 _3923_ (.A(_1908_),
    .B(_1905_),
    .C(_1909_),
    .Y(_0127_));
 sg13g2_xnor2_1 _3924_ (.Y(_1910_),
    .A(_1705_),
    .B(_1908_));
 sg13g2_nor2_1 _3925_ (.A(_1650_),
    .B(_1910_),
    .Y(_0128_));
 sg13g2_and3_1 _3926_ (.X(_1911_),
    .A(_1895_),
    .B(_1732_),
    .C(_1896_));
 sg13g2_buf_1 _3927_ (.A(_1911_),
    .X(_1912_));
 sg13g2_nor2b_1 _3928_ (.A(_1907_),
    .B_N(_1705_),
    .Y(_1913_));
 sg13g2_xnor2_1 _3929_ (.Y(_1914_),
    .A(_0029_),
    .B(_1913_));
 sg13g2_nand2_1 _3930_ (.Y(_1915_),
    .A(_1912_),
    .B(_1914_));
 sg13g2_o21ai_1 _3931_ (.B1(_1915_),
    .Y(_0129_),
    .A1(_1707_),
    .A2(_1865_));
 sg13g2_nand2_1 _3932_ (.Y(_1916_),
    .A(_1913_),
    .B(_1706_));
 sg13g2_nor2_1 _3933_ (.A(_1916_),
    .B(_1863_),
    .Y(_1917_));
 sg13g2_xnor2_1 _3934_ (.Y(_1918_),
    .A(net72),
    .B(_1917_));
 sg13g2_nor2_1 _3935_ (.A(_1650_),
    .B(_1918_),
    .Y(_0130_));
 sg13g2_nand2_1 _3936_ (.Y(_1919_),
    .A(_1917_),
    .B(_1702_));
 sg13g2_nor2_2 _3937_ (.A(_1703_),
    .B(_1916_),
    .Y(_1920_));
 sg13g2_a221oi_1 _3938_ (.B2(_1920_),
    .C1(_1905_),
    .B1(_1896_),
    .A1(_1723_),
    .Y(_0131_),
    .A2(_1919_));
 sg13g2_xnor2_1 _3939_ (.Y(_1921_),
    .A(_0030_),
    .B(_1920_));
 sg13g2_nand2_1 _3940_ (.Y(_1922_),
    .A(_1912_),
    .B(_1921_));
 sg13g2_o21ai_1 _3941_ (.B1(_1922_),
    .Y(_0132_),
    .A1(_1699_),
    .A2(_1865_));
 sg13g2_a21o_1 _3942_ (.A2(_1698_),
    .A1(_1920_),
    .B1(_1894_),
    .X(_1923_));
 sg13g2_nand3_1 _3943_ (.B(_1698_),
    .C(_1894_),
    .A(_1920_),
    .Y(_1924_));
 sg13g2_nand3_1 _3944_ (.B(_1923_),
    .C(_1924_),
    .A(_1912_),
    .Y(_1925_));
 sg13g2_o21ai_1 _3945_ (.B1(_1925_),
    .Y(_0133_),
    .A1(_1729_),
    .A2(_1864_));
 sg13g2_and2_1 _3946_ (.A(_0004_),
    .B(_0003_),
    .X(_0057_));
 sg13g2_nand2_1 _3947_ (.Y(_1926_),
    .A(_1586_),
    .B(_0055_));
 sg13g2_inv_1 _3948_ (.Y(_0058_),
    .A(_1926_));
 sg13g2_buf_1 _3949_ (.A(net67),
    .X(_1927_));
 sg13g2_nand2_1 _3950_ (.Y(_1928_),
    .A(\counter[7] ),
    .B(\counter[6] ));
 sg13g2_nor4_1 _3951_ (.A(_1599_),
    .B(_1600_),
    .C(_1928_),
    .D(_1607_),
    .Y(_1929_));
 sg13g2_nor2_1 _3952_ (.A(\counter[10] ),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_nor2_1 _3953_ (.A(_1598_),
    .B(_1613_),
    .Y(_1931_));
 sg13g2_nor3_1 _3954_ (.A(net53),
    .B(_1930_),
    .C(_1931_),
    .Y(_0059_));
 sg13g2_nor2_1 _3955_ (.A(\counter[11] ),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_nor3_1 _3956_ (.A(net53),
    .B(_1614_),
    .C(_1932_),
    .Y(_0060_));
 sg13g2_nor2_1 _3957_ (.A(_1573_),
    .B(_1614_),
    .Y(_1933_));
 sg13g2_inv_1 _3958_ (.Y(_1934_),
    .A(_1615_));
 sg13g2_nor3_1 _3959_ (.A(net53),
    .B(_1933_),
    .C(_1934_),
    .Y(_0061_));
 sg13g2_nor2_1 _3960_ (.A(_1572_),
    .B(_1934_),
    .Y(_1935_));
 sg13g2_nor3_1 _3961_ (.A(net53),
    .B(_1616_),
    .C(_1935_),
    .Y(_0062_));
 sg13g2_nand4_1 _3962_ (.B(\counter[10] ),
    .C(_1572_),
    .A(\counter[11] ),
    .Y(_1936_),
    .D(_1573_));
 sg13g2_nand2b_1 _3963_ (.Y(_1937_),
    .B(_1929_),
    .A_N(_1936_));
 sg13g2_inv_1 _3964_ (.Y(_1938_),
    .A(_1937_));
 sg13g2_nor2_1 _3965_ (.A(_1574_),
    .B(_1938_),
    .Y(_1939_));
 sg13g2_nand2_1 _3966_ (.Y(_1940_),
    .A(_1938_),
    .B(_1574_));
 sg13g2_inv_1 _3967_ (.Y(_1941_),
    .A(_1940_));
 sg13g2_nor3_1 _3968_ (.A(net53),
    .B(_1939_),
    .C(_1941_),
    .Y(_0063_));
 sg13g2_nor2_1 _3969_ (.A(\counter[15] ),
    .B(_1941_),
    .Y(_1942_));
 sg13g2_inv_1 _3970_ (.Y(_1943_),
    .A(_1617_));
 sg13g2_nor3_1 _3971_ (.A(net53),
    .B(_1942_),
    .C(_1943_),
    .Y(_0064_));
 sg13g2_nor2_1 _3972_ (.A(\counter[16] ),
    .B(_1943_),
    .Y(_1944_));
 sg13g2_nor3_1 _3973_ (.A(net53),
    .B(_1618_),
    .C(_1944_),
    .Y(_0065_));
 sg13g2_nor2_1 _3974_ (.A(\counter[17] ),
    .B(_1618_),
    .Y(_1945_));
 sg13g2_inv_1 _3975_ (.Y(_1946_),
    .A(_1619_));
 sg13g2_nor3_1 _3976_ (.A(net53),
    .B(_1945_),
    .C(_1946_),
    .Y(_0066_));
 sg13g2_nor2_1 _3977_ (.A(\counter[18] ),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_nor3_1 _3978_ (.A(_1927_),
    .B(_1620_),
    .C(_1947_),
    .Y(_0067_));
 sg13g2_buf_1 _3979_ (.A(net67),
    .X(_1948_));
 sg13g2_nor2_1 _3980_ (.A(\counter[19] ),
    .B(_1620_),
    .Y(_1949_));
 sg13g2_inv_1 _3981_ (.Y(_1950_),
    .A(_1621_));
 sg13g2_nor3_1 _3982_ (.A(net52),
    .B(_1949_),
    .C(_1950_),
    .Y(_0068_));
 sg13g2_inv_1 _3983_ (.Y(_1951_),
    .A(_1603_));
 sg13g2_nor3_1 _3984_ (.A(net52),
    .B(_1568_),
    .C(_1951_),
    .Y(_0069_));
 sg13g2_nor2_1 _3985_ (.A(\counter[20] ),
    .B(_1950_),
    .Y(_1952_));
 sg13g2_nor3_1 _3986_ (.A(net52),
    .B(_1622_),
    .C(_1952_),
    .Y(_0070_));
 sg13g2_nor2_1 _3987_ (.A(\counter[21] ),
    .B(_1622_),
    .Y(_1953_));
 sg13g2_nor3_1 _3988_ (.A(net52),
    .B(_1953_),
    .C(_1624_),
    .Y(_0071_));
 sg13g2_nor2_1 _3989_ (.A(\counter[22] ),
    .B(_1624_),
    .Y(_1954_));
 sg13g2_nor2b_1 _3990_ (.A(_1625_),
    .B_N(\counter[22] ),
    .Y(_1955_));
 sg13g2_nor3_1 _3991_ (.A(net52),
    .B(_1954_),
    .C(_1955_),
    .Y(_0072_));
 sg13g2_nor2_1 _3992_ (.A(_1591_),
    .B(_1625_),
    .Y(_1956_));
 sg13g2_nor2_1 _3993_ (.A(\counter[23] ),
    .B(_1955_),
    .Y(_1957_));
 sg13g2_nor3_1 _3994_ (.A(net52),
    .B(_1956_),
    .C(_1957_),
    .Y(_0073_));
 sg13g2_nor2_1 _3995_ (.A(\counter[24] ),
    .B(_1956_),
    .Y(_1958_));
 sg13g2_nand2_1 _3996_ (.Y(_1959_),
    .A(_1956_),
    .B(\counter[24] ));
 sg13g2_inv_1 _3997_ (.Y(_1960_),
    .A(_1959_));
 sg13g2_nor3_1 _3998_ (.A(_1948_),
    .B(_1958_),
    .C(_1960_),
    .Y(_0074_));
 sg13g2_a221oi_1 _3999_ (.B2(_1589_),
    .C1(_1927_),
    .B1(_1959_),
    .A1(_1592_),
    .Y(_0075_),
    .A2(_1624_));
 sg13g2_nor2_1 _4000_ (.A(_1562_),
    .B(_1626_),
    .Y(_1961_));
 sg13g2_nor3_1 _4001_ (.A(_1948_),
    .B(_1961_),
    .C(_1632_),
    .Y(_0076_));
 sg13g2_nor2_1 _4002_ (.A(\counter[2] ),
    .B(_1951_),
    .Y(_1962_));
 sg13g2_nor3_1 _4003_ (.A(net52),
    .B(_1604_),
    .C(_1962_),
    .Y(_0080_));
 sg13g2_nor2b_1 _4004_ (.A(_1630_),
    .B_N(\counter[30] ),
    .Y(_1963_));
 sg13g2_nor2_1 _4005_ (.A(\counter[30] ),
    .B(_1631_),
    .Y(_1964_));
 sg13g2_nor3_1 _4006_ (.A(net52),
    .B(_1963_),
    .C(_1964_),
    .Y(_0081_));
 sg13g2_o21ai_1 _4007_ (.B1(_1586_),
    .Y(_1965_),
    .A1(\counter[31] ),
    .A2(_1963_));
 sg13g2_a21oi_1 _4008_ (.A1(\counter[31] ),
    .A2(_1963_),
    .Y(_0082_),
    .B1(_1965_));
 sg13g2_nor2_1 _4009_ (.A(\counter[3] ),
    .B(_1604_),
    .Y(_1966_));
 sg13g2_nor3_1 _4010_ (.A(net67),
    .B(_1966_),
    .C(_1639_),
    .Y(_0083_));
 sg13g2_nor2_1 _4011_ (.A(_1565_),
    .B(_1605_),
    .Y(_1967_));
 sg13g2_nor2_1 _4012_ (.A(\counter[4] ),
    .B(_1639_),
    .Y(_1968_));
 sg13g2_nor3_1 _4013_ (.A(net67),
    .B(_1967_),
    .C(_1968_),
    .Y(_0084_));
 sg13g2_nor2_1 _4014_ (.A(\counter[5] ),
    .B(_1967_),
    .Y(_1969_));
 sg13g2_nor3_1 _4015_ (.A(net67),
    .B(_1606_),
    .C(_1969_),
    .Y(_0085_));
 sg13g2_nor2_1 _4016_ (.A(\counter[6] ),
    .B(_1606_),
    .Y(_1970_));
 sg13g2_nor3_1 _4017_ (.A(_1588_),
    .B(_1970_),
    .C(_1608_),
    .Y(_0086_));
 sg13g2_nor2_1 _4018_ (.A(\counter[7] ),
    .B(_1608_),
    .Y(_1971_));
 sg13g2_inv_1 _4019_ (.Y(_1972_),
    .A(_1609_));
 sg13g2_nor3_1 _4020_ (.A(_1588_),
    .B(_1971_),
    .C(_1972_),
    .Y(_0087_));
 sg13g2_nor2_1 _4021_ (.A(\counter[8] ),
    .B(_1972_),
    .Y(_1973_));
 sg13g2_nor3_1 _4022_ (.A(net67),
    .B(_1610_),
    .C(_1973_),
    .Y(_0088_));
 sg13g2_nor2_1 _4023_ (.A(\counter[9] ),
    .B(_1610_),
    .Y(_1974_));
 sg13g2_nor3_1 _4024_ (.A(net67),
    .B(_1974_),
    .C(_1612_),
    .Y(_0089_));
 sg13g2_inv_1 _4025_ (.Y(_1975_),
    .A(_0056_));
 sg13g2_o21ai_1 _4026_ (.B1(_1578_),
    .Y(_1976_),
    .A1(\i_project.controller_0.mode_ramp_base[0] ),
    .A2(_1903_));
 sg13g2_a21oi_1 _4027_ (.A1(_1975_),
    .A2(_1903_),
    .Y(_0101_),
    .B1(_1976_));
 sg13g2_buf_1 _4028_ (.A(_1789_),
    .X(_1977_));
 sg13g2_buf_2 _4029_ (.A(\i_project.controller_0.mode_ramp_base[7] ),
    .X(_1978_));
 sg13g2_inv_1 _4030_ (.Y(_1979_),
    .A(_1978_));
 sg13g2_buf_8 _4031_ (.A(\i_project.controller_0.mode_ramp_base[6] ),
    .X(_1980_));
 sg13g2_inv_1 _4032_ (.Y(_1981_),
    .A(net70));
 sg13g2_buf_8 _4033_ (.A(\i_project.controller_0.mode_ramp_base[5] ),
    .X(_1982_));
 sg13g2_inv_1 _4034_ (.Y(_1983_),
    .A(_1982_));
 sg13g2_buf_1 _4035_ (.A(\i_project.controller_0.mode_ramp_base[4] ),
    .X(_1984_));
 sg13g2_buf_2 _4036_ (.A(_1984_),
    .X(_1985_));
 sg13g2_inv_1 _4037_ (.Y(_1986_),
    .A(net59));
 sg13g2_buf_1 _4038_ (.A(\i_project.controller_0.mode_ramp_base[3] ),
    .X(_1987_));
 sg13g2_inv_1 _4039_ (.Y(_1988_),
    .A(net69));
 sg13g2_buf_2 _4040_ (.A(\i_project.controller_0.mode_ramp_base[1] ),
    .X(_1989_));
 sg13g2_inv_1 _4041_ (.Y(_1990_),
    .A(_1989_));
 sg13g2_inv_1 _4042_ (.Y(_1991_),
    .A(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_nor3_1 _4043_ (.A(_1990_),
    .B(_1991_),
    .C(_1904_),
    .Y(_1992_));
 sg13g2_buf_2 _4044_ (.A(\i_project.controller_0.mode_ramp_base[2] ),
    .X(_1993_));
 sg13g2_nand2_1 _4045_ (.Y(_1994_),
    .A(_1992_),
    .B(_1993_));
 sg13g2_nor2_1 _4046_ (.A(_1988_),
    .B(_1994_),
    .Y(_1995_));
 sg13g2_inv_1 _4047_ (.Y(_1996_),
    .A(_1995_));
 sg13g2_nor2_1 _4048_ (.A(_1986_),
    .B(_1996_),
    .Y(_1997_));
 sg13g2_inv_1 _4049_ (.Y(_1998_),
    .A(_1997_));
 sg13g2_nor2_1 _4050_ (.A(_1983_),
    .B(_1998_),
    .Y(_1999_));
 sg13g2_inv_1 _4051_ (.Y(_2000_),
    .A(_1999_));
 sg13g2_nor3_1 _4052_ (.A(_1979_),
    .B(_1981_),
    .C(_2000_),
    .Y(_2001_));
 sg13g2_buf_2 _4053_ (.A(\i_project.controller_0.t[8] ),
    .X(_2002_));
 sg13g2_nand2_1 _4054_ (.Y(_2003_),
    .A(_2001_),
    .B(_2002_));
 sg13g2_buf_1 _4055_ (.A(\i_project.controller_0.t[9] ),
    .X(_2004_));
 sg13g2_nor2b_1 _4056_ (.A(_2003_),
    .B_N(_2004_),
    .Y(_2005_));
 sg13g2_nor2_1 _4057_ (.A(\i_project.controller_0.t[10] ),
    .B(_2005_),
    .Y(_2006_));
 sg13g2_and2_1 _4058_ (.A(_2005_),
    .B(\i_project.controller_0.t[10] ),
    .X(_2007_));
 sg13g2_buf_1 _4059_ (.A(_2007_),
    .X(_2008_));
 sg13g2_nor3_1 _4060_ (.A(net51),
    .B(_2006_),
    .C(_2008_),
    .Y(_0102_));
 sg13g2_buf_1 _4061_ (.A(\i_project.controller_0.t[11] ),
    .X(_2009_));
 sg13g2_o21ai_1 _4062_ (.B1(net68),
    .Y(_2010_),
    .A1(_2009_),
    .A2(_2008_));
 sg13g2_a21oi_1 _4063_ (.A1(_2009_),
    .A2(_2008_),
    .Y(_0103_),
    .B1(_2010_));
 sg13g2_a21oi_1 _4064_ (.A1(_1903_),
    .A2(\i_project.controller_0.mode_ramp_base[0] ),
    .Y(_2011_),
    .B1(_1989_));
 sg13g2_nor3_1 _4065_ (.A(net51),
    .B(_2011_),
    .C(_1992_),
    .Y(_0104_));
 sg13g2_nor2_1 _4066_ (.A(_1993_),
    .B(_1992_),
    .Y(_2012_));
 sg13g2_inv_1 _4067_ (.Y(_2013_),
    .A(_1994_));
 sg13g2_nor3_1 _4068_ (.A(net51),
    .B(_2012_),
    .C(_2013_),
    .Y(_0105_));
 sg13g2_nor2_1 _4069_ (.A(net69),
    .B(_2013_),
    .Y(_2014_));
 sg13g2_nor3_1 _4070_ (.A(net51),
    .B(_1995_),
    .C(_2014_),
    .Y(_0106_));
 sg13g2_nor2_1 _4071_ (.A(net59),
    .B(_1995_),
    .Y(_2015_));
 sg13g2_nor3_1 _4072_ (.A(net51),
    .B(_2015_),
    .C(_1997_),
    .Y(_0107_));
 sg13g2_buf_1 _4073_ (.A(_1982_),
    .X(_2016_));
 sg13g2_nor2_1 _4074_ (.A(net58),
    .B(_1997_),
    .Y(_2017_));
 sg13g2_nor3_1 _4075_ (.A(net51),
    .B(_2017_),
    .C(_1999_),
    .Y(_0108_));
 sg13g2_nor2_1 _4076_ (.A(net70),
    .B(_1999_),
    .Y(_2018_));
 sg13g2_nor2_1 _4077_ (.A(_1981_),
    .B(_2000_),
    .Y(_2019_));
 sg13g2_nor3_1 _4078_ (.A(net51),
    .B(_2018_),
    .C(_2019_),
    .Y(_0109_));
 sg13g2_nor2_1 _4079_ (.A(_1978_),
    .B(_2019_),
    .Y(_2020_));
 sg13g2_nor3_1 _4080_ (.A(net51),
    .B(_2001_),
    .C(_2020_),
    .Y(_0110_));
 sg13g2_nor2_1 _4081_ (.A(_2002_),
    .B(_2001_),
    .Y(_2021_));
 sg13g2_inv_1 _4082_ (.Y(_2022_),
    .A(_2003_));
 sg13g2_nor3_1 _4083_ (.A(_1977_),
    .B(_2021_),
    .C(_2022_),
    .Y(_0111_));
 sg13g2_nor2_1 _4084_ (.A(_2004_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_nor3_1 _4085_ (.A(_1977_),
    .B(_2005_),
    .C(_2023_),
    .Y(_0112_));
 sg13g2_nand2_1 _4086_ (.Y(_2024_),
    .A(net74),
    .B(net4));
 sg13g2_inv_1 _4087_ (.Y(_0143_),
    .A(_2024_));
 sg13g2_nor3_2 _4088_ (.A(_1757_),
    .B(_1792_),
    .C(_1771_),
    .Y(_2025_));
 sg13g2_buf_8 _4089_ (.A(_2025_),
    .X(_2026_));
 sg13g2_inv_4 _4090_ (.A(net48),
    .Y(_2027_));
 sg13g2_xnor2_1 _4091_ (.Y(_2028_),
    .A(_1673_),
    .B(\i_project.controller_0.mode_ramp_base[6] ));
 sg13g2_xnor2_1 _4092_ (.Y(_2029_),
    .A(_1671_),
    .B(_1982_));
 sg13g2_nand2_1 _4093_ (.Y(_2030_),
    .A(_1666_),
    .B(_1987_));
 sg13g2_xnor2_1 _4094_ (.Y(_2031_),
    .A(\i_project.controller_0.h[1] ),
    .B(_1984_));
 sg13g2_nand2_1 _4095_ (.Y(_2032_),
    .A(net73),
    .B(_1984_));
 sg13g2_o21ai_1 _4096_ (.B1(_2032_),
    .Y(_2033_),
    .A1(_2030_),
    .A2(_2031_));
 sg13g2_buf_1 _4097_ (.A(_2033_),
    .X(_2034_));
 sg13g2_nand2b_1 _4098_ (.Y(_2035_),
    .B(_2034_),
    .A_N(_2029_));
 sg13g2_nand2_1 _4099_ (.Y(_2036_),
    .A(_1671_),
    .B(_1982_));
 sg13g2_nand2_1 _4100_ (.Y(_2037_),
    .A(_2035_),
    .B(_2036_));
 sg13g2_xnor2_1 _4101_ (.Y(_2038_),
    .A(_2028_),
    .B(_2037_));
 sg13g2_inv_2 _4102_ (.Y(_2039_),
    .A(_1713_));
 sg13g2_nand2_1 _4103_ (.Y(_2040_),
    .A(_2039_),
    .B(_1780_));
 sg13g2_nand2_1 _4104_ (.Y(_2041_),
    .A(_1713_),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _4105_ (.Y(_2042_),
    .A(_2040_),
    .B(_2041_));
 sg13g2_xor2_1 _4106_ (.B(_1776_),
    .A(_1716_),
    .X(_2043_));
 sg13g2_xor2_1 _4107_ (.B(\i_project.controller_0.voffset[2] ),
    .A(_1712_),
    .X(_2044_));
 sg13g2_nand2_2 _4108_ (.Y(_2045_),
    .A(_1715_),
    .B(\i_project.controller_0.voffset[0] ));
 sg13g2_inv_2 _4109_ (.Y(_2046_),
    .A(_2045_));
 sg13g2_nand3_1 _4110_ (.B(_2044_),
    .C(_2046_),
    .A(_2043_),
    .Y(_2047_));
 sg13g2_nand2_1 _4111_ (.Y(_2048_),
    .A(_1716_),
    .B(_1776_));
 sg13g2_nor2_1 _4112_ (.A(_1712_),
    .B(\i_project.controller_0.voffset[2] ),
    .Y(_2049_));
 sg13g2_nand2_1 _4113_ (.Y(_2050_),
    .A(_1712_),
    .B(\i_project.controller_0.voffset[2] ));
 sg13g2_o21ai_1 _4114_ (.B1(_2050_),
    .Y(_2051_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_inv_2 _4115_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_nand2_1 _4116_ (.Y(_2053_),
    .A(_2047_),
    .B(_2052_));
 sg13g2_nand2b_1 _4117_ (.Y(_2054_),
    .B(_2053_),
    .A_N(_2042_));
 sg13g2_nand3_1 _4118_ (.B(_2042_),
    .C(_2052_),
    .A(_2047_),
    .Y(_2055_));
 sg13g2_nand2_1 _4119_ (.Y(_2056_),
    .A(_2054_),
    .B(_2055_));
 sg13g2_buf_8 _4120_ (.A(_2056_),
    .X(_2057_));
 sg13g2_xnor2_1 _4121_ (.Y(_2058_),
    .A(_1980_),
    .B(_2057_));
 sg13g2_nand2_1 _4122_ (.Y(_2059_),
    .A(_2043_),
    .B(_2046_));
 sg13g2_xnor2_1 _4123_ (.Y(_2060_),
    .A(_1716_),
    .B(_1776_));
 sg13g2_nand2_1 _4124_ (.Y(_2061_),
    .A(_2060_),
    .B(_2045_));
 sg13g2_nand2_2 _4125_ (.Y(_2062_),
    .A(_2059_),
    .B(_2061_));
 sg13g2_nand2_1 _4126_ (.Y(_2063_),
    .A(_2062_),
    .B(_0043_));
 sg13g2_nand2_1 _4127_ (.Y(_2064_),
    .A(_1886_),
    .B(_1739_));
 sg13g2_nand2_1 _4128_ (.Y(_2065_),
    .A(_2064_),
    .B(_2045_));
 sg13g2_buf_2 _4129_ (.A(_2065_),
    .X(_2066_));
 sg13g2_nor2_1 _4130_ (.A(_1988_),
    .B(_2066_),
    .Y(_2067_));
 sg13g2_buf_8 _4131_ (.A(_2062_),
    .X(_2068_));
 sg13g2_nor2_1 _4132_ (.A(_0043_),
    .B(net36),
    .Y(_2069_));
 sg13g2_a21oi_1 _4133_ (.A1(_2063_),
    .A2(_2067_),
    .Y(_2070_),
    .B1(_2069_));
 sg13g2_inv_1 _4134_ (.Y(_2071_),
    .A(_2070_));
 sg13g2_nor2_1 _4135_ (.A(_1716_),
    .B(_1776_),
    .Y(_2072_));
 sg13g2_inv_1 _4136_ (.Y(_2073_),
    .A(_2072_));
 sg13g2_inv_1 _4137_ (.Y(_2074_),
    .A(_2048_));
 sg13g2_a21oi_1 _4138_ (.A1(_2073_),
    .A2(_2046_),
    .Y(_2075_),
    .B1(_2074_));
 sg13g2_nand2_1 _4139_ (.Y(_2076_),
    .A(_1721_),
    .B(_1778_));
 sg13g2_nand2_2 _4140_ (.Y(_2077_),
    .A(_2076_),
    .B(_2050_));
 sg13g2_nand2_1 _4141_ (.Y(_2078_),
    .A(_2075_),
    .B(_2077_));
 sg13g2_o21ai_1 _4142_ (.B1(_2048_),
    .Y(_2079_),
    .A1(_2045_),
    .A2(_2072_));
 sg13g2_buf_2 _4143_ (.A(_2079_),
    .X(_2080_));
 sg13g2_nand2_1 _4144_ (.Y(_2081_),
    .A(_2080_),
    .B(_2044_));
 sg13g2_nand2_1 _4145_ (.Y(_2082_),
    .A(_2078_),
    .B(_2081_));
 sg13g2_buf_2 _4146_ (.A(_2082_),
    .X(_2083_));
 sg13g2_nand2_1 _4147_ (.Y(_2084_),
    .A(_2083_),
    .B(_1982_));
 sg13g2_nand3_1 _4148_ (.B(_2081_),
    .C(_1983_),
    .A(_2078_),
    .Y(_2085_));
 sg13g2_nand2_1 _4149_ (.Y(_2086_),
    .A(_2084_),
    .B(_2085_));
 sg13g2_nand2_1 _4150_ (.Y(_2087_),
    .A(_2071_),
    .B(_2086_));
 sg13g2_xnor2_1 _4151_ (.Y(_2088_),
    .A(_2077_),
    .B(_2080_));
 sg13g2_buf_8 _4152_ (.A(_2088_),
    .X(_2089_));
 sg13g2_inv_1 _4153_ (.Y(_2090_),
    .A(_0042_));
 sg13g2_nand2_1 _4154_ (.Y(_2091_),
    .A(_2089_),
    .B(_2090_));
 sg13g2_nand2_1 _4155_ (.Y(_2092_),
    .A(_2087_),
    .B(_2091_));
 sg13g2_inv_1 _4156_ (.Y(_2093_),
    .A(_2092_));
 sg13g2_nand2b_1 _4157_ (.Y(_2094_),
    .B(_2093_),
    .A_N(_2058_));
 sg13g2_nand2_1 _4158_ (.Y(_2095_),
    .A(_2092_),
    .B(_2058_));
 sg13g2_nand2_1 _4159_ (.Y(_2096_),
    .A(_2094_),
    .B(_2095_));
 sg13g2_xnor2_1 _4160_ (.Y(_2097_),
    .A(_2038_),
    .B(_2096_));
 sg13g2_buf_8 _4161_ (.A(_2057_),
    .X(_2098_));
 sg13g2_xnor2_1 _4162_ (.Y(_2099_),
    .A(_1674_),
    .B(_2098_));
 sg13g2_nor3_1 _4163_ (.A(_1760_),
    .B(_0027_),
    .C(_1794_),
    .Y(_2100_));
 sg13g2_buf_1 _4164_ (.A(_2100_),
    .X(_2101_));
 sg13g2_a21oi_1 _4165_ (.A1(_2099_),
    .A2(net47),
    .Y(_2102_),
    .B1(net48));
 sg13g2_inv_1 _4166_ (.Y(_2103_),
    .A(_2102_));
 sg13g2_o21ai_1 _4167_ (.B1(_2103_),
    .Y(_2104_),
    .A1(net41),
    .A2(_2097_));
 sg13g2_xnor2_1 _4168_ (.Y(_2105_),
    .A(_1859_),
    .B(_2083_));
 sg13g2_inv_1 _4169_ (.Y(_2106_),
    .A(_2105_));
 sg13g2_nor3_1 _4170_ (.A(_1757_),
    .B(_1760_),
    .C(_1771_),
    .Y(_2107_));
 sg13g2_buf_1 _4171_ (.A(_2107_),
    .X(_2108_));
 sg13g2_buf_1 _4172_ (.A(net50),
    .X(_2109_));
 sg13g2_nor3_1 _4173_ (.A(_1760_),
    .B(_1794_),
    .C(_1762_),
    .Y(_2110_));
 sg13g2_buf_2 _4174_ (.A(_2110_),
    .X(_2111_));
 sg13g2_buf_8 _4175_ (.A(_2111_),
    .X(_2112_));
 sg13g2_buf_1 _4176_ (.A(net40),
    .X(_2113_));
 sg13g2_a21oi_1 _4177_ (.A1(_2106_),
    .A2(_2109_),
    .Y(_2114_),
    .B1(net35));
 sg13g2_nand2_1 _4178_ (.Y(_2115_),
    .A(_2104_),
    .B(_2114_));
 sg13g2_nor3_2 _4179_ (.A(_1757_),
    .B(_1792_),
    .C(_1762_),
    .Y(_2116_));
 sg13g2_buf_8 _4180_ (.A(_2116_),
    .X(_2117_));
 sg13g2_buf_1 _4181_ (.A(_2117_),
    .X(_2118_));
 sg13g2_inv_1 _4182_ (.Y(_2119_),
    .A(net39));
 sg13g2_nor2_1 _4183_ (.A(_1698_),
    .B(_1700_),
    .Y(_2120_));
 sg13g2_inv_1 _4184_ (.Y(_2121_),
    .A(_2120_));
 sg13g2_nand2_1 _4185_ (.Y(_2122_),
    .A(_1580_),
    .B(_0054_));
 sg13g2_a21oi_1 _4186_ (.A1(_1579_),
    .A2(_0038_),
    .Y(_2123_),
    .B1(_1582_));
 sg13g2_nand2_1 _4187_ (.Y(_2124_),
    .A(_1741_),
    .B(_1579_));
 sg13g2_o21ai_1 _4188_ (.B1(_2124_),
    .Y(_2125_),
    .A1(_1579_),
    .A2(_0037_));
 sg13g2_a22oi_1 _4189_ (.Y(_2126_),
    .B1(_1582_),
    .B2(_2125_),
    .A2(_2123_),
    .A1(_2122_));
 sg13g2_nand2_1 _4190_ (.Y(_2127_),
    .A(_2121_),
    .B(_1850_));
 sg13g2_o21ai_1 _4191_ (.B1(_2127_),
    .Y(_2128_),
    .A1(_2121_),
    .A2(_2126_));
 sg13g2_buf_1 _4192_ (.A(_2128_),
    .X(_2129_));
 sg13g2_buf_1 _4193_ (.A(_2129_),
    .X(_2130_));
 sg13g2_buf_1 _4194_ (.A(net29),
    .X(_2131_));
 sg13g2_buf_1 _4195_ (.A(_1579_),
    .X(_2132_));
 sg13g2_nand2_1 _4196_ (.Y(_2133_),
    .A(net57),
    .B(_0051_));
 sg13g2_inv_1 _4197_ (.Y(_2134_),
    .A(_2133_));
 sg13g2_a21oi_1 _4198_ (.A1(_1580_),
    .A2(_0053_),
    .Y(_2135_),
    .B1(_2134_));
 sg13g2_inv_1 _4199_ (.Y(_2136_),
    .A(_2135_));
 sg13g2_nand2_1 _4200_ (.Y(_2137_),
    .A(_2125_),
    .B(net55));
 sg13g2_o21ai_1 _4201_ (.B1(_2137_),
    .Y(_2138_),
    .A1(net55),
    .A2(_2136_));
 sg13g2_inv_1 _4202_ (.Y(_2139_),
    .A(_2138_));
 sg13g2_inv_1 _4203_ (.Y(_2140_),
    .A(net40));
 sg13g2_a21oi_1 _4204_ (.A1(net29),
    .A2(_2139_),
    .Y(_2141_),
    .B1(_2140_));
 sg13g2_o21ai_1 _4205_ (.B1(_2141_),
    .Y(_2142_),
    .A1(net25),
    .A2(_2139_));
 sg13g2_nand3_1 _4206_ (.B(net34),
    .C(_2142_),
    .A(_2115_),
    .Y(_2143_));
 sg13g2_buf_1 _4207_ (.A(net39),
    .X(_2144_));
 sg13g2_nand2_1 _4208_ (.Y(_2145_),
    .A(_1696_),
    .B(_1680_));
 sg13g2_buf_2 _4209_ (.A(_2145_),
    .X(_2146_));
 sg13g2_inv_4 _4210_ (.A(_2146_),
    .Y(_2147_));
 sg13g2_buf_1 _4211_ (.A(net28),
    .X(_2148_));
 sg13g2_a21oi_1 _4212_ (.A1(_2138_),
    .A2(_2144_),
    .Y(_2149_),
    .B1(_2148_));
 sg13g2_xnor2_1 _4213_ (.Y(_2150_),
    .A(net72),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_xnor2_1 _4214_ (.Y(_2151_),
    .A(_1706_),
    .B(_1783_));
 sg13g2_nor2_1 _4215_ (.A(_2150_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_xnor2_1 _4216_ (.Y(_2153_),
    .A(_1705_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _4217_ (.A(_2153_),
    .B(_2042_),
    .Y(_2154_));
 sg13g2_and2_1 _4218_ (.A(_2152_),
    .B(_2154_),
    .X(_2155_));
 sg13g2_nand2_1 _4219_ (.Y(_2156_),
    .A(_2053_),
    .B(_2155_));
 sg13g2_nand2_1 _4220_ (.Y(_2157_),
    .A(_1705_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _4221_ (.A(_1705_),
    .B(\i_project.controller_0.voffset[4] ),
    .Y(_2158_));
 sg13g2_a21oi_1 _4222_ (.A1(_2041_),
    .A2(_2157_),
    .Y(_2159_),
    .B1(_2158_));
 sg13g2_nand2_1 _4223_ (.Y(_2160_),
    .A(_1706_),
    .B(_1783_));
 sg13g2_nor2_1 _4224_ (.A(net72),
    .B(\i_project.controller_0.voffset[6] ),
    .Y(_2161_));
 sg13g2_nand2_1 _4225_ (.Y(_2162_),
    .A(net72),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_o21ai_1 _4226_ (.B1(_2162_),
    .Y(_2163_),
    .A1(_2160_),
    .A2(_2161_));
 sg13g2_a21oi_1 _4227_ (.A1(_2152_),
    .A2(_2159_),
    .Y(_2164_),
    .B1(_2163_));
 sg13g2_nand2_1 _4228_ (.Y(_2165_),
    .A(_2156_),
    .B(_2164_));
 sg13g2_nor2_1 _4229_ (.A(_1701_),
    .B(\i_project.controller_0.voffset[7] ),
    .Y(_2166_));
 sg13g2_nand2_1 _4230_ (.Y(_2167_),
    .A(_1701_),
    .B(\i_project.controller_0.voffset[7] ));
 sg13g2_inv_1 _4231_ (.Y(_2168_),
    .A(_2167_));
 sg13g2_nor2_1 _4232_ (.A(_2166_),
    .B(_2168_),
    .Y(_2169_));
 sg13g2_nand2_1 _4233_ (.Y(_2170_),
    .A(_2165_),
    .B(_2169_));
 sg13g2_nand2b_1 _4234_ (.Y(_2171_),
    .B(_2168_),
    .A_N(_0030_));
 sg13g2_o21ai_1 _4235_ (.B1(_2171_),
    .Y(_2172_),
    .A1(_1699_),
    .A2(_2170_));
 sg13g2_nand2b_1 _4236_ (.Y(_2173_),
    .B(_1700_),
    .A_N(_2172_));
 sg13g2_inv_1 _4237_ (.Y(_2174_),
    .A(_1666_));
 sg13g2_nand2_1 _4238_ (.Y(_2175_),
    .A(_2172_),
    .B(_1729_));
 sg13g2_nand3_1 _4239_ (.B(_2174_),
    .C(_2175_),
    .A(_2173_),
    .Y(_2176_));
 sg13g2_nor2_1 _4240_ (.A(_2077_),
    .B(_2042_),
    .Y(_2177_));
 sg13g2_nand2_1 _4241_ (.Y(_2178_),
    .A(_2177_),
    .B(_2080_));
 sg13g2_inv_1 _4242_ (.Y(_2179_),
    .A(_2050_));
 sg13g2_inv_1 _4243_ (.Y(_2180_),
    .A(_2041_));
 sg13g2_a21oi_1 _4244_ (.A1(_2040_),
    .A2(_2179_),
    .Y(_2181_),
    .B1(_2180_));
 sg13g2_nand2_1 _4245_ (.Y(_2182_),
    .A(_2178_),
    .B(_2181_));
 sg13g2_nor2_1 _4246_ (.A(_2153_),
    .B(_2151_),
    .Y(_2183_));
 sg13g2_inv_1 _4247_ (.Y(_2184_),
    .A(_2169_));
 sg13g2_nor2_1 _4248_ (.A(_2150_),
    .B(_2184_),
    .Y(_2185_));
 sg13g2_nand3_1 _4249_ (.B(_2183_),
    .C(_2185_),
    .A(_2182_),
    .Y(_2186_));
 sg13g2_o21ai_1 _4250_ (.B1(_2160_),
    .Y(_2187_),
    .A1(_2157_),
    .A2(_2151_));
 sg13g2_o21ai_1 _4251_ (.B1(_2167_),
    .Y(_2188_),
    .A1(_2162_),
    .A2(_2166_));
 sg13g2_a21oi_1 _4252_ (.A1(_2187_),
    .A2(_2185_),
    .Y(_2189_),
    .B1(_2188_));
 sg13g2_nand2_1 _4253_ (.Y(_2190_),
    .A(_2186_),
    .B(_2189_));
 sg13g2_xnor2_1 _4254_ (.Y(_2191_),
    .A(_1698_),
    .B(_2190_));
 sg13g2_nand2_1 _4255_ (.Y(_2192_),
    .A(_2191_),
    .B(net64));
 sg13g2_nor2_1 _4256_ (.A(_0038_),
    .B(_0037_),
    .Y(_2193_));
 sg13g2_nand3_1 _4257_ (.B(_2192_),
    .C(_2193_),
    .A(_2176_),
    .Y(_2194_));
 sg13g2_nand2_1 _4258_ (.Y(_2195_),
    .A(_2194_),
    .B(_1745_));
 sg13g2_inv_1 _4259_ (.Y(_2196_),
    .A(_2157_));
 sg13g2_nor2_1 _4260_ (.A(_2158_),
    .B(_2196_),
    .Y(_2197_));
 sg13g2_nand2_1 _4261_ (.Y(_2198_),
    .A(_2182_),
    .B(_2197_));
 sg13g2_nand3_1 _4262_ (.B(_2181_),
    .C(_2153_),
    .A(_2178_),
    .Y(_2199_));
 sg13g2_nand2_1 _4263_ (.Y(_2200_),
    .A(_2198_),
    .B(_2199_));
 sg13g2_buf_8 _4264_ (.A(_2200_),
    .X(_0145_));
 sg13g2_a21oi_1 _4265_ (.A1(_2051_),
    .A2(_2154_),
    .Y(_0146_),
    .B1(_2159_));
 sg13g2_nor2_1 _4266_ (.A(_2060_),
    .B(_2077_),
    .Y(_0147_));
 sg13g2_nand3_1 _4267_ (.B(_0147_),
    .C(_2046_),
    .A(_2154_),
    .Y(_0148_));
 sg13g2_nand2_1 _4268_ (.Y(_0149_),
    .A(_0146_),
    .B(_0148_));
 sg13g2_xor2_1 _4269_ (.B(_1783_),
    .A(_1706_),
    .X(_0150_));
 sg13g2_nand2_1 _4270_ (.Y(_0151_),
    .A(_0149_),
    .B(_0150_));
 sg13g2_nand3_1 _4271_ (.B(_0148_),
    .C(_2151_),
    .A(_0146_),
    .Y(_0152_));
 sg13g2_nand2_1 _4272_ (.Y(_0153_),
    .A(_0151_),
    .B(_0152_));
 sg13g2_buf_8 _4273_ (.A(_0153_),
    .X(_0154_));
 sg13g2_a22oi_1 _4274_ (.Y(_0155_),
    .B1(_1670_),
    .B2(_0154_),
    .A2(net20),
    .A1(_1866_));
 sg13g2_nand2_1 _4275_ (.Y(_0156_),
    .A(_2197_),
    .B(_0150_));
 sg13g2_nor2_1 _4276_ (.A(_0156_),
    .B(_2181_),
    .Y(_0157_));
 sg13g2_nor2_1 _4277_ (.A(_2187_),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_nand3_1 _4278_ (.B(_2080_),
    .C(_2183_),
    .A(_2177_),
    .Y(_0159_));
 sg13g2_nand2_1 _4279_ (.Y(_0160_),
    .A(_0158_),
    .B(_0159_));
 sg13g2_nand2b_1 _4280_ (.Y(_0161_),
    .B(_0160_),
    .A_N(_2150_));
 sg13g2_nand3_1 _4281_ (.B(_0159_),
    .C(_2150_),
    .A(_0158_),
    .Y(_0162_));
 sg13g2_nand2_2 _4282_ (.Y(_0163_),
    .A(_0161_),
    .B(_0162_));
 sg13g2_buf_8 _4283_ (.A(_0163_),
    .X(_0164_));
 sg13g2_nand3_1 _4284_ (.B(_1669_),
    .C(net64),
    .A(net18),
    .Y(_0165_));
 sg13g2_nand3_1 _4285_ (.B(_2184_),
    .C(_2164_),
    .A(_2156_),
    .Y(_0166_));
 sg13g2_nand2_1 _4286_ (.Y(_0167_),
    .A(_2170_),
    .B(_0166_));
 sg13g2_buf_2 _4287_ (.A(_0167_),
    .X(_0168_));
 sg13g2_nand2_1 _4288_ (.Y(_0169_),
    .A(_0168_),
    .B(_1682_));
 sg13g2_nand3_1 _4289_ (.B(_0165_),
    .C(_0169_),
    .A(_0155_),
    .Y(_0170_));
 sg13g2_a21oi_1 _4290_ (.A1(_2089_),
    .A2(net64),
    .Y(_0171_),
    .B1(_1668_));
 sg13g2_o21ai_1 _4291_ (.B1(_0171_),
    .Y(_0172_),
    .A1(net64),
    .A2(_2098_));
 sg13g2_a22oi_1 _4292_ (.Y(_0173_),
    .B1(_1670_),
    .B2(_2068_),
    .A2(_2066_),
    .A1(_1866_));
 sg13g2_a21oi_1 _4293_ (.A1(_0172_),
    .A2(_0173_),
    .Y(_0174_),
    .B1(_1691_));
 sg13g2_a21oi_1 _4294_ (.A1(_0170_),
    .A2(_1746_),
    .Y(_0175_),
    .B1(_0174_));
 sg13g2_a21oi_2 _4295_ (.B1(_2146_),
    .Y(_0176_),
    .A2(_0175_),
    .A1(_2195_));
 sg13g2_a21oi_1 _4296_ (.A1(_2143_),
    .A2(_2149_),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_buf_1 _4297_ (.A(\depth[1] ),
    .X(_0178_));
 sg13g2_buf_1 _4298_ (.A(\depth[0] ),
    .X(_0179_));
 sg13g2_nand2_1 _4299_ (.Y(_0180_),
    .A(_0178_),
    .B(_0179_));
 sg13g2_nor2_1 _4300_ (.A(_0046_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_inv_1 _4301_ (.Y(_0182_),
    .A(_0178_));
 sg13g2_inv_1 _4302_ (.Y(_0183_),
    .A(\depth[2] ));
 sg13g2_nor3_1 _4303_ (.A(_0179_),
    .B(_0182_),
    .C(_0183_),
    .Y(_0184_));
 sg13g2_nor2_1 _4304_ (.A(_0181_),
    .B(_0184_),
    .Y(_0185_));
 sg13g2_inv_1 _4305_ (.Y(_0186_),
    .A(_0185_));
 sg13g2_inv_1 _4306_ (.Y(_0187_),
    .A(_0179_));
 sg13g2_nor3_2 _4307_ (.A(_0178_),
    .B(_0187_),
    .C(_0183_),
    .Y(_0188_));
 sg13g2_nand3b_1 _4308_ (.B(_1725_),
    .C(_1889_),
    .Y(_0189_),
    .A_N(net72));
 sg13g2_nand3_1 _4309_ (.B(_1701_),
    .C(_1730_),
    .A(_0189_),
    .Y(_0190_));
 sg13g2_nand4_1 _4310_ (.B(_1708_),
    .C(_1717_),
    .A(_1704_),
    .Y(_0191_),
    .D(_1889_));
 sg13g2_inv_1 _4311_ (.Y(_0192_),
    .A(_0029_));
 sg13g2_a21oi_1 _4312_ (.A1(_1704_),
    .A2(_0192_),
    .Y(_0193_),
    .B1(_1700_));
 sg13g2_nand2_1 _4313_ (.Y(_0194_),
    .A(_0191_),
    .B(_0193_));
 sg13g2_nand3_1 _4314_ (.B(_1728_),
    .C(_2121_),
    .A(_0194_),
    .Y(_0195_));
 sg13g2_nand3_1 _4315_ (.B(_0190_),
    .C(_0195_),
    .A(_1755_),
    .Y(_0196_));
 sg13g2_inv_4 _4316_ (.A(_1764_),
    .Y(_0197_));
 sg13g2_nand2_1 _4317_ (.Y(_0198_),
    .A(_0196_),
    .B(_0197_));
 sg13g2_buf_2 _4318_ (.A(_0198_),
    .X(_0199_));
 sg13g2_o21ai_1 _4319_ (.B1(_0199_),
    .Y(_0200_),
    .A1(_0186_),
    .A2(_0188_));
 sg13g2_a21oi_1 _4320_ (.A1(_0018_),
    .A2(_1765_),
    .Y(_0201_),
    .B1(_0200_));
 sg13g2_o21ai_1 _4321_ (.B1(_0201_),
    .Y(_0202_),
    .A1(net49),
    .A2(_0177_));
 sg13g2_inv_1 _4322_ (.Y(_0203_),
    .A(_0046_));
 sg13g2_a21oi_1 _4323_ (.A1(_0182_),
    .A2(_0187_),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_inv_1 _4324_ (.Y(_0205_),
    .A(_0180_));
 sg13g2_nor2_1 _4325_ (.A(\depth[2] ),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_inv_1 _4326_ (.Y(_0207_),
    .A(_0206_));
 sg13g2_nor2_1 _4327_ (.A(_0204_),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_buf_8 _4328_ (.A(_0208_),
    .X(_0209_));
 sg13g2_inv_1 _4329_ (.Y(_0210_),
    .A(_0209_));
 sg13g2_nand2_1 _4330_ (.Y(_0211_),
    .A(_0202_),
    .B(_0210_));
 sg13g2_nor3_1 _4331_ (.A(_0179_),
    .B(_0182_),
    .C(_0203_),
    .Y(_0212_));
 sg13g2_buf_2 _4332_ (.A(_0212_),
    .X(_0213_));
 sg13g2_inv_2 _4333_ (.Y(_0214_),
    .A(_0213_));
 sg13g2_xor2_1 _4334_ (.B(_2004_),
    .A(_1662_),
    .X(_0215_));
 sg13g2_nand2_1 _4335_ (.Y(_0216_),
    .A(net62),
    .B(net70));
 sg13g2_o21ai_1 _4336_ (.B1(_0216_),
    .Y(_0217_),
    .A1(_2036_),
    .A2(_2028_));
 sg13g2_xnor2_1 _4337_ (.Y(_0218_),
    .A(_1654_),
    .B(_2002_));
 sg13g2_xnor2_1 _4338_ (.Y(_0219_),
    .A(_1651_),
    .B(_1978_));
 sg13g2_nor2_1 _4339_ (.A(_0218_),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_nand2_1 _4340_ (.Y(_0221_),
    .A(_1651_),
    .B(_1978_));
 sg13g2_nand2_1 _4341_ (.Y(_0222_),
    .A(_1654_),
    .B(_2002_));
 sg13g2_o21ai_1 _4342_ (.B1(_0222_),
    .Y(_0223_),
    .A1(_0221_),
    .A2(_0218_));
 sg13g2_a21oi_1 _4343_ (.A1(_0217_),
    .A2(_0220_),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_nor2_1 _4344_ (.A(_2028_),
    .B(_2029_),
    .Y(_0225_));
 sg13g2_nand3_1 _4345_ (.B(_0225_),
    .C(_0220_),
    .A(_2034_),
    .Y(_0226_));
 sg13g2_nand2_1 _4346_ (.Y(_0227_),
    .A(_0224_),
    .B(_0226_));
 sg13g2_xnor2_1 _4347_ (.Y(_0228_),
    .A(_0215_),
    .B(_0227_));
 sg13g2_buf_1 _4348_ (.A(_0020_),
    .X(_0229_));
 sg13g2_inv_1 _4349_ (.Y(_0230_),
    .A(_0229_));
 sg13g2_xnor2_1 _4350_ (.Y(_0231_),
    .A(_0230_),
    .B(_0163_));
 sg13g2_xnor2_1 _4351_ (.Y(_0232_),
    .A(_0228_),
    .B(_0231_));
 sg13g2_inv_1 _4352_ (.Y(_0233_),
    .A(net22));
 sg13g2_inv_1 _4353_ (.Y(_0234_),
    .A(_0041_));
 sg13g2_nand2_1 _4354_ (.Y(_0235_),
    .A(_0233_),
    .B(_0234_));
 sg13g2_nand2_1 _4355_ (.Y(_0236_),
    .A(_2095_),
    .B(_0235_));
 sg13g2_inv_1 _4356_ (.Y(_0237_),
    .A(_2002_));
 sg13g2_nand2_1 _4357_ (.Y(_0238_),
    .A(_0149_),
    .B(_2151_));
 sg13g2_nand3_1 _4358_ (.B(_0148_),
    .C(_0150_),
    .A(_0146_),
    .Y(_0239_));
 sg13g2_nand2_2 _4359_ (.Y(_0240_),
    .A(_0238_),
    .B(_0239_));
 sg13g2_xnor2_1 _4360_ (.Y(_0241_),
    .A(_0237_),
    .B(_0240_));
 sg13g2_buf_1 _4361_ (.A(_0040_),
    .X(_0242_));
 sg13g2_nor2_2 _4362_ (.A(_0242_),
    .B(net20),
    .Y(_0243_));
 sg13g2_inv_1 _4363_ (.Y(_0244_),
    .A(_0242_));
 sg13g2_xnor2_1 _4364_ (.Y(_0245_),
    .A(_2153_),
    .B(_2182_));
 sg13g2_nor2_1 _4365_ (.A(_0244_),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_nor2_2 _4366_ (.A(_0243_),
    .B(_0246_),
    .Y(_0247_));
 sg13g2_nand3_1 _4367_ (.B(_0241_),
    .C(_0247_),
    .A(_0236_),
    .Y(_0248_));
 sg13g2_nand2_1 _4368_ (.Y(_0249_),
    .A(net19),
    .B(_0039_));
 sg13g2_nor2_1 _4369_ (.A(_0039_),
    .B(net19),
    .Y(_0250_));
 sg13g2_a21oi_1 _4370_ (.A1(_0249_),
    .A2(_0243_),
    .Y(_0251_),
    .B1(_0250_));
 sg13g2_nand2_1 _4371_ (.Y(_0252_),
    .A(_0248_),
    .B(_0251_));
 sg13g2_nand2b_1 _4372_ (.Y(_0253_),
    .B(_0252_),
    .A_N(_0232_));
 sg13g2_nand3_1 _4373_ (.B(_0232_),
    .C(_0251_),
    .A(_0248_),
    .Y(_0254_));
 sg13g2_nand3_1 _4374_ (.B(_0254_),
    .C(net48),
    .A(_0253_),
    .Y(_0255_));
 sg13g2_xnor2_1 _4375_ (.Y(_0256_),
    .A(_1684_),
    .B(_0164_));
 sg13g2_a21oi_1 _4376_ (.A1(_0256_),
    .A2(_2101_),
    .Y(_0257_),
    .B1(_2025_));
 sg13g2_inv_1 _4377_ (.Y(_0258_),
    .A(_0257_));
 sg13g2_nand2_1 _4378_ (.Y(_0259_),
    .A(_0255_),
    .B(_0258_));
 sg13g2_xnor2_1 _4379_ (.Y(_0260_),
    .A(_1694_),
    .B(net19));
 sg13g2_inv_1 _4380_ (.Y(_0261_),
    .A(_0260_));
 sg13g2_a21oi_1 _4381_ (.A1(_0261_),
    .A2(_2108_),
    .Y(_0262_),
    .B1(_2112_));
 sg13g2_nand2_1 _4382_ (.Y(_0263_),
    .A(_0259_),
    .B(_0262_));
 sg13g2_nor2b_1 _4383_ (.A(net57),
    .B_N(_0051_),
    .Y(_0264_));
 sg13g2_a21oi_1 _4384_ (.A1(net57),
    .A2(_0048_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_nand2_1 _4385_ (.Y(_0266_),
    .A(_0024_),
    .B(_2132_));
 sg13g2_o21ai_1 _4386_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_2132_),
    .A2(_1750_));
 sg13g2_nor2_1 _4387_ (.A(net55),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_a21o_1 _4388_ (.A2(_0265_),
    .A1(net55),
    .B1(_0268_),
    .X(_0269_));
 sg13g2_buf_1 _4389_ (.A(_0269_),
    .X(_0270_));
 sg13g2_xnor2_1 _4390_ (.Y(_0271_),
    .A(_0270_),
    .B(_2130_));
 sg13g2_a21oi_1 _4391_ (.A1(_0271_),
    .A2(net40),
    .Y(_0272_),
    .B1(_2117_));
 sg13g2_nand2_1 _4392_ (.Y(_0273_),
    .A(_0263_),
    .B(_0272_));
 sg13g2_a21oi_1 _4393_ (.A1(_0270_),
    .A2(net39),
    .Y(_0274_),
    .B1(_2147_));
 sg13g2_nand2_1 _4394_ (.Y(_0275_),
    .A(_0273_),
    .B(_0274_));
 sg13g2_inv_4 _4395_ (.A(_0176_),
    .Y(_0276_));
 sg13g2_nand2_1 _4396_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_buf_8 _4397_ (.A(_0197_),
    .X(_0278_));
 sg13g2_nand2_1 _4398_ (.Y(_0279_),
    .A(_0277_),
    .B(net38));
 sg13g2_nand2_1 _4399_ (.Y(_0280_),
    .A(_1764_),
    .B(_0050_));
 sg13g2_buf_1 _4400_ (.A(_0280_),
    .X(_0281_));
 sg13g2_nand3_1 _4401_ (.B(_0199_),
    .C(_0281_),
    .A(_0279_),
    .Y(_0282_));
 sg13g2_nor2_1 _4402_ (.A(_0214_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_nor2_1 _4403_ (.A(_0211_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_nand2_1 _4404_ (.Y(_0285_),
    .A(_0227_),
    .B(_0215_));
 sg13g2_nand2_1 _4405_ (.Y(_0286_),
    .A(_1662_),
    .B(_2004_));
 sg13g2_nand2_1 _4406_ (.Y(_0287_),
    .A(_0285_),
    .B(_0286_));
 sg13g2_nand2_1 _4407_ (.Y(_0288_),
    .A(_0168_),
    .B(_0019_));
 sg13g2_inv_1 _4408_ (.Y(_0289_),
    .A(_0019_));
 sg13g2_nand3_1 _4409_ (.B(_0166_),
    .C(_0289_),
    .A(_2170_),
    .Y(_0290_));
 sg13g2_buf_1 _4410_ (.A(_0290_),
    .X(_0291_));
 sg13g2_nor2_1 _4411_ (.A(net60),
    .B(\i_project.controller_0.t[10] ),
    .Y(_0292_));
 sg13g2_nand2_1 _4412_ (.Y(_0293_),
    .A(_1663_),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_nor2b_1 _4413_ (.A(_0292_),
    .B_N(_0293_),
    .Y(_0294_));
 sg13g2_nand3_1 _4414_ (.B(_0291_),
    .C(_0294_),
    .A(_0288_),
    .Y(_0295_));
 sg13g2_nand2_1 _4415_ (.Y(_0296_),
    .A(_0168_),
    .B(_0289_));
 sg13g2_nand3_1 _4416_ (.B(_0166_),
    .C(_0019_),
    .A(_2170_),
    .Y(_0297_));
 sg13g2_inv_1 _4417_ (.Y(_0298_),
    .A(_0294_));
 sg13g2_nand3_1 _4418_ (.B(_0297_),
    .C(_0298_),
    .A(_0296_),
    .Y(_0299_));
 sg13g2_nand2_1 _4419_ (.Y(_0300_),
    .A(_0295_),
    .B(_0299_));
 sg13g2_xnor2_1 _4420_ (.Y(_0301_),
    .A(_0287_),
    .B(_0300_));
 sg13g2_nand2_1 _4421_ (.Y(_0302_),
    .A(_0247_),
    .B(_2058_));
 sg13g2_nand2_1 _4422_ (.Y(_0303_),
    .A(_0231_),
    .B(_0241_));
 sg13g2_nor3_1 _4423_ (.A(_2093_),
    .B(_0302_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_inv_1 _4424_ (.Y(_0305_),
    .A(_0304_));
 sg13g2_inv_1 _4425_ (.Y(_0306_),
    .A(_0243_));
 sg13g2_o21ai_1 _4426_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_0235_),
    .A2(_0246_));
 sg13g2_dfrbp_1 _4427_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net83),
    .D(_0000_),
    .Q_N(_2255_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _4428_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net84),
    .D(_0001_),
    .Q_N(_2256_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _4429_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0002_),
    .Q_N(_2254_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4430_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net86),
    .D(_0057_),
    .Q_N(_2257_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _4431_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net87),
    .D(_0003_),
    .Q_N(_2253_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4432_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_0004_),
    .Q_N(_2252_),
    .Q(_0144_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4427__83 (.L_HI(net83));
 sg13g2_buf_1 _4435_ (.A(net89),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4436_ (.A(net90),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4437_ (.A(net91),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4438_ (.A(net92),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4439_ (.A(net93),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4440_ (.A(net94),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4441_ (.A(net95),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4442_ (.A(net96),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4443_ (.A(net75),
    .X(uio_out[0]));
 sg13g2_buf_1 _4444_ (.A(net76),
    .X(uio_out[1]));
 sg13g2_buf_1 _4445_ (.A(net77),
    .X(uio_out[2]));
 sg13g2_buf_1 _4446_ (.A(net78),
    .X(uio_out[3]));
 sg13g2_buf_1 _4447_ (.A(net79),
    .X(uio_out[4]));
 sg13g2_buf_1 _4448_ (.A(net80),
    .X(uio_out[5]));
 sg13g2_buf_1 _4449_ (.A(net81),
    .X(uio_out[6]));
 sg13g2_buf_1 _4450_ (.A(net82),
    .X(uio_out[7]));
 sg13g2_buf_1 _4451_ (.A(\i_project.controller_0.vga_sync.o_vsync ),
    .X(net11));
 sg13g2_buf_1 _4452_ (.A(hsync),
    .X(net15));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net97),
    .D(_0058_),
    .Q_N(_0055_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[10]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net98),
    .D(_0059_),
    .Q_N(_2251_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 \counter[11]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net99),
    .D(_0060_),
    .Q_N(_2250_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 \counter[12]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(_0061_),
    .Q_N(_2249_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 \counter[13]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net101),
    .D(_0062_),
    .Q_N(_2248_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 \counter[14]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(_0063_),
    .Q_N(_2247_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 \counter[15]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_0064_),
    .Q_N(_2246_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 \counter[16]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net104),
    .D(_0065_),
    .Q_N(_2245_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 \counter[17]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net105),
    .D(_0066_),
    .Q_N(_2244_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 \counter[18]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net106),
    .D(_0067_),
    .Q_N(_2243_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 \counter[19]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net107),
    .D(_0068_),
    .Q_N(_2242_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net108),
    .D(_0069_),
    .Q_N(_2241_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[20]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net109),
    .D(_0070_),
    .Q_N(_2240_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 \counter[21]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_2239_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 \counter[22]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net111),
    .D(_0072_),
    .Q_N(_2238_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 \counter[23]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net112),
    .D(_0073_),
    .Q_N(_2237_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 \counter[24]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net113),
    .D(_0074_),
    .Q_N(_2236_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 \counter[25]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net114),
    .D(_0075_),
    .Q_N(_2235_),
    .Q(\counter[25] ));
 sg13g2_dfrbp_1 \counter[26]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net115),
    .D(_0076_),
    .Q_N(_2234_),
    .Q(\counter[26] ));
 sg13g2_dfrbp_1 \counter[27]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net116),
    .D(_0077_),
    .Q_N(_2233_),
    .Q(\counter[27] ));
 sg13g2_dfrbp_1 \counter[28]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net117),
    .D(_0078_),
    .Q_N(_2232_),
    .Q(\counter[28] ));
 sg13g2_dfrbp_1 \counter[29]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net118),
    .D(_0079_),
    .Q_N(_2231_),
    .Q(\counter[29] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net119),
    .D(_0080_),
    .Q_N(_2230_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[30]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net120),
    .D(_0081_),
    .Q_N(_2229_),
    .Q(\counter[30] ));
 sg13g2_dfrbp_1 \counter[31]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net121),
    .D(_0082_),
    .Q_N(_2228_),
    .Q(\counter[31] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net122),
    .D(_0083_),
    .Q_N(_2227_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net123),
    .D(_0084_),
    .Q_N(_2226_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net124),
    .D(_0085_),
    .Q_N(_2225_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net125),
    .D(_0086_),
    .Q_N(_2224_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net126),
    .D(_0087_),
    .Q_N(_2223_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net127),
    .D(_0088_),
    .Q_N(_2222_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net128),
    .D(_0089_),
    .Q_N(_2258_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \depth[0]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net129),
    .D(_0005_),
    .Q_N(_2259_),
    .Q(\depth[0] ));
 sg13g2_dfrbp_1 \depth[1]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_0006_),
    .Q_N(_2260_),
    .Q(\depth[1] ));
 sg13g2_dfrbp_1 \depth[2]$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(_0007_),
    .Q_N(_0046_),
    .Q(\depth[2] ));
 sg13g2_dfrbp_1 \dither_threshold[0]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net132),
    .D(_0090_),
    .Q_N(_0022_),
    .Q(\dither_threshold[0] ));
 sg13g2_dfrbp_1 \dither_threshold[1]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_0091_),
    .Q_N(_0031_),
    .Q(\dither_threshold[1] ));
 sg13g2_dfrbp_1 \dither_threshold[2]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0092_),
    .Q_N(_2221_),
    .Q(\dither_threshold[2] ));
 sg13g2_dfrbp_1 \dither_threshold[3]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net135),
    .D(_0093_),
    .Q_N(_0032_),
    .Q(\dither_threshold[3] ));
 sg13g2_dfrbp_1 \dither_threshold[4]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net136),
    .D(_0094_),
    .Q_N(_0033_),
    .Q(\dither_threshold[4] ));
 sg13g2_dfrbp_1 \dither_threshold[5]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net137),
    .D(_0095_),
    .Q_N(_0034_),
    .Q(\dither_threshold[5] ));
 sg13g2_dfrbp_1 \dither_threshold[6]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net138),
    .D(_0096_),
    .Q_N(_0035_),
    .Q(\dither_threshold[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[2]$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net139),
    .D(_0003_),
    .Q_N(_2220_),
    .Q(\i_project.controller_0.divider[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[3]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net140),
    .D(_0004_),
    .Q_N(_2219_),
    .Q(\i_project.controller_0.divider[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[4]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(_0097_),
    .Q_N(_2218_),
    .Q(\i_project.controller_0.mode[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[5]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net142),
    .D(_0098_),
    .Q_N(_2217_),
    .Q(\i_project.controller_0.mode[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[6]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net143),
    .D(_0099_),
    .Q_N(_0027_),
    .Q(\i_project.controller_0.mode[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[7]$_DFFE_PN_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net144),
    .D(_0100_),
    .Q_N(_0025_),
    .Q(\i_project.controller_0.vga_sync.mode ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[0]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net145),
    .D(_0101_),
    .Q_N(_0056_),
    .Q(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[10]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net146),
    .D(_0102_),
    .Q_N(_0019_),
    .Q(\i_project.controller_0.t[10] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[11]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net147),
    .D(_0103_),
    .Q_N(_2216_),
    .Q(\i_project.controller_0.t[11] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[1]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net148),
    .D(_0104_),
    .Q_N(_0021_),
    .Q(\i_project.controller_0.mode_ramp_base[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[2]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net149),
    .D(_0105_),
    .Q_N(_0045_),
    .Q(\i_project.controller_0.mode_ramp_base[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[3]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net150),
    .D(_0106_),
    .Q_N(_0044_),
    .Q(\i_project.controller_0.mode_ramp_base[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[4]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net151),
    .D(_0107_),
    .Q_N(_0043_),
    .Q(\i_project.controller_0.mode_ramp_base[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[5]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net152),
    .D(_0108_),
    .Q_N(_0042_),
    .Q(\i_project.controller_0.mode_ramp_base[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[6]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net153),
    .D(_0109_),
    .Q_N(_0041_),
    .Q(\i_project.controller_0.mode_ramp_base[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[7]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net154),
    .D(_0110_),
    .Q_N(_0040_),
    .Q(\i_project.controller_0.mode_ramp_base[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[8]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net155),
    .D(_0111_),
    .Q_N(_0039_),
    .Q(\i_project.controller_0.t[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[9]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net156),
    .D(_0112_),
    .Q_N(_0020_),
    .Q(\i_project.controller_0.t[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net157),
    .D(_0113_),
    .Q_N(_0054_),
    .Q(\i_project.controller_0.h[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net158),
    .D(_0114_),
    .Q_N(_0038_),
    .Q(\i_project.controller_0.h[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net159),
    .D(_0115_),
    .Q_N(_0037_),
    .Q(\i_project.controller_0.h[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net160),
    .D(_0116_),
    .Q_N(_0023_),
    .Q(\i_project.controller_0.h[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net161),
    .D(_0117_),
    .Q_N(_0053_),
    .Q(\i_project.controller_0.h[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net162),
    .D(_0118_),
    .Q_N(_0051_),
    .Q(\i_project.controller_0.h[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net163),
    .D(_0119_),
    .Q_N(_0048_),
    .Q(\i_project.controller_0.h[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net164),
    .D(_0120_),
    .Q_N(_0026_),
    .Q(\i_project.controller_0.h[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net165),
    .D(_0121_),
    .Q_N(_0024_),
    .Q(\i_project.controller_0.h[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net166),
    .D(_0122_),
    .Q_N(_0049_),
    .Q(\i_project.controller_0.h[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hsync$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net167),
    .D(_0123_),
    .Q_N(hsync),
    .Q(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net168),
    .D(_0124_),
    .Q_N(_2215_),
    .Q(\i_project.controller_0.v[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net169),
    .D(_0125_),
    .Q_N(_2214_),
    .Q(\i_project.controller_0.v[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net170),
    .D(_0126_),
    .Q_N(_2213_),
    .Q(\i_project.controller_0.v[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net171),
    .D(_0127_),
    .Q_N(_2212_),
    .Q(\i_project.controller_0.v[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net172),
    .D(_0128_),
    .Q_N(_2211_),
    .Q(\i_project.controller_0.v[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net173),
    .D(_0129_),
    .Q_N(_0029_),
    .Q(\i_project.controller_0.v[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net174),
    .D(_0130_),
    .Q_N(_2210_),
    .Q(\i_project.controller_0.v[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net175),
    .D(_0131_),
    .Q_N(_2209_),
    .Q(\i_project.controller_0.v[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net176),
    .D(_0132_),
    .Q_N(_0030_),
    .Q(\i_project.controller_0.v[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net177),
    .D(_0133_),
    .Q_N(_0028_),
    .Q(\i_project.controller_0.v[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vsync$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net178),
    .D(_0134_),
    .Q_N(_2208_),
    .Q(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[0]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net179),
    .D(_0135_),
    .Q_N(_2207_),
    .Q(\i_project.controller_0.voffset[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[1]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net180),
    .D(_0136_),
    .Q_N(_2206_),
    .Q(\i_project.controller_0.voffset[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[2]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net181),
    .D(_0137_),
    .Q_N(_2205_),
    .Q(\i_project.controller_0.voffset[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net182),
    .D(_0138_),
    .Q_N(_2204_),
    .Q(\i_project.controller_0.voffset[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net183),
    .D(_0139_),
    .Q_N(_2203_),
    .Q(\i_project.controller_0.voffset[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[5]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net184),
    .D(_0140_),
    .Q_N(_2202_),
    .Q(\i_project.controller_0.voffset[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[6]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net185),
    .D(_0141_),
    .Q_N(_2201_),
    .Q(\i_project.controller_0.voffset[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[7]$_SDFFCE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net186),
    .D(_0142_),
    .Q_N(_2261_),
    .Q(\i_project.controller_0.voffset[7] ));
 sg13g2_dfrbp_1 \project_rst_n$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net187),
    .D(_0008_),
    .Q_N(_2262_),
    .Q(\i_project.controller_0.rst_n ));
 sg13g2_dfrbp_1 \project_ui_in[2]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net188),
    .D(\counter[30] ),
    .Q_N(_0018_),
    .Q(\i_project.controller_0.grey_pass[10] ));
 sg13g2_dfrbp_1 \project_ui_in[3]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net189),
    .D(\counter[31] ),
    .Q_N(_0017_),
    .Q(\i_project.controller_0.grey_pass[11] ));
 sg13g2_dfrbp_1 \project_ui_in[4]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net190),
    .D(_0009_),
    .Q_N(_0052_),
    .Q(\i_project.controller_0.grey_pass[12] ));
 sg13g2_dfrbp_1 \project_ui_in[5]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net191),
    .D(_0010_),
    .Q_N(_0050_),
    .Q(\i_project.controller_0.grey_pass[13] ));
 sg13g2_dfrbp_1 \project_ui_in[6]$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net192),
    .D(_0011_),
    .Q_N(_0047_),
    .Q(\i_project.controller_0.grey_pass[14] ));
 sg13g2_dfrbp_1 \project_ui_in[7]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net193),
    .D(_0143_),
    .Q_N(_0036_),
    .Q(\i_project.controller_0.grey_pass[15] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout16 (.A(_0470_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0408_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0164_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0154_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0145_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1865_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_2098_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0210_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_2148_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_2131_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0422_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0405_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2147_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2130_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0434_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0430_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0418_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2144_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2119_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2113_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2068_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0281_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0278_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_2118_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2112_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2027_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0786_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0410_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0359_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2117_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2109_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2101_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2026_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1765_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2108_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1977_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1948_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1927_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1785_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1584_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0400_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2132_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2016_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1985_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1685_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1684_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1674_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1672_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1667_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1655_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1652_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1588_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1578_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1987_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1980_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1711_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1702_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1668_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1647_),
    .X(net74));
 sg13g2_tielo _4443__75 (.L_LO(net75));
 sg13g2_tielo _4444__76 (.L_LO(net76));
 sg13g2_tielo _4445__77 (.L_LO(net77));
 sg13g2_tielo _4446__78 (.L_LO(net78));
 sg13g2_tielo _4447__79 (.L_LO(net79));
 sg13g2_tielo _4448__80 (.L_LO(net80));
 sg13g2_tielo _4449__81 (.L_LO(net81));
 sg13g2_tielo _4450__82 (.L_LO(net82));
 sg13g2_tiehi _4428__84 (.L_HI(net84));
 sg13g2_tiehi _4429__85 (.L_HI(net85));
 sg13g2_tiehi _4430__86 (.L_HI(net86));
 sg13g2_tiehi _4431__87 (.L_HI(net87));
 sg13g2_tiehi _4432__88 (.L_HI(net88));
 sg13g2_tiehi _4435__89 (.L_HI(net89));
 sg13g2_tiehi _4436__90 (.L_HI(net90));
 sg13g2_tiehi _4437__91 (.L_HI(net91));
 sg13g2_tiehi _4438__92 (.L_HI(net92));
 sg13g2_tiehi _4439__93 (.L_HI(net93));
 sg13g2_tiehi _4440__94 (.L_HI(net94));
 sg13g2_tiehi _4441__95 (.L_HI(net95));
 sg13g2_tiehi _4442__96 (.L_HI(net96));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \counter[10]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \counter[11]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \counter[12]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \counter[13]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter[14]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[15]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[16]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[17]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[18]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[19]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[20]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[21]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \counter[22]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \counter[23]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \counter[24]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \counter[25]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \counter[26]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \counter[27]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \counter[28]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \counter[29]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \counter[30]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \counter[31]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \depth[0]$_DFF_P__129  (.L_HI(net129));
 sg13g2_tiehi \depth[1]$_DFF_P__130  (.L_HI(net130));
 sg13g2_tiehi \depth[2]$_DFF_P__131  (.L_HI(net131));
 sg13g2_tiehi \dither_threshold[0]$_SDFFE_PP0P__132  (.L_HI(net132));
 sg13g2_tiehi \dither_threshold[1]$_SDFF_PP0__133  (.L_HI(net133));
 sg13g2_tiehi \dither_threshold[2]$_SDFF_PP0__134  (.L_HI(net134));
 sg13g2_tiehi \dither_threshold[3]$_SDFF_PP0__135  (.L_HI(net135));
 sg13g2_tiehi \dither_threshold[4]$_SDFF_PP0__136  (.L_HI(net136));
 sg13g2_tiehi \dither_threshold[5]$_SDFF_PP0__137  (.L_HI(net137));
 sg13g2_tiehi \dither_threshold[6]$_SDFF_PP0__138  (.L_HI(net138));
 sg13g2_tiehi \i_project.controller_0.mode_params[2]$_DFFE_PN__139  (.L_HI(net139));
 sg13g2_tiehi \i_project.controller_0.mode_params[3]$_DFFE_PN__140  (.L_HI(net140));
 sg13g2_tiehi \i_project.controller_0.mode_params[4]$_DFFE_PN__141  (.L_HI(net141));
 sg13g2_tiehi \i_project.controller_0.mode_params[5]$_DFFE_PN__142  (.L_HI(net142));
 sg13g2_tiehi \i_project.controller_0.mode_params[6]$_DFFE_PN__143  (.L_HI(net143));
 sg13g2_tiehi \i_project.controller_0.mode_params[7]$_DFFE_PN__144  (.L_HI(net144));
 sg13g2_tiehi \i_project.controller_0.t[0]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \i_project.controller_0.t[10]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \i_project.controller_0.t[11]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \i_project.controller_0.t[1]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \i_project.controller_0.t[2]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \i_project.controller_0.t[3]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \i_project.controller_0.t[4]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \i_project.controller_0.t[5]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \i_project.controller_0.t[6]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \i_project.controller_0.t[7]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \i_project.controller_0.t[8]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \i_project.controller_0.t[9]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0__157  (.L_HI(net157));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0__158  (.L_HI(net158));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0__159  (.L_HI(net159));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0__161  (.L_HI(net161));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0__162  (.L_HI(net162));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0__163  (.L_HI(net163));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0__164  (.L_HI(net164));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hsync$_DFFE_PP__167  (.L_HI(net167));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P__168  (.L_HI(net168));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P__169  (.L_HI(net169));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P__170  (.L_HI(net170));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vsync$_DFFE_PP__178  (.L_HI(net178));
 sg13g2_tiehi \i_project.controller_0.voffset[0]$_DFFE_PP__179  (.L_HI(net179));
 sg13g2_tiehi \i_project.controller_0.voffset[1]$_DFFE_PP__180  (.L_HI(net180));
 sg13g2_tiehi \i_project.controller_0.voffset[2]$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \i_project.controller_0.voffset[3]$_SDFFCE_PP0P__182  (.L_HI(net182));
 sg13g2_tiehi \i_project.controller_0.voffset[4]$_SDFFCE_PP0P__183  (.L_HI(net183));
 sg13g2_tiehi \i_project.controller_0.voffset[5]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \i_project.controller_0.voffset[6]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \i_project.controller_0.voffset[7]$_SDFFCE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \project_rst_n$_DFF_P__187  (.L_HI(net187));
 sg13g2_tiehi \project_ui_in[2]$_DFF_P__188  (.L_HI(net188));
 sg13g2_tiehi \project_ui_in[3]$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \project_ui_in[4]$_DFF_P__190  (.L_HI(net190));
 sg13g2_tiehi \project_ui_in[5]$_DFF_P__191  (.L_HI(net191));
 sg13g2_tiehi \project_ui_in[6]$_DFF_P__192  (.L_HI(net192));
 sg13g2_tiehi \project_ui_in[7]$_SDFF_PN0__193  (.L_HI(net193));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_fill_2 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_30 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_4 FILLER_0_77 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_fill_2 FILLER_0_96 ();
 sg13g2_fill_2 FILLER_0_102 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_154 ();
 sg13g2_fill_1 FILLER_0_159 ();
 sg13g2_fill_1 FILLER_0_195 ();
 sg13g2_fill_2 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_fill_2 FILLER_0_287 ();
 sg13g2_fill_1 FILLER_0_306 ();
 sg13g2_fill_1 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_4 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_23 ();
 sg13g2_fill_1 FILLER_1_40 ();
 sg13g2_decap_4 FILLER_1_53 ();
 sg13g2_fill_1 FILLER_1_57 ();
 sg13g2_fill_2 FILLER_1_78 ();
 sg13g2_fill_2 FILLER_1_87 ();
 sg13g2_fill_1 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_129 ();
 sg13g2_decap_4 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_fill_2 FILLER_1_161 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_176 ();
 sg13g2_fill_1 FILLER_1_198 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_212 ();
 sg13g2_fill_1 FILLER_1_221 ();
 sg13g2_fill_2 FILLER_1_226 ();
 sg13g2_fill_2 FILLER_1_233 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_fill_2 FILLER_1_245 ();
 sg13g2_fill_1 FILLER_1_251 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_fill_1 FILLER_1_262 ();
 sg13g2_fill_2 FILLER_1_286 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_312 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_1 FILLER_1_332 ();
 sg13g2_fill_2 FILLER_1_339 ();
 sg13g2_decap_4 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_fill_2 FILLER_1_366 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_23 ();
 sg13g2_fill_1 FILLER_2_36 ();
 sg13g2_fill_1 FILLER_2_41 ();
 sg13g2_fill_1 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_58 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_fill_1 FILLER_2_65 ();
 sg13g2_decap_4 FILLER_2_83 ();
 sg13g2_fill_2 FILLER_2_96 ();
 sg13g2_fill_1 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_151 ();
 sg13g2_fill_1 FILLER_2_158 ();
 sg13g2_fill_2 FILLER_2_167 ();
 sg13g2_fill_1 FILLER_2_173 ();
 sg13g2_fill_1 FILLER_2_178 ();
 sg13g2_fill_1 FILLER_2_182 ();
 sg13g2_fill_2 FILLER_2_195 ();
 sg13g2_fill_1 FILLER_2_197 ();
 sg13g2_decap_4 FILLER_2_201 ();
 sg13g2_decap_4 FILLER_2_221 ();
 sg13g2_fill_1 FILLER_2_236 ();
 sg13g2_decap_4 FILLER_2_253 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_fill_2 FILLER_2_279 ();
 sg13g2_fill_2 FILLER_2_286 ();
 sg13g2_decap_4 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_306 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_fill_2 FILLER_2_319 ();
 sg13g2_fill_1 FILLER_2_321 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_331 ();
 sg13g2_fill_2 FILLER_2_355 ();
 sg13g2_decap_4 FILLER_2_365 ();
 sg13g2_fill_1 FILLER_2_378 ();
 sg13g2_decap_4 FILLER_2_383 ();
 sg13g2_fill_1 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_fill_2 FILLER_2_403 ();
 sg13g2_decap_4 FILLER_2_409 ();
 sg13g2_fill_1 FILLER_2_413 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_9 ();
 sg13g2_fill_2 FILLER_3_54 ();
 sg13g2_fill_1 FILLER_3_56 ();
 sg13g2_fill_1 FILLER_3_115 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_fill_1 FILLER_3_151 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_178 ();
 sg13g2_fill_2 FILLER_3_201 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_fill_1 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_285 ();
 sg13g2_fill_2 FILLER_3_299 ();
 sg13g2_decap_4 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_309 ();
 sg13g2_fill_1 FILLER_3_317 ();
 sg13g2_fill_1 FILLER_3_327 ();
 sg13g2_fill_1 FILLER_3_357 ();
 sg13g2_decap_4 FILLER_3_386 ();
 sg13g2_decap_4 FILLER_3_394 ();
 sg13g2_fill_2 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_412 ();
 sg13g2_fill_1 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_22 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_decap_4 FILLER_4_34 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_fill_1 FILLER_4_51 ();
 sg13g2_fill_2 FILLER_4_83 ();
 sg13g2_fill_2 FILLER_4_93 ();
 sg13g2_fill_2 FILLER_4_98 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_fill_2 FILLER_4_113 ();
 sg13g2_fill_2 FILLER_4_118 ();
 sg13g2_fill_2 FILLER_4_124 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_fill_1 FILLER_4_155 ();
 sg13g2_fill_1 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_174 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_211 ();
 sg13g2_fill_1 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_248 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_decap_4 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_263 ();
 sg13g2_fill_2 FILLER_4_299 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_fill_1 FILLER_4_360 ();
 sg13g2_fill_2 FILLER_4_397 ();
 sg13g2_fill_1 FILLER_4_399 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_12 ();
 sg13g2_fill_1 FILLER_5_17 ();
 sg13g2_fill_1 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_2 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_37 ();
 sg13g2_fill_2 FILLER_5_57 ();
 sg13g2_fill_2 FILLER_5_76 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_128 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_fill_1 FILLER_5_185 ();
 sg13g2_fill_2 FILLER_5_205 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_decap_4 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_4 FILLER_5_307 ();
 sg13g2_decap_4 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_349 ();
 sg13g2_decap_4 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_fill_1 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_49 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_64 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_102 ();
 sg13g2_fill_1 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_118 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_170 ();
 sg13g2_fill_2 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_fill_1 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_fill_2 FILLER_6_310 ();
 sg13g2_fill_2 FILLER_6_350 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_fill_1 FILLER_6_383 ();
 sg13g2_fill_1 FILLER_6_416 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_27 ();
 sg13g2_fill_1 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_83 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_109 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_139 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_decap_4 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_4 FILLER_7_242 ();
 sg13g2_fill_1 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_decap_4 FILLER_7_293 ();
 sg13g2_decap_4 FILLER_7_320 ();
 sg13g2_fill_1 FILLER_7_324 ();
 sg13g2_fill_2 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_44 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_fill_2 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_68 ();
 sg13g2_decap_4 FILLER_8_77 ();
 sg13g2_fill_2 FILLER_8_81 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_2 FILLER_8_125 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_241 ();
 sg13g2_fill_2 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_259 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_271 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_decap_4 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_348 ();
 sg13g2_fill_2 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_decap_4 FILLER_8_362 ();
 sg13g2_fill_2 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_8_372 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_19 ();
 sg13g2_decap_4 FILLER_9_38 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_4 FILLER_9_81 ();
 sg13g2_decap_4 FILLER_9_89 ();
 sg13g2_fill_1 FILLER_9_93 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_138 ();
 sg13g2_fill_2 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_4 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_2 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_fill_2 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_fill_2 FILLER_9_337 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_fill_2 FILLER_9_393 ();
 sg13g2_fill_2 FILLER_9_402 ();
 sg13g2_fill_2 FILLER_10_32 ();
 sg13g2_fill_2 FILLER_10_52 ();
 sg13g2_fill_1 FILLER_10_54 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_decap_4 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_226 ();
 sg13g2_fill_1 FILLER_10_230 ();
 sg13g2_decap_4 FILLER_10_236 ();
 sg13g2_fill_1 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_4 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_188 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_fill_1 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_365 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_34 ();
 sg13g2_fill_2 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_4 FILLER_12_113 ();
 sg13g2_fill_1 FILLER_12_117 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_160 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_2 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_decap_4 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_390 ();
 sg13g2_fill_1 FILLER_12_409 ();
 sg13g2_fill_2 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_419 ();
 sg13g2_decap_4 FILLER_12_426 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_43 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_122 ();
 sg13g2_fill_2 FILLER_13_128 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_310 ();
 sg13g2_fill_2 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_decap_4 FILLER_13_349 ();
 sg13g2_decap_4 FILLER_13_356 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_369 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_396 ();
 sg13g2_fill_1 FILLER_13_407 ();
 sg13g2_fill_1 FILLER_13_415 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_53 ();
 sg13g2_decap_4 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_62 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_2 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_fill_2 FILLER_14_197 ();
 sg13g2_decap_4 FILLER_14_223 ();
 sg13g2_fill_2 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_decap_4 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_38 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_122 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_decap_4 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_fill_2 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_363 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_18 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_47 ();
 sg13g2_decap_4 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_60 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_2 FILLER_16_193 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_fill_1 FILLER_16_421 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_6 ();
 sg13g2_fill_1 FILLER_17_13 ();
 sg13g2_fill_1 FILLER_17_22 ();
 sg13g2_fill_1 FILLER_17_50 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_fill_1 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_17_412 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_2 FILLER_18_83 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_341 ();
 sg13g2_fill_1 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_fill_2 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_13 ();
 sg13g2_fill_1 FILLER_20_15 ();
 sg13g2_fill_2 FILLER_20_20 ();
 sg13g2_fill_1 FILLER_20_22 ();
 sg13g2_fill_2 FILLER_20_50 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_decap_4 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_153 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_4 FILLER_20_190 ();
 sg13g2_decap_4 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_4 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_fill_1 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_decap_4 FILLER_21_37 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_4 FILLER_21_93 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_218 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_394 ();
 sg13g2_decap_4 FILLER_21_418 ();
 sg13g2_fill_2 FILLER_21_422 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_decap_4 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_1 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_decap_4 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_129 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_decap_8 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_decap_4 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_decap_4 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_374 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_15 ();
 sg13g2_decap_8 FILLER_23_22 ();
 sg13g2_decap_8 FILLER_23_29 ();
 sg13g2_decap_8 FILLER_23_36 ();
 sg13g2_decap_8 FILLER_23_47 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_422 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_67 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_4 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_decap_4 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_394 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_decap_4 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_decap_4 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_416 ();
 sg13g2_fill_2 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_26_3 ();
 sg13g2_fill_2 FILLER_26_19 ();
 sg13g2_decap_4 FILLER_26_32 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_decap_8 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_193 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_decap_4 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_397 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_11 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_decap_4 FILLER_27_186 ();
 sg13g2_decap_4 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_57 ();
 sg13g2_decap_4 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_79 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_decap_8 FILLER_28_93 ();
 sg13g2_decap_8 FILLER_28_100 ();
 sg13g2_decap_4 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_409 ();
 sg13g2_fill_2 FILLER_28_415 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_15 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_4 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_4 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_38 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_60 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_397 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_decap_4 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_78 ();
 sg13g2_decap_8 FILLER_31_97 ();
 sg13g2_decap_4 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_32_3 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_decap_4 FILLER_32_183 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_decap_4 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_121 ();
 sg13g2_fill_1 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_11 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_71 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_decap_4 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_421 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_fill_1 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_51 ();
 sg13g2_fill_1 FILLER_36_66 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_138 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_43 ();
 sg13g2_fill_1 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_1 FILLER_38_50 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_decap_4 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_402 ();
endmodule
