module tt_um_MichaelBell_canon (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire clknet_0_clk;
 wire net180;
 wire \crotchet[0] ;
 wire \crotchet[1] ;
 wire \crotchet[2] ;
 wire \crotchet[3] ;
 wire \crotchet[4] ;
 wire \crotchet[5] ;
 wire \crotchet[6] ;
 wire \i_display.colour[0] ;
 wire \i_display.colour[1] ;
 wire \i_display.colour[2] ;
 wire \i_display.colour[3] ;
 wire \i_display.colour[4] ;
 wire \i_display.colour[5] ;
 wire \i_display.frame[0] ;
 wire \i_display.frame[1] ;
 wire \i_display.frame[2] ;
 wire \i_display.frame[3] ;
 wire \i_display.frame[4] ;
 wire \i_display.frame[5] ;
 wire \i_display.frame[6] ;
 wire \i_display.frame[7] ;
 wire \i_display.frame[8] ;
 wire \i_display.frame[9] ;
 wire \i_display.frame_crotchet[0] ;
 wire \i_display.frame_crotchet[1] ;
 wire \i_display.frame_crotchet[2] ;
 wire \i_display.frame_crotchet[3] ;
 wire \i_display.frame_crotchet[4] ;
 wire \i_display.frame_crotchet[5] ;
 wire \i_display.frame_crotchet[6] ;
 wire \i_display.hsync ;
 wire \i_display.i_vga.hblank ;
 wire \i_display.i_vga.hblank_tmp ;
 wire \i_display.i_vga.hsync_tmp ;
 wire \i_display.i_vga.low_count[0] ;
 wire \i_display.i_vga.low_count[1] ;
 wire \i_display.i_vga.low_count[2] ;
 wire \i_display.i_vga.low_count[3] ;
 wire \i_display.i_vga.low_count[4] ;
 wire \i_display.i_vga.low_count[5] ;
 wire \i_display.i_vga.low_count[6] ;
 wire \i_display.i_vga.low_count[7] ;
 wire \i_display.i_vga.low_count[8] ;
 wire \i_display.i_vga.low_count[9] ;
 wire \i_display.i_vga.timing_ver.blank ;
 wire \i_display.i_vga.timing_ver.counter[0] ;
 wire \i_display.i_vga.timing_ver.counter[10] ;
 wire \i_display.i_vga.timing_ver.counter[1] ;
 wire \i_display.i_vga.timing_ver.counter[2] ;
 wire \i_display.i_vga.timing_ver.counter[3] ;
 wire \i_display.i_vga.timing_ver.counter[4] ;
 wire \i_display.i_vga.timing_ver.counter[5] ;
 wire \i_display.i_vga.timing_ver.counter[6] ;
 wire \i_display.i_vga.timing_ver.counter[7] ;
 wire \i_display.i_vga.timing_ver.counter[8] ;
 wire \i_display.i_vga.timing_ver.counter[9] ;
 wire \i_display.i_vga.timing_ver.sync ;
 wire \i_display.i_vga.timing_ver.sync_tmp ;
 wire \i_display.i_vga.vblank ;
 wire \i_display.in_line ;
 wire \i_display.x_idx[0] ;
 wire \i_display.x_idx[1] ;
 wire \i_display.x_idx[2] ;
 wire \i_display.x_idx[3] ;
 wire \i_display.x_idx[4] ;
 wire \i_display.x_idx[5] ;
 wire \i_display.x_idx[6] ;
 wire \i_display.x_idx[7] ;
 wire \i_display.x_idx[8] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-1] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-2] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-3] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-4] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-5] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[0] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[1] ;
 wire \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[2] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[0] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[1] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[2] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[3] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[4] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[5] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[6] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[7] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[8] ;
 wire \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[9] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[2] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[5] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[6] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7] ;
 wire \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8] ;
 wire \i_music.count[10] ;
 wire \i_music.count[11] ;
 wire \i_music.count[12] ;
 wire \i_music.count[13] ;
 wire \i_music.count[14] ;
 wire \i_music.count[15] ;
 wire \i_music.count[16] ;
 wire \i_music.count[17] ;
 wire \i_music.count[18] ;
 wire \i_music.count[19] ;
 wire \i_music.count[20] ;
 wire \i_music.count[21] ;
 wire \i_music.count[22] ;
 wire \i_music.count[23] ;
 wire \i_music.count[24] ;
 wire \i_music.i_pwm.count[0] ;
 wire \i_music.i_pwm.count[1] ;
 wire \i_music.i_pwm.count[2] ;
 wire \i_music.i_pwm.count[3] ;
 wire \i_music.i_pwm.count[4] ;
 wire \i_music.i_pwm.count[5] ;
 wire \i_music.i_pwm.count[6] ;
 wire \i_music.i_pwm.count[7] ;
 wire \i_music.i_pwm.pwm ;
 wire \i_music.i_pwm.sample[0] ;
 wire \i_music.i_pwm.sample[1] ;
 wire \i_music.i_pwm.sample[2] ;
 wire \i_music.i_pwm.sample[3] ;
 wire \i_music.i_pwm.sample[4] ;
 wire \i_music.i_pwm.sample[5] ;
 wire \i_music.i_pwm.sample[6] ;
 wire \i_music.i_pwm.sample[7] ;
 wire \i_music.i_sample.sample_acc[0] ;
 wire \i_music.i_sample.sample_acc[1] ;
 wire \i_music.i_sample.sample_acc[2] ;
 wire \i_music.i_sample.sample_acc[3] ;
 wire \i_music.i_sample.sample_acc[4] ;
 wire \i_music.i_sample.sample_acc[5] ;
 wire \i_music.i_sample.sample_acc[6] ;
 wire \i_music.i_sample.sample_acc[7] ;
 wire \i_music.i_sample.sample_acc[8] ;
 wire \i_music.i_sample.sample_idx[0] ;
 wire \i_music.i_sample.sample_idx[1] ;
 wire \i_music.i_sample.sample_idx[2] ;
 wire \i_music.i_sample.sample_idx[3] ;
 wire \i_music.i_sample.sample_idx[4] ;
 wire \i_music.i_sample.sample_idx[5] ;
 wire \i_music.i_sample.sample_idx[6] ;
 wire \i_music.i_sample.sample_idx[7] ;
 wire \i_music.i_sample.t1.CG.GCLK ;
 wire \i_music.i_sample.t1.genblk1[0].state.D ;
 wire \i_music.i_sample.t1.genblk1[0].state.Q ;
 wire \i_music.i_sample.t1.genblk1[10].state.D ;
 wire \i_music.i_sample.t1.genblk1[10].state.Q ;
 wire \i_music.i_sample.t1.genblk1[11].state.D ;
 wire \i_music.i_sample.t1.genblk1[11].state.Q ;
 wire \i_music.i_sample.t1.genblk1[12].state.D ;
 wire \i_music.i_sample.t1.genblk1[12].state.Q ;
 wire \i_music.i_sample.t1.genblk1[13].state.D ;
 wire \i_music.i_sample.t1.genblk1[13].state.Q ;
 wire \i_music.i_sample.t1.genblk1[14].state.D ;
 wire \i_music.i_sample.t1.genblk1[14].state.Q ;
 wire \i_music.i_sample.t1.genblk1[15].state.D ;
 wire \i_music.i_sample.t1.genblk1[15].state.Q ;
 wire \i_music.i_sample.t1.genblk1[16].state.D ;
 wire \i_music.i_sample.t1.genblk1[16].state.Q ;
 wire \i_music.i_sample.t1.genblk1[17].state.D ;
 wire \i_music.i_sample.t1.genblk1[17].state.Q ;
 wire \i_music.i_sample.t1.genblk1[18].state.D ;
 wire \i_music.i_sample.t1.genblk1[18].state.Q ;
 wire \i_music.i_sample.t1.genblk1[1].state.D ;
 wire \i_music.i_sample.t1.genblk1[1].state.Q ;
 wire \i_music.i_sample.t1.genblk1[2].state.D ;
 wire \i_music.i_sample.t1.genblk1[2].state.Q ;
 wire \i_music.i_sample.t1.genblk1[3].state.D ;
 wire \i_music.i_sample.t1.genblk1[3].state.Q ;
 wire \i_music.i_sample.t1.genblk1[4].state.D ;
 wire \i_music.i_sample.t1.genblk1[4].state.Q ;
 wire \i_music.i_sample.t1.genblk1[5].state.D ;
 wire \i_music.i_sample.t1.genblk1[5].state.Q ;
 wire \i_music.i_sample.t1.genblk1[6].state.D ;
 wire \i_music.i_sample.t1.genblk1[6].state.Q ;
 wire \i_music.i_sample.t1.genblk1[7].state.D ;
 wire \i_music.i_sample.t1.genblk1[7].state.Q ;
 wire \i_music.i_sample.t1.genblk1[8].state.D ;
 wire \i_music.i_sample.t1.genblk1[8].state.Q ;
 wire \i_music.i_sample.t1.genblk1[9].state.D ;
 wire \i_music.i_sample.t1.genblk1[9].state.Q ;
 wire \i_music.i_sample.t2.CG.GCLK ;
 wire \i_music.i_sample.t2.genblk1[0].state.Q ;
 wire \i_music.i_sample.t2.genblk1[10].state.Q ;
 wire \i_music.i_sample.t2.genblk1[11].state.Q ;
 wire \i_music.i_sample.t2.genblk1[12].state.Q ;
 wire \i_music.i_sample.t2.genblk1[13].state.Q ;
 wire \i_music.i_sample.t2.genblk1[14].state.Q ;
 wire \i_music.i_sample.t2.genblk1[15].state.Q ;
 wire \i_music.i_sample.t2.genblk1[16].state.Q ;
 wire \i_music.i_sample.t2.genblk1[17].state.Q ;
 wire \i_music.i_sample.t2.genblk1[1].state.Q ;
 wire \i_music.i_sample.t2.genblk1[2].state.Q ;
 wire \i_music.i_sample.t2.genblk1[3].state.Q ;
 wire \i_music.i_sample.t2.genblk1[4].state.Q ;
 wire \i_music.i_sample.t2.genblk1[5].state.Q ;
 wire \i_music.i_sample.t2.genblk1[6].state.Q ;
 wire \i_music.i_sample.t2.genblk1[7].state.Q ;
 wire \i_music.i_sample.t2.genblk1[8].state.Q ;
 wire \i_music.i_sample.t2.genblk1[9].state.Q ;
 wire \i_music.i_sample.t3.CG.GCLK ;
 wire \i_music.i_sample.t3.genblk1[0].state.Q ;
 wire \i_music.i_sample.t3.genblk1[10].state.Q ;
 wire \i_music.i_sample.t3.genblk1[11].state.Q ;
 wire \i_music.i_sample.t3.genblk1[12].state.Q ;
 wire \i_music.i_sample.t3.genblk1[13].state.Q ;
 wire \i_music.i_sample.t3.genblk1[14].state.Q ;
 wire \i_music.i_sample.t3.genblk1[15].state.Q ;
 wire \i_music.i_sample.t3.genblk1[16].state.Q ;
 wire \i_music.i_sample.t3.genblk1[17].state.Q ;
 wire \i_music.i_sample.t3.genblk1[1].state.Q ;
 wire \i_music.i_sample.t3.genblk1[2].state.Q ;
 wire \i_music.i_sample.t3.genblk1[3].state.Q ;
 wire \i_music.i_sample.t3.genblk1[4].state.Q ;
 wire \i_music.i_sample.t3.genblk1[5].state.Q ;
 wire \i_music.i_sample.t3.genblk1[6].state.Q ;
 wire \i_music.i_sample.t3.genblk1[7].state.Q ;
 wire \i_music.i_sample.t3.genblk1[8].state.Q ;
 wire \i_music.i_sample.t3.genblk1[9].state.Q ;
 wire \i_music.i_sample.t4.CG.GCLK ;
 wire \i_music.i_sample.t4.genblk1[0].state.Q ;
 wire \i_music.i_sample.t4.genblk1[10].state.Q ;
 wire \i_music.i_sample.t4.genblk1[11].state.Q ;
 wire \i_music.i_sample.t4.genblk1[12].state.Q ;
 wire \i_music.i_sample.t4.genblk1[13].state.Q ;
 wire \i_music.i_sample.t4.genblk1[14].state.Q ;
 wire \i_music.i_sample.t4.genblk1[15].state.Q ;
 wire \i_music.i_sample.t4.genblk1[16].state.Q ;
 wire \i_music.i_sample.t4.genblk1[17].state.Q ;
 wire \i_music.i_sample.t4.genblk1[1].state.Q ;
 wire \i_music.i_sample.t4.genblk1[2].state.Q ;
 wire \i_music.i_sample.t4.genblk1[3].state.Q ;
 wire \i_music.i_sample.t4.genblk1[4].state.Q ;
 wire \i_music.i_sample.t4.genblk1[5].state.Q ;
 wire \i_music.i_sample.t4.genblk1[6].state.Q ;
 wire \i_music.i_sample.t4.genblk1[7].state.Q ;
 wire \i_music.i_sample.t4.genblk1[8].state.Q ;
 wire \i_music.i_sample.t4.genblk1[9].state.Q ;
 wire \i_music.i_sample.thresh[0] ;
 wire \i_music.i_sample.thresh[10] ;
 wire \i_music.i_sample.thresh[1] ;
 wire \i_music.i_sample.thresh[2] ;
 wire \i_music.i_sample.thresh[3] ;
 wire \i_music.i_sample.thresh[4] ;
 wire \i_music.i_sample.thresh[5] ;
 wire \i_music.i_sample.thresh[6] ;
 wire \i_music.i_sample.thresh[7] ;
 wire \i_music.i_sample.thresh[8] ;
 wire \i_music.i_sample.thresh[9] ;
 wire \i_music.violin_note_idx[1][0] ;
 wire \i_music.violin_note_idx[1][1] ;
 wire \i_music.violin_note_idx[1][2] ;
 wire \i_music.violin_note_idx[1][3] ;
 wire \i_music.violin_note_idx[1][4] ;
 wire \i_music.violin_note_idx[1][5] ;
 wire \i_music.violin_note_idx[1][6] ;
 wire \i_music.violin_note_idx[1][7] ;
 wire \i_music.violin_note_idx[1][8] ;
 wire \i_music.violin_note_idx[2][0] ;
 wire \i_music.violin_note_idx[2][1] ;
 wire \i_music.violin_note_idx[2][2] ;
 wire \i_music.violin_note_idx[2][3] ;
 wire \i_music.violin_note_idx[2][4] ;
 wire \i_music.violin_note_idx[2][5] ;
 wire \i_music.violin_note_idx[2][6] ;
 wire \i_music.violin_note_idx[2][7] ;
 wire \i_music.violin_note_idx[2][8] ;
 wire \i_music.violin_note_idx[3][0] ;
 wire \i_music.violin_note_idx[3][1] ;
 wire \i_music.violin_note_idx[3][2] ;
 wire \i_music.violin_note_idx[3][3] ;
 wire \i_music.violin_note_idx[3][4] ;
 wire \i_music.violin_note_idx[3][5] ;
 wire \i_music.violin_note_idx[3][6] ;
 wire \i_music.violin_note_idx[3][7] ;
 wire \i_music.violin_note_idx[3][8] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire clknet_level_0_1_10_clk;
 wire clknet_level_1_1_11_clk;
 wire clknet_level_2_1_12_clk;
 wire clknet_level_0_1_23_clk;
 wire clknet_level_1_1_24_clk;
 wire clknet_level_2_1_25_clk;
 wire clknet_level_0_1_36_clk;
 wire clknet_level_1_1_37_clk;
 wire clknet_level_2_1_38_clk;
 wire clknet_level_0_1_49_clk;
 wire clknet_level_1_1_410_clk;
 wire clknet_level_2_1_411_clk;
 wire clknet_level_0_1_512_clk;
 wire clknet_level_1_1_513_clk;
 wire clknet_level_2_1_514_clk;
 wire clknet_level_0_1_615_clk;
 wire clknet_level_1_1_616_clk;
 wire clknet_level_2_1_617_clk;
 wire clknet_level_0_1_718_clk;
 wire clknet_level_1_1_719_clk;
 wire clknet_level_2_1_720_clk;
 wire clknet_level_0_1_821_clk;
 wire clknet_level_1_1_822_clk;
 wire clknet_level_2_1_823_clk;
 wire clknet_level_0_1_924_clk;
 wire clknet_level_1_1_925_clk;
 wire clknet_level_2_1_926_clk;
 wire clknet_level_0_1_1027_clk;
 wire clknet_level_1_1_1028_clk;
 wire clknet_level_2_1_1029_clk;
 wire clknet_level_0_1_1130_clk;
 wire clknet_level_1_1_1131_clk;
 wire clknet_level_2_1_1132_clk;
 wire clknet_level_0_1_1233_clk;
 wire clknet_level_1_1_1234_clk;
 wire clknet_level_2_1_1235_clk;
 wire clknet_level_0_1_1336_clk;
 wire clknet_level_1_1_1337_clk;
 wire clknet_level_2_1_1338_clk;
 wire clknet_level_0_1_1439_clk;
 wire clknet_level_1_1_1440_clk;
 wire clknet_level_2_1_1441_clk;
 wire clknet_level_0_1_1542_clk;
 wire clknet_level_1_1_1543_clk;
 wire clknet_level_2_1_1544_clk;
 wire clknet_level_0_1_1645_clk;
 wire clknet_level_1_1_1646_clk;
 wire clknet_level_2_1_1647_clk;
 wire clknet_level_0_1_1748_clk;
 wire clknet_level_1_1_1749_clk;
 wire clknet_level_2_1_1750_clk;
 wire clknet_level_0_1_1851_clk;
 wire clknet_level_1_1_1852_clk;
 wire clknet_level_2_1_1853_clk;
 wire clknet_level_0_1_1954_clk;
 wire clknet_level_1_1_1955_clk;
 wire clknet_level_2_1_1956_clk;
 wire clknet_level_0_1_2057_clk;
 wire clknet_level_1_1_2058_clk;
 wire clknet_level_2_1_2059_clk;
 wire clknet_level_0_1_2160_clk;
 wire clknet_level_1_1_2161_clk;
 wire clknet_level_2_1_2162_clk;
 wire clknet_level_0_1_2263_clk;
 wire clknet_level_1_1_2264_clk;
 wire clknet_level_2_1_2265_clk;
 wire clknet_level_0_1_2366_clk;
 wire clknet_level_1_1_2367_clk;
 wire clknet_level_2_1_2368_clk;
 wire clknet_level_0_1_2469_clk;
 wire clknet_level_1_1_2470_clk;
 wire clknet_level_2_1_2471_clk;
 wire clknet_level_0_1_2572_clk;
 wire clknet_level_1_1_2573_clk;
 wire clknet_level_2_1_2574_clk;
 wire clknet_level_0_1_2675_clk;
 wire clknet_level_1_1_2676_clk;
 wire clknet_level_2_1_2677_clk;
 wire clknet_level_0_1_2778_clk;
 wire clknet_level_1_1_2779_clk;
 wire clknet_level_2_1_2780_clk;
 wire clknet_level_0_1_2881_clk;
 wire clknet_level_1_1_2882_clk;
 wire clknet_level_2_1_2883_clk;
 wire clknet_level_0_1_2984_clk;
 wire clknet_level_1_1_2985_clk;
 wire clknet_level_2_1_2986_clk;
 wire clknet_level_0_1_3087_clk;
 wire clknet_level_1_1_3088_clk;
 wire clknet_level_2_1_3089_clk;
 wire clknet_level_0_1_3190_clk;
 wire clknet_level_1_1_3191_clk;
 wire clknet_level_2_1_3192_clk;
 wire clknet_level_0_1_3293_clk;
 wire clknet_level_1_1_3294_clk;
 wire clknet_level_2_1_3295_clk;
 wire \clknet_0_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ;
 wire \clknet_0_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ;
 wire \clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ;

 sg13g2_buf_1 _4706_ (.A(rst_n),
    .X(_4140_));
 sg13g2_inv_1 _4707_ (.Y(_4141_),
    .A(net165));
 sg13g2_buf_8 _4708_ (.A(\i_display.x_idx[1] ),
    .X(_4142_));
 sg13g2_buf_8 _4709_ (.A(\i_display.x_idx[3] ),
    .X(_4143_));
 sg13g2_buf_8 _4710_ (.A(_4143_),
    .X(_4144_));
 sg13g2_inv_8 _4711_ (.Y(_4145_),
    .A(net155));
 sg13g2_buf_8 _4712_ (.A(\i_display.x_idx[2] ),
    .X(_4146_));
 sg13g2_nand2_1 _4713_ (.Y(_4147_),
    .A(_4145_),
    .B(net163));
 sg13g2_buf_8 _4714_ (.A(_4147_),
    .X(_4148_));
 sg13g2_nor2_1 _4715_ (.A(net164),
    .B(_4148_),
    .Y(_4149_));
 sg13g2_buf_2 _4716_ (.A(_0089_),
    .X(_4150_));
 sg13g2_inv_2 _4717_ (.Y(_4151_),
    .A(_4150_));
 sg13g2_buf_16 _4718_ (.X(_4152_),
    .A(\i_display.x_idx[4] ));
 sg13g2_inv_16 _4719_ (.A(_4152_),
    .Y(_4153_));
 sg13g2_buf_8 _4720_ (.A(\i_display.x_idx[5] ),
    .X(_4154_));
 sg13g2_nand2_1 _4721_ (.Y(_4155_),
    .A(_4153_),
    .B(_4154_));
 sg13g2_nor2_1 _4722_ (.A(_4151_),
    .B(_4155_),
    .Y(_4156_));
 sg13g2_buf_8 _4723_ (.A(\i_display.x_idx[7] ),
    .X(_4157_));
 sg13g2_buf_1 _4724_ (.A(\i_display.x_idx[6] ),
    .X(_4158_));
 sg13g2_nand2_1 _4725_ (.Y(_4159_),
    .A(_4157_),
    .B(net162));
 sg13g2_buf_2 _4726_ (.A(_4159_),
    .X(_4160_));
 sg13g2_inv_2 _4727_ (.Y(_4161_),
    .A(_4160_));
 sg13g2_nand3_1 _4728_ (.B(_4156_),
    .C(_4161_),
    .A(_4149_),
    .Y(_4162_));
 sg13g2_buf_8 _4729_ (.A(_4152_),
    .X(_4163_));
 sg13g2_nor2_1 _4730_ (.A(net154),
    .B(_4154_),
    .Y(_4164_));
 sg13g2_nand2_1 _4731_ (.Y(_4165_),
    .A(_4164_),
    .B(_4150_));
 sg13g2_nor2_1 _4732_ (.A(_4160_),
    .B(_4165_),
    .Y(_4166_));
 sg13g2_buf_8 _4733_ (.A(\i_display.x_idx[0] ),
    .X(_4167_));
 sg13g2_inv_4 _4734_ (.A(net163),
    .Y(_4168_));
 sg13g2_nor2_1 _4735_ (.A(_4167_),
    .B(_4168_),
    .Y(_4169_));
 sg13g2_inv_1 _4736_ (.Y(_4170_),
    .A(_4169_));
 sg13g2_nor2b_1 _4737_ (.A(_4170_),
    .B_N(net164),
    .Y(_4171_));
 sg13g2_nand2_1 _4738_ (.Y(_4172_),
    .A(_4166_),
    .B(_4171_));
 sg13g2_nand3_1 _4739_ (.B(_4144_),
    .C(_4150_),
    .A(_4168_),
    .Y(_4173_));
 sg13g2_inv_4 _4740_ (.A(_4167_),
    .Y(_4174_));
 sg13g2_nor2_2 _4741_ (.A(_4142_),
    .B(_4174_),
    .Y(_4175_));
 sg13g2_nor2b_1 _4742_ (.A(_4173_),
    .B_N(_4175_),
    .Y(_4176_));
 sg13g2_nand2_2 _4743_ (.Y(_4177_),
    .A(net154),
    .B(_4154_));
 sg13g2_nor2_1 _4744_ (.A(_4160_),
    .B(_4177_),
    .Y(_4178_));
 sg13g2_nand2_1 _4745_ (.Y(_4179_),
    .A(_4176_),
    .B(_4178_));
 sg13g2_nand3_1 _4746_ (.B(_4172_),
    .C(_4179_),
    .A(_4162_),
    .Y(_4180_));
 sg13g2_nor2_2 _4747_ (.A(net163),
    .B(_4143_),
    .Y(_4181_));
 sg13g2_nor2_1 _4748_ (.A(net164),
    .B(_4181_),
    .Y(_4182_));
 sg13g2_nand2_1 _4749_ (.Y(_4183_),
    .A(_4156_),
    .B(_4182_));
 sg13g2_a21oi_1 _4750_ (.A1(net164),
    .A2(net163),
    .Y(_4184_),
    .B1(net155));
 sg13g2_nor2_1 _4751_ (.A(_4151_),
    .B(_4177_),
    .Y(_4185_));
 sg13g2_nand2_1 _4752_ (.Y(_4186_),
    .A(_4184_),
    .B(_4185_));
 sg13g2_nand2_1 _4753_ (.Y(_4187_),
    .A(_4183_),
    .B(_4186_));
 sg13g2_inv_8 _4754_ (.Y(_4188_),
    .A(_4157_));
 sg13g2_nor2_2 _4755_ (.A(net162),
    .B(_4188_),
    .Y(_4189_));
 sg13g2_nand2_1 _4756_ (.Y(_4190_),
    .A(_4187_),
    .B(_4189_));
 sg13g2_inv_4 _4757_ (.A(_4175_),
    .Y(_4191_));
 sg13g2_nor2_1 _4758_ (.A(_4168_),
    .B(_4191_),
    .Y(_4192_));
 sg13g2_nand2_1 _4759_ (.Y(_4193_),
    .A(_4166_),
    .B(_4192_));
 sg13g2_nand2_1 _4760_ (.Y(_4194_),
    .A(_4190_),
    .B(_4193_));
 sg13g2_nor2_1 _4761_ (.A(_4180_),
    .B(_4194_),
    .Y(_4195_));
 sg13g2_nand2_1 _4762_ (.Y(_4196_),
    .A(net164),
    .B(_4167_));
 sg13g2_nand2b_1 _4763_ (.Y(_4197_),
    .B(_4181_),
    .A_N(_4196_));
 sg13g2_inv_1 _4764_ (.Y(_4198_),
    .A(_4148_));
 sg13g2_nand2_1 _4765_ (.Y(_4199_),
    .A(_4198_),
    .B(_4175_));
 sg13g2_nand2_1 _4766_ (.Y(_4200_),
    .A(_4197_),
    .B(_4199_));
 sg13g2_nor2_2 _4767_ (.A(_4154_),
    .B(_4153_),
    .Y(_4201_));
 sg13g2_inv_2 _4768_ (.Y(_4202_),
    .A(_4201_));
 sg13g2_nor2_1 _4769_ (.A(_4157_),
    .B(net162),
    .Y(_4203_));
 sg13g2_buf_8 _4770_ (.A(_4203_),
    .X(_4204_));
 sg13g2_nand2_1 _4771_ (.Y(_4205_),
    .A(_4204_),
    .B(_4150_));
 sg13g2_nor2_2 _4772_ (.A(_4202_),
    .B(_4205_),
    .Y(_4206_));
 sg13g2_nand2_1 _4773_ (.Y(_4207_),
    .A(_4200_),
    .B(_4206_));
 sg13g2_inv_1 _4774_ (.Y(_4208_),
    .A(_4204_));
 sg13g2_nor2_2 _4775_ (.A(_4208_),
    .B(_4165_),
    .Y(_4209_));
 sg13g2_nand2_2 _4776_ (.Y(_4210_),
    .A(\i_display.x_idx[2] ),
    .B(_4143_));
 sg13g2_nor2_1 _4777_ (.A(_4210_),
    .B(_4191_),
    .Y(_4211_));
 sg13g2_nand2_1 _4778_ (.Y(_4212_),
    .A(_4209_),
    .B(_4211_));
 sg13g2_nand2_1 _4779_ (.Y(_4213_),
    .A(_4207_),
    .B(_4212_));
 sg13g2_nor3_1 _4780_ (.A(net164),
    .B(_4154_),
    .C(_4148_),
    .Y(_4214_));
 sg13g2_nand2_1 _4781_ (.Y(_4215_),
    .A(_4167_),
    .B(_4163_));
 sg13g2_inv_1 _4782_ (.Y(_4216_),
    .A(_4215_));
 sg13g2_inv_4 _4783_ (.A(_4189_),
    .Y(_4217_));
 sg13g2_nor2_1 _4784_ (.A(_4151_),
    .B(_4217_),
    .Y(_4218_));
 sg13g2_nand3_1 _4785_ (.B(_4216_),
    .C(_4218_),
    .A(_4214_),
    .Y(_4219_));
 sg13g2_nand3_1 _4786_ (.B(_4142_),
    .C(net163),
    .A(_4145_),
    .Y(_4220_));
 sg13g2_nor2b_1 _4787_ (.A(_4220_),
    .B_N(_4201_),
    .Y(_4221_));
 sg13g2_nand3_1 _4788_ (.B(_4174_),
    .C(_4218_),
    .A(_4221_),
    .Y(_4222_));
 sg13g2_nand2_1 _4789_ (.Y(_4223_),
    .A(_4219_),
    .B(_4222_));
 sg13g2_nor2_1 _4790_ (.A(_4213_),
    .B(_4223_),
    .Y(_4224_));
 sg13g2_buf_1 _4791_ (.A(\i_display.i_vga.low_count[6] ),
    .X(_4225_));
 sg13g2_nor2_1 _4792_ (.A(\i_display.i_vga.low_count[7] ),
    .B(_4225_),
    .Y(_4226_));
 sg13g2_inv_1 _4793_ (.Y(_4227_),
    .A(_4226_));
 sg13g2_nor2_1 _4794_ (.A(\i_display.i_vga.low_count[5] ),
    .B(_4227_),
    .Y(_4228_));
 sg13g2_inv_2 _4795_ (.Y(_4229_),
    .A(_4228_));
 sg13g2_buf_1 _4796_ (.A(\i_display.i_vga.low_count[2] ),
    .X(_4230_));
 sg13g2_inv_1 _4797_ (.Y(_4231_),
    .A(_4230_));
 sg13g2_buf_1 _4798_ (.A(\i_display.i_vga.low_count[0] ),
    .X(_4232_));
 sg13g2_buf_8 _4799_ (.A(\i_display.i_vga.low_count[1] ),
    .X(_4233_));
 sg13g2_nand2_1 _4800_ (.Y(_4234_),
    .A(_4232_),
    .B(_4233_));
 sg13g2_nor2_1 _4801_ (.A(_4231_),
    .B(_4234_),
    .Y(_4235_));
 sg13g2_buf_1 _4802_ (.A(\i_display.i_vga.low_count[8] ),
    .X(_4236_));
 sg13g2_buf_1 _4803_ (.A(\i_display.i_vga.low_count[9] ),
    .X(_4237_));
 sg13g2_buf_2 _4804_ (.A(\i_display.i_vga.low_count[4] ),
    .X(_4238_));
 sg13g2_buf_2 _4805_ (.A(\i_display.i_vga.low_count[3] ),
    .X(_4239_));
 sg13g2_nand2_1 _4806_ (.Y(_4240_),
    .A(_4238_),
    .B(_4239_));
 sg13g2_inv_1 _4807_ (.Y(_4241_),
    .A(_4240_));
 sg13g2_nand4_1 _4808_ (.B(_4236_),
    .C(_4237_),
    .A(_4235_),
    .Y(_4242_),
    .D(_4241_));
 sg13g2_nor2_1 _4809_ (.A(_4229_),
    .B(_4242_),
    .Y(_4243_));
 sg13g2_nor2_1 _4810_ (.A(\i_display.hsync ),
    .B(_4243_),
    .Y(_4244_));
 sg13g2_buf_8 _4811_ (.A(_4244_),
    .X(_4245_));
 sg13g2_nand2_1 _4812_ (.Y(_4246_),
    .A(_4175_),
    .B(_4181_));
 sg13g2_nand2b_1 _4813_ (.Y(_4247_),
    .B(_4206_),
    .A_N(_4246_));
 sg13g2_nand2_1 _4814_ (.Y(_4248_),
    .A(_4204_),
    .B(_4164_));
 sg13g2_nand2b_1 _4815_ (.Y(_4249_),
    .B(_4176_),
    .A_N(_4248_));
 sg13g2_nand2_1 _4816_ (.Y(_4250_),
    .A(_4247_),
    .B(_4249_));
 sg13g2_nor2_1 _4817_ (.A(_4208_),
    .B(_4202_),
    .Y(_4251_));
 sg13g2_nand3_1 _4818_ (.B(_4211_),
    .C(_4150_),
    .A(_4251_),
    .Y(_4252_));
 sg13g2_inv_1 _4819_ (.Y(_4253_),
    .A(_4210_));
 sg13g2_nor2_1 _4820_ (.A(net164),
    .B(_4167_),
    .Y(_4254_));
 sg13g2_buf_2 _4821_ (.A(_4254_),
    .X(_4255_));
 sg13g2_nand2_1 _4822_ (.Y(_4256_),
    .A(_4253_),
    .B(_4255_));
 sg13g2_inv_1 _4823_ (.Y(_4257_),
    .A(_4256_));
 sg13g2_nand2_2 _4824_ (.Y(_4258_),
    .A(_4188_),
    .B(net162));
 sg13g2_nor2_1 _4825_ (.A(_4177_),
    .B(_4258_),
    .Y(_4259_));
 sg13g2_nand3_1 _4826_ (.B(_4259_),
    .C(_4150_),
    .A(_4257_),
    .Y(_4260_));
 sg13g2_nand2_1 _4827_ (.Y(_4261_),
    .A(_4252_),
    .B(_4260_));
 sg13g2_nor2_1 _4828_ (.A(_4250_),
    .B(_4261_),
    .Y(_4262_));
 sg13g2_nand4_1 _4829_ (.B(_4224_),
    .C(_4245_),
    .A(_4195_),
    .Y(_4263_),
    .D(_4262_));
 sg13g2_buf_1 _4830_ (.A(_4263_),
    .X(_4264_));
 sg13g2_buf_1 _4831_ (.A(_0092_),
    .X(_4265_));
 sg13g2_inv_1 _4832_ (.Y(_4266_),
    .A(_4265_));
 sg13g2_inv_8 _4833_ (.Y(_4267_),
    .A(_4245_));
 sg13g2_nand2_2 _4834_ (.Y(_4268_),
    .A(_4267_),
    .B(_0093_));
 sg13g2_nand3_1 _4835_ (.B(_4266_),
    .C(_4268_),
    .A(_4264_),
    .Y(_4269_));
 sg13g2_nand2_1 _4836_ (.Y(_4270_),
    .A(_4221_),
    .B(_4218_));
 sg13g2_nor2_1 _4837_ (.A(_4174_),
    .B(_4270_),
    .Y(_4271_));
 sg13g2_nor3_1 _4838_ (.A(_4271_),
    .B(_4250_),
    .C(_4261_),
    .Y(_4272_));
 sg13g2_inv_4 _4839_ (.A(_4255_),
    .Y(_4273_));
 sg13g2_nor2_1 _4840_ (.A(_4145_),
    .B(_4273_),
    .Y(_4274_));
 sg13g2_nand2_1 _4841_ (.Y(_4275_),
    .A(_4209_),
    .B(_4274_));
 sg13g2_inv_1 _4842_ (.Y(_4276_),
    .A(_4181_));
 sg13g2_nor2_1 _4843_ (.A(_4276_),
    .B(_4273_),
    .Y(_4277_));
 sg13g2_nand2_1 _4844_ (.Y(_4278_),
    .A(_4206_),
    .B(_4277_));
 sg13g2_nand3_1 _4845_ (.B(_4275_),
    .C(_4278_),
    .A(_4212_),
    .Y(_4279_));
 sg13g2_nor2_1 _4846_ (.A(_4180_),
    .B(_4279_),
    .Y(_4280_));
 sg13g2_nand3_1 _4847_ (.B(_4280_),
    .C(_4245_),
    .A(_4272_),
    .Y(_4281_));
 sg13g2_buf_8 _4848_ (.A(_4281_),
    .X(_4282_));
 sg13g2_inv_1 _4849_ (.Y(_4283_),
    .A(_0090_));
 sg13g2_nand2_2 _4850_ (.Y(_4284_),
    .A(_4267_),
    .B(_0091_));
 sg13g2_nand3_1 _4851_ (.B(_4283_),
    .C(_4284_),
    .A(_4282_),
    .Y(_4285_));
 sg13g2_buf_2 _4852_ (.A(_4285_),
    .X(_4286_));
 sg13g2_nand2_1 _4853_ (.Y(_4287_),
    .A(_4269_),
    .B(_4286_));
 sg13g2_buf_2 _4854_ (.A(_0094_),
    .X(_4288_));
 sg13g2_buf_8 _4855_ (.A(_4245_),
    .X(_4289_));
 sg13g2_nor2b_1 _4856_ (.A(net102),
    .B_N(_0095_),
    .Y(_4290_));
 sg13g2_nand3_1 _4857_ (.B(_4161_),
    .C(_4185_),
    .A(_4277_),
    .Y(_4291_));
 sg13g2_nand2_1 _4858_ (.Y(_4292_),
    .A(_4291_),
    .B(_4270_));
 sg13g2_nor2_1 _4859_ (.A(_4148_),
    .B(_4273_),
    .Y(_4293_));
 sg13g2_buf_1 _4860_ (.A(net164),
    .X(_4294_));
 sg13g2_nand2_1 _4861_ (.Y(_4295_),
    .A(_4174_),
    .B(_4294_));
 sg13g2_nor2_1 _4862_ (.A(_4295_),
    .B(_4276_),
    .Y(_4296_));
 sg13g2_nor2_1 _4863_ (.A(_4293_),
    .B(_4296_),
    .Y(_4297_));
 sg13g2_inv_1 _4864_ (.Y(_4298_),
    .A(_4211_));
 sg13g2_nand3_1 _4865_ (.B(_4204_),
    .C(_4150_),
    .A(_4201_),
    .Y(_4299_));
 sg13g2_a21oi_1 _4866_ (.A1(_4297_),
    .A2(_4298_),
    .Y(_4300_),
    .B1(_4299_));
 sg13g2_nor2_1 _4867_ (.A(_4292_),
    .B(_4300_),
    .Y(_4301_));
 sg13g2_inv_1 _4868_ (.Y(_4302_),
    .A(_4149_));
 sg13g2_inv_1 _4869_ (.Y(_4303_),
    .A(_4209_));
 sg13g2_nor2_1 _4870_ (.A(_4302_),
    .B(_4303_),
    .Y(_4304_));
 sg13g2_a21oi_1 _4871_ (.A1(_4200_),
    .A2(_4206_),
    .Y(_4305_),
    .B1(_4304_));
 sg13g2_and3_1 _4872_ (.X(_4306_),
    .A(_4301_),
    .B(net102),
    .C(_4305_));
 sg13g2_nor2_2 _4873_ (.A(_4290_),
    .B(_4306_),
    .Y(_4307_));
 sg13g2_inv_4 _4874_ (.A(_4307_),
    .Y(_4308_));
 sg13g2_nor2_1 _4875_ (.A(_4288_),
    .B(_4308_),
    .Y(_4309_));
 sg13g2_nor2_1 _4876_ (.A(_4286_),
    .B(_4269_),
    .Y(_4310_));
 sg13g2_a21oi_1 _4877_ (.A1(_4287_),
    .A2(_4309_),
    .Y(_4311_),
    .B1(_4310_));
 sg13g2_inv_1 _4878_ (.Y(_4312_),
    .A(_4311_));
 sg13g2_buf_1 _4879_ (.A(_0099_),
    .X(_4313_));
 sg13g2_nor2_1 _4880_ (.A(_4246_),
    .B(_4299_),
    .Y(_4314_));
 sg13g2_nor3_1 _4881_ (.A(_4191_),
    .B(_4173_),
    .C(_4248_),
    .Y(_4315_));
 sg13g2_nor2_1 _4882_ (.A(_4314_),
    .B(_4315_),
    .Y(_4316_));
 sg13g2_nor2_1 _4883_ (.A(_4256_),
    .B(_4299_),
    .Y(_4317_));
 sg13g2_inv_1 _4884_ (.Y(_4318_),
    .A(_4317_));
 sg13g2_nand2_1 _4885_ (.Y(_4319_),
    .A(_4316_),
    .B(_4318_));
 sg13g2_nor2b_1 _4886_ (.A(_4319_),
    .B_N(_4207_),
    .Y(_4320_));
 sg13g2_nand2_1 _4887_ (.Y(_4321_),
    .A(_4162_),
    .B(_4179_));
 sg13g2_inv_1 _4888_ (.Y(_4322_),
    .A(_4321_));
 sg13g2_a22oi_1 _4889_ (.Y(_4323_),
    .B1(_4209_),
    .B2(_4192_),
    .A2(_4211_),
    .A1(_4206_));
 sg13g2_nand4_1 _4890_ (.B(net102),
    .C(_4322_),
    .A(_4320_),
    .Y(_4324_),
    .D(_4323_));
 sg13g2_buf_8 _4891_ (.A(_4267_),
    .X(_4325_));
 sg13g2_nand2_1 _4892_ (.Y(_4326_),
    .A(_4325_),
    .B(_0098_));
 sg13g2_nand2_1 _4893_ (.Y(_4327_),
    .A(_4324_),
    .B(_4326_));
 sg13g2_buf_8 _4894_ (.A(_4327_),
    .X(_4328_));
 sg13g2_nor2_1 _4895_ (.A(net161),
    .B(net82),
    .Y(_4329_));
 sg13g2_inv_1 _4896_ (.Y(_4330_),
    .A(_4190_));
 sg13g2_nand2_1 _4897_ (.Y(_4331_),
    .A(_4316_),
    .B(_4179_));
 sg13g2_nor3_1 _4898_ (.A(_4330_),
    .B(_4292_),
    .C(_4331_),
    .Y(_4332_));
 sg13g2_nand2_1 _4899_ (.Y(_4333_),
    .A(_4275_),
    .B(_4278_));
 sg13g2_nor2_1 _4900_ (.A(_4304_),
    .B(_4333_),
    .Y(_4334_));
 sg13g2_nand3_1 _4901_ (.B(net102),
    .C(_4334_),
    .A(_4332_),
    .Y(_4335_));
 sg13g2_buf_1 _4902_ (.A(_4335_),
    .X(_4336_));
 sg13g2_inv_1 _4903_ (.Y(_4337_),
    .A(_0100_));
 sg13g2_nor2_1 _4904_ (.A(_4337_),
    .B(_4289_),
    .Y(_4338_));
 sg13g2_inv_1 _4905_ (.Y(_4339_),
    .A(_4338_));
 sg13g2_nand2_1 _4906_ (.Y(_4340_),
    .A(_4336_),
    .B(_4339_));
 sg13g2_inv_2 _4907_ (.Y(_4341_),
    .A(_4340_));
 sg13g2_buf_2 _4908_ (.A(_0028_),
    .X(_4342_));
 sg13g2_inv_1 _4909_ (.Y(_4343_),
    .A(_4342_));
 sg13g2_nand2_1 _4910_ (.Y(_4344_),
    .A(_4341_),
    .B(_4343_));
 sg13g2_xor2_1 _4911_ (.B(_4344_),
    .A(_4329_),
    .X(_4345_));
 sg13g2_inv_1 _4912_ (.Y(_4346_),
    .A(_4345_));
 sg13g2_nand2_1 _4913_ (.Y(_4347_),
    .A(_4312_),
    .B(_4346_));
 sg13g2_nand2_1 _4914_ (.Y(_4348_),
    .A(_4311_),
    .B(_4345_));
 sg13g2_nand2_1 _4915_ (.Y(_4349_),
    .A(_4347_),
    .B(_4348_));
 sg13g2_buf_2 _4916_ (.A(_0097_),
    .X(_4350_));
 sg13g2_inv_1 _4917_ (.Y(_4351_),
    .A(_4350_));
 sg13g2_nand3_1 _4918_ (.B(_4351_),
    .C(_4339_),
    .A(_4336_),
    .Y(_4352_));
 sg13g2_buf_1 _4919_ (.A(_4352_),
    .X(_4353_));
 sg13g2_inv_1 _4920_ (.Y(_4354_),
    .A(_4329_));
 sg13g2_nor2_1 _4921_ (.A(_4353_),
    .B(_4354_),
    .Y(_4355_));
 sg13g2_inv_1 _4922_ (.Y(_4356_),
    .A(_4355_));
 sg13g2_nand2_1 _4923_ (.Y(_4357_),
    .A(_4349_),
    .B(_4356_));
 sg13g2_nand3_1 _4924_ (.B(_4348_),
    .C(_4355_),
    .A(_4347_),
    .Y(_4358_));
 sg13g2_nand2_1 _4925_ (.Y(_4359_),
    .A(_4357_),
    .B(_4358_));
 sg13g2_nand3_1 _4926_ (.B(_4318_),
    .C(_4260_),
    .A(_4316_),
    .Y(_4360_));
 sg13g2_nand2_1 _4927_ (.Y(_4361_),
    .A(_4209_),
    .B(_4293_));
 sg13g2_nor2b_1 _4928_ (.A(_4333_),
    .B_N(_4361_),
    .Y(_4362_));
 sg13g2_nor2b_1 _4929_ (.A(_4360_),
    .B_N(_4362_),
    .Y(_4363_));
 sg13g2_a22oi_1 _4930_ (.Y(_4364_),
    .B1(_4166_),
    .B2(_4192_),
    .A2(_4178_),
    .A1(_4176_));
 sg13g2_nand3_1 _4931_ (.B(_4289_),
    .C(_4364_),
    .A(_4363_),
    .Y(_4365_));
 sg13g2_nand2_1 _4932_ (.Y(_4366_),
    .A(_4267_),
    .B(_0088_));
 sg13g2_nand2_1 _4933_ (.Y(_4367_),
    .A(_4365_),
    .B(_4366_));
 sg13g2_buf_8 _4934_ (.A(_4367_),
    .X(_4368_));
 sg13g2_nor2_1 _4935_ (.A(_0090_),
    .B(net84),
    .Y(_4369_));
 sg13g2_inv_1 _4936_ (.Y(_4370_),
    .A(_0027_));
 sg13g2_nor2_2 _4937_ (.A(_4370_),
    .B(_4245_),
    .Y(_4371_));
 sg13g2_inv_1 _4938_ (.Y(_4372_),
    .A(_4194_));
 sg13g2_nand2_1 _4939_ (.Y(_4373_),
    .A(_4214_),
    .B(_4218_));
 sg13g2_nand2_1 _4940_ (.Y(_4374_),
    .A(_4373_),
    .B(_4270_));
 sg13g2_nor2_1 _4941_ (.A(_4374_),
    .B(_4321_),
    .Y(_4375_));
 sg13g2_nand2_1 _4942_ (.Y(_4376_),
    .A(_4372_),
    .B(_4375_));
 sg13g2_inv_1 _4943_ (.Y(_4377_),
    .A(_4185_));
 sg13g2_nor3_1 _4944_ (.A(_4258_),
    .B(_4256_),
    .C(_4377_),
    .Y(_4378_));
 sg13g2_nor3_1 _4945_ (.A(_4317_),
    .B(_4378_),
    .C(_4250_),
    .Y(_4379_));
 sg13g2_nand2_1 _4946_ (.Y(_4380_),
    .A(_4379_),
    .B(_4362_));
 sg13g2_nor3_2 _4947_ (.A(_4325_),
    .B(_4376_),
    .C(_4380_),
    .Y(_4381_));
 sg13g2_nor2_1 _4948_ (.A(_4371_),
    .B(_4381_),
    .Y(_4382_));
 sg13g2_inv_1 _4949_ (.Y(_4383_),
    .A(_0096_));
 sg13g2_nand2_1 _4950_ (.Y(_4384_),
    .A(_4382_),
    .B(_4383_));
 sg13g2_xnor2_1 _4951_ (.Y(_4385_),
    .A(_4369_),
    .B(_4384_));
 sg13g2_nand2_1 _4952_ (.Y(_4386_),
    .A(_4264_),
    .B(_4268_));
 sg13g2_buf_2 _4953_ (.A(_4386_),
    .X(_4387_));
 sg13g2_nor2b_1 _4954_ (.A(_4387_),
    .B_N(_4266_),
    .Y(_4388_));
 sg13g2_nand2_1 _4955_ (.Y(_4389_),
    .A(_4282_),
    .B(_4284_));
 sg13g2_buf_8 _4956_ (.A(_4389_),
    .X(_4390_));
 sg13g2_nor2_2 _4957_ (.A(_4288_),
    .B(_4390_),
    .Y(_4391_));
 sg13g2_nand2_1 _4958_ (.Y(_4392_),
    .A(_4388_),
    .B(_4391_));
 sg13g2_inv_1 _4959_ (.Y(_4393_),
    .A(_4288_));
 sg13g2_nand3_1 _4960_ (.B(_4393_),
    .C(_4268_),
    .A(_4264_),
    .Y(_4394_));
 sg13g2_nand3_1 _4961_ (.B(_4266_),
    .C(_4284_),
    .A(_4282_),
    .Y(_4395_));
 sg13g2_nand2_1 _4962_ (.Y(_4396_),
    .A(_4394_),
    .B(_4395_));
 sg13g2_nand2_1 _4963_ (.Y(_4397_),
    .A(_4392_),
    .B(_4396_));
 sg13g2_nor2_1 _4964_ (.A(_4350_),
    .B(_4308_),
    .Y(_4398_));
 sg13g2_inv_1 _4965_ (.Y(_4399_),
    .A(_4398_));
 sg13g2_nand2_1 _4966_ (.Y(_4400_),
    .A(_4397_),
    .B(_4399_));
 sg13g2_nand3_1 _4967_ (.B(_4396_),
    .C(_4398_),
    .A(_4392_),
    .Y(_4401_));
 sg13g2_nand2_1 _4968_ (.Y(_4402_),
    .A(_4400_),
    .B(_4401_));
 sg13g2_nand2b_1 _4969_ (.Y(_4403_),
    .B(_4402_),
    .A_N(_4385_));
 sg13g2_nand3_1 _4970_ (.B(_4401_),
    .C(_4385_),
    .A(_4400_),
    .Y(_4404_));
 sg13g2_buf_1 _4971_ (.A(_4404_),
    .X(_4405_));
 sg13g2_nand2_1 _4972_ (.Y(_4406_),
    .A(_4403_),
    .B(_4405_));
 sg13g2_inv_1 _4973_ (.Y(_4407_),
    .A(_4286_));
 sg13g2_nand2_1 _4974_ (.Y(_4408_),
    .A(_4388_),
    .B(_4407_));
 sg13g2_nand2_1 _4975_ (.Y(_4409_),
    .A(_4408_),
    .B(_4287_));
 sg13g2_inv_1 _4976_ (.Y(_4410_),
    .A(_4309_));
 sg13g2_nand2_1 _4977_ (.Y(_4411_),
    .A(_4409_),
    .B(_4410_));
 sg13g2_nand3_1 _4978_ (.B(_4287_),
    .C(_4309_),
    .A(_4408_),
    .Y(_4412_));
 sg13g2_buf_2 _4979_ (.A(\i_display.frame[0] ),
    .X(_4413_));
 sg13g2_inv_1 _4980_ (.Y(_4414_),
    .A(_4413_));
 sg13g2_nor2_1 _4981_ (.A(_4414_),
    .B(net84),
    .Y(_4415_));
 sg13g2_nand3_1 _4982_ (.B(_4412_),
    .C(_4415_),
    .A(_4411_),
    .Y(_4416_));
 sg13g2_inv_1 _4983_ (.Y(_4417_),
    .A(_4416_));
 sg13g2_nand2_1 _4984_ (.Y(_4418_),
    .A(_4406_),
    .B(_4417_));
 sg13g2_nand3_1 _4985_ (.B(_4405_),
    .C(_4416_),
    .A(_4403_),
    .Y(_4419_));
 sg13g2_nand2_1 _4986_ (.Y(_4420_),
    .A(_4418_),
    .B(_4419_));
 sg13g2_nand2b_1 _4987_ (.Y(_4421_),
    .B(_4420_),
    .A_N(_4359_));
 sg13g2_nand3_1 _4988_ (.B(_4418_),
    .C(_4419_),
    .A(_4359_),
    .Y(_4422_));
 sg13g2_nand2_1 _4989_ (.Y(_4423_),
    .A(_4421_),
    .B(_4422_));
 sg13g2_nor3_1 _4990_ (.A(_4288_),
    .B(net82),
    .C(_4353_),
    .Y(_4424_));
 sg13g2_nor2_1 _4991_ (.A(_4350_),
    .B(_4327_),
    .Y(_4425_));
 sg13g2_nor2_1 _4992_ (.A(net161),
    .B(_4340_),
    .Y(_4426_));
 sg13g2_xor2_1 _4993_ (.B(_4426_),
    .A(_4425_),
    .X(_4427_));
 sg13g2_nand3_1 _4994_ (.B(_4283_),
    .C(_4268_),
    .A(_4264_),
    .Y(_4428_));
 sg13g2_nand3_1 _4995_ (.B(_4383_),
    .C(_4284_),
    .A(_4282_),
    .Y(_4429_));
 sg13g2_nand2_1 _4996_ (.Y(_4430_),
    .A(_4428_),
    .B(_4429_));
 sg13g2_buf_2 _4997_ (.A(\i_display.frame[2] ),
    .X(_4431_));
 sg13g2_inv_2 _4998_ (.Y(_4432_),
    .A(_4431_));
 sg13g2_nor2_1 _4999_ (.A(_4432_),
    .B(_4308_),
    .Y(_4433_));
 sg13g2_nand3_1 _5000_ (.B(_4383_),
    .C(_4268_),
    .A(_4264_),
    .Y(_4434_));
 sg13g2_buf_1 _5001_ (.A(_4434_),
    .X(_4435_));
 sg13g2_nor2_1 _5002_ (.A(_4286_),
    .B(_4435_),
    .Y(_4436_));
 sg13g2_a21oi_2 _5003_ (.B1(_4436_),
    .Y(_4437_),
    .A2(_4433_),
    .A1(_4430_));
 sg13g2_xor2_1 _5004_ (.B(_4437_),
    .A(_4427_),
    .X(_4438_));
 sg13g2_nand2b_1 _5005_ (.Y(_4439_),
    .B(_4438_),
    .A_N(_4424_));
 sg13g2_xnor2_1 _5006_ (.Y(_4440_),
    .A(_4427_),
    .B(_4437_));
 sg13g2_nand2_1 _5007_ (.Y(_4441_),
    .A(_4440_),
    .B(_4424_));
 sg13g2_nand2_1 _5008_ (.Y(_4442_),
    .A(_4411_),
    .B(_4412_));
 sg13g2_nand2_1 _5009_ (.Y(_4443_),
    .A(_4442_),
    .B(_4415_));
 sg13g2_inv_1 _5010_ (.Y(_4444_),
    .A(_4415_));
 sg13g2_nand3_1 _5011_ (.B(_4412_),
    .C(_4444_),
    .A(_4411_),
    .Y(_4445_));
 sg13g2_nand2_1 _5012_ (.Y(_4446_),
    .A(_4443_),
    .B(_4445_));
 sg13g2_nand3_1 _5013_ (.B(_4441_),
    .C(_4446_),
    .A(_4439_),
    .Y(_4447_));
 sg13g2_buf_2 _5014_ (.A(_4447_),
    .X(_4448_));
 sg13g2_nand2_1 _5015_ (.Y(_4449_),
    .A(_4423_),
    .B(_4448_));
 sg13g2_inv_1 _5016_ (.Y(_4450_),
    .A(_4448_));
 sg13g2_nand3_1 _5017_ (.B(_4422_),
    .C(_4450_),
    .A(_4421_),
    .Y(_4451_));
 sg13g2_nor2b_1 _5018_ (.A(_4437_),
    .B_N(_4427_),
    .Y(_4452_));
 sg13g2_a21oi_1 _5019_ (.A1(_4440_),
    .A2(_4424_),
    .Y(_4453_),
    .B1(_4452_));
 sg13g2_inv_1 _5020_ (.Y(_4454_),
    .A(_4453_));
 sg13g2_nand3_1 _5021_ (.B(_4451_),
    .C(_4454_),
    .A(_4449_),
    .Y(_4455_));
 sg13g2_nand2_1 _5022_ (.Y(_4456_),
    .A(_4423_),
    .B(_4450_));
 sg13g2_nand3_1 _5023_ (.B(_4422_),
    .C(_4448_),
    .A(_4421_),
    .Y(_4457_));
 sg13g2_nand3_1 _5024_ (.B(_4457_),
    .C(_4453_),
    .A(_4456_),
    .Y(_4458_));
 sg13g2_nand2_1 _5025_ (.Y(_4459_),
    .A(_4439_),
    .B(_4441_));
 sg13g2_nand2b_1 _5026_ (.Y(_4460_),
    .B(_4459_),
    .A_N(_4446_));
 sg13g2_nand2_1 _5027_ (.Y(_4461_),
    .A(_4460_),
    .B(_4448_));
 sg13g2_buf_1 _5028_ (.A(\i_display.frame[3] ),
    .X(_4462_));
 sg13g2_buf_1 _5029_ (.A(_4462_),
    .X(_4463_));
 sg13g2_nand2_1 _5030_ (.Y(_4464_),
    .A(_4341_),
    .B(net152));
 sg13g2_nor2_1 _5031_ (.A(_4432_),
    .B(net82),
    .Y(_4465_));
 sg13g2_nor2b_2 _5032_ (.A(_4464_),
    .B_N(_4465_),
    .Y(_4466_));
 sg13g2_nand2_1 _5033_ (.Y(_4467_),
    .A(_4307_),
    .B(_4283_));
 sg13g2_or2_1 _5034_ (.X(_4468_),
    .B(_4435_),
    .A(_4467_));
 sg13g2_nor2_1 _5035_ (.A(_4288_),
    .B(net82),
    .Y(_4469_));
 sg13g2_xor2_1 _5036_ (.B(_4469_),
    .A(_4353_),
    .X(_4470_));
 sg13g2_xnor2_1 _5037_ (.Y(_4471_),
    .A(_4468_),
    .B(_4470_));
 sg13g2_xnor2_1 _5038_ (.Y(_4472_),
    .A(_4466_),
    .B(_4471_));
 sg13g2_o21ai_1 _5039_ (.B1(_4430_),
    .Y(_4473_),
    .A1(_4286_),
    .A2(_4435_));
 sg13g2_xnor2_1 _5040_ (.Y(_4474_),
    .A(_4433_),
    .B(_4473_));
 sg13g2_nand2_1 _5041_ (.Y(_4475_),
    .A(_4472_),
    .B(_4474_));
 sg13g2_nand2_1 _5042_ (.Y(_4476_),
    .A(_4461_),
    .B(_4475_));
 sg13g2_nor2_1 _5043_ (.A(_4468_),
    .B(_4470_),
    .Y(_4477_));
 sg13g2_nand2b_1 _5044_ (.Y(_4478_),
    .B(_4466_),
    .A_N(_4471_));
 sg13g2_nor2b_1 _5045_ (.A(_4477_),
    .B_N(_4478_),
    .Y(_4479_));
 sg13g2_inv_1 _5046_ (.Y(_4480_),
    .A(_4479_));
 sg13g2_xor2_1 _5047_ (.B(_4471_),
    .A(_4466_),
    .X(_4481_));
 sg13g2_nor2b_1 _5048_ (.A(_4481_),
    .B_N(_4474_),
    .Y(_4482_));
 sg13g2_nand3_1 _5049_ (.B(_4448_),
    .C(_4482_),
    .A(_4460_),
    .Y(_4483_));
 sg13g2_inv_1 _5050_ (.Y(_4484_),
    .A(_4483_));
 sg13g2_a21oi_1 _5051_ (.A1(_4476_),
    .A2(_4480_),
    .Y(_4485_),
    .B1(_4484_));
 sg13g2_inv_1 _5052_ (.Y(_4486_),
    .A(_4485_));
 sg13g2_a21oi_1 _5053_ (.A1(_4455_),
    .A2(_4458_),
    .Y(_4487_),
    .B1(_4486_));
 sg13g2_nand3_1 _5054_ (.B(_4483_),
    .C(_4480_),
    .A(_4476_),
    .Y(_4488_));
 sg13g2_nand2_1 _5055_ (.Y(_4489_),
    .A(_4461_),
    .B(_4482_));
 sg13g2_nand3_1 _5056_ (.B(_4448_),
    .C(_4475_),
    .A(_4460_),
    .Y(_4490_));
 sg13g2_nand3_1 _5057_ (.B(_4490_),
    .C(_4479_),
    .A(_4489_),
    .Y(_4491_));
 sg13g2_nand2_1 _5058_ (.Y(_4492_),
    .A(_4488_),
    .B(_4491_));
 sg13g2_nor2_1 _5059_ (.A(_4265_),
    .B(_4340_),
    .Y(_4493_));
 sg13g2_buf_1 _5060_ (.A(\i_display.frame[1] ),
    .X(_4494_));
 sg13g2_inv_1 _5061_ (.Y(_4495_),
    .A(net160));
 sg13g2_nor2_1 _5062_ (.A(_4495_),
    .B(net82),
    .Y(_4496_));
 sg13g2_nand2_1 _5063_ (.Y(_4497_),
    .A(_4493_),
    .B(_4496_));
 sg13g2_xnor2_1 _5064_ (.Y(_4498_),
    .A(_4465_),
    .B(_4464_));
 sg13g2_nor2b_1 _5065_ (.A(_4497_),
    .B_N(_4498_),
    .Y(_4499_));
 sg13g2_inv_1 _5066_ (.Y(_4500_),
    .A(_4499_));
 sg13g2_xnor2_1 _5067_ (.Y(_4501_),
    .A(_4497_),
    .B(_4498_));
 sg13g2_xor2_1 _5068_ (.B(_4435_),
    .A(_4467_),
    .X(_4502_));
 sg13g2_and2_1 _5069_ (.A(_4501_),
    .B(_4502_),
    .X(_4503_));
 sg13g2_inv_1 _5070_ (.Y(_4504_),
    .A(_4503_));
 sg13g2_xnor2_1 _5071_ (.Y(_4505_),
    .A(_4474_),
    .B(_4472_));
 sg13g2_a21oi_1 _5072_ (.A1(_4500_),
    .A2(_4504_),
    .Y(_4506_),
    .B1(_4505_));
 sg13g2_inv_1 _5073_ (.Y(_4507_),
    .A(_4506_));
 sg13g2_nand2_1 _5074_ (.Y(_4508_),
    .A(_4492_),
    .B(_4507_));
 sg13g2_nor4_1 _5075_ (.A(_4414_),
    .B(_0090_),
    .C(net82),
    .D(_4340_),
    .Y(_4509_));
 sg13g2_nand3_1 _5076_ (.B(_4383_),
    .C(_4307_),
    .A(_4509_),
    .Y(_4510_));
 sg13g2_xnor2_1 _5077_ (.Y(_4511_),
    .A(_4496_),
    .B(_4493_));
 sg13g2_a21oi_1 _5078_ (.A1(_4383_),
    .A2(_4307_),
    .Y(_4512_),
    .B1(_4509_));
 sg13g2_a21oi_1 _5079_ (.A1(_4510_),
    .A2(_4511_),
    .Y(_4513_),
    .B1(_4512_));
 sg13g2_o21ai_1 _5080_ (.B1(_4513_),
    .Y(_4514_),
    .A1(_4502_),
    .A2(_4501_));
 sg13g2_nor2_1 _5081_ (.A(_4500_),
    .B(_4505_),
    .Y(_4515_));
 sg13g2_nor2b_1 _5082_ (.A(_4499_),
    .B_N(_4505_),
    .Y(_4516_));
 sg13g2_nor4_2 _5083_ (.A(_4503_),
    .B(_4514_),
    .C(_4515_),
    .Y(_4517_),
    .D(_4516_));
 sg13g2_nor2_1 _5084_ (.A(_4507_),
    .B(_4492_),
    .Y(_4518_));
 sg13g2_a21oi_2 _5085_ (.B1(_4518_),
    .Y(_4519_),
    .A2(_4517_),
    .A1(_4508_));
 sg13g2_nand3_1 _5086_ (.B(_4458_),
    .C(_4486_),
    .A(_4455_),
    .Y(_4520_));
 sg13g2_o21ai_1 _5087_ (.B1(_4520_),
    .Y(_4521_),
    .A1(_4487_),
    .A2(_4519_));
 sg13g2_buf_1 _5088_ (.A(_4521_),
    .X(_4522_));
 sg13g2_inv_1 _5089_ (.Y(_4523_),
    .A(_4451_));
 sg13g2_a21oi_1 _5090_ (.A1(_4449_),
    .A2(_4454_),
    .Y(_4524_),
    .B1(_4523_));
 sg13g2_inv_1 _5091_ (.Y(_4525_),
    .A(_4524_));
 sg13g2_o21ai_1 _5092_ (.B1(_4421_),
    .Y(_4526_),
    .A1(_4416_),
    .A2(_4406_));
 sg13g2_nor3_1 _5093_ (.A(_4495_),
    .B(_4371_),
    .C(_4381_),
    .Y(_4527_));
 sg13g2_nand3_1 _5094_ (.B(_4275_),
    .C(_4278_),
    .A(_4361_),
    .Y(_4528_));
 sg13g2_nor2_1 _5095_ (.A(_4528_),
    .B(_4319_),
    .Y(_4529_));
 sg13g2_nor2_1 _5096_ (.A(_4292_),
    .B(_4194_),
    .Y(_4530_));
 sg13g2_nand3_1 _5097_ (.B(_4530_),
    .C(_4245_),
    .A(_4529_),
    .Y(_4531_));
 sg13g2_nand2_1 _5098_ (.Y(_4532_),
    .A(_4267_),
    .B(_0035_));
 sg13g2_nand2_1 _5099_ (.Y(_4533_),
    .A(_4531_),
    .B(_4532_));
 sg13g2_buf_8 _5100_ (.A(_4533_),
    .X(_4534_));
 sg13g2_nor2_1 _5101_ (.A(_4413_),
    .B(net83),
    .Y(_4535_));
 sg13g2_inv_1 _5102_ (.Y(_4536_),
    .A(_4535_));
 sg13g2_nand2_1 _5103_ (.Y(_4537_),
    .A(_4527_),
    .B(_4536_));
 sg13g2_inv_1 _5104_ (.Y(_4538_),
    .A(_4375_));
 sg13g2_nor2_1 _5105_ (.A(_4194_),
    .B(_4538_),
    .Y(_4539_));
 sg13g2_nand3_1 _5106_ (.B(_4245_),
    .C(_4539_),
    .A(_4363_),
    .Y(_4540_));
 sg13g2_buf_8 _5107_ (.A(_4540_),
    .X(_4541_));
 sg13g2_inv_4 _5108_ (.A(_4371_),
    .Y(_4542_));
 sg13g2_nand3_1 _5109_ (.B(net160),
    .C(_4542_),
    .A(_4541_),
    .Y(_4543_));
 sg13g2_nand2_1 _5110_ (.Y(_4544_),
    .A(_4543_),
    .B(_4535_));
 sg13g2_nand2_1 _5111_ (.Y(_4545_),
    .A(_4537_),
    .B(_4544_));
 sg13g2_nor2_1 _5112_ (.A(_4432_),
    .B(net84),
    .Y(_4546_));
 sg13g2_nand2_1 _5113_ (.Y(_4547_),
    .A(_4545_),
    .B(_4546_));
 sg13g2_inv_1 _5114_ (.Y(_4548_),
    .A(_4546_));
 sg13g2_nand3_1 _5115_ (.B(_4544_),
    .C(_4548_),
    .A(_4537_),
    .Y(_4549_));
 sg13g2_nand2_1 _5116_ (.Y(_4550_),
    .A(_4547_),
    .B(_4549_));
 sg13g2_nor2b_1 _5117_ (.A(_4384_),
    .B_N(_4369_),
    .Y(_4551_));
 sg13g2_inv_1 _5118_ (.Y(_4552_),
    .A(_4551_));
 sg13g2_nand2_1 _5119_ (.Y(_4553_),
    .A(_4550_),
    .B(_4552_));
 sg13g2_nand3_1 _5120_ (.B(_4549_),
    .C(_4551_),
    .A(_4547_),
    .Y(_4554_));
 sg13g2_nor2_2 _5121_ (.A(net161),
    .B(_4308_),
    .Y(_4555_));
 sg13g2_buf_1 _5122_ (.A(\i_display.frame[4] ),
    .X(_4556_));
 sg13g2_inv_1 _5123_ (.Y(_4557_),
    .A(_4556_));
 sg13g2_nor2_1 _5124_ (.A(_4557_),
    .B(_4387_),
    .Y(_4558_));
 sg13g2_xnor2_1 _5125_ (.Y(_4559_),
    .A(_4391_),
    .B(_4558_));
 sg13g2_xnor2_1 _5126_ (.Y(_4560_),
    .A(_4555_),
    .B(_4559_));
 sg13g2_nand3_1 _5127_ (.B(_4554_),
    .C(_4560_),
    .A(_4553_),
    .Y(_4561_));
 sg13g2_nand2_1 _5128_ (.Y(_4562_),
    .A(_4550_),
    .B(_4551_));
 sg13g2_nand3_1 _5129_ (.B(_4549_),
    .C(_4552_),
    .A(_4547_),
    .Y(_4563_));
 sg13g2_xor2_1 _5130_ (.B(_4559_),
    .A(_4555_),
    .X(_4564_));
 sg13g2_nand3_1 _5131_ (.B(_4563_),
    .C(_4564_),
    .A(_4562_),
    .Y(_4565_));
 sg13g2_nand2_1 _5132_ (.Y(_4566_),
    .A(_4561_),
    .B(_4565_));
 sg13g2_nand2_1 _5133_ (.Y(_4567_),
    .A(_4566_),
    .B(_4405_));
 sg13g2_inv_1 _5134_ (.Y(_4568_),
    .A(_4405_));
 sg13g2_nand3_1 _5135_ (.B(_4565_),
    .C(_4568_),
    .A(_4561_),
    .Y(_4569_));
 sg13g2_nor2_1 _5136_ (.A(_4342_),
    .B(net82),
    .Y(_4570_));
 sg13g2_inv_1 _5137_ (.Y(_4571_),
    .A(_4313_));
 sg13g2_nand3_1 _5138_ (.B(_4571_),
    .C(_4341_),
    .A(_4570_),
    .Y(_4572_));
 sg13g2_inv_1 _5139_ (.Y(_4573_),
    .A(_4572_));
 sg13g2_a22oi_1 _5140_ (.Y(_4574_),
    .B1(_4398_),
    .B2(_4396_),
    .A2(_4388_),
    .A1(_4391_));
 sg13g2_buf_2 _5141_ (.A(_0036_),
    .X(_4575_));
 sg13g2_inv_1 _5142_ (.Y(_4576_),
    .A(_4575_));
 sg13g2_nand3_1 _5143_ (.B(_4576_),
    .C(_4339_),
    .A(_4336_),
    .Y(_4577_));
 sg13g2_buf_1 _5144_ (.A(_4577_),
    .X(_4578_));
 sg13g2_inv_1 _5145_ (.Y(_4579_),
    .A(_4578_));
 sg13g2_nand2_1 _5146_ (.Y(_4580_),
    .A(_4579_),
    .B(_4570_));
 sg13g2_nand3_1 _5147_ (.B(_4343_),
    .C(_4326_),
    .A(_4324_),
    .Y(_4581_));
 sg13g2_nand2_1 _5148_ (.Y(_4582_),
    .A(_4578_),
    .B(_4581_));
 sg13g2_nand2_1 _5149_ (.Y(_4583_),
    .A(_4580_),
    .B(_4582_));
 sg13g2_nand2_1 _5150_ (.Y(_4584_),
    .A(_4583_),
    .B(net83));
 sg13g2_inv_1 _5151_ (.Y(_4585_),
    .A(net83));
 sg13g2_nand3_1 _5152_ (.B(_4582_),
    .C(_4585_),
    .A(_4580_),
    .Y(_4586_));
 sg13g2_nand2_1 _5153_ (.Y(_4587_),
    .A(_4584_),
    .B(_4586_));
 sg13g2_xnor2_1 _5154_ (.Y(_4588_),
    .A(_4574_),
    .B(_4587_));
 sg13g2_xnor2_1 _5155_ (.Y(_4589_),
    .A(_4573_),
    .B(_4588_));
 sg13g2_nand3_1 _5156_ (.B(_4569_),
    .C(_4589_),
    .A(_4567_),
    .Y(_4590_));
 sg13g2_nand2_1 _5157_ (.Y(_4591_),
    .A(_4566_),
    .B(_4568_));
 sg13g2_nand3_1 _5158_ (.B(_4565_),
    .C(_4405_),
    .A(_4561_),
    .Y(_4592_));
 sg13g2_xnor2_1 _5159_ (.Y(_4593_),
    .A(_4572_),
    .B(_4588_));
 sg13g2_nand3_1 _5160_ (.B(_4592_),
    .C(_4593_),
    .A(_4591_),
    .Y(_4594_));
 sg13g2_nand2_1 _5161_ (.Y(_4595_),
    .A(_4590_),
    .B(_4594_));
 sg13g2_nand2b_1 _5162_ (.Y(_4596_),
    .B(_4595_),
    .A_N(_4526_));
 sg13g2_nand3_1 _5163_ (.B(_4526_),
    .C(_4594_),
    .A(_4590_),
    .Y(_4597_));
 sg13g2_nand2_1 _5164_ (.Y(_4598_),
    .A(_4596_),
    .B(_4597_));
 sg13g2_inv_1 _5165_ (.Y(_4599_),
    .A(_4347_));
 sg13g2_inv_1 _5166_ (.Y(_4600_),
    .A(_4358_));
 sg13g2_nor2_1 _5167_ (.A(_4599_),
    .B(_4600_),
    .Y(_4601_));
 sg13g2_nand2_1 _5168_ (.Y(_0260_),
    .A(_4598_),
    .B(_4601_));
 sg13g2_inv_1 _5169_ (.Y(_0261_),
    .A(_4601_));
 sg13g2_nand3_1 _5170_ (.B(_4597_),
    .C(_0261_),
    .A(_4596_),
    .Y(_0262_));
 sg13g2_nand2_1 _5171_ (.Y(_0263_),
    .A(_0260_),
    .B(_0262_));
 sg13g2_xnor2_1 _5172_ (.Y(_0264_),
    .A(_4525_),
    .B(_0263_));
 sg13g2_nand2_1 _5173_ (.Y(_0265_),
    .A(_4522_),
    .B(_0264_));
 sg13g2_nand3_1 _5174_ (.B(_0262_),
    .C(_4525_),
    .A(_0260_),
    .Y(_0266_));
 sg13g2_buf_1 _5175_ (.A(_0266_),
    .X(_0267_));
 sg13g2_nand2_1 _5176_ (.Y(_0268_),
    .A(_0265_),
    .B(_0267_));
 sg13g2_inv_1 _5177_ (.Y(_0269_),
    .A(_4554_));
 sg13g2_a21oi_2 _5178_ (.B1(_0269_),
    .Y(_0270_),
    .A2(_4560_),
    .A1(_4553_));
 sg13g2_nand2_1 _5179_ (.Y(_0271_),
    .A(_4543_),
    .B(_4536_));
 sg13g2_nor2_1 _5180_ (.A(_4536_),
    .B(_4543_),
    .Y(_0272_));
 sg13g2_a21oi_2 _5181_ (.B1(_0272_),
    .Y(_0273_),
    .A2(_4546_),
    .A1(_0271_));
 sg13g2_nor3_1 _5182_ (.A(_4432_),
    .B(_4371_),
    .C(_4381_),
    .Y(_0274_));
 sg13g2_nor2_1 _5183_ (.A(net160),
    .B(net83),
    .Y(_0275_));
 sg13g2_nand2_1 _5184_ (.Y(_0276_),
    .A(_0274_),
    .B(_0275_));
 sg13g2_nand3_1 _5185_ (.B(_4431_),
    .C(_4542_),
    .A(_4541_),
    .Y(_0277_));
 sg13g2_inv_2 _5186_ (.Y(_0278_),
    .A(_0275_));
 sg13g2_nand2_1 _5187_ (.Y(_0279_),
    .A(_0277_),
    .B(_0278_));
 sg13g2_inv_1 _5188_ (.Y(_0280_),
    .A(_4462_));
 sg13g2_nor2_1 _5189_ (.A(_0280_),
    .B(net84),
    .Y(_0281_));
 sg13g2_nand3_1 _5190_ (.B(_0279_),
    .C(_0281_),
    .A(_0276_),
    .Y(_0282_));
 sg13g2_nand2_1 _5191_ (.Y(_0283_),
    .A(_0274_),
    .B(_0278_));
 sg13g2_nand2_1 _5192_ (.Y(_0284_),
    .A(_0277_),
    .B(_0275_));
 sg13g2_inv_1 _5193_ (.Y(_0285_),
    .A(_0281_));
 sg13g2_nand3_1 _5194_ (.B(_0284_),
    .C(_0285_),
    .A(_0283_),
    .Y(_0286_));
 sg13g2_nand2_1 _5195_ (.Y(_0287_),
    .A(_0282_),
    .B(_0286_));
 sg13g2_nand2b_1 _5196_ (.Y(_0288_),
    .B(_0287_),
    .A_N(_0273_));
 sg13g2_nand3_1 _5197_ (.B(_0282_),
    .C(_0286_),
    .A(_0273_),
    .Y(_0289_));
 sg13g2_nand2_1 _5198_ (.Y(_0290_),
    .A(_0288_),
    .B(_0289_));
 sg13g2_nor2_2 _5199_ (.A(_4342_),
    .B(_4308_),
    .Y(_0291_));
 sg13g2_nor2_1 _5200_ (.A(_4350_),
    .B(_4390_),
    .Y(_0292_));
 sg13g2_nor2_1 _5201_ (.A(net161),
    .B(_4387_),
    .Y(_0293_));
 sg13g2_xnor2_1 _5202_ (.Y(_0294_),
    .A(_0292_),
    .B(_0293_));
 sg13g2_xnor2_1 _5203_ (.Y(_0295_),
    .A(_0291_),
    .B(_0294_));
 sg13g2_nand2_1 _5204_ (.Y(_0296_),
    .A(_0290_),
    .B(_0295_));
 sg13g2_xor2_1 _5205_ (.B(_0294_),
    .A(_0291_),
    .X(_0297_));
 sg13g2_nand3_1 _5206_ (.B(_0289_),
    .C(_0297_),
    .A(_0288_),
    .Y(_0298_));
 sg13g2_nand2_1 _5207_ (.Y(_0299_),
    .A(_0296_),
    .B(_0298_));
 sg13g2_nand2b_1 _5208_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_0270_));
 sg13g2_nand3_1 _5209_ (.B(_0270_),
    .C(_0298_),
    .A(_0296_),
    .Y(_0301_));
 sg13g2_nand2_1 _5210_ (.Y(_0302_),
    .A(_0300_),
    .B(_0301_));
 sg13g2_inv_1 _5211_ (.Y(_0303_),
    .A(_4580_));
 sg13g2_inv_1 _5212_ (.Y(_0304_),
    .A(_4586_));
 sg13g2_nor2_1 _5213_ (.A(_0303_),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_buf_1 _5214_ (.A(_0038_),
    .X(_0306_));
 sg13g2_nor2_1 _5215_ (.A(_0306_),
    .B(_4328_),
    .Y(_0307_));
 sg13g2_inv_1 _5216_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_nor2_2 _5217_ (.A(_4578_),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_inv_1 _5218_ (.Y(_0310_),
    .A(_0306_));
 sg13g2_nor2_1 _5219_ (.A(_4575_),
    .B(net82),
    .Y(_0311_));
 sg13g2_a21oi_1 _5220_ (.A1(_4341_),
    .A2(_0310_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_nor2_1 _5221_ (.A(_0309_),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_nor2b_1 _5222_ (.A(_4559_),
    .B_N(_4555_),
    .Y(_0314_));
 sg13g2_nand2_1 _5223_ (.Y(_0315_),
    .A(_4558_),
    .B(_4391_));
 sg13g2_nor2b_1 _5224_ (.A(_0314_),
    .B_N(_0315_),
    .Y(_0316_));
 sg13g2_xnor2_1 _5225_ (.Y(_0317_),
    .A(_0313_),
    .B(_0316_));
 sg13g2_xnor2_1 _5226_ (.Y(_0318_),
    .A(_0305_),
    .B(_0317_));
 sg13g2_nand2_1 _5227_ (.Y(_0319_),
    .A(_0302_),
    .B(_0318_));
 sg13g2_inv_1 _5228_ (.Y(_0320_),
    .A(_0305_));
 sg13g2_xnor2_1 _5229_ (.Y(_0321_),
    .A(_0320_),
    .B(_0317_));
 sg13g2_nand3_1 _5230_ (.B(_0301_),
    .C(_0321_),
    .A(_0300_),
    .Y(_0322_));
 sg13g2_nand2_1 _5231_ (.Y(_0323_),
    .A(_0319_),
    .B(_0322_));
 sg13g2_inv_1 _5232_ (.Y(_0324_),
    .A(_4569_));
 sg13g2_a21oi_2 _5233_ (.B1(_0324_),
    .Y(_0325_),
    .A2(_4589_),
    .A1(_4567_));
 sg13g2_nand2_1 _5234_ (.Y(_0326_),
    .A(_0323_),
    .B(_0325_));
 sg13g2_nor2_1 _5235_ (.A(_4574_),
    .B(_4587_),
    .Y(_0327_));
 sg13g2_nand2b_1 _5236_ (.Y(_0328_),
    .B(_4573_),
    .A_N(_4588_));
 sg13g2_nor2b_1 _5237_ (.A(_0327_),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_inv_1 _5238_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nor2_1 _5239_ (.A(_0325_),
    .B(_0323_),
    .Y(_0331_));
 sg13g2_a21oi_1 _5240_ (.A1(_0326_),
    .A2(_0330_),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_inv_1 _5241_ (.Y(_0333_),
    .A(_0332_));
 sg13g2_nand2_1 _5242_ (.Y(_0334_),
    .A(_0299_),
    .B(_0270_));
 sg13g2_nor2_1 _5243_ (.A(_0270_),
    .B(_0299_),
    .Y(_0335_));
 sg13g2_a21oi_2 _5244_ (.B1(_0335_),
    .Y(_0336_),
    .A2(_0318_),
    .A1(_0334_));
 sg13g2_nand2_1 _5245_ (.Y(_0337_),
    .A(_0287_),
    .B(_0273_));
 sg13g2_nor2_1 _5246_ (.A(_0273_),
    .B(_0287_),
    .Y(_0338_));
 sg13g2_a21oi_2 _5247_ (.B1(_0338_),
    .Y(_0339_),
    .A2(_0295_),
    .A1(_0337_));
 sg13g2_nor2_1 _5248_ (.A(_4575_),
    .B(_4308_),
    .Y(_0340_));
 sg13g2_nor2_1 _5249_ (.A(net161),
    .B(_4390_),
    .Y(_0341_));
 sg13g2_nor2_1 _5250_ (.A(_4342_),
    .B(_4387_),
    .Y(_0342_));
 sg13g2_xnor2_1 _5251_ (.Y(_0343_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_xnor2_1 _5252_ (.Y(_0344_),
    .A(_0340_),
    .B(_0343_));
 sg13g2_nor2_1 _5253_ (.A(_0278_),
    .B(_0277_),
    .Y(_0345_));
 sg13g2_a21oi_2 _5254_ (.B1(_0345_),
    .Y(_0346_),
    .A2(_0281_),
    .A1(_0279_));
 sg13g2_nor2_1 _5255_ (.A(_4431_),
    .B(net83),
    .Y(_0347_));
 sg13g2_nor3_1 _5256_ (.A(_0280_),
    .B(_4371_),
    .C(_4381_),
    .Y(_0348_));
 sg13g2_nand2b_1 _5257_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0347_));
 sg13g2_nand3_1 _5258_ (.B(_4462_),
    .C(_4542_),
    .A(_4541_),
    .Y(_0350_));
 sg13g2_nand2_1 _5259_ (.Y(_0351_),
    .A(_0350_),
    .B(_0347_));
 sg13g2_nand2_1 _5260_ (.Y(_0352_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_nor2_1 _5261_ (.A(_4557_),
    .B(net84),
    .Y(_0353_));
 sg13g2_nand2_1 _5262_ (.Y(_0354_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_inv_1 _5263_ (.Y(_0355_),
    .A(_0353_));
 sg13g2_nand3_1 _5264_ (.B(_0351_),
    .C(_0355_),
    .A(_0349_),
    .Y(_0356_));
 sg13g2_nand2_1 _5265_ (.Y(_0357_),
    .A(_0354_),
    .B(_0356_));
 sg13g2_nand2b_1 _5266_ (.Y(_0358_),
    .B(_0357_),
    .A_N(_0346_));
 sg13g2_nand3_1 _5267_ (.B(_0356_),
    .C(_0346_),
    .A(_0354_),
    .Y(_0359_));
 sg13g2_nand3b_1 _5268_ (.B(_0358_),
    .C(_0359_),
    .Y(_0360_),
    .A_N(_0344_));
 sg13g2_nand2_1 _5269_ (.Y(_0361_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_nand2_1 _5270_ (.Y(_0362_),
    .A(_0361_),
    .B(_0344_));
 sg13g2_nand2_1 _5271_ (.Y(_0363_),
    .A(_0360_),
    .B(_0362_));
 sg13g2_nand2b_1 _5272_ (.Y(_0364_),
    .B(_0363_),
    .A_N(_0339_));
 sg13g2_nand3_1 _5273_ (.B(_0362_),
    .C(_0339_),
    .A(_0360_),
    .Y(_0365_));
 sg13g2_nand2_1 _5274_ (.Y(_0366_),
    .A(_0364_),
    .B(_0365_));
 sg13g2_inv_1 _5275_ (.Y(_0367_),
    .A(_0040_));
 sg13g2_nand2_1 _5276_ (.Y(_0368_),
    .A(_4341_),
    .B(_0367_));
 sg13g2_xnor2_1 _5277_ (.Y(_0369_),
    .A(_0307_),
    .B(_0368_));
 sg13g2_nor2b_1 _5278_ (.A(_0294_),
    .B_N(_0291_),
    .Y(_0370_));
 sg13g2_nand2_1 _5279_ (.Y(_0371_),
    .A(_0293_),
    .B(_0292_));
 sg13g2_nor2b_1 _5280_ (.A(_0370_),
    .B_N(_0371_),
    .Y(_0372_));
 sg13g2_xnor2_1 _5281_ (.Y(_0373_),
    .A(_0369_),
    .B(_0372_));
 sg13g2_xor2_1 _5282_ (.B(_0373_),
    .A(_0309_),
    .X(_0374_));
 sg13g2_nand2_1 _5283_ (.Y(_0375_),
    .A(_0366_),
    .B(_0374_));
 sg13g2_xnor2_1 _5284_ (.Y(_0376_),
    .A(_0309_),
    .B(_0373_));
 sg13g2_nand3_1 _5285_ (.B(_0365_),
    .C(_0376_),
    .A(_0364_),
    .Y(_0377_));
 sg13g2_nand2_1 _5286_ (.Y(_0378_),
    .A(_0375_),
    .B(_0377_));
 sg13g2_nand2b_1 _5287_ (.Y(_0379_),
    .B(_0378_),
    .A_N(_0336_));
 sg13g2_nand3_1 _5288_ (.B(_0377_),
    .C(_0336_),
    .A(_0375_),
    .Y(_0380_));
 sg13g2_nand2_1 _5289_ (.Y(_0381_),
    .A(_0379_),
    .B(_0380_));
 sg13g2_nor2b_1 _5290_ (.A(_0316_),
    .B_N(_0313_),
    .Y(_0382_));
 sg13g2_a21oi_1 _5291_ (.A1(_0317_),
    .A2(_0320_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_inv_1 _5292_ (.Y(_0384_),
    .A(_0383_));
 sg13g2_nand2_1 _5293_ (.Y(_0385_),
    .A(_0381_),
    .B(_0384_));
 sg13g2_nand3_1 _5294_ (.B(_0380_),
    .C(_0383_),
    .A(_0379_),
    .Y(_0386_));
 sg13g2_nand2_1 _5295_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_xnor2_1 _5296_ (.Y(_0388_),
    .A(_0333_),
    .B(_0387_));
 sg13g2_inv_1 _5297_ (.Y(_0389_),
    .A(_4597_));
 sg13g2_a21oi_2 _5298_ (.B1(_0389_),
    .Y(_0390_),
    .A2(_0261_),
    .A1(_4596_));
 sg13g2_nand2b_1 _5299_ (.Y(_0391_),
    .B(_0323_),
    .A_N(_0325_));
 sg13g2_nand3_1 _5300_ (.B(_0322_),
    .C(_0325_),
    .A(_0319_),
    .Y(_0392_));
 sg13g2_nand2_1 _5301_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_nand2_1 _5302_ (.Y(_0394_),
    .A(_0393_),
    .B(_0330_));
 sg13g2_nand3_1 _5303_ (.B(_0392_),
    .C(_0329_),
    .A(_0391_),
    .Y(_0395_));
 sg13g2_nand2_1 _5304_ (.Y(_0396_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_nor2_1 _5305_ (.A(_0390_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_inv_2 _5306_ (.Y(_0398_),
    .A(_0390_));
 sg13g2_a21oi_1 _5307_ (.A1(_0394_),
    .A2(_0395_),
    .Y(_0399_),
    .B1(_0398_));
 sg13g2_nor2_1 _5308_ (.A(_0397_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_nand2_1 _5309_ (.Y(_0401_),
    .A(_0388_),
    .B(_0400_));
 sg13g2_inv_1 _5310_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_nand2_1 _5311_ (.Y(_0403_),
    .A(_0268_),
    .B(_0402_));
 sg13g2_nand2_1 _5312_ (.Y(_0404_),
    .A(_0387_),
    .B(_0332_));
 sg13g2_nand2_1 _5313_ (.Y(_0405_),
    .A(_0404_),
    .B(_0397_));
 sg13g2_nand3_1 _5314_ (.B(_0385_),
    .C(_0386_),
    .A(_0333_),
    .Y(_0406_));
 sg13g2_nand2_1 _5315_ (.Y(_0407_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_inv_1 _5316_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nand2_1 _5317_ (.Y(_0409_),
    .A(_0403_),
    .B(_0408_));
 sg13g2_buf_1 _5318_ (.A(\i_display.frame[6] ),
    .X(_0410_));
 sg13g2_inv_1 _5319_ (.Y(_0411_),
    .A(net159));
 sg13g2_nor2_1 _5320_ (.A(_0411_),
    .B(net84),
    .Y(_0412_));
 sg13g2_buf_1 _5321_ (.A(\i_display.frame[5] ),
    .X(_0413_));
 sg13g2_inv_1 _5322_ (.Y(_0414_),
    .A(net158));
 sg13g2_nand2_1 _5323_ (.Y(_0415_),
    .A(_4541_),
    .B(_4542_));
 sg13g2_nor2_1 _5324_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nor2_1 _5325_ (.A(_4556_),
    .B(net83),
    .Y(_0417_));
 sg13g2_inv_1 _5326_ (.Y(_0418_),
    .A(_0417_));
 sg13g2_nand2_1 _5327_ (.Y(_0419_),
    .A(_0416_),
    .B(_0418_));
 sg13g2_nand3_1 _5328_ (.B(net158),
    .C(_4542_),
    .A(_4541_),
    .Y(_0420_));
 sg13g2_nand2_1 _5329_ (.Y(_0421_),
    .A(_0420_),
    .B(_0417_));
 sg13g2_nand3b_1 _5330_ (.B(_0419_),
    .C(_0421_),
    .Y(_0422_),
    .A_N(_0412_));
 sg13g2_nand2_1 _5331_ (.Y(_0423_),
    .A(_0419_),
    .B(_0421_));
 sg13g2_nand2_1 _5332_ (.Y(_0424_),
    .A(_0423_),
    .B(_0412_));
 sg13g2_nand2_1 _5333_ (.Y(_0425_),
    .A(_0422_),
    .B(_0424_));
 sg13g2_nand3_1 _5334_ (.B(_4556_),
    .C(_4542_),
    .A(_4541_),
    .Y(_0426_));
 sg13g2_nor2_1 _5335_ (.A(net152),
    .B(net83),
    .Y(_0427_));
 sg13g2_inv_2 _5336_ (.Y(_0428_),
    .A(_0427_));
 sg13g2_nand2_1 _5337_ (.Y(_0429_),
    .A(_0426_),
    .B(_0428_));
 sg13g2_nor2_1 _5338_ (.A(_0414_),
    .B(net84),
    .Y(_0430_));
 sg13g2_nor2_1 _5339_ (.A(_0428_),
    .B(_0426_),
    .Y(_0431_));
 sg13g2_a21oi_1 _5340_ (.A1(_0429_),
    .A2(_0430_),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_nand2_1 _5341_ (.Y(_0433_),
    .A(_0425_),
    .B(_0432_));
 sg13g2_inv_1 _5342_ (.Y(_0434_),
    .A(_0432_));
 sg13g2_nand3_1 _5343_ (.B(_0422_),
    .C(_0424_),
    .A(_0434_),
    .Y(_0435_));
 sg13g2_inv_1 _5344_ (.Y(_0436_),
    .A(\i_display.frame[9] ));
 sg13g2_nor2_1 _5345_ (.A(_0436_),
    .B(_4308_),
    .Y(_0437_));
 sg13g2_nand3_1 _5346_ (.B(_4576_),
    .C(_4284_),
    .A(_4282_),
    .Y(_0438_));
 sg13g2_buf_1 _5347_ (.A(_0438_),
    .X(_0439_));
 sg13g2_buf_1 _5348_ (.A(\i_display.frame[8] ),
    .X(_0440_));
 sg13g2_inv_1 _5349_ (.Y(_0441_),
    .A(_0440_));
 sg13g2_nor2_1 _5350_ (.A(_0441_),
    .B(_4387_),
    .Y(_0442_));
 sg13g2_xor2_1 _5351_ (.B(_0442_),
    .A(_0439_),
    .X(_0443_));
 sg13g2_xnor2_1 _5352_ (.Y(_0444_),
    .A(_0437_),
    .B(_0443_));
 sg13g2_nand3_1 _5353_ (.B(_0435_),
    .C(_0444_),
    .A(_0433_),
    .Y(_0445_));
 sg13g2_nand2_1 _5354_ (.Y(_0446_),
    .A(_0425_),
    .B(_0434_));
 sg13g2_nand3_1 _5355_ (.B(_0424_),
    .C(_0432_),
    .A(_0422_),
    .Y(_0447_));
 sg13g2_inv_1 _5356_ (.Y(_0448_),
    .A(_0444_));
 sg13g2_nand3_1 _5357_ (.B(_0447_),
    .C(_0448_),
    .A(_0446_),
    .Y(_0449_));
 sg13g2_nand2_1 _5358_ (.Y(_0450_),
    .A(_0445_),
    .B(_0449_));
 sg13g2_nor2_1 _5359_ (.A(_4557_),
    .B(_0415_),
    .Y(_0451_));
 sg13g2_nand2_1 _5360_ (.Y(_0452_),
    .A(_0451_),
    .B(_0427_));
 sg13g2_nand2_1 _5361_ (.Y(_0453_),
    .A(_0452_),
    .B(_0429_));
 sg13g2_inv_1 _5362_ (.Y(_0454_),
    .A(_0430_));
 sg13g2_nand2_1 _5363_ (.Y(_0455_),
    .A(_0453_),
    .B(_0454_));
 sg13g2_nand3_1 _5364_ (.B(_0429_),
    .C(_0430_),
    .A(_0452_),
    .Y(_0456_));
 sg13g2_nand2_1 _5365_ (.Y(_0457_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_nand2b_1 _5366_ (.Y(_0458_),
    .B(_0350_),
    .A_N(_0347_));
 sg13g2_nor2b_1 _5367_ (.A(_0350_),
    .B_N(_0347_),
    .Y(_0459_));
 sg13g2_a21oi_2 _5368_ (.B1(_0459_),
    .Y(_0460_),
    .A2(_0353_),
    .A1(_0458_));
 sg13g2_nand2_1 _5369_ (.Y(_0461_),
    .A(_0457_),
    .B(_0460_));
 sg13g2_nor2_1 _5370_ (.A(_0441_),
    .B(_4308_),
    .Y(_0462_));
 sg13g2_nor2_1 _5371_ (.A(_4342_),
    .B(_4390_),
    .Y(_0463_));
 sg13g2_buf_2 _5372_ (.A(\i_display.frame[7] ),
    .X(_0464_));
 sg13g2_inv_1 _5373_ (.Y(_0465_),
    .A(_0464_));
 sg13g2_nor2_1 _5374_ (.A(_0465_),
    .B(_4387_),
    .Y(_0466_));
 sg13g2_xnor2_1 _5375_ (.Y(_0467_),
    .A(_0463_),
    .B(_0466_));
 sg13g2_xnor2_1 _5376_ (.Y(_0468_),
    .A(_0462_),
    .B(_0467_));
 sg13g2_nor2_1 _5377_ (.A(_0460_),
    .B(_0457_),
    .Y(_0469_));
 sg13g2_a21oi_1 _5378_ (.A1(_0461_),
    .A2(_0468_),
    .Y(_0470_),
    .B1(_0469_));
 sg13g2_nand2_1 _5379_ (.Y(_0471_),
    .A(_0450_),
    .B(_0470_));
 sg13g2_and2_1 _5380_ (.A(_0466_),
    .B(_0463_),
    .X(_0472_));
 sg13g2_nor2b_1 _5381_ (.A(_0467_),
    .B_N(_0462_),
    .Y(_0473_));
 sg13g2_nor2_1 _5382_ (.A(_0472_),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_inv_1 _5383_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_inv_1 _5384_ (.Y(_0476_),
    .A(_0470_));
 sg13g2_nand3_1 _5385_ (.B(_0445_),
    .C(_0449_),
    .A(_0476_),
    .Y(_0477_));
 sg13g2_inv_1 _5386_ (.Y(_0478_),
    .A(_0477_));
 sg13g2_a21oi_1 _5387_ (.A1(_0471_),
    .A2(_0475_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_o21ai_1 _5388_ (.B1(_0439_),
    .Y(_0480_),
    .A1(_0441_),
    .A2(_4387_));
 sg13g2_nor3_1 _5389_ (.A(_0441_),
    .B(_4387_),
    .C(_0439_),
    .Y(_0481_));
 sg13g2_a21oi_1 _5390_ (.A1(_0480_),
    .A2(_0437_),
    .Y(_0482_),
    .B1(_0481_));
 sg13g2_nor2_1 _5391_ (.A(_0306_),
    .B(_4390_),
    .Y(_0483_));
 sg13g2_nand3_1 _5392_ (.B(_0367_),
    .C(_4268_),
    .A(_4264_),
    .Y(_0484_));
 sg13g2_xnor2_1 _5393_ (.Y(_0485_),
    .A(_0483_),
    .B(_0484_));
 sg13g2_nor2_1 _5394_ (.A(_0465_),
    .B(_4368_),
    .Y(_0486_));
 sg13g2_nor2_1 _5395_ (.A(net158),
    .B(net83),
    .Y(_0487_));
 sg13g2_inv_1 _5396_ (.Y(_0488_),
    .A(_0487_));
 sg13g2_nand2_1 _5397_ (.Y(_0489_),
    .A(_4382_),
    .B(net159));
 sg13g2_nor2_1 _5398_ (.A(_0488_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_nand2_1 _5399_ (.Y(_0491_),
    .A(_0489_),
    .B(_0488_));
 sg13g2_nand2b_1 _5400_ (.Y(_0492_),
    .B(_0491_),
    .A_N(_0490_));
 sg13g2_nand2b_1 _5401_ (.Y(_0493_),
    .B(_0492_),
    .A_N(_0486_));
 sg13g2_nand3b_1 _5402_ (.B(_0486_),
    .C(_0491_),
    .Y(_0494_),
    .A_N(_0490_));
 sg13g2_nand2_1 _5403_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_nand2_1 _5404_ (.Y(_0496_),
    .A(_0420_),
    .B(_0418_));
 sg13g2_nor2_1 _5405_ (.A(_0418_),
    .B(_0420_),
    .Y(_0497_));
 sg13g2_a21oi_1 _5406_ (.A1(_0496_),
    .A2(_0412_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_nand2_1 _5407_ (.Y(_0499_),
    .A(_0495_),
    .B(_0498_));
 sg13g2_inv_1 _5408_ (.Y(_0500_),
    .A(_0498_));
 sg13g2_nand3_1 _5409_ (.B(_0494_),
    .C(_0500_),
    .A(_0493_),
    .Y(_0501_));
 sg13g2_nand2_1 _5410_ (.Y(_0502_),
    .A(_0499_),
    .B(_0501_));
 sg13g2_nand2b_1 _5411_ (.Y(_0503_),
    .B(_0502_),
    .A_N(_0485_));
 sg13g2_nand3_1 _5412_ (.B(_0501_),
    .C(_0485_),
    .A(_0499_),
    .Y(_0504_));
 sg13g2_nand2_1 _5413_ (.Y(_0505_),
    .A(_0503_),
    .B(_0504_));
 sg13g2_inv_1 _5414_ (.Y(_0506_),
    .A(_0435_));
 sg13g2_a21oi_1 _5415_ (.A1(_0433_),
    .A2(_0444_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_nand2_1 _5416_ (.Y(_0508_),
    .A(_0505_),
    .B(_0507_));
 sg13g2_inv_1 _5417_ (.Y(_0509_),
    .A(_0507_));
 sg13g2_nand3_1 _5418_ (.B(_0504_),
    .C(_0509_),
    .A(_0503_),
    .Y(_0510_));
 sg13g2_nand2_1 _5419_ (.Y(_0511_),
    .A(_0508_),
    .B(_0510_));
 sg13g2_xnor2_1 _5420_ (.Y(_0512_),
    .A(_0482_),
    .B(_0511_));
 sg13g2_xor2_1 _5421_ (.B(_0512_),
    .A(_0479_),
    .X(_0513_));
 sg13g2_nand3_1 _5422_ (.B(_0471_),
    .C(_0475_),
    .A(_0477_),
    .Y(_0514_));
 sg13g2_nand2_1 _5423_ (.Y(_0515_),
    .A(_0450_),
    .B(_0476_));
 sg13g2_nand3_1 _5424_ (.B(_0449_),
    .C(_0470_),
    .A(_0445_),
    .Y(_0516_));
 sg13g2_nand3_1 _5425_ (.B(_0516_),
    .C(_0474_),
    .A(_0515_),
    .Y(_0517_));
 sg13g2_nand2_1 _5426_ (.Y(_0518_),
    .A(_0514_),
    .B(_0517_));
 sg13g2_nand2b_1 _5427_ (.Y(_0519_),
    .B(_0457_),
    .A_N(_0460_));
 sg13g2_nand3_1 _5428_ (.B(_0455_),
    .C(_0456_),
    .A(_0460_),
    .Y(_0520_));
 sg13g2_nand3b_1 _5429_ (.B(_0519_),
    .C(_0520_),
    .Y(_0521_),
    .A_N(_0468_));
 sg13g2_nand2_1 _5430_ (.Y(_0522_),
    .A(_0519_),
    .B(_0520_));
 sg13g2_nand2_1 _5431_ (.Y(_0523_),
    .A(_0522_),
    .B(_0468_));
 sg13g2_nand2_1 _5432_ (.Y(_0524_),
    .A(_0521_),
    .B(_0523_));
 sg13g2_nand2_1 _5433_ (.Y(_0525_),
    .A(_0357_),
    .B(_0346_));
 sg13g2_nor2_1 _5434_ (.A(_0346_),
    .B(_0357_),
    .Y(_0526_));
 sg13g2_a21oi_2 _5435_ (.B1(_0526_),
    .Y(_0527_),
    .A2(_0344_),
    .A1(_0525_));
 sg13g2_nand2_1 _5436_ (.Y(_0528_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_nor2_1 _5437_ (.A(_0368_),
    .B(_0308_),
    .Y(_0529_));
 sg13g2_nor2_1 _5438_ (.A(_0436_),
    .B(_4328_),
    .Y(_0530_));
 sg13g2_or2_1 _5439_ (.X(_0531_),
    .B(_0342_),
    .A(_0341_));
 sg13g2_a22oi_1 _5440_ (.Y(_0532_),
    .B1(_0340_),
    .B2(_0531_),
    .A2(_0463_),
    .A1(_0293_));
 sg13g2_xnor2_1 _5441_ (.Y(_0533_),
    .A(_0530_),
    .B(_0532_));
 sg13g2_xnor2_1 _5442_ (.Y(_0534_),
    .A(_0529_),
    .B(_0533_));
 sg13g2_inv_1 _5443_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_nor2_1 _5444_ (.A(_0527_),
    .B(_0524_),
    .Y(_0536_));
 sg13g2_a21oi_2 _5445_ (.B1(_0536_),
    .Y(_0537_),
    .A2(_0535_),
    .A1(_0528_));
 sg13g2_nand2_1 _5446_ (.Y(_0538_),
    .A(_0518_),
    .B(_0537_));
 sg13g2_nor2b_1 _5447_ (.A(_0532_),
    .B_N(_0530_),
    .Y(_0539_));
 sg13g2_a21oi_1 _5448_ (.A1(_0533_),
    .A2(_0529_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_inv_1 _5449_ (.Y(_0541_),
    .A(_0540_));
 sg13g2_nor2_1 _5450_ (.A(_0537_),
    .B(_0518_),
    .Y(_0542_));
 sg13g2_a21oi_1 _5451_ (.A1(_0538_),
    .A2(_0541_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_nand2b_1 _5452_ (.Y(_0544_),
    .B(_0543_),
    .A_N(_0513_));
 sg13g2_nand2b_1 _5453_ (.Y(_0545_),
    .B(_0513_),
    .A_N(_0543_));
 sg13g2_nand2_2 _5454_ (.Y(_0546_),
    .A(_0544_),
    .B(_0545_));
 sg13g2_inv_1 _5455_ (.Y(_0547_),
    .A(_0482_));
 sg13g2_inv_1 _5456_ (.Y(_0548_),
    .A(_0510_));
 sg13g2_a21oi_1 _5457_ (.A1(_0508_),
    .A2(_0547_),
    .Y(_0549_),
    .B1(_0548_));
 sg13g2_nor2b_1 _5458_ (.A(_0484_),
    .B_N(_0483_),
    .Y(_0550_));
 sg13g2_and2_1 _5459_ (.A(_0504_),
    .B(_0501_),
    .X(_0551_));
 sg13g2_buf_1 _5460_ (.A(_0551_),
    .X(_0552_));
 sg13g2_nor2_1 _5461_ (.A(_0436_),
    .B(_4390_),
    .Y(_0553_));
 sg13g2_a21oi_1 _5462_ (.A1(_0491_),
    .A2(_0486_),
    .Y(_0554_),
    .B1(_0490_));
 sg13g2_nor2_1 _5463_ (.A(_0441_),
    .B(_4368_),
    .Y(_0555_));
 sg13g2_nor2_1 _5464_ (.A(net159),
    .B(_4534_),
    .Y(_0556_));
 sg13g2_nand2_1 _5465_ (.Y(_0557_),
    .A(_4382_),
    .B(_0464_));
 sg13g2_xnor2_1 _5466_ (.Y(_0558_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_xnor2_1 _5467_ (.Y(_0559_),
    .A(_0555_),
    .B(_0558_));
 sg13g2_nor2_1 _5468_ (.A(_0554_),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_nand2_1 _5469_ (.Y(_0561_),
    .A(_0559_),
    .B(_0554_));
 sg13g2_nor2b_1 _5470_ (.A(_0560_),
    .B_N(_0561_),
    .Y(_0562_));
 sg13g2_xnor2_1 _5471_ (.Y(_0563_),
    .A(_0553_),
    .B(_0562_));
 sg13g2_xnor2_1 _5472_ (.Y(_0564_),
    .A(_0552_),
    .B(_0563_));
 sg13g2_xnor2_1 _5473_ (.Y(_0565_),
    .A(_0550_),
    .B(_0564_));
 sg13g2_xor2_1 _5474_ (.B(_0565_),
    .A(_0549_),
    .X(_0566_));
 sg13g2_nor2_1 _5475_ (.A(_0479_),
    .B(_0512_),
    .Y(_0567_));
 sg13g2_nand2b_1 _5476_ (.Y(_0568_),
    .B(_0567_),
    .A_N(_0566_));
 sg13g2_nand2b_1 _5477_ (.Y(_0569_),
    .B(_0566_),
    .A_N(_0567_));
 sg13g2_nand2_1 _5478_ (.Y(_0570_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_buf_2 _5479_ (.A(_0570_),
    .X(_0571_));
 sg13g2_nand2_1 _5480_ (.Y(_0572_),
    .A(_0378_),
    .B(_0336_));
 sg13g2_nor2_1 _5481_ (.A(_0336_),
    .B(_0378_),
    .Y(_0573_));
 sg13g2_a21oi_2 _5482_ (.B1(_0573_),
    .Y(_0574_),
    .A2(_0384_),
    .A1(_0572_));
 sg13g2_nand2_1 _5483_ (.Y(_0575_),
    .A(_0363_),
    .B(_0339_));
 sg13g2_nor2_1 _5484_ (.A(_0339_),
    .B(_0363_),
    .Y(_0576_));
 sg13g2_a21oi_2 _5485_ (.B1(_0576_),
    .Y(_0577_),
    .A2(_0374_),
    .A1(_0575_));
 sg13g2_nand2b_1 _5486_ (.Y(_0578_),
    .B(_0524_),
    .A_N(_0527_));
 sg13g2_nand3_1 _5487_ (.B(_0523_),
    .C(_0527_),
    .A(_0521_),
    .Y(_0579_));
 sg13g2_nand2_1 _5488_ (.Y(_0580_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_nand2_1 _5489_ (.Y(_0581_),
    .A(_0580_),
    .B(_0535_));
 sg13g2_nand3_1 _5490_ (.B(_0579_),
    .C(_0534_),
    .A(_0578_),
    .Y(_0582_));
 sg13g2_nand2_1 _5491_ (.Y(_0583_),
    .A(_0581_),
    .B(_0582_));
 sg13g2_nand2b_1 _5492_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0577_));
 sg13g2_nand3_1 _5493_ (.B(_0577_),
    .C(_0582_),
    .A(_0581_),
    .Y(_0585_));
 sg13g2_nand2_1 _5494_ (.Y(_0586_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_nor2b_1 _5495_ (.A(_0372_),
    .B_N(_0369_),
    .Y(_0587_));
 sg13g2_a21oi_1 _5496_ (.A1(_0373_),
    .A2(_0309_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_inv_1 _5497_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_nand2_1 _5498_ (.Y(_0590_),
    .A(_0586_),
    .B(_0589_));
 sg13g2_nand3_1 _5499_ (.B(_0585_),
    .C(_0588_),
    .A(_0584_),
    .Y(_0591_));
 sg13g2_nand2_2 _5500_ (.Y(_0592_),
    .A(_0590_),
    .B(_0591_));
 sg13g2_xor2_1 _5501_ (.B(_0592_),
    .A(_0574_),
    .X(_0593_));
 sg13g2_nand2_1 _5502_ (.Y(_0594_),
    .A(_0583_),
    .B(_0577_));
 sg13g2_nor2_1 _5503_ (.A(_0577_),
    .B(_0583_),
    .Y(_0595_));
 sg13g2_a21oi_1 _5504_ (.A1(_0594_),
    .A2(_0589_),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_inv_1 _5505_ (.Y(_0597_),
    .A(_0596_));
 sg13g2_nand3_1 _5506_ (.B(_0514_),
    .C(_0517_),
    .A(_0537_),
    .Y(_0598_));
 sg13g2_inv_1 _5507_ (.Y(_0599_),
    .A(_0537_));
 sg13g2_nand2_1 _5508_ (.Y(_0600_),
    .A(_0518_),
    .B(_0599_));
 sg13g2_nand2_1 _5509_ (.Y(_0601_),
    .A(_0598_),
    .B(_0600_));
 sg13g2_nand2_1 _5510_ (.Y(_0602_),
    .A(_0601_),
    .B(_0541_));
 sg13g2_nand3_1 _5511_ (.B(_0598_),
    .C(_0540_),
    .A(_0600_),
    .Y(_0603_));
 sg13g2_nand2_1 _5512_ (.Y(_0604_),
    .A(_0602_),
    .B(_0603_));
 sg13g2_xnor2_1 _5513_ (.Y(_0605_),
    .A(_0597_),
    .B(_0604_));
 sg13g2_nand2_1 _5514_ (.Y(_0606_),
    .A(_0593_),
    .B(_0605_));
 sg13g2_nor3_1 _5515_ (.A(_0546_),
    .B(_0571_),
    .C(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _5516_ (.Y(_0608_),
    .A(_0409_),
    .B(_0607_));
 sg13g2_nor2_1 _5517_ (.A(_0574_),
    .B(_0592_),
    .Y(_0609_));
 sg13g2_nand2_1 _5518_ (.Y(_0610_),
    .A(_0604_),
    .B(_0596_));
 sg13g2_nand2_1 _5519_ (.Y(_0611_),
    .A(_0609_),
    .B(_0610_));
 sg13g2_nand3_1 _5520_ (.B(_0602_),
    .C(_0603_),
    .A(_0597_),
    .Y(_0612_));
 sg13g2_nand2_1 _5521_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_nor2_1 _5522_ (.A(_0546_),
    .B(_0571_),
    .Y(_0614_));
 sg13g2_o21ai_1 _5523_ (.B1(_0568_),
    .Y(_0615_),
    .A1(_0545_),
    .A2(_0571_));
 sg13g2_a21oi_1 _5524_ (.A1(_0613_),
    .A2(_0614_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_nand2_1 _5525_ (.Y(_0617_),
    .A(_0608_),
    .B(_0616_));
 sg13g2_nor2b_1 _5526_ (.A(_0557_),
    .B_N(_0556_),
    .Y(_0618_));
 sg13g2_a21oi_1 _5527_ (.A1(_0558_),
    .A2(_0555_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nor2_1 _5528_ (.A(_0436_),
    .B(net84),
    .Y(_0620_));
 sg13g2_nor2_1 _5529_ (.A(_0464_),
    .B(_4534_),
    .Y(_0621_));
 sg13g2_nand2_1 _5530_ (.Y(_0622_),
    .A(_4382_),
    .B(_0440_));
 sg13g2_xnor2_1 _5531_ (.Y(_0623_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_xnor2_1 _5532_ (.Y(_0624_),
    .A(_0620_),
    .B(_0623_));
 sg13g2_xor2_1 _5533_ (.B(_0624_),
    .A(_0619_),
    .X(_0625_));
 sg13g2_a21oi_1 _5534_ (.A1(_0561_),
    .A2(_0553_),
    .Y(_0626_),
    .B1(_0560_));
 sg13g2_xor2_1 _5535_ (.B(_0626_),
    .A(_0625_),
    .X(_0627_));
 sg13g2_nand2_1 _5536_ (.Y(_0628_),
    .A(_0563_),
    .B(_0552_));
 sg13g2_nor2_1 _5537_ (.A(_0552_),
    .B(_0563_),
    .Y(_0629_));
 sg13g2_a21oi_1 _5538_ (.A1(_0628_),
    .A2(_0550_),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_xnor2_1 _5539_ (.Y(_0631_),
    .A(_0627_),
    .B(_0630_));
 sg13g2_nand2b_1 _5540_ (.Y(_0632_),
    .B(_0565_),
    .A_N(_0549_));
 sg13g2_nor2_1 _5541_ (.A(_0631_),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_nand2_1 _5542_ (.Y(_0634_),
    .A(_0632_),
    .B(_0631_));
 sg13g2_inv_1 _5543_ (.Y(_0635_),
    .A(_0634_));
 sg13g2_nor2_1 _5544_ (.A(_0633_),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_inv_1 _5545_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_nand2_1 _5546_ (.Y(_0638_),
    .A(_0617_),
    .B(_0637_));
 sg13g2_nand3_1 _5547_ (.B(_0616_),
    .C(_0636_),
    .A(_0608_),
    .Y(_0639_));
 sg13g2_buf_1 _5548_ (.A(net92),
    .X(_0640_));
 sg13g2_inv_1 _5549_ (.Y(_0641_),
    .A(_4277_));
 sg13g2_nand2_1 _5550_ (.Y(_0642_),
    .A(_0641_),
    .B(net154));
 sg13g2_nor2_1 _5551_ (.A(net153),
    .B(_4168_),
    .Y(_0643_));
 sg13g2_nand2_1 _5552_ (.Y(_0644_),
    .A(_4273_),
    .B(_4153_));
 sg13g2_nor2_1 _5553_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_inv_1 _5554_ (.Y(_0646_),
    .A(_0642_));
 sg13g2_buf_1 _5555_ (.A(_4154_),
    .X(_0647_));
 sg13g2_inv_1 _5556_ (.Y(_0648_),
    .A(net151));
 sg13g2_buf_1 _5557_ (.A(_0648_),
    .X(_0649_));
 sg13g2_o21ai_1 _5558_ (.B1(net132),
    .Y(_0650_),
    .A1(_0645_),
    .A2(_0646_));
 sg13g2_a21oi_1 _5559_ (.A1(_4169_),
    .A2(_0642_),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_inv_1 _5560_ (.Y(_0652_),
    .A(_0651_));
 sg13g2_nor2_1 _5561_ (.A(net153),
    .B(net163),
    .Y(_0653_));
 sg13g2_buf_1 _5562_ (.A(_0033_),
    .X(_0654_));
 sg13g2_inv_1 _5563_ (.Y(_0655_),
    .A(_0654_));
 sg13g2_a21oi_1 _5564_ (.A1(_0653_),
    .A2(_0655_),
    .Y(_0656_),
    .B1(_4153_));
 sg13g2_nor2_1 _5565_ (.A(net154),
    .B(_4149_),
    .Y(_0657_));
 sg13g2_o21ai_1 _5566_ (.B1(net151),
    .Y(_0658_),
    .A1(_0656_),
    .A2(_0657_));
 sg13g2_a21o_1 _5567_ (.A2(_0658_),
    .A1(_0652_),
    .B1(_4160_),
    .X(_0659_));
 sg13g2_inv_1 _5568_ (.Y(_0660_),
    .A(_0032_));
 sg13g2_o21ai_1 _5569_ (.B1(_4302_),
    .Y(_0661_),
    .A1(_4153_),
    .A2(_0660_));
 sg13g2_a21oi_1 _5570_ (.A1(_0661_),
    .A2(_0648_),
    .Y(_0662_),
    .B1(_4217_));
 sg13g2_buf_1 _5571_ (.A(net154),
    .X(_0663_));
 sg13g2_nor2_1 _5572_ (.A(_0034_),
    .B(_4191_),
    .Y(_0664_));
 sg13g2_inv_1 _5573_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_nor3_1 _5574_ (.A(_0663_),
    .B(_0654_),
    .C(_0665_),
    .Y(_0666_));
 sg13g2_buf_1 _5575_ (.A(net151),
    .X(_0667_));
 sg13g2_nand2_1 _5576_ (.Y(_0668_),
    .A(_0666_),
    .B(net140));
 sg13g2_nor2_1 _5577_ (.A(_4146_),
    .B(_4145_),
    .Y(_0669_));
 sg13g2_nor2_1 _5578_ (.A(_0669_),
    .B(_4198_),
    .Y(_0670_));
 sg13g2_nor2_1 _5579_ (.A(net153),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_buf_1 _5580_ (.A(_4153_),
    .X(_0672_));
 sg13g2_o21ai_1 _5581_ (.B1(net139),
    .Y(_0673_),
    .A1(_4145_),
    .A2(_4273_));
 sg13g2_inv_1 _5582_ (.Y(_0674_),
    .A(_0034_));
 sg13g2_nand2_2 _5583_ (.Y(_0675_),
    .A(_4274_),
    .B(_0674_));
 sg13g2_nor2_2 _5584_ (.A(net139),
    .B(_4184_),
    .Y(_0676_));
 sg13g2_nand2_1 _5585_ (.Y(_0677_),
    .A(_0675_),
    .B(_0676_));
 sg13g2_o21ai_1 _5586_ (.B1(_0677_),
    .Y(_0678_),
    .A1(_0671_),
    .A2(_0673_));
 sg13g2_nand2_1 _5587_ (.Y(_0679_),
    .A(_0678_),
    .B(net140));
 sg13g2_nor2_1 _5588_ (.A(_4163_),
    .B(_4182_),
    .Y(_0680_));
 sg13g2_nor3_1 _5589_ (.A(net139),
    .B(_4181_),
    .C(_0643_),
    .Y(_0681_));
 sg13g2_o21ai_1 _5590_ (.B1(_0648_),
    .Y(_0682_),
    .A1(_0680_),
    .A2(_0681_));
 sg13g2_nor2_1 _5591_ (.A(net162),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_inv_1 _5592_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_a21oi_1 _5593_ (.A1(net139),
    .A2(_4167_),
    .Y(_0685_),
    .B1(net153));
 sg13g2_inv_1 _5594_ (.Y(_0686_),
    .A(net162));
 sg13g2_nor2_1 _5595_ (.A(net151),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_nor2b_1 _5596_ (.A(_0685_),
    .B_N(_0687_),
    .Y(_0688_));
 sg13g2_nor2_1 _5597_ (.A(net153),
    .B(_4145_),
    .Y(_0689_));
 sg13g2_nand2_1 _5598_ (.Y(_0690_),
    .A(_0689_),
    .B(net163));
 sg13g2_nand2_1 _5599_ (.Y(_0691_),
    .A(_0688_),
    .B(_0690_));
 sg13g2_nand3_1 _5600_ (.B(_0684_),
    .C(_0691_),
    .A(_0679_),
    .Y(_0692_));
 sg13g2_nor2_1 _5601_ (.A(_4151_),
    .B(net92),
    .Y(_0693_));
 sg13g2_buf_2 _5602_ (.A(_0693_),
    .X(_0694_));
 sg13g2_inv_1 _5603_ (.Y(_0695_),
    .A(_0694_));
 sg13g2_a221oi_1 _5604_ (.B2(_4188_),
    .C1(_0695_),
    .B1(_0692_),
    .A1(_0662_),
    .Y(_0696_),
    .A2(_0668_));
 sg13g2_a22oi_1 _5605_ (.Y(_0697_),
    .B1(_0659_),
    .B2(_0696_),
    .A2(net86),
    .A1(_0046_));
 sg13g2_inv_1 _5606_ (.Y(_0698_),
    .A(_0697_));
 sg13g2_nand3_1 _5607_ (.B(_0639_),
    .C(_0698_),
    .A(_0638_),
    .Y(_0699_));
 sg13g2_buf_1 _5608_ (.A(_0699_),
    .X(_0700_));
 sg13g2_nand2_1 _5609_ (.Y(_0701_),
    .A(_0617_),
    .B(_0636_));
 sg13g2_nand3_1 _5610_ (.B(_0616_),
    .C(_0637_),
    .A(_0608_),
    .Y(_0702_));
 sg13g2_nand3_1 _5611_ (.B(_0702_),
    .C(_0697_),
    .A(_0701_),
    .Y(_0703_));
 sg13g2_buf_1 _5612_ (.A(net102),
    .X(_0704_));
 sg13g2_buf_1 _5613_ (.A(net91),
    .X(_0705_));
 sg13g2_buf_2 _5614_ (.A(\i_display.i_vga.vblank ),
    .X(_0706_));
 sg13g2_nor2_2 _5615_ (.A(_0706_),
    .B(\i_display.i_vga.hblank ),
    .Y(_0707_));
 sg13g2_inv_4 _5616_ (.A(_0707_),
    .Y(_0708_));
 sg13g2_buf_1 _5617_ (.A(_0708_),
    .X(_0709_));
 sg13g2_nor2_1 _5618_ (.A(_0047_),
    .B(net131),
    .Y(_0710_));
 sg13g2_buf_1 _5619_ (.A(_0706_),
    .X(_0711_));
 sg13g2_inv_1 _5620_ (.Y(_0712_),
    .A(\i_display.i_vga.timing_ver.counter[9] ));
 sg13g2_nor2_1 _5621_ (.A(net150),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_inv_1 _5622_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_nor2_1 _5623_ (.A(_0714_),
    .B(net85),
    .Y(_0715_));
 sg13g2_a21o_1 _5624_ (.A2(_0710_),
    .A1(net85),
    .B1(_0715_),
    .X(_0716_));
 sg13g2_nand3_1 _5625_ (.B(_0703_),
    .C(_0716_),
    .A(_0700_),
    .Y(_0717_));
 sg13g2_nand3_1 _5626_ (.B(_0702_),
    .C(_0698_),
    .A(_0701_),
    .Y(_0718_));
 sg13g2_nand3_1 _5627_ (.B(_0639_),
    .C(_0697_),
    .A(_0638_),
    .Y(_0719_));
 sg13g2_inv_1 _5628_ (.Y(_0720_),
    .A(_0716_));
 sg13g2_nand3_1 _5629_ (.B(_0719_),
    .C(_0720_),
    .A(_0718_),
    .Y(_0721_));
 sg13g2_nand2_1 _5630_ (.Y(_0722_),
    .A(_0717_),
    .B(_0721_));
 sg13g2_xnor2_1 _5631_ (.Y(_0723_),
    .A(_0574_),
    .B(_0592_));
 sg13g2_nand2_1 _5632_ (.Y(_0724_),
    .A(_0409_),
    .B(_0723_));
 sg13g2_nand3_1 _5633_ (.B(_0593_),
    .C(_0408_),
    .A(_0403_),
    .Y(_0725_));
 sg13g2_inv_1 _5634_ (.Y(_0726_),
    .A(_4155_));
 sg13g2_nand2_1 _5635_ (.Y(_0727_),
    .A(_0664_),
    .B(_4145_));
 sg13g2_nor2_1 _5636_ (.A(_4255_),
    .B(_0689_),
    .Y(_0728_));
 sg13g2_inv_1 _5637_ (.Y(_0729_),
    .A(_0728_));
 sg13g2_a21oi_1 _5638_ (.A1(_0729_),
    .A2(_4168_),
    .Y(_0730_),
    .B1(_4177_));
 sg13g2_a21o_1 _5639_ (.A2(_0727_),
    .A1(_0726_),
    .B1(_0730_),
    .X(_0731_));
 sg13g2_o21ai_1 _5640_ (.B1(_4161_),
    .Y(_0732_),
    .A1(_0731_),
    .A2(_0651_));
 sg13g2_nor2_1 _5641_ (.A(_0034_),
    .B(_4273_),
    .Y(_0733_));
 sg13g2_inv_1 _5642_ (.Y(_0734_),
    .A(_0733_));
 sg13g2_nor2_1 _5643_ (.A(net155),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_nor2_1 _5644_ (.A(net141),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_inv_1 _5645_ (.Y(_0737_),
    .A(_0736_));
 sg13g2_o21ai_1 _5646_ (.B1(net141),
    .Y(_0738_),
    .A1(net140),
    .A2(_4148_));
 sg13g2_nand2_1 _5647_ (.Y(_0739_),
    .A(_0737_),
    .B(_0738_));
 sg13g2_a21oi_1 _5648_ (.A1(_0733_),
    .A2(_0655_),
    .Y(_0740_),
    .B1(net139));
 sg13g2_o21ai_1 _5649_ (.B1(net140),
    .Y(_0741_),
    .A1(_0740_),
    .A2(_0736_));
 sg13g2_nand2_1 _5650_ (.Y(_0742_),
    .A(_4273_),
    .B(_4145_));
 sg13g2_nor2_1 _5651_ (.A(_0653_),
    .B(_4255_),
    .Y(_0743_));
 sg13g2_inv_1 _5652_ (.Y(_0744_),
    .A(_0743_));
 sg13g2_o21ai_1 _5653_ (.B1(_0744_),
    .Y(_0745_),
    .A1(net141),
    .A2(_0742_));
 sg13g2_nand2_1 _5654_ (.Y(_0746_),
    .A(_0745_),
    .B(_0687_));
 sg13g2_nand3_1 _5655_ (.B(_0684_),
    .C(_0746_),
    .A(_0741_),
    .Y(_0747_));
 sg13g2_a221oi_1 _5656_ (.B2(_4188_),
    .C1(_0695_),
    .B1(_0747_),
    .A1(_4189_),
    .Y(_0748_),
    .A2(_0739_));
 sg13g2_a22oi_1 _5657_ (.Y(_0749_),
    .B1(_0732_),
    .B2(_0748_),
    .A2(net92),
    .A1(_0042_));
 sg13g2_inv_1 _5658_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nand3_1 _5659_ (.B(_0725_),
    .C(_0750_),
    .A(_0724_),
    .Y(_0751_));
 sg13g2_buf_1 _5660_ (.A(_0751_),
    .X(_0752_));
 sg13g2_nand2_1 _5661_ (.Y(_0753_),
    .A(_0409_),
    .B(_0593_));
 sg13g2_nand3_1 _5662_ (.B(_0723_),
    .C(_0408_),
    .A(_0403_),
    .Y(_0754_));
 sg13g2_nand3_1 _5663_ (.B(_0754_),
    .C(_0749_),
    .A(_0753_),
    .Y(_0755_));
 sg13g2_nand2_1 _5664_ (.Y(_0756_),
    .A(_0752_),
    .B(_0755_));
 sg13g2_nand3b_1 _5665_ (.B(_0690_),
    .C(_0727_),
    .Y(_0757_),
    .A_N(_0673_));
 sg13g2_o21ai_1 _5666_ (.B1(_0675_),
    .Y(_0758_),
    .A1(_4216_),
    .A2(_0676_));
 sg13g2_a21oi_1 _5667_ (.A1(_0757_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(net132));
 sg13g2_a22oi_1 _5668_ (.Y(_0760_),
    .B1(net155),
    .B2(_4216_),
    .A2(net141),
    .A1(net153));
 sg13g2_o21ai_1 _5669_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_4149_),
    .A2(_0644_));
 sg13g2_a21o_1 _5670_ (.A2(_0761_),
    .A1(_0687_),
    .B1(_0683_),
    .X(_0762_));
 sg13g2_o21ai_1 _5671_ (.B1(_4188_),
    .Y(_0763_),
    .A1(_0759_),
    .A2(_0762_));
 sg13g2_a21oi_1 _5672_ (.A1(net153),
    .A2(net139),
    .Y(_0764_),
    .B1(_4148_));
 sg13g2_a21oi_1 _5673_ (.A1(_0764_),
    .A2(net132),
    .Y(_0765_),
    .B1(_4217_));
 sg13g2_nor2_1 _5674_ (.A(_4216_),
    .B(_0676_),
    .Y(_0766_));
 sg13g2_nand3_1 _5675_ (.B(net140),
    .C(_0766_),
    .A(_0757_),
    .Y(_0767_));
 sg13g2_nor2_1 _5676_ (.A(_4155_),
    .B(_0735_),
    .Y(_0768_));
 sg13g2_nor2_1 _5677_ (.A(_0730_),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_nand2_1 _5678_ (.Y(_0770_),
    .A(_0652_),
    .B(_0769_));
 sg13g2_a221oi_1 _5679_ (.B2(_4161_),
    .C1(_0695_),
    .B1(_0770_),
    .A1(_0765_),
    .Y(_0771_),
    .A2(_0767_));
 sg13g2_a22oi_1 _5680_ (.Y(_0772_),
    .B1(_0763_),
    .B2(_0771_),
    .A2(net86),
    .A1(_0043_));
 sg13g2_nand2_1 _5681_ (.Y(_0773_),
    .A(_0406_),
    .B(_0404_));
 sg13g2_nor2_1 _5682_ (.A(_0773_),
    .B(_0723_),
    .Y(_0774_));
 sg13g2_nand3_1 _5683_ (.B(_0394_),
    .C(_0395_),
    .A(_0398_),
    .Y(_0775_));
 sg13g2_a21oi_1 _5684_ (.A1(_0775_),
    .A2(_0267_),
    .Y(_0776_),
    .B1(_0399_));
 sg13g2_nor2_1 _5685_ (.A(_0332_),
    .B(_0387_),
    .Y(_0777_));
 sg13g2_nor2_1 _5686_ (.A(_0777_),
    .B(_0609_),
    .Y(_0778_));
 sg13g2_nand2_1 _5687_ (.Y(_0779_),
    .A(_0592_),
    .B(_0574_));
 sg13g2_nor2b_1 _5688_ (.A(_0778_),
    .B_N(_0779_),
    .Y(_0780_));
 sg13g2_a21oi_1 _5689_ (.A1(_0774_),
    .A2(_0776_),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_nand2_1 _5690_ (.Y(_0782_),
    .A(_0263_),
    .B(_4524_));
 sg13g2_nand2_1 _5691_ (.Y(_0783_),
    .A(_0782_),
    .B(_0267_));
 sg13g2_nand2_1 _5692_ (.Y(_0784_),
    .A(_0396_),
    .B(_0390_));
 sg13g2_nand2_1 _5693_ (.Y(_0785_),
    .A(_0775_),
    .B(_0784_));
 sg13g2_nor2_1 _5694_ (.A(_0783_),
    .B(_0785_),
    .Y(_0786_));
 sg13g2_nand3_1 _5695_ (.B(_0786_),
    .C(_4522_),
    .A(_0774_),
    .Y(_0787_));
 sg13g2_nand2_1 _5696_ (.Y(_0788_),
    .A(_0781_),
    .B(_0787_));
 sg13g2_nand2_1 _5697_ (.Y(_0789_),
    .A(_0788_),
    .B(_0605_));
 sg13g2_nand2_1 _5698_ (.Y(_0790_),
    .A(_0612_),
    .B(_0610_));
 sg13g2_nand3_1 _5699_ (.B(_0787_),
    .C(_0790_),
    .A(_0781_),
    .Y(_0791_));
 sg13g2_nand2_1 _5700_ (.Y(_0792_),
    .A(_0789_),
    .B(_0791_));
 sg13g2_nand2b_1 _5701_ (.Y(_0793_),
    .B(_0792_),
    .A_N(_0772_));
 sg13g2_nand3_1 _5702_ (.B(_0791_),
    .C(_0772_),
    .A(_0789_),
    .Y(_0794_));
 sg13g2_nand2_1 _5703_ (.Y(_0795_),
    .A(_0793_),
    .B(_0794_));
 sg13g2_nor2_1 _5704_ (.A(_0756_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_nor2_1 _5705_ (.A(net155),
    .B(net154),
    .Y(_0797_));
 sg13g2_a21oi_1 _5706_ (.A1(_0734_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(_0645_));
 sg13g2_buf_1 _5707_ (.A(_0031_),
    .X(_0799_));
 sg13g2_inv_1 _5708_ (.Y(_0800_),
    .A(_0799_));
 sg13g2_nand3_1 _5709_ (.B(_0798_),
    .C(_0800_),
    .A(_0758_),
    .Y(_0801_));
 sg13g2_nand3_1 _5710_ (.B(_0798_),
    .C(net151),
    .A(_0758_),
    .Y(_0802_));
 sg13g2_a21oi_1 _5711_ (.A1(_4255_),
    .A2(_0648_),
    .Y(_0803_),
    .B1(_4258_));
 sg13g2_a22oi_1 _5712_ (.Y(_0804_),
    .B1(_0802_),
    .B2(_0803_),
    .A2(_4204_),
    .A1(_0801_));
 sg13g2_a21oi_1 _5713_ (.A1(_0642_),
    .A2(_0644_),
    .Y(_0805_),
    .B1(net151));
 sg13g2_o21ai_1 _5714_ (.B1(_0805_),
    .Y(_0806_),
    .A1(_4170_),
    .A2(_0646_));
 sg13g2_a21o_1 _5715_ (.A2(_0658_),
    .A1(_0806_),
    .B1(_0686_),
    .X(_0807_));
 sg13g2_nand4_1 _5716_ (.B(net151),
    .C(_0766_),
    .A(_0807_),
    .Y(_0808_),
    .D(_0798_));
 sg13g2_inv_1 _5717_ (.Y(_0809_),
    .A(_0662_));
 sg13g2_o21ai_1 _5718_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_4188_),
    .A2(_0807_));
 sg13g2_a21oi_1 _5719_ (.A1(_0808_),
    .A2(_0810_),
    .Y(_0811_),
    .B1(_0695_));
 sg13g2_a22oi_1 _5720_ (.Y(_0812_),
    .B1(_0804_),
    .B2(_0811_),
    .A2(net92),
    .A1(_0029_));
 sg13g2_inv_1 _5721_ (.Y(_0813_),
    .A(_4519_));
 sg13g2_inv_1 _5722_ (.Y(_0814_),
    .A(_4520_));
 sg13g2_nor2_1 _5723_ (.A(_4487_),
    .B(_0814_),
    .Y(_0815_));
 sg13g2_nand2_1 _5724_ (.Y(_0816_),
    .A(_0813_),
    .B(_0815_));
 sg13g2_nand2_1 _5725_ (.Y(_0817_),
    .A(_4455_),
    .B(_4458_));
 sg13g2_nand2_1 _5726_ (.Y(_0818_),
    .A(_0817_),
    .B(_4485_));
 sg13g2_nand2_1 _5727_ (.Y(_0819_),
    .A(_0818_),
    .B(_4520_));
 sg13g2_nand2_1 _5728_ (.Y(_0820_),
    .A(_4519_),
    .B(_0819_));
 sg13g2_nand2_1 _5729_ (.Y(_0821_),
    .A(_0816_),
    .B(_0820_));
 sg13g2_nand2b_1 _5730_ (.Y(_0822_),
    .B(_0821_),
    .A_N(_0812_));
 sg13g2_nand2b_1 _5731_ (.Y(_0823_),
    .B(_4508_),
    .A_N(_4518_));
 sg13g2_xor2_1 _5732_ (.B(_0823_),
    .A(_4517_),
    .X(_0824_));
 sg13g2_nor2_1 _5733_ (.A(_0101_),
    .B(net92),
    .Y(_0825_));
 sg13g2_nor2b_1 _5734_ (.A(_0824_),
    .B_N(_0825_),
    .Y(_0826_));
 sg13g2_nand3_1 _5735_ (.B(_0820_),
    .C(_0812_),
    .A(_0816_),
    .Y(_0827_));
 sg13g2_inv_1 _5736_ (.Y(_0828_),
    .A(_0827_));
 sg13g2_a21oi_1 _5737_ (.A1(_0822_),
    .A2(_0826_),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_inv_2 _5738_ (.Y(_0830_),
    .A(_0829_));
 sg13g2_a21oi_1 _5739_ (.A1(net151),
    .A2(_0656_),
    .Y(_0831_),
    .B1(_0768_));
 sg13g2_a21o_1 _5740_ (.A2(_0831_),
    .A1(_0806_),
    .B1(_4160_),
    .X(_0832_));
 sg13g2_a21oi_1 _5741_ (.A1(net154),
    .A2(_0653_),
    .Y(_0833_),
    .B1(_0676_));
 sg13g2_a21oi_1 _5742_ (.A1(net155),
    .A2(_0654_),
    .Y(_0834_),
    .B1(net154));
 sg13g2_nand2_1 _5743_ (.Y(_0835_),
    .A(_0665_),
    .B(_0834_));
 sg13g2_a21oi_1 _5744_ (.A1(_0833_),
    .A2(_0835_),
    .Y(_0836_),
    .B1(_0649_));
 sg13g2_inv_1 _5745_ (.Y(_0837_),
    .A(_0735_));
 sg13g2_a22oi_1 _5746_ (.Y(_0838_),
    .B1(_4164_),
    .B2(_0837_),
    .A2(_4201_),
    .A1(_4302_));
 sg13g2_nand2b_1 _5747_ (.Y(_0839_),
    .B(_0838_),
    .A_N(_0836_));
 sg13g2_inv_1 _5748_ (.Y(_0840_),
    .A(_0675_));
 sg13g2_o21ai_1 _5749_ (.B1(_0835_),
    .Y(_0841_),
    .A1(_0840_),
    .A2(_0833_));
 sg13g2_nand2b_1 _5750_ (.Y(_0842_),
    .B(_0647_),
    .A_N(_0841_));
 sg13g2_nor2_1 _5751_ (.A(_4255_),
    .B(_0643_),
    .Y(_0843_));
 sg13g2_inv_1 _5752_ (.Y(_0844_),
    .A(_0843_));
 sg13g2_a21oi_1 _5753_ (.A1(_0844_),
    .A2(_0649_),
    .Y(_0845_),
    .B1(_4258_));
 sg13g2_nor2_1 _5754_ (.A(_0799_),
    .B(_0841_),
    .Y(_0846_));
 sg13g2_o21ai_1 _5755_ (.B1(_0694_),
    .Y(_0847_),
    .A1(_4208_),
    .A2(_0846_));
 sg13g2_a221oi_1 _5756_ (.B2(_0845_),
    .C1(_0847_),
    .B1(_0842_),
    .A1(_4189_),
    .Y(_0848_),
    .A2(_0839_));
 sg13g2_a22oi_1 _5757_ (.Y(_0849_),
    .B1(_0832_),
    .B2(_0848_),
    .A2(net92),
    .A1(_0037_));
 sg13g2_nor2_1 _5758_ (.A(_0819_),
    .B(_4519_),
    .Y(_0850_));
 sg13g2_nor2_1 _5759_ (.A(_0814_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_nand2_1 _5760_ (.Y(_0852_),
    .A(_0851_),
    .B(_0783_));
 sg13g2_nand2_1 _5761_ (.Y(_0853_),
    .A(_0265_),
    .B(_0852_));
 sg13g2_nand2b_1 _5762_ (.Y(_0854_),
    .B(_0853_),
    .A_N(_0849_));
 sg13g2_nand3_1 _5763_ (.B(_0852_),
    .C(_0849_),
    .A(_0265_),
    .Y(_0855_));
 sg13g2_inv_1 _5764_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_a21oi_1 _5765_ (.A1(_0830_),
    .A2(_0854_),
    .Y(_0857_),
    .B1(_0856_));
 sg13g2_nand2_1 _5766_ (.Y(_0858_),
    .A(_0268_),
    .B(_0785_));
 sg13g2_nand3_1 _5767_ (.B(_0267_),
    .C(_0400_),
    .A(_0265_),
    .Y(_0859_));
 sg13g2_nand2_1 _5768_ (.Y(_0860_),
    .A(_0858_),
    .B(_0859_));
 sg13g2_nand3_1 _5769_ (.B(_0660_),
    .C(_0655_),
    .A(_0733_),
    .Y(_0861_));
 sg13g2_o21ai_1 _5770_ (.B1(_4204_),
    .Y(_0862_),
    .A1(_0799_),
    .A2(_0861_));
 sg13g2_a21oi_1 _5771_ (.A1(_0729_),
    .A2(net132),
    .Y(_0863_),
    .B1(_4258_));
 sg13g2_o21ai_1 _5772_ (.B1(_0863_),
    .Y(_0864_),
    .A1(net132),
    .A2(_0861_));
 sg13g2_nand2_1 _5773_ (.Y(_0865_),
    .A(_0862_),
    .B(_0864_));
 sg13g2_nor2_1 _5774_ (.A(_0865_),
    .B(_0810_),
    .Y(_0866_));
 sg13g2_a22oi_1 _5775_ (.Y(_0867_),
    .B1(_0694_),
    .B2(_0866_),
    .A2(net92),
    .A1(_0039_));
 sg13g2_nand2_1 _5776_ (.Y(_0868_),
    .A(_0860_),
    .B(_0867_));
 sg13g2_inv_1 _5777_ (.Y(_0869_),
    .A(_0867_));
 sg13g2_nand3_1 _5778_ (.B(_0859_),
    .C(_0869_),
    .A(_0858_),
    .Y(_0870_));
 sg13g2_nand2_1 _5779_ (.Y(_0871_),
    .A(_0868_),
    .B(_0870_));
 sg13g2_nor2_1 _5780_ (.A(_0857_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_a21oi_1 _5781_ (.A1(_0744_),
    .A2(_0655_),
    .Y(_0873_),
    .B1(net141));
 sg13g2_o21ai_1 _5782_ (.B1(_0647_),
    .Y(_0874_),
    .A1(_0676_),
    .A2(_0873_));
 sg13g2_a21oi_1 _5783_ (.A1(_0874_),
    .A2(_0838_),
    .Y(_0875_),
    .B1(_4217_));
 sg13g2_a21oi_1 _5784_ (.A1(_0650_),
    .A2(_0831_),
    .Y(_0876_),
    .B1(_4160_));
 sg13g2_nor2b_1 _5785_ (.A(_0873_),
    .B_N(_0677_),
    .Y(_0877_));
 sg13g2_nor2_1 _5786_ (.A(net132),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_nor3_1 _5787_ (.A(_0683_),
    .B(_0688_),
    .C(_0878_),
    .Y(_0879_));
 sg13g2_nor2_1 _5788_ (.A(_4157_),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_or3_1 _5789_ (.A(_0875_),
    .B(_0876_),
    .C(_0880_),
    .X(_0881_));
 sg13g2_inv_1 _5790_ (.Y(_0882_),
    .A(_0881_));
 sg13g2_a22oi_1 _5791_ (.Y(_0883_),
    .B1(_0694_),
    .B2(_0882_),
    .A2(net92),
    .A1(_0041_));
 sg13g2_nand2_1 _5792_ (.Y(_0884_),
    .A(_0786_),
    .B(_4522_));
 sg13g2_inv_2 _5793_ (.Y(_0885_),
    .A(_0776_));
 sg13g2_nand2_1 _5794_ (.Y(_0886_),
    .A(_0884_),
    .B(_0885_));
 sg13g2_nand2_1 _5795_ (.Y(_0887_),
    .A(_0886_),
    .B(_0388_));
 sg13g2_nand3_1 _5796_ (.B(_0773_),
    .C(_0885_),
    .A(_0884_),
    .Y(_0888_));
 sg13g2_nand2_1 _5797_ (.Y(_0889_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_xnor2_1 _5798_ (.Y(_0890_),
    .A(_0883_),
    .B(_0889_));
 sg13g2_nand2_1 _5799_ (.Y(_0891_),
    .A(_0872_),
    .B(_0890_));
 sg13g2_nand2_1 _5800_ (.Y(_0892_),
    .A(_0886_),
    .B(_0773_));
 sg13g2_nand3_1 _5801_ (.B(_0388_),
    .C(_0885_),
    .A(_0884_),
    .Y(_0893_));
 sg13g2_inv_1 _5802_ (.Y(_0894_),
    .A(_0883_));
 sg13g2_nand3_1 _5803_ (.B(_0893_),
    .C(_0894_),
    .A(_0892_),
    .Y(_0895_));
 sg13g2_inv_1 _5804_ (.Y(_0896_),
    .A(_0868_));
 sg13g2_nor2_1 _5805_ (.A(_0894_),
    .B(_0889_),
    .Y(_0897_));
 sg13g2_a21oi_1 _5806_ (.A1(_0895_),
    .A2(_0896_),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nand2_1 _5807_ (.Y(_0899_),
    .A(_0891_),
    .B(_0898_));
 sg13g2_nand2_1 _5808_ (.Y(_0900_),
    .A(_0796_),
    .B(_0899_));
 sg13g2_inv_1 _5809_ (.Y(_0901_),
    .A(_0755_));
 sg13g2_inv_1 _5810_ (.Y(_0902_),
    .A(_0794_));
 sg13g2_a21oi_1 _5811_ (.A1(_0901_),
    .A2(_0793_),
    .Y(_0903_),
    .B1(_0902_));
 sg13g2_nand2_1 _5812_ (.Y(_0904_),
    .A(_0900_),
    .B(_0903_));
 sg13g2_nand3_1 _5813_ (.B(_4168_),
    .C(_0660_),
    .A(_0729_),
    .Y(_0905_));
 sg13g2_a21o_1 _5814_ (.A2(_0905_),
    .A1(net140),
    .B1(_0805_),
    .X(_0906_));
 sg13g2_inv_1 _5815_ (.Y(_0907_),
    .A(_4258_));
 sg13g2_a21oi_1 _5816_ (.A1(_0744_),
    .A2(_0742_),
    .Y(_0908_),
    .B1(net141));
 sg13g2_a21oi_1 _5817_ (.A1(net141),
    .A2(_0843_),
    .Y(_0909_),
    .B1(_0908_));
 sg13g2_nor4_1 _5818_ (.A(net153),
    .B(net163),
    .C(net155),
    .D(_0672_),
    .Y(_0910_));
 sg13g2_a21oi_1 _5819_ (.A1(_0672_),
    .A2(_0689_),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_nand3_1 _5820_ (.B(net140),
    .C(_0675_),
    .A(_0911_),
    .Y(_0912_));
 sg13g2_o21ai_1 _5821_ (.B1(_0912_),
    .Y(_0913_),
    .A1(net140),
    .A2(_0909_));
 sg13g2_a22oi_1 _5822_ (.Y(_0914_),
    .B1(_0907_),
    .B2(_0913_),
    .A2(_4161_),
    .A1(_0906_));
 sg13g2_a21oi_1 _5823_ (.A1(_0911_),
    .A2(_0675_),
    .Y(_0915_),
    .B1(_0799_));
 sg13g2_nand2b_1 _5824_ (.Y(_0916_),
    .B(_4204_),
    .A_N(_0915_));
 sg13g2_o21ai_1 _5825_ (.B1(_0765_),
    .Y(_0917_),
    .A1(net132),
    .A2(_0911_));
 sg13g2_nand3_1 _5826_ (.B(_0916_),
    .C(_0917_),
    .A(_0914_),
    .Y(_0918_));
 sg13g2_inv_1 _5827_ (.Y(_0919_),
    .A(_0918_));
 sg13g2_a22oi_1 _5828_ (.Y(_0920_),
    .B1(_0694_),
    .B2(_0919_),
    .A2(net86),
    .A1(_0044_));
 sg13g2_nor2_1 _5829_ (.A(_0401_),
    .B(_0606_),
    .Y(_0921_));
 sg13g2_nand2_1 _5830_ (.Y(_0922_),
    .A(_0921_),
    .B(_0268_));
 sg13g2_nor2_1 _5831_ (.A(_0790_),
    .B(_0723_),
    .Y(_0923_));
 sg13g2_a21oi_1 _5832_ (.A1(_0923_),
    .A2(_0407_),
    .Y(_0924_),
    .B1(_0613_));
 sg13g2_nand2_1 _5833_ (.Y(_0925_),
    .A(_0922_),
    .B(_0924_));
 sg13g2_nand2_1 _5834_ (.Y(_0926_),
    .A(_0925_),
    .B(_0546_));
 sg13g2_inv_2 _5835_ (.Y(_0927_),
    .A(_0546_));
 sg13g2_nand3_1 _5836_ (.B(_0924_),
    .C(_0927_),
    .A(_0922_),
    .Y(_0928_));
 sg13g2_nand3b_1 _5837_ (.B(_0926_),
    .C(_0928_),
    .Y(_0929_),
    .A_N(_0920_));
 sg13g2_nand2_1 _5838_ (.Y(_0930_),
    .A(_0925_),
    .B(_0927_));
 sg13g2_nand3_1 _5839_ (.B(_0924_),
    .C(_0546_),
    .A(_0922_),
    .Y(_0931_));
 sg13g2_nand3_1 _5840_ (.B(_0931_),
    .C(_0920_),
    .A(_0930_),
    .Y(_0932_));
 sg13g2_nand2_1 _5841_ (.Y(_0933_),
    .A(_0929_),
    .B(_0932_));
 sg13g2_a21oi_1 _5842_ (.A1(net155),
    .A2(_0664_),
    .Y(_0934_),
    .B1(_0735_));
 sg13g2_a21oi_1 _5843_ (.A1(_0934_),
    .A2(net139),
    .Y(_0935_),
    .B1(_0740_));
 sg13g2_nor2b_1 _5844_ (.A(_4255_),
    .B_N(_4164_),
    .Y(_0936_));
 sg13g2_inv_1 _5845_ (.Y(_0937_),
    .A(_0671_));
 sg13g2_a22oi_1 _5846_ (.Y(_0938_),
    .B1(_0936_),
    .B2(_0937_),
    .A2(_0728_),
    .A1(_4201_));
 sg13g2_o21ai_1 _5847_ (.B1(_0938_),
    .Y(_0939_),
    .A1(net132),
    .A2(_0935_));
 sg13g2_nand2_1 _5848_ (.Y(_0940_),
    .A(_0939_),
    .B(_0907_));
 sg13g2_nand2_1 _5849_ (.Y(_0941_),
    .A(_0935_),
    .B(_0800_));
 sg13g2_nand3_1 _5850_ (.B(_0660_),
    .C(_0655_),
    .A(_0653_),
    .Y(_0942_));
 sg13g2_a21o_1 _5851_ (.A2(_0942_),
    .A1(_0667_),
    .B1(_0805_),
    .X(_0943_));
 sg13g2_nor2_1 _5852_ (.A(_4155_),
    .B(_0934_),
    .Y(_0944_));
 sg13g2_o21ai_1 _5853_ (.B1(_0694_),
    .Y(_0945_),
    .A1(_0809_),
    .A2(_0944_));
 sg13g2_a221oi_1 _5854_ (.B2(_0943_),
    .C1(_0945_),
    .B1(_4161_),
    .A1(_0941_),
    .Y(_0946_),
    .A2(_4204_));
 sg13g2_a22oi_1 _5855_ (.Y(_0947_),
    .B1(_0940_),
    .B2(_0946_),
    .A2(net86),
    .A1(_0045_));
 sg13g2_a21oi_1 _5856_ (.A1(_0818_),
    .A2(_4518_),
    .Y(_0948_),
    .B1(_0814_));
 sg13g2_nand2b_1 _5857_ (.Y(_0949_),
    .B(_0786_),
    .A_N(_0948_));
 sg13g2_nand2_1 _5858_ (.Y(_0950_),
    .A(_0949_),
    .B(_0885_));
 sg13g2_nand2_1 _5859_ (.Y(_0951_),
    .A(_0605_),
    .B(_0927_));
 sg13g2_inv_1 _5860_ (.Y(_0952_),
    .A(_0774_));
 sg13g2_nor2_1 _5861_ (.A(_0951_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_nor2_1 _5862_ (.A(_0546_),
    .B(_0790_),
    .Y(_0954_));
 sg13g2_nand2_1 _5863_ (.Y(_0955_),
    .A(_0780_),
    .B(_0954_));
 sg13g2_nand2_1 _5864_ (.Y(_0956_),
    .A(_0612_),
    .B(_0545_));
 sg13g2_nand2_1 _5865_ (.Y(_0957_),
    .A(_0956_),
    .B(_0544_));
 sg13g2_nand2_1 _5866_ (.Y(_0958_),
    .A(_0955_),
    .B(_0957_));
 sg13g2_a21oi_1 _5867_ (.A1(_0950_),
    .A2(_0953_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nand2b_1 _5868_ (.Y(_0960_),
    .B(_0815_),
    .A_N(_0823_));
 sg13g2_nor3_1 _5869_ (.A(_0960_),
    .B(_0783_),
    .C(_0785_),
    .Y(_0961_));
 sg13g2_nand3_1 _5870_ (.B(_4517_),
    .C(_0961_),
    .A(_0953_),
    .Y(_0962_));
 sg13g2_nand2_1 _5871_ (.Y(_0963_),
    .A(_0959_),
    .B(_0962_));
 sg13g2_nand2_1 _5872_ (.Y(_0964_),
    .A(_0963_),
    .B(_0571_));
 sg13g2_inv_1 _5873_ (.Y(_0965_),
    .A(_0571_));
 sg13g2_nand3_1 _5874_ (.B(_0965_),
    .C(_0962_),
    .A(_0959_),
    .Y(_0966_));
 sg13g2_nand3b_1 _5875_ (.B(_0964_),
    .C(_0966_),
    .Y(_0967_),
    .A_N(_0947_));
 sg13g2_nand2_1 _5876_ (.Y(_0968_),
    .A(_0963_),
    .B(_0965_));
 sg13g2_nand3_1 _5877_ (.B(_0571_),
    .C(_0962_),
    .A(_0959_),
    .Y(_0969_));
 sg13g2_nand3_1 _5878_ (.B(_0969_),
    .C(_0947_),
    .A(_0968_),
    .Y(_0970_));
 sg13g2_buf_1 _5879_ (.A(_0970_),
    .X(_0971_));
 sg13g2_nand2_1 _5880_ (.Y(_0972_),
    .A(_0967_),
    .B(_0971_));
 sg13g2_nor2_1 _5881_ (.A(_0933_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_nand2_1 _5882_ (.Y(_0974_),
    .A(_0904_),
    .B(_0973_));
 sg13g2_nand2_1 _5883_ (.Y(_0975_),
    .A(_0971_),
    .B(_0932_));
 sg13g2_nand2_1 _5884_ (.Y(_0976_),
    .A(_0975_),
    .B(_0967_));
 sg13g2_nand2_1 _5885_ (.Y(_0977_),
    .A(_0974_),
    .B(_0976_));
 sg13g2_nand2b_1 _5886_ (.Y(_0978_),
    .B(_0977_),
    .A_N(_0722_));
 sg13g2_nand3_1 _5887_ (.B(_0722_),
    .C(_0976_),
    .A(_0974_),
    .Y(_0979_));
 sg13g2_nand2_1 _5888_ (.Y(_0980_),
    .A(_0707_),
    .B(_4236_));
 sg13g2_inv_1 _5889_ (.Y(_0981_),
    .A(\i_display.i_vga.timing_ver.counter[8] ));
 sg13g2_nor2_2 _5890_ (.A(net150),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_nor2_1 _5891_ (.A(_0982_),
    .B(net85),
    .Y(_0983_));
 sg13g2_a21oi_1 _5892_ (.A1(net85),
    .A2(_0980_),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_xor2_1 _5893_ (.B(_0972_),
    .A(_0984_),
    .X(_0985_));
 sg13g2_nand2_1 _5894_ (.Y(_0986_),
    .A(_0830_),
    .B(_0854_));
 sg13g2_nand2_1 _5895_ (.Y(_0987_),
    .A(_0986_),
    .B(_0855_));
 sg13g2_nand2_1 _5896_ (.Y(_0988_),
    .A(_0987_),
    .B(_0870_));
 sg13g2_nand2_1 _5897_ (.Y(_0989_),
    .A(_0988_),
    .B(_0868_));
 sg13g2_nand2_1 _5898_ (.Y(_0990_),
    .A(_0989_),
    .B(_0890_));
 sg13g2_nor2_1 _5899_ (.A(_0897_),
    .B(_0901_),
    .Y(_0991_));
 sg13g2_nand2_1 _5900_ (.Y(_0992_),
    .A(_0990_),
    .B(_0991_));
 sg13g2_nor2_1 _5901_ (.A(_0795_),
    .B(_0933_),
    .Y(_0993_));
 sg13g2_nand3_1 _5902_ (.B(_0993_),
    .C(_0752_),
    .A(_0992_),
    .Y(_0994_));
 sg13g2_inv_1 _5903_ (.Y(_0995_),
    .A(_0929_));
 sg13g2_a21oi_1 _5904_ (.A1(_0932_),
    .A2(_0794_),
    .Y(_0996_),
    .B1(_0995_));
 sg13g2_inv_1 _5905_ (.Y(_0997_),
    .A(_0996_));
 sg13g2_nand2_1 _5906_ (.Y(_0998_),
    .A(_0994_),
    .B(_0997_));
 sg13g2_xnor2_1 _5907_ (.Y(_0999_),
    .A(_0985_),
    .B(_0998_));
 sg13g2_a21oi_1 _5908_ (.A1(_0978_),
    .A2(_0979_),
    .Y(_1000_),
    .B1(_0999_));
 sg13g2_inv_1 _5909_ (.Y(_1001_),
    .A(\i_display.i_vga.low_count[7] ));
 sg13g2_nor2_1 _5910_ (.A(_1001_),
    .B(net131),
    .Y(_1002_));
 sg13g2_buf_1 _5911_ (.A(\i_display.i_vga.timing_ver.counter[7] ),
    .X(_1003_));
 sg13g2_inv_1 _5912_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_nor2_1 _5913_ (.A(net150),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_nor2b_1 _5914_ (.A(net85),
    .B_N(_1005_),
    .Y(_1006_));
 sg13g2_a21oi_1 _5915_ (.A1(net85),
    .A2(_1002_),
    .Y(_1007_),
    .B1(_1006_));
 sg13g2_xnor2_1 _5916_ (.Y(_1008_),
    .A(_1007_),
    .B(_0933_));
 sg13g2_xnor2_1 _5917_ (.Y(_1009_),
    .A(_1008_),
    .B(_0904_));
 sg13g2_inv_1 _5918_ (.Y(_1010_),
    .A(_4238_));
 sg13g2_nor2_2 _5919_ (.A(_1010_),
    .B(_0708_),
    .Y(_1011_));
 sg13g2_inv_1 _5920_ (.Y(_1012_),
    .A(_1011_));
 sg13g2_buf_2 _5921_ (.A(\i_display.i_vga.timing_ver.counter[4] ),
    .X(_1013_));
 sg13g2_inv_1 _5922_ (.Y(_1014_),
    .A(_1013_));
 sg13g2_nor2_1 _5923_ (.A(net150),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_nor2_1 _5924_ (.A(_1015_),
    .B(_0705_),
    .Y(_1016_));
 sg13g2_a21oi_1 _5925_ (.A1(net85),
    .A2(_1012_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_xnor2_1 _5926_ (.Y(_1018_),
    .A(_0890_),
    .B(_0989_));
 sg13g2_nor2_1 _5927_ (.A(_1017_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_inv_1 _5928_ (.Y(_1020_),
    .A(\i_display.i_vga.low_count[5] ));
 sg13g2_nor2_1 _5929_ (.A(_1020_),
    .B(_0708_),
    .Y(_1021_));
 sg13g2_inv_1 _5930_ (.Y(_1022_),
    .A(_1021_));
 sg13g2_buf_1 _5931_ (.A(\i_display.i_vga.timing_ver.counter[5] ),
    .X(_1023_));
 sg13g2_inv_1 _5932_ (.Y(_1024_),
    .A(_1023_));
 sg13g2_nor2_2 _5933_ (.A(_0706_),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_nor2_1 _5934_ (.A(_1025_),
    .B(_0704_),
    .Y(_1026_));
 sg13g2_a21o_1 _5935_ (.A2(_1022_),
    .A1(net91),
    .B1(_1026_),
    .X(_1027_));
 sg13g2_nand2_1 _5936_ (.Y(_1028_),
    .A(_0756_),
    .B(_1027_));
 sg13g2_inv_1 _5937_ (.Y(_1029_),
    .A(_1027_));
 sg13g2_nand3_1 _5938_ (.B(_0755_),
    .C(_1029_),
    .A(_0752_),
    .Y(_1030_));
 sg13g2_nand2_1 _5939_ (.Y(_1031_),
    .A(_1028_),
    .B(_1030_));
 sg13g2_a22oi_1 _5940_ (.Y(_1032_),
    .B1(_0899_),
    .B2(_1031_),
    .A2(_1017_),
    .A1(_1018_));
 sg13g2_nand2b_1 _5941_ (.Y(_1033_),
    .B(_1032_),
    .A_N(_1019_));
 sg13g2_nand2_1 _5942_ (.Y(_1034_),
    .A(_0895_),
    .B(_0896_));
 sg13g2_inv_1 _5943_ (.Y(_1035_),
    .A(_0897_));
 sg13g2_nand2_1 _5944_ (.Y(_1036_),
    .A(_1034_),
    .B(_1035_));
 sg13g2_a21oi_1 _5945_ (.A1(_0872_),
    .A2(_0890_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_nor2b_1 _5946_ (.A(_1031_),
    .B_N(_1037_),
    .Y(_1038_));
 sg13g2_nor2_2 _5947_ (.A(_4231_),
    .B(_0708_),
    .Y(_1039_));
 sg13g2_inv_1 _5948_ (.Y(_1040_),
    .A(_1039_));
 sg13g2_buf_1 _5949_ (.A(\i_display.i_vga.timing_ver.counter[2] ),
    .X(_1041_));
 sg13g2_inv_1 _5950_ (.Y(_1042_),
    .A(_1041_));
 sg13g2_nor2_2 _5951_ (.A(_0711_),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_nor2_1 _5952_ (.A(_1043_),
    .B(net91),
    .Y(_1044_));
 sg13g2_a21oi_1 _5953_ (.A1(net91),
    .A2(_1040_),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_nand2_1 _5954_ (.Y(_1046_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_xnor2_1 _5955_ (.Y(_1047_),
    .A(_0829_),
    .B(_1046_));
 sg13g2_nor2_1 _5956_ (.A(_1045_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_nand2_1 _5957_ (.Y(_1049_),
    .A(_1047_),
    .B(_1045_));
 sg13g2_inv_1 _5958_ (.Y(_1050_),
    .A(_4232_));
 sg13g2_nor2_2 _5959_ (.A(_1050_),
    .B(_0708_),
    .Y(_1051_));
 sg13g2_inv_1 _5960_ (.Y(_1052_),
    .A(_1051_));
 sg13g2_buf_1 _5961_ (.A(\i_display.i_vga.timing_ver.counter[0] ),
    .X(_1053_));
 sg13g2_inv_1 _5962_ (.Y(_1054_),
    .A(_1053_));
 sg13g2_nor2_2 _5963_ (.A(net150),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_nor2_1 _5964_ (.A(_1055_),
    .B(net91),
    .Y(_1056_));
 sg13g2_a21oi_1 _5965_ (.A1(net91),
    .A2(_1052_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_xnor2_1 _5966_ (.Y(_1058_),
    .A(_0825_),
    .B(_0824_));
 sg13g2_xor2_1 _5967_ (.B(_1058_),
    .A(_1057_),
    .X(_1059_));
 sg13g2_nand2_1 _5968_ (.Y(_1060_),
    .A(_0822_),
    .B(_0827_));
 sg13g2_inv_1 _5969_ (.Y(_1061_),
    .A(_0826_));
 sg13g2_nand2_1 _5970_ (.Y(_1062_),
    .A(_1060_),
    .B(_1061_));
 sg13g2_nand3_1 _5971_ (.B(_0827_),
    .C(_0826_),
    .A(_0822_),
    .Y(_1063_));
 sg13g2_nand2_1 _5972_ (.Y(_1064_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_nand2_1 _5973_ (.Y(_1065_),
    .A(_0707_),
    .B(_4233_));
 sg13g2_inv_1 _5974_ (.Y(_1066_),
    .A(_1065_));
 sg13g2_buf_1 _5975_ (.A(\i_display.i_vga.timing_ver.counter[1] ),
    .X(_1067_));
 sg13g2_inv_1 _5976_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_nor2_2 _5977_ (.A(net150),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_inv_1 _5978_ (.Y(_1070_),
    .A(_1069_));
 sg13g2_nor2_1 _5979_ (.A(_1070_),
    .B(net102),
    .Y(_1071_));
 sg13g2_a21o_1 _5980_ (.A2(_1066_),
    .A1(net102),
    .B1(_1071_),
    .X(_1072_));
 sg13g2_nand2_1 _5981_ (.Y(_1073_),
    .A(_1064_),
    .B(_1072_));
 sg13g2_inv_1 _5982_ (.Y(_1074_),
    .A(_1072_));
 sg13g2_nand3_1 _5983_ (.B(_1063_),
    .C(_1074_),
    .A(_1062_),
    .Y(_1075_));
 sg13g2_nand2_1 _5984_ (.Y(_1076_),
    .A(_1073_),
    .B(_1075_));
 sg13g2_nor2_1 _5985_ (.A(_1059_),
    .B(_1076_),
    .Y(_1077_));
 sg13g2_nand2_1 _5986_ (.Y(_1078_),
    .A(_1049_),
    .B(_1077_));
 sg13g2_nor2_1 _5987_ (.A(_1048_),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_inv_1 _5988_ (.Y(_1080_),
    .A(_4239_));
 sg13g2_nor2_1 _5989_ (.A(_1080_),
    .B(_0708_),
    .Y(_1081_));
 sg13g2_inv_1 _5990_ (.Y(_1082_),
    .A(_1081_));
 sg13g2_buf_1 _5991_ (.A(\i_display.i_vga.timing_ver.counter[3] ),
    .X(_1083_));
 sg13g2_inv_1 _5992_ (.Y(_1084_),
    .A(_1083_));
 sg13g2_nor2_2 _5993_ (.A(_0711_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nor2_1 _5994_ (.A(_1085_),
    .B(net91),
    .Y(_1086_));
 sg13g2_a21oi_1 _5995_ (.A1(net91),
    .A2(_1082_),
    .Y(_1087_),
    .B1(_1086_));
 sg13g2_nand2b_1 _5996_ (.Y(_1088_),
    .B(_0871_),
    .A_N(_1087_));
 sg13g2_nand3_1 _5997_ (.B(_0870_),
    .C(_1087_),
    .A(_0868_),
    .Y(_1089_));
 sg13g2_nand3_1 _5998_ (.B(_1089_),
    .C(_0857_),
    .A(_1088_),
    .Y(_1090_));
 sg13g2_nand2_1 _5999_ (.Y(_1091_),
    .A(_1088_),
    .B(_1089_));
 sg13g2_nand2_1 _6000_ (.Y(_1092_),
    .A(_1091_),
    .B(_0987_));
 sg13g2_nand3_1 _6001_ (.B(_1090_),
    .C(_1092_),
    .A(_1079_),
    .Y(_1093_));
 sg13g2_nor2_1 _6002_ (.A(_1038_),
    .B(_1093_),
    .Y(_1094_));
 sg13g2_inv_1 _6003_ (.Y(_1095_),
    .A(_4225_));
 sg13g2_nor2_1 _6004_ (.A(_1095_),
    .B(_0708_),
    .Y(_1096_));
 sg13g2_inv_1 _6005_ (.Y(_1097_),
    .A(_1096_));
 sg13g2_inv_1 _6006_ (.Y(_1098_),
    .A(\i_display.i_vga.timing_ver.counter[6] ));
 sg13g2_nor2_2 _6007_ (.A(_0706_),
    .B(_1098_),
    .Y(_1099_));
 sg13g2_nor2_1 _6008_ (.A(_1099_),
    .B(_0705_),
    .Y(_1100_));
 sg13g2_a21oi_1 _6009_ (.A1(net85),
    .A2(_1097_),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_xor2_1 _6010_ (.B(_0795_),
    .A(_1101_),
    .X(_1102_));
 sg13g2_inv_2 _6011_ (.Y(_1103_),
    .A(_1102_));
 sg13g2_nand2_1 _6012_ (.Y(_1104_),
    .A(_0992_),
    .B(_0752_));
 sg13g2_nand2_1 _6013_ (.Y(_1105_),
    .A(_1103_),
    .B(_1104_));
 sg13g2_inv_1 _6014_ (.Y(_1106_),
    .A(_1104_));
 sg13g2_nand2_1 _6015_ (.Y(_1107_),
    .A(_1106_),
    .B(_1102_));
 sg13g2_nand3_1 _6016_ (.B(_1105_),
    .C(_1107_),
    .A(_1094_),
    .Y(_1108_));
 sg13g2_nor3_1 _6017_ (.A(_1009_),
    .B(_1033_),
    .C(_1108_),
    .Y(_1109_));
 sg13g2_nand2_1 _6018_ (.Y(_1110_),
    .A(_0703_),
    .B(_0971_));
 sg13g2_a21oi_1 _6019_ (.A1(_1110_),
    .A2(_0700_),
    .Y(_1111_),
    .B1(_0996_));
 sg13g2_nand2_1 _6020_ (.Y(_1112_),
    .A(_1111_),
    .B(_0994_));
 sg13g2_nand2_1 _6021_ (.Y(_1113_),
    .A(_0700_),
    .B(_0703_));
 sg13g2_nand2_1 _6022_ (.Y(_1114_),
    .A(_1110_),
    .B(_0700_));
 sg13g2_o21ai_1 _6023_ (.B1(_1114_),
    .Y(_1115_),
    .A1(_1113_),
    .A2(_0972_));
 sg13g2_nand2_1 _6024_ (.Y(_1116_),
    .A(_1112_),
    .B(_1115_));
 sg13g2_nor2_1 _6025_ (.A(_0637_),
    .B(_0568_),
    .Y(_1117_));
 sg13g2_nor3_1 _6026_ (.A(_0571_),
    .B(_0637_),
    .C(_0957_),
    .Y(_1118_));
 sg13g2_nor3_1 _6027_ (.A(_0571_),
    .B(_0637_),
    .C(_0951_),
    .Y(_1119_));
 sg13g2_nor2b_1 _6028_ (.A(_0781_),
    .B_N(_1119_),
    .Y(_1120_));
 sg13g2_nor4_1 _6029_ (.A(_0633_),
    .B(_1117_),
    .C(_1118_),
    .D(_1120_),
    .Y(_1121_));
 sg13g2_nand4_1 _6030_ (.B(_4522_),
    .C(_0774_),
    .A(_1119_),
    .Y(_1122_),
    .D(_0786_));
 sg13g2_nor2b_1 _6031_ (.A(_0626_),
    .B_N(_0625_),
    .Y(_1123_));
 sg13g2_nor2_1 _6032_ (.A(_0619_),
    .B(_0624_),
    .Y(_1124_));
 sg13g2_nand2_1 _6033_ (.Y(_1125_),
    .A(_4585_),
    .B(_0306_));
 sg13g2_nor2_1 _6034_ (.A(_0436_),
    .B(_0415_),
    .Y(_1126_));
 sg13g2_xnor2_1 _6035_ (.Y(_1127_),
    .A(_1125_),
    .B(_1126_));
 sg13g2_nor2b_1 _6036_ (.A(_0622_),
    .B_N(_0621_),
    .Y(_1128_));
 sg13g2_a21oi_1 _6037_ (.A1(_0623_),
    .A2(_0620_),
    .Y(_1129_),
    .B1(_1128_));
 sg13g2_xnor2_1 _6038_ (.Y(_1130_),
    .A(_1127_),
    .B(_1129_));
 sg13g2_xnor2_1 _6039_ (.Y(_1131_),
    .A(_1124_),
    .B(_1130_));
 sg13g2_xor2_1 _6040_ (.B(_1131_),
    .A(_1123_),
    .X(_1132_));
 sg13g2_inv_1 _6041_ (.Y(_1133_),
    .A(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[9] ));
 sg13g2_nor4_1 _6042_ (.A(net162),
    .B(_0799_),
    .C(_4151_),
    .D(_0030_),
    .Y(_1134_));
 sg13g2_nand3_1 _6043_ (.B(_0666_),
    .C(_1134_),
    .A(net102),
    .Y(_1135_));
 sg13g2_o21ai_1 _6044_ (.B1(_1135_),
    .Y(_1136_),
    .A1(_1133_),
    .A2(_0704_));
 sg13g2_nor2_1 _6045_ (.A(_0627_),
    .B(_0630_),
    .Y(_1137_));
 sg13g2_xnor2_1 _6046_ (.Y(_1138_),
    .A(_1136_),
    .B(_1137_));
 sg13g2_xnor2_1 _6047_ (.Y(_1139_),
    .A(_1132_),
    .B(_1138_));
 sg13g2_a21oi_1 _6048_ (.A1(_1121_),
    .A2(_1122_),
    .Y(_1140_),
    .B1(_1139_));
 sg13g2_nand3_1 _6049_ (.B(_1122_),
    .C(_1139_),
    .A(_1121_),
    .Y(_1141_));
 sg13g2_nor2b_1 _6050_ (.A(_1140_),
    .B_N(_1141_),
    .Y(_1142_));
 sg13g2_inv_1 _6051_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_nand2_1 _6052_ (.Y(_1144_),
    .A(_1116_),
    .B(_1143_));
 sg13g2_nand3_1 _6053_ (.B(_1115_),
    .C(_1142_),
    .A(_1112_),
    .Y(_1145_));
 sg13g2_nand2_1 _6054_ (.Y(_1146_),
    .A(_1144_),
    .B(_1145_));
 sg13g2_nand3_1 _6055_ (.B(_1109_),
    .C(_1146_),
    .A(_1000_),
    .Y(_1147_));
 sg13g2_nand2_1 _6056_ (.Y(_1148_),
    .A(_1023_),
    .B(\i_display.i_vga.timing_ver.counter[6] ));
 sg13g2_nor3_1 _6057_ (.A(_1013_),
    .B(_1004_),
    .C(_1148_),
    .Y(_1149_));
 sg13g2_inv_1 _6058_ (.Y(_1150_),
    .A(\i_display.i_vga.timing_ver.counter[10] ));
 sg13g2_nor3_2 _6059_ (.A(_0712_),
    .B(_0981_),
    .C(_1150_),
    .Y(_1151_));
 sg13g2_nor2_1 _6060_ (.A(_1067_),
    .B(_1054_),
    .Y(_1152_));
 sg13g2_nor2_1 _6061_ (.A(_1041_),
    .B(_1084_),
    .Y(_1153_));
 sg13g2_nand4_1 _6062_ (.B(_1151_),
    .C(_1152_),
    .A(_1149_),
    .Y(_1154_),
    .D(_1153_));
 sg13g2_inv_1 _6063_ (.Y(_1155_),
    .A(_4237_));
 sg13g2_inv_1 _6064_ (.Y(_1156_),
    .A(_4233_));
 sg13g2_buf_1 _6065_ (.A(_1156_),
    .X(_1157_));
 sg13g2_buf_1 _6066_ (.A(net138),
    .X(_1158_));
 sg13g2_nor4_1 _6067_ (.A(_1155_),
    .B(_1050_),
    .C(_4231_),
    .D(_1158_),
    .Y(_1159_));
 sg13g2_inv_1 _6068_ (.Y(_1160_),
    .A(_4236_));
 sg13g2_nor4_1 _6069_ (.A(\i_display.i_vga.low_count[7] ),
    .B(_4225_),
    .C(_1160_),
    .D(\i_display.i_vga.low_count[5] ),
    .Y(_1161_));
 sg13g2_nand3_1 _6070_ (.B(_4241_),
    .C(_1161_),
    .A(_1159_),
    .Y(_1162_));
 sg13g2_buf_1 _6071_ (.A(_1162_),
    .X(_1163_));
 sg13g2_mux2_1 _6072_ (.A0(_1154_),
    .A1(\i_display.hsync ),
    .S(_1163_),
    .X(_1164_));
 sg13g2_nand2_1 _6073_ (.Y(_1165_),
    .A(_1147_),
    .B(_1164_));
 sg13g2_nand2_1 _6074_ (.Y(_1166_),
    .A(_1165_),
    .B(_0640_));
 sg13g2_buf_1 _6075_ (.A(_1166_),
    .X(_1167_));
 sg13g2_nand2_1 _6076_ (.Y(_1168_),
    .A(net27),
    .B(_0032_));
 sg13g2_nand2_1 _6077_ (.Y(_1169_),
    .A(_1149_),
    .B(_1153_));
 sg13g2_nand2_1 _6078_ (.Y(_1170_),
    .A(_1151_),
    .B(_1152_));
 sg13g2_inv_1 _6079_ (.Y(_1171_),
    .A(_4243_));
 sg13g2_nor3_1 _6080_ (.A(_1169_),
    .B(_1170_),
    .C(_1171_),
    .Y(_1172_));
 sg13g2_inv_1 _6081_ (.Y(_1173_),
    .A(_1172_));
 sg13g2_xnor2_1 _6082_ (.Y(_1174_),
    .A(net141),
    .B(_4210_));
 sg13g2_xnor2_1 _6083_ (.Y(_1175_),
    .A(net8),
    .B(\crotchet[6] ));
 sg13g2_buf_2 _6084_ (.A(_1175_),
    .X(_1176_));
 sg13g2_xnor2_1 _6085_ (.Y(_1177_),
    .A(net6),
    .B(\crotchet[4] ));
 sg13g2_buf_1 _6086_ (.A(_1177_),
    .X(_1178_));
 sg13g2_xnor2_1 _6087_ (.Y(_1179_),
    .A(net7),
    .B(\crotchet[5] ));
 sg13g2_buf_1 _6088_ (.A(_1179_),
    .X(_1180_));
 sg13g2_inv_1 _6089_ (.Y(_1181_),
    .A(net148));
 sg13g2_nor3_1 _6090_ (.A(_1176_),
    .B(net149),
    .C(_1181_),
    .Y(_1182_));
 sg13g2_nor2_1 _6091_ (.A(net148),
    .B(net149),
    .Y(_1183_));
 sg13g2_inv_1 _6092_ (.Y(_1184_),
    .A(_1183_));
 sg13g2_buf_1 _6093_ (.A(\crotchet[0] ),
    .X(_1185_));
 sg13g2_buf_1 _6094_ (.A(\crotchet[1] ),
    .X(_1186_));
 sg13g2_xnor2_1 _6095_ (.Y(_1187_),
    .A(net3),
    .B(_1186_));
 sg13g2_inv_1 _6096_ (.Y(_1188_),
    .A(_1187_));
 sg13g2_nor2_1 _6097_ (.A(_1185_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_inv_1 _6098_ (.Y(_1190_),
    .A(_1189_));
 sg13g2_buf_1 _6099_ (.A(\crotchet[3] ),
    .X(_1191_));
 sg13g2_xnor2_1 _6100_ (.Y(_1192_),
    .A(net5),
    .B(_1191_));
 sg13g2_buf_1 _6101_ (.A(_1192_),
    .X(_1193_));
 sg13g2_inv_1 _6102_ (.Y(_1194_),
    .A(net137));
 sg13g2_buf_1 _6103_ (.A(\crotchet[2] ),
    .X(_1195_));
 sg13g2_xnor2_1 _6104_ (.Y(_1196_),
    .A(net4),
    .B(_1195_));
 sg13g2_buf_2 _6105_ (.A(_1196_),
    .X(_1197_));
 sg13g2_inv_2 _6106_ (.Y(_1198_),
    .A(_1197_));
 sg13g2_nor2_1 _6107_ (.A(_1194_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_inv_1 _6108_ (.Y(_1200_),
    .A(_1199_));
 sg13g2_nor2_1 _6109_ (.A(_1190_),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_inv_2 _6110_ (.Y(_1202_),
    .A(_1176_));
 sg13g2_xor2_1 _6111_ (.B(net149),
    .A(net148),
    .X(_1203_));
 sg13g2_nor2_1 _6112_ (.A(_1202_),
    .B(_1203_),
    .Y(_1204_));
 sg13g2_inv_1 _6113_ (.Y(_1205_),
    .A(_1204_));
 sg13g2_a21oi_1 _6114_ (.A1(_1184_),
    .A2(_1201_),
    .Y(_1206_),
    .B1(_1205_));
 sg13g2_nor2_1 _6115_ (.A(net137),
    .B(_1198_),
    .Y(_1207_));
 sg13g2_inv_1 _6116_ (.Y(_1208_),
    .A(_1207_));
 sg13g2_o21ai_1 _6117_ (.B1(_1208_),
    .Y(_1209_),
    .A1(_1182_),
    .A2(_1206_));
 sg13g2_nor2_1 _6118_ (.A(net137),
    .B(net149),
    .Y(_1210_));
 sg13g2_a21oi_1 _6119_ (.A1(_1210_),
    .A2(_1198_),
    .Y(_1211_),
    .B1(net148));
 sg13g2_inv_1 _6120_ (.Y(_1212_),
    .A(_1211_));
 sg13g2_nand2_1 _6121_ (.Y(_1213_),
    .A(net137),
    .B(net149));
 sg13g2_nor2b_1 _6122_ (.A(_1212_),
    .B_N(_1213_),
    .Y(_1214_));
 sg13g2_nor2_1 _6123_ (.A(_1197_),
    .B(_1194_),
    .Y(_1215_));
 sg13g2_nor2_1 _6124_ (.A(_1181_),
    .B(_1210_),
    .Y(_1216_));
 sg13g2_o21ai_1 _6125_ (.B1(_1216_),
    .Y(_1217_),
    .A1(_1207_),
    .A2(_1215_));
 sg13g2_nand2b_1 _6126_ (.Y(_1218_),
    .B(_1217_),
    .A_N(_1214_));
 sg13g2_a21oi_1 _6127_ (.A1(_1218_),
    .A2(_1202_),
    .Y(_1219_),
    .B1(_1173_));
 sg13g2_a22oi_1 _6128_ (.Y(_1220_),
    .B1(_1209_),
    .B2(_1219_),
    .A2(_1174_),
    .A1(_1173_));
 sg13g2_nand3_1 _6129_ (.B(net86),
    .C(_1220_),
    .A(_1165_),
    .Y(_1221_));
 sg13g2_nand2_1 _6130_ (.Y(_1222_),
    .A(_1168_),
    .B(_1221_));
 sg13g2_buf_2 _6131_ (.A(_1222_),
    .X(_1223_));
 sg13g2_nor2_1 _6132_ (.A(_4141_),
    .B(_1223_),
    .Y(_1224_));
 sg13g2_buf_1 _6133_ (.A(_1224_),
    .X(_1225_));
 sg13g2_inv_4 _6134_ (.A(net23),
    .Y(_1226_));
 sg13g2_nand4_1 _6135_ (.B(_1109_),
    .C(_1146_),
    .A(_1000_),
    .Y(_1227_),
    .D(net86));
 sg13g2_inv_1 _6136_ (.Y(_1228_),
    .A(_1152_));
 sg13g2_inv_1 _6137_ (.Y(_1229_),
    .A(_1148_));
 sg13g2_nand3_1 _6138_ (.B(_1003_),
    .C(_1229_),
    .A(_1151_),
    .Y(_1230_));
 sg13g2_nor3_1 _6139_ (.A(_1041_),
    .B(_1013_),
    .C(_1084_),
    .Y(_1231_));
 sg13g2_nand2b_1 _6140_ (.Y(_1232_),
    .B(_1231_),
    .A_N(_1230_));
 sg13g2_nand2_1 _6141_ (.Y(_1233_),
    .A(_4236_),
    .B(_4237_));
 sg13g2_nand2_1 _6142_ (.Y(_1234_),
    .A(_4235_),
    .B(_4239_));
 sg13g2_nor2_1 _6143_ (.A(_1010_),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_inv_1 _6144_ (.Y(_1236_),
    .A(_1235_));
 sg13g2_nor3_1 _6145_ (.A(_4229_),
    .B(_1233_),
    .C(_1236_),
    .Y(_1237_));
 sg13g2_inv_1 _6146_ (.Y(_1238_),
    .A(_1237_));
 sg13g2_nor3_1 _6147_ (.A(_1228_),
    .B(_1232_),
    .C(_1238_),
    .Y(_1239_));
 sg13g2_inv_1 _6148_ (.Y(_1240_),
    .A(_1239_));
 sg13g2_nand2_1 _6149_ (.Y(_1241_),
    .A(_1227_),
    .B(net90));
 sg13g2_buf_8 _6150_ (.A(_1241_),
    .X(_1242_));
 sg13g2_inv_1 _6151_ (.Y(_1243_),
    .A(_0670_));
 sg13g2_o21ai_1 _6152_ (.B1(_1206_),
    .Y(_1244_),
    .A1(net137),
    .A2(_1188_));
 sg13g2_nand2b_1 _6153_ (.Y(_1245_),
    .B(_1181_),
    .A_N(_1214_));
 sg13g2_nand2_1 _6154_ (.Y(_1246_),
    .A(_1197_),
    .B(net149));
 sg13g2_nor2_1 _6155_ (.A(_1194_),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_nor2_1 _6156_ (.A(_1176_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_a21oi_1 _6157_ (.A1(_1245_),
    .A2(_1248_),
    .Y(_1249_),
    .B1(net90));
 sg13g2_a22oi_1 _6158_ (.Y(_1250_),
    .B1(_1244_),
    .B2(_1249_),
    .A2(_1243_),
    .A1(net90));
 sg13g2_inv_1 _6159_ (.Y(_1251_),
    .A(_1250_));
 sg13g2_nand2_1 _6160_ (.Y(_1252_),
    .A(net28),
    .B(_1251_));
 sg13g2_nand3_1 _6161_ (.B(_0655_),
    .C(net90),
    .A(_1227_),
    .Y(_1253_));
 sg13g2_nand2_1 _6162_ (.Y(_1254_),
    .A(_1252_),
    .B(_1253_));
 sg13g2_nand2_1 _6163_ (.Y(_1255_),
    .A(_1254_),
    .B(net165));
 sg13g2_buf_2 _6164_ (.A(_1255_),
    .X(_1256_));
 sg13g2_nand2_1 _6165_ (.Y(_1257_),
    .A(net19),
    .B(_1256_));
 sg13g2_nor2_1 _6166_ (.A(_1154_),
    .B(_1163_),
    .Y(_1258_));
 sg13g2_inv_1 _6167_ (.Y(_1259_),
    .A(_1258_));
 sg13g2_nor2_1 _6168_ (.A(_4210_),
    .B(_4177_),
    .Y(_1260_));
 sg13g2_nand2_1 _6169_ (.Y(_1261_),
    .A(_1260_),
    .B(net162));
 sg13g2_xnor2_1 _6170_ (.Y(_1262_),
    .A(_0030_),
    .B(_1261_));
 sg13g2_inv_1 _6171_ (.Y(_1263_),
    .A(net149));
 sg13g2_nor3_1 _6172_ (.A(_1202_),
    .B(_1181_),
    .C(_1263_),
    .Y(_1264_));
 sg13g2_a221oi_1 _6173_ (.B2(_1248_),
    .C1(net90),
    .B1(_1212_),
    .A1(_1201_),
    .Y(_1265_),
    .A2(_1264_));
 sg13g2_a21oi_1 _6174_ (.A1(_1259_),
    .A2(_1262_),
    .Y(_1266_),
    .B1(_1265_));
 sg13g2_nand2_1 _6175_ (.Y(_1267_),
    .A(net28),
    .B(_1266_));
 sg13g2_o21ai_1 _6176_ (.B1(_1267_),
    .Y(_1268_),
    .A1(_0030_),
    .A2(net28));
 sg13g2_nand2_1 _6177_ (.Y(_1269_),
    .A(_1268_),
    .B(net165));
 sg13g2_buf_2 _6178_ (.A(_1269_),
    .X(_1270_));
 sg13g2_inv_4 _6179_ (.A(_1270_),
    .Y(_1271_));
 sg13g2_nor2_1 _6180_ (.A(net139),
    .B(_4210_),
    .Y(_1272_));
 sg13g2_xnor2_1 _6181_ (.Y(_1273_),
    .A(_0800_),
    .B(_1272_));
 sg13g2_xnor2_1 _6182_ (.Y(_1274_),
    .A(_1198_),
    .B(_1189_));
 sg13g2_o21ai_1 _6183_ (.B1(_1216_),
    .Y(_1275_),
    .A1(_1213_),
    .A2(_1274_));
 sg13g2_inv_1 _6184_ (.Y(_1276_),
    .A(_1215_));
 sg13g2_a21oi_1 _6185_ (.A1(_1276_),
    .A2(_1183_),
    .Y(_1277_),
    .B1(_1202_));
 sg13g2_nand2_1 _6186_ (.Y(_1278_),
    .A(_1275_),
    .B(_1277_));
 sg13g2_nor2_1 _6187_ (.A(net148),
    .B(_1263_),
    .Y(_1279_));
 sg13g2_a21oi_1 _6188_ (.A1(_1263_),
    .A2(net137),
    .Y(_1280_),
    .B1(_1197_));
 sg13g2_a22oi_1 _6189_ (.Y(_1281_),
    .B1(net148),
    .B2(_1280_),
    .A2(_1279_),
    .A1(_1207_));
 sg13g2_a21oi_1 _6190_ (.A1(_1202_),
    .A2(_1281_),
    .Y(_1282_),
    .B1(net90));
 sg13g2_a22oi_1 _6191_ (.Y(_1283_),
    .B1(_1278_),
    .B2(_1282_),
    .A2(_1273_),
    .A1(_1259_));
 sg13g2_nand2_1 _6192_ (.Y(_1284_),
    .A(net28),
    .B(_1283_));
 sg13g2_o21ai_1 _6193_ (.B1(_1284_),
    .Y(_1285_),
    .A1(_0799_),
    .A2(_1242_));
 sg13g2_nand2_1 _6194_ (.Y(_1286_),
    .A(_1285_),
    .B(net165));
 sg13g2_buf_8 _6195_ (.A(_1286_),
    .X(_1287_));
 sg13g2_inv_1 _6196_ (.Y(_1288_),
    .A(net28));
 sg13g2_inv_1 _6197_ (.Y(_1289_),
    .A(_0087_));
 sg13g2_nand2_1 _6198_ (.Y(_1290_),
    .A(_1288_),
    .B(_1289_));
 sg13g2_xnor2_1 _6199_ (.Y(_1291_),
    .A(_1289_),
    .B(_1260_));
 sg13g2_inv_1 _6200_ (.Y(_1292_),
    .A(_1210_));
 sg13g2_a21oi_1 _6201_ (.A1(_1292_),
    .A2(_1246_),
    .Y(_1293_),
    .B1(_1176_));
 sg13g2_nand3_1 _6202_ (.B(_1197_),
    .C(net149),
    .A(_1189_),
    .Y(_1294_));
 sg13g2_nand2_1 _6203_ (.Y(_1295_),
    .A(_1294_),
    .B(net137));
 sg13g2_a221oi_1 _6204_ (.B2(_1204_),
    .C1(_1240_),
    .B1(_1295_),
    .A1(_1293_),
    .Y(_1296_),
    .A2(_1212_));
 sg13g2_a21oi_1 _6205_ (.A1(_1259_),
    .A2(_1291_),
    .Y(_1297_),
    .B1(_1296_));
 sg13g2_nand2_1 _6206_ (.Y(_1298_),
    .A(_1242_),
    .B(_1297_));
 sg13g2_nand2_1 _6207_ (.Y(_1299_),
    .A(_1290_),
    .B(_1298_));
 sg13g2_nand2_1 _6208_ (.Y(_1300_),
    .A(_1299_),
    .B(net165));
 sg13g2_buf_8 _6209_ (.A(_1300_),
    .X(_1301_));
 sg13g2_nand2_2 _6210_ (.Y(_1302_),
    .A(_1287_),
    .B(_1301_));
 sg13g2_nor2_2 _6211_ (.A(net26),
    .B(_1302_),
    .Y(_1303_));
 sg13g2_inv_2 _6212_ (.Y(_1304_),
    .A(_1303_));
 sg13g2_nor2_1 _6213_ (.A(_1285_),
    .B(_1301_),
    .Y(_1305_));
 sg13g2_buf_1 _6214_ (.A(_1305_),
    .X(_1306_));
 sg13g2_nand3_1 _6215_ (.B(_1223_),
    .C(_1271_),
    .A(net18),
    .Y(_1307_));
 sg13g2_o21ai_1 _6216_ (.B1(_1307_),
    .Y(_0011_),
    .A1(_1257_),
    .A2(_1304_));
 sg13g2_buf_1 _6217_ (.A(_4141_),
    .X(_1308_));
 sg13g2_nand2_1 _6218_ (.Y(_1309_),
    .A(net27),
    .B(_0654_));
 sg13g2_nand3_1 _6219_ (.B(net86),
    .C(_1250_),
    .A(_1165_),
    .Y(_1310_));
 sg13g2_nand2_2 _6220_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_nor2_1 _6221_ (.A(net147),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_buf_8 _6222_ (.A(_1312_),
    .X(_1313_));
 sg13g2_buf_8 _6223_ (.A(_1287_),
    .X(_1314_));
 sg13g2_nor3_1 _6224_ (.A(_1313_),
    .B(net19),
    .C(net25),
    .Y(_1315_));
 sg13g2_inv_1 _6225_ (.Y(_1316_),
    .A(_0053_));
 sg13g2_o21ai_1 _6226_ (.B1(_1206_),
    .Y(_1317_),
    .A1(_1316_),
    .A2(net137));
 sg13g2_a22oi_1 _6227_ (.Y(_1318_),
    .B1(_1317_),
    .B2(_1249_),
    .A2(net90),
    .A1(_4168_));
 sg13g2_nand2b_1 _6228_ (.Y(_1319_),
    .B(net28),
    .A_N(_1318_));
 sg13g2_nand3_1 _6229_ (.B(_0674_),
    .C(net90),
    .A(_1227_),
    .Y(_1320_));
 sg13g2_nand2_1 _6230_ (.Y(_1321_),
    .A(_1319_),
    .B(_1320_));
 sg13g2_nand3_1 _6231_ (.B(_1321_),
    .C(net165),
    .A(_1223_),
    .Y(_1322_));
 sg13g2_buf_1 _6232_ (.A(_1322_),
    .X(_1323_));
 sg13g2_inv_1 _6233_ (.Y(_1324_),
    .A(_1323_));
 sg13g2_nand2_1 _6234_ (.Y(_1325_),
    .A(_1324_),
    .B(_1314_));
 sg13g2_nor2b_1 _6235_ (.A(_1315_),
    .B_N(_1325_),
    .Y(_1326_));
 sg13g2_nor2_2 _6236_ (.A(_1301_),
    .B(_1270_),
    .Y(_1327_));
 sg13g2_inv_1 _6237_ (.Y(_1328_),
    .A(_1327_));
 sg13g2_nand2_1 _6238_ (.Y(_1329_),
    .A(_1321_),
    .B(net165));
 sg13g2_buf_8 _6239_ (.A(_1329_),
    .X(_1330_));
 sg13g2_nand3_1 _6240_ (.B(net19),
    .C(_1330_),
    .A(_1287_),
    .Y(_1331_));
 sg13g2_buf_2 _6241_ (.A(_1331_),
    .X(_1332_));
 sg13g2_buf_1 _6242_ (.A(_1301_),
    .X(_1333_));
 sg13g2_a21oi_1 _6243_ (.A1(_1332_),
    .A2(net22),
    .Y(_1334_),
    .B1(net26));
 sg13g2_nor2_2 _6244_ (.A(_1311_),
    .B(_1330_),
    .Y(_1335_));
 sg13g2_nand2_1 _6245_ (.Y(_1336_),
    .A(_1335_),
    .B(net23));
 sg13g2_inv_16 _6246_ (.A(_1287_),
    .Y(_1337_));
 sg13g2_nand2_1 _6247_ (.Y(_1338_),
    .A(_1336_),
    .B(_1337_));
 sg13g2_nand2_1 _6248_ (.Y(_1339_),
    .A(net27),
    .B(_0034_));
 sg13g2_nand3_1 _6249_ (.B(net86),
    .C(_1318_),
    .A(_1165_),
    .Y(_1340_));
 sg13g2_nand2_1 _6250_ (.Y(_1341_),
    .A(_1339_),
    .B(_1340_));
 sg13g2_nor2_1 _6251_ (.A(net147),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_a21oi_1 _6252_ (.A1(net25),
    .A2(_1342_),
    .Y(_1343_),
    .B1(net22));
 sg13g2_nand2_1 _6253_ (.Y(_1344_),
    .A(_1338_),
    .B(_1343_));
 sg13g2_nand2_1 _6254_ (.Y(_1345_),
    .A(_1334_),
    .B(_1344_));
 sg13g2_o21ai_1 _6255_ (.B1(_1345_),
    .Y(_0012_),
    .A1(_1326_),
    .A2(_1328_));
 sg13g2_nand2_1 _6256_ (.Y(_1346_),
    .A(_1287_),
    .B(_1313_));
 sg13g2_nand2_1 _6257_ (.Y(_1347_),
    .A(_1338_),
    .B(_1346_));
 sg13g2_inv_4 _6258_ (.A(_1301_),
    .Y(_1348_));
 sg13g2_nand2_1 _6259_ (.Y(_1349_),
    .A(_1347_),
    .B(net21));
 sg13g2_nand3_1 _6260_ (.B(_1223_),
    .C(_1341_),
    .A(_1313_),
    .Y(_1350_));
 sg13g2_buf_1 _6261_ (.A(_1350_),
    .X(_1351_));
 sg13g2_nand2_2 _6262_ (.Y(_1352_),
    .A(_1342_),
    .B(_1256_));
 sg13g2_a21o_1 _6263_ (.A2(_1352_),
    .A1(_1351_),
    .B1(_1302_),
    .X(_1353_));
 sg13g2_nand2_1 _6264_ (.Y(_1354_),
    .A(_1349_),
    .B(_1353_));
 sg13g2_buf_1 _6265_ (.A(_1270_),
    .X(_1355_));
 sg13g2_nand2_1 _6266_ (.Y(_1356_),
    .A(_1354_),
    .B(net24));
 sg13g2_nor2_1 _6267_ (.A(_1223_),
    .B(_1330_),
    .Y(_1357_));
 sg13g2_inv_1 _6268_ (.Y(_1358_),
    .A(_1357_));
 sg13g2_nand3_1 _6269_ (.B(_1256_),
    .C(_1337_),
    .A(_1358_),
    .Y(_1359_));
 sg13g2_nand2_1 _6270_ (.Y(_1360_),
    .A(_1359_),
    .B(_1325_));
 sg13g2_nor3_1 _6271_ (.A(_1254_),
    .B(_1270_),
    .C(_1302_),
    .Y(_1361_));
 sg13g2_a21oi_1 _6272_ (.A1(_1360_),
    .A2(_1327_),
    .Y(_1362_),
    .B1(_1361_));
 sg13g2_nand2_1 _6273_ (.Y(_0013_),
    .A(_1356_),
    .B(_1362_));
 sg13g2_inv_1 _6274_ (.Y(_1363_),
    .A(_1223_));
 sg13g2_nand2_2 _6275_ (.Y(_1364_),
    .A(_1313_),
    .B(_1363_));
 sg13g2_nor2_1 _6276_ (.A(_1341_),
    .B(_1364_),
    .Y(_1365_));
 sg13g2_buf_8 _6277_ (.A(_1337_),
    .X(_1366_));
 sg13g2_a21oi_1 _6278_ (.A1(_1365_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(_1333_));
 sg13g2_nand2_1 _6279_ (.Y(_1368_),
    .A(net19),
    .B(_1330_));
 sg13g2_nand3_1 _6280_ (.B(_1358_),
    .C(net25),
    .A(_1368_),
    .Y(_1369_));
 sg13g2_nand3_1 _6281_ (.B(net24),
    .C(_1369_),
    .A(_1367_),
    .Y(_1370_));
 sg13g2_nand2_1 _6282_ (.Y(_1371_),
    .A(_1360_),
    .B(_1327_));
 sg13g2_nand2_1 _6283_ (.Y(_1372_),
    .A(_1352_),
    .B(_1226_));
 sg13g2_nand3_1 _6284_ (.B(_1364_),
    .C(_1372_),
    .A(_1303_),
    .Y(_1373_));
 sg13g2_nand3_1 _6285_ (.B(_1371_),
    .C(_1373_),
    .A(_1370_),
    .Y(_0014_));
 sg13g2_nor2_1 _6286_ (.A(_1254_),
    .B(_1330_),
    .Y(_1374_));
 sg13g2_nand2_1 _6287_ (.Y(_1375_),
    .A(_1374_),
    .B(net23));
 sg13g2_nand2_1 _6288_ (.Y(_1376_),
    .A(_1375_),
    .B(_1257_));
 sg13g2_nand2_1 _6289_ (.Y(_1377_),
    .A(_1376_),
    .B(net20));
 sg13g2_nand2_1 _6290_ (.Y(_1378_),
    .A(_1377_),
    .B(_1332_));
 sg13g2_nand2_1 _6291_ (.Y(_1379_),
    .A(_1378_),
    .B(_1327_));
 sg13g2_buf_1 _6292_ (.A(net165),
    .X(_1380_));
 sg13g2_nand3_1 _6293_ (.B(_1254_),
    .C(net157),
    .A(_1341_),
    .Y(_1381_));
 sg13g2_nand2_1 _6294_ (.Y(_1382_),
    .A(_1352_),
    .B(_1381_));
 sg13g2_nand2_1 _6295_ (.Y(_1383_),
    .A(_1382_),
    .B(_1225_));
 sg13g2_nand2_1 _6296_ (.Y(_1384_),
    .A(_1383_),
    .B(_1257_));
 sg13g2_nand3_1 _6297_ (.B(net24),
    .C(net18),
    .A(_1384_),
    .Y(_1385_));
 sg13g2_a21o_1 _6298_ (.A2(_1375_),
    .A1(_1351_),
    .B1(_1304_),
    .X(_1386_));
 sg13g2_nand3_1 _6299_ (.B(_1385_),
    .C(_1386_),
    .A(_1379_),
    .Y(_0015_));
 sg13g2_nand2_1 _6300_ (.Y(_1387_),
    .A(_1330_),
    .B(_1256_));
 sg13g2_nor2_1 _6301_ (.A(net19),
    .B(_1387_),
    .Y(_1388_));
 sg13g2_nand2_1 _6302_ (.Y(_1389_),
    .A(_1388_),
    .B(net20));
 sg13g2_a21oi_1 _6303_ (.A1(_1389_),
    .A2(_1332_),
    .Y(_1390_),
    .B1(_1328_));
 sg13g2_nand4_1 _6304_ (.B(net18),
    .C(_1355_),
    .A(_1358_),
    .Y(_1391_),
    .D(_1364_));
 sg13g2_nor2_1 _6305_ (.A(net23),
    .B(_1335_),
    .Y(_1392_));
 sg13g2_a21oi_1 _6306_ (.A1(_1303_),
    .A2(_1392_),
    .Y(_1393_),
    .B1(_1361_));
 sg13g2_nand3b_1 _6307_ (.B(_1391_),
    .C(_1393_),
    .Y(_0016_),
    .A_N(_1390_));
 sg13g2_a22oi_1 _6308_ (.Y(_1394_),
    .B1(_1355_),
    .B2(_1367_),
    .A2(_1392_),
    .A1(_1303_));
 sg13g2_nand2_1 _6309_ (.Y(_0017_),
    .A(_1394_),
    .B(_1379_));
 sg13g2_o21ai_1 _6310_ (.B1(_1332_),
    .Y(_1395_),
    .A1(_1314_),
    .A2(_1375_));
 sg13g2_nand2_1 _6311_ (.Y(_1396_),
    .A(_1395_),
    .B(_1327_));
 sg13g2_nand2_1 _6312_ (.Y(_0018_),
    .A(_1396_),
    .B(_1393_));
 sg13g2_nand2_1 _6313_ (.Y(_1397_),
    .A(_1358_),
    .B(_1381_));
 sg13g2_nand2_1 _6314_ (.Y(_1398_),
    .A(_1397_),
    .B(net20));
 sg13g2_nor2_1 _6315_ (.A(net21),
    .B(_1364_),
    .Y(_1399_));
 sg13g2_a21oi_2 _6316_ (.B1(net26),
    .Y(_1400_),
    .A2(net25),
    .A1(_1399_));
 sg13g2_nand2_1 _6317_ (.Y(_1401_),
    .A(_1302_),
    .B(net26));
 sg13g2_a21oi_1 _6318_ (.A1(_1397_),
    .A2(net22),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_nand3_1 _6319_ (.B(net21),
    .C(_1332_),
    .A(_1359_),
    .Y(_1403_));
 sg13g2_a22oi_1 _6320_ (.Y(_0002_),
    .B1(_1402_),
    .B2(_1403_),
    .A2(_1400_),
    .A1(_1398_));
 sg13g2_nand3_1 _6321_ (.B(_1381_),
    .C(_1226_),
    .A(_1352_),
    .Y(_1404_));
 sg13g2_nand2_1 _6322_ (.Y(_1405_),
    .A(_1404_),
    .B(_1337_));
 sg13g2_nand2_1 _6323_ (.Y(_1406_),
    .A(_1352_),
    .B(net25));
 sg13g2_nand2_1 _6324_ (.Y(_1407_),
    .A(_1405_),
    .B(_1406_));
 sg13g2_nand2_1 _6325_ (.Y(_1408_),
    .A(_1407_),
    .B(net22));
 sg13g2_inv_4 _6326_ (.A(_1387_),
    .Y(_1409_));
 sg13g2_a21oi_1 _6327_ (.A1(_1409_),
    .A2(net20),
    .Y(_1410_),
    .B1(_1333_));
 sg13g2_nand3_1 _6328_ (.B(_1223_),
    .C(_1313_),
    .A(net25),
    .Y(_1411_));
 sg13g2_a21oi_1 _6329_ (.A1(_1410_),
    .A2(_1411_),
    .Y(_1412_),
    .B1(net24));
 sg13g2_o21ai_1 _6330_ (.B1(net18),
    .Y(_1413_),
    .A1(_1374_),
    .A2(_1324_));
 sg13g2_nand2_1 _6331_ (.Y(_1414_),
    .A(_1400_),
    .B(_1413_));
 sg13g2_nor2b_1 _6332_ (.A(_1414_),
    .B_N(_1405_),
    .Y(_1415_));
 sg13g2_a21oi_1 _6333_ (.A1(_1408_),
    .A2(_1412_),
    .Y(_0003_),
    .B1(_1415_));
 sg13g2_nand2_1 _6334_ (.Y(_1416_),
    .A(_1323_),
    .B(_1256_));
 sg13g2_nand2_1 _6335_ (.Y(_1417_),
    .A(_1416_),
    .B(_1337_));
 sg13g2_nand2_1 _6336_ (.Y(_1418_),
    .A(_1287_),
    .B(net23));
 sg13g2_nand2_1 _6337_ (.Y(_1419_),
    .A(_1417_),
    .B(_1418_));
 sg13g2_nand2_1 _6338_ (.Y(_1420_),
    .A(_1419_),
    .B(net21));
 sg13g2_nand2_1 _6339_ (.Y(_1421_),
    .A(_1351_),
    .B(_1337_));
 sg13g2_nand2_1 _6340_ (.Y(_1422_),
    .A(_1421_),
    .B(_1346_));
 sg13g2_nand2_1 _6341_ (.Y(_1423_),
    .A(_1422_),
    .B(net22));
 sg13g2_nand2_1 _6342_ (.Y(_1424_),
    .A(_1420_),
    .B(_1423_));
 sg13g2_nand2_1 _6343_ (.Y(_1425_),
    .A(_1424_),
    .B(net26));
 sg13g2_inv_1 _6344_ (.Y(_1426_),
    .A(_1351_));
 sg13g2_a21oi_1 _6345_ (.A1(_1335_),
    .A2(net19),
    .Y(_1427_),
    .B1(_1409_));
 sg13g2_a22oi_1 _6346_ (.Y(_1428_),
    .B1(net18),
    .B2(_1427_),
    .A2(net20),
    .A1(_1426_));
 sg13g2_nand2_1 _6347_ (.Y(_1429_),
    .A(_1428_),
    .B(net24));
 sg13g2_nand2_1 _6348_ (.Y(_0004_),
    .A(_1425_),
    .B(_1429_));
 sg13g2_o21ai_1 _6349_ (.B1(_1301_),
    .Y(_1430_),
    .A1(net23),
    .A2(_1287_));
 sg13g2_inv_1 _6350_ (.Y(_1431_),
    .A(_1306_));
 sg13g2_a21oi_1 _6351_ (.A1(_1372_),
    .A2(_1375_),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_nand2_1 _6352_ (.Y(_1433_),
    .A(net20),
    .B(net23));
 sg13g2_nand2_1 _6353_ (.Y(_1434_),
    .A(_1400_),
    .B(_1433_));
 sg13g2_nor2_1 _6354_ (.A(_1432_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_a21oi_1 _6355_ (.A1(_1412_),
    .A2(_1430_),
    .Y(_0005_),
    .B1(_1435_));
 sg13g2_o21ai_1 _6356_ (.B1(_1256_),
    .Y(_1436_),
    .A1(net23),
    .A2(net25));
 sg13g2_nand2_1 _6357_ (.Y(_1437_),
    .A(_1436_),
    .B(net22));
 sg13g2_nand2_1 _6358_ (.Y(_1438_),
    .A(_1420_),
    .B(_1437_));
 sg13g2_nand2_1 _6359_ (.Y(_1439_),
    .A(_1438_),
    .B(net26));
 sg13g2_a21oi_1 _6360_ (.A1(net18),
    .A2(_1416_),
    .Y(_1440_),
    .B1(_1315_));
 sg13g2_nand2_1 _6361_ (.Y(_1441_),
    .A(_1440_),
    .B(net24));
 sg13g2_nand2_1 _6362_ (.Y(_0006_),
    .A(_1439_),
    .B(_1441_));
 sg13g2_a22oi_1 _6363_ (.Y(_1442_),
    .B1(net20),
    .B2(_1388_),
    .A2(_1256_),
    .A1(net19));
 sg13g2_nand2_1 _6364_ (.Y(_1443_),
    .A(_1442_),
    .B(net21));
 sg13g2_nand2_1 _6365_ (.Y(_1444_),
    .A(_1337_),
    .B(_1323_));
 sg13g2_nand2_1 _6366_ (.Y(_1445_),
    .A(_1444_),
    .B(_1406_));
 sg13g2_inv_1 _6367_ (.Y(_1446_),
    .A(_1299_));
 sg13g2_a21oi_1 _6368_ (.A1(_1445_),
    .A2(_1446_),
    .Y(_1447_),
    .B1(net24));
 sg13g2_nand2_1 _6369_ (.Y(_1448_),
    .A(_1400_),
    .B(_1444_));
 sg13g2_nand2_1 _6370_ (.Y(_1449_),
    .A(_1409_),
    .B(net19));
 sg13g2_nand3_1 _6371_ (.B(net18),
    .C(_1364_),
    .A(_1449_),
    .Y(_1450_));
 sg13g2_nor2b_1 _6372_ (.A(_1448_),
    .B_N(_1450_),
    .Y(_1451_));
 sg13g2_a21oi_1 _6373_ (.A1(_1443_),
    .A2(_1447_),
    .Y(_0007_),
    .B1(_1451_));
 sg13g2_a21oi_1 _6374_ (.A1(_1383_),
    .A2(_1323_),
    .Y(_1452_),
    .B1(_1431_));
 sg13g2_nand2_1 _6375_ (.Y(_1453_),
    .A(_1427_),
    .B(net20));
 sg13g2_nand2_1 _6376_ (.Y(_1454_),
    .A(_1400_),
    .B(_1453_));
 sg13g2_nor2_1 _6377_ (.A(_1452_),
    .B(_1454_),
    .Y(_1455_));
 sg13g2_nor2_1 _6378_ (.A(net21),
    .B(_1453_),
    .Y(_1456_));
 sg13g2_a21oi_1 _6379_ (.A1(_1285_),
    .A2(_1311_),
    .Y(_1457_),
    .B1(_1446_));
 sg13g2_nor2_1 _6380_ (.A(_1409_),
    .B(_1302_),
    .Y(_1458_));
 sg13g2_nor3_1 _6381_ (.A(_1270_),
    .B(_1457_),
    .C(_1458_),
    .Y(_1459_));
 sg13g2_nor2b_1 _6382_ (.A(_1456_),
    .B_N(_1459_),
    .Y(_1460_));
 sg13g2_nor2_1 _6383_ (.A(_1455_),
    .B(_1460_),
    .Y(_0008_));
 sg13g2_nand2_1 _6384_ (.Y(_1461_),
    .A(_1430_),
    .B(_1270_));
 sg13g2_a21oi_1 _6385_ (.A1(_1446_),
    .A2(_1335_),
    .Y(_1462_),
    .B1(_1461_));
 sg13g2_nor2_1 _6386_ (.A(_1357_),
    .B(_1346_),
    .Y(_1463_));
 sg13g2_nor2_1 _6387_ (.A(net25),
    .B(_1392_),
    .Y(_1464_));
 sg13g2_o21ai_1 _6388_ (.B1(_1348_),
    .Y(_1465_),
    .A1(_1463_),
    .A2(_1464_));
 sg13g2_nand3_1 _6389_ (.B(net26),
    .C(net22),
    .A(_1346_),
    .Y(_1466_));
 sg13g2_nand4_1 _6390_ (.B(net26),
    .C(_1311_),
    .A(_1418_),
    .Y(_1467_),
    .D(net21));
 sg13g2_o21ai_1 _6391_ (.B1(_1467_),
    .Y(_1468_),
    .A1(_1464_),
    .A2(_1466_));
 sg13g2_a21oi_1 _6392_ (.A1(_1462_),
    .A2(_1465_),
    .Y(_0009_),
    .B1(_1468_));
 sg13g2_nor2_1 _6393_ (.A(_1364_),
    .B(net18),
    .Y(_1469_));
 sg13g2_nor3_1 _6394_ (.A(net22),
    .B(_1335_),
    .C(_1418_),
    .Y(_1470_));
 sg13g2_nor2_1 _6395_ (.A(_1469_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_nor2_1 _6396_ (.A(_1399_),
    .B(_1401_),
    .Y(_1472_));
 sg13g2_o21ai_1 _6397_ (.B1(_1366_),
    .Y(_1473_),
    .A1(_1313_),
    .A2(_1357_));
 sg13g2_nand2_1 _6398_ (.Y(_1474_),
    .A(_1473_),
    .B(_1418_));
 sg13g2_nand2_1 _6399_ (.Y(_1475_),
    .A(_1474_),
    .B(net21));
 sg13g2_a22oi_1 _6400_ (.Y(_0010_),
    .B1(_1472_),
    .B2(_1475_),
    .A2(_1471_),
    .A1(net24));
 sg13g2_inv_1 _6401_ (.Y(_1476_),
    .A(_0054_));
 sg13g2_nor2_1 _6402_ (.A(net147),
    .B(_1173_),
    .Y(_1477_));
 sg13g2_inv_1 _6403_ (.Y(_1478_),
    .A(_1477_));
 sg13g2_nor2_1 _6404_ (.A(_1178_),
    .B(_1478_),
    .Y(_1479_));
 sg13g2_a21oi_1 _6405_ (.A1(_1476_),
    .A2(_1478_),
    .Y(_0000_),
    .B1(_1479_));
 sg13g2_inv_1 _6406_ (.Y(_0001_),
    .A(_0000_));
 sg13g2_nor2_2 _6407_ (.A(_4232_),
    .B(net138),
    .Y(_1480_));
 sg13g2_buf_8 _6408_ (.A(_1480_),
    .X(_1481_));
 sg13g2_buf_1 _6409_ (.A(net124),
    .X(_1482_));
 sg13g2_buf_1 _6410_ (.A(net116),
    .X(_1483_));
 sg13g2_nor2_1 _6411_ (.A(_4233_),
    .B(_1050_),
    .Y(_1484_));
 sg13g2_buf_2 _6412_ (.A(_1484_),
    .X(_1485_));
 sg13g2_buf_1 _6413_ (.A(_1485_),
    .X(_1486_));
 sg13g2_a22oi_1 _6414_ (.Y(_1487_),
    .B1(\i_music.i_sample.t3.genblk1[8].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t4.genblk1[8].state.Q ),
    .A1(net112));
 sg13g2_buf_1 _6415_ (.A(_4232_),
    .X(_1488_));
 sg13g2_buf_1 _6416_ (.A(_4233_),
    .X(_1489_));
 sg13g2_nor2_1 _6417_ (.A(_1488_),
    .B(_1489_),
    .Y(_1490_));
 sg13g2_buf_1 _6418_ (.A(_1490_),
    .X(_1491_));
 sg13g2_buf_1 _6419_ (.A(_1491_),
    .X(_1492_));
 sg13g2_buf_1 _6420_ (.A(net122),
    .X(_1493_));
 sg13g2_buf_1 _6421_ (.A(net115),
    .X(_1494_));
 sg13g2_buf_1 _6422_ (.A(net111),
    .X(_1495_));
 sg13g2_buf_1 _6423_ (.A(net108),
    .X(_1496_));
 sg13g2_nand2_1 _6424_ (.Y(_1497_),
    .A(_1496_),
    .B(\i_music.i_sample.t2.genblk1[8].state.Q ));
 sg13g2_inv_1 _6425_ (.Y(_1498_),
    .A(_4234_));
 sg13g2_buf_1 _6426_ (.A(_1498_),
    .X(_1499_));
 sg13g2_buf_1 _6427_ (.A(net129),
    .X(_1500_));
 sg13g2_buf_1 _6428_ (.A(_1500_),
    .X(_1501_));
 sg13g2_nand2_1 _6429_ (.Y(_1502_),
    .A(_1501_),
    .B(\i_music.i_sample.t1.genblk1[8].state.Q ));
 sg13g2_nand3_1 _6430_ (.B(_1497_),
    .C(_1502_),
    .A(_1487_),
    .Y(_0249_));
 sg13g2_a22oi_1 _6431_ (.Y(_1503_),
    .B1(\i_music.i_sample.t3.genblk1[9].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t4.genblk1[9].state.Q ),
    .A1(net112));
 sg13g2_nand2_1 _6432_ (.Y(_1504_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[9].state.Q ));
 sg13g2_nand2_1 _6433_ (.Y(_1505_),
    .A(_1501_),
    .B(\i_music.i_sample.t1.genblk1[9].state.Q ));
 sg13g2_nand3_1 _6434_ (.B(_1504_),
    .C(_1505_),
    .A(_1503_),
    .Y(_0251_));
 sg13g2_a22oi_1 _6435_ (.Y(_1506_),
    .B1(\i_music.i_sample.t3.genblk1[10].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t4.genblk1[10].state.Q ),
    .A1(net112));
 sg13g2_nand2_1 _6436_ (.Y(_1507_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[10].state.Q ));
 sg13g2_nand2_1 _6437_ (.Y(_1508_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[10].state.Q ));
 sg13g2_nand3_1 _6438_ (.B(_1507_),
    .C(_1508_),
    .A(_1506_),
    .Y(_0252_));
 sg13g2_a22oi_1 _6439_ (.Y(_1509_),
    .B1(\i_music.i_sample.t3.genblk1[11].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t4.genblk1[11].state.Q ),
    .A1(net112));
 sg13g2_nand2_1 _6440_ (.Y(_1510_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[11].state.Q ));
 sg13g2_nand2_1 _6441_ (.Y(_1511_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[11].state.Q ));
 sg13g2_nand3_1 _6442_ (.B(_1510_),
    .C(_1511_),
    .A(_1509_),
    .Y(_0253_));
 sg13g2_a22oi_1 _6443_ (.Y(_1512_),
    .B1(\i_music.i_sample.t3.genblk1[12].state.Q ),
    .B2(_1486_),
    .A2(\i_music.i_sample.t4.genblk1[12].state.Q ),
    .A1(net112));
 sg13g2_nand2_1 _6444_ (.Y(_1513_),
    .A(_1496_),
    .B(\i_music.i_sample.t2.genblk1[12].state.Q ));
 sg13g2_nand2_1 _6445_ (.Y(_1514_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[12].state.Q ));
 sg13g2_nand3_1 _6446_ (.B(_1513_),
    .C(_1514_),
    .A(_1512_),
    .Y(_0254_));
 sg13g2_a22oi_1 _6447_ (.Y(_1515_),
    .B1(\i_music.i_sample.t3.genblk1[13].state.Q ),
    .B2(_1486_),
    .A2(\i_music.i_sample.t4.genblk1[13].state.Q ),
    .A1(net116));
 sg13g2_nand2_1 _6448_ (.Y(_1516_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[13].state.Q ));
 sg13g2_nand2_1 _6449_ (.Y(_1517_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[13].state.Q ));
 sg13g2_nand3_1 _6450_ (.B(_1516_),
    .C(_1517_),
    .A(_1515_),
    .Y(_0255_));
 sg13g2_a22oi_1 _6451_ (.Y(_1518_),
    .B1(\i_music.i_sample.t3.genblk1[14].state.Q ),
    .B2(_1485_),
    .A2(\i_music.i_sample.t4.genblk1[14].state.Q ),
    .A1(net116));
 sg13g2_nand2_1 _6452_ (.Y(_1519_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[14].state.Q ));
 sg13g2_nand2_1 _6453_ (.Y(_1520_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[14].state.Q ));
 sg13g2_nand3_1 _6454_ (.B(_1519_),
    .C(_1520_),
    .A(_1518_),
    .Y(_0256_));
 sg13g2_a22oi_1 _6455_ (.Y(_1521_),
    .B1(\i_music.i_sample.t3.genblk1[15].state.Q ),
    .B2(_1485_),
    .A2(\i_music.i_sample.t4.genblk1[15].state.Q ),
    .A1(net116));
 sg13g2_nand2_1 _6456_ (.Y(_1522_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[15].state.Q ));
 sg13g2_nand2_1 _6457_ (.Y(_1523_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[15].state.Q ));
 sg13g2_nand3_1 _6458_ (.B(_1522_),
    .C(_1523_),
    .A(_1521_),
    .Y(_0257_));
 sg13g2_a22oi_1 _6459_ (.Y(_1524_),
    .B1(\i_music.i_sample.t3.genblk1[16].state.Q ),
    .B2(_1485_),
    .A2(\i_music.i_sample.t4.genblk1[16].state.Q ),
    .A1(_1482_));
 sg13g2_nand2_1 _6460_ (.Y(_1525_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[16].state.Q ));
 sg13g2_nand2_1 _6461_ (.Y(_1526_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[16].state.Q ));
 sg13g2_nand3_1 _6462_ (.B(_1525_),
    .C(_1526_),
    .A(_1524_),
    .Y(_0258_));
 sg13g2_a22oi_1 _6463_ (.Y(_1527_),
    .B1(\i_music.i_sample.t3.genblk1[17].state.Q ),
    .B2(_1485_),
    .A2(\i_music.i_sample.t4.genblk1[17].state.Q ),
    .A1(net116));
 sg13g2_nand2_1 _6464_ (.Y(_1528_),
    .A(net101),
    .B(\i_music.i_sample.t2.genblk1[17].state.Q ));
 sg13g2_nand2_1 _6465_ (.Y(_1529_),
    .A(net121),
    .B(\i_music.i_sample.t1.genblk1[17].state.Q ));
 sg13g2_nand3_1 _6466_ (.B(_1528_),
    .C(_1529_),
    .A(_1527_),
    .Y(_0259_));
 sg13g2_buf_1 _6467_ (.A(_4234_),
    .X(_1530_));
 sg13g2_nor2b_1 _6468_ (.A(net136),
    .B_N(\i_music.i_sample.t1.genblk1[18].state.Q ),
    .Y(_0250_));
 sg13g2_buf_1 _6469_ (.A(\i_music.i_sample.t1.genblk1[0].state.Q ),
    .X(_1531_));
 sg13g2_inv_1 _6470_ (.Y(_1532_),
    .A(net80));
 sg13g2_o21ai_1 _6471_ (.B1(net145),
    .Y(_1533_),
    .A1(net146),
    .A2(\i_music.i_sample.t4.genblk1[0].state.Q ));
 sg13g2_buf_1 _6472_ (.A(net108),
    .X(_1534_));
 sg13g2_a22oi_1 _6473_ (.Y(_1535_),
    .B1(\i_music.i_sample.t3.genblk1[0].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t2.genblk1[0].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6474_ (.Y(_0241_),
    .B1(_1533_),
    .B2(_1535_),
    .A2(net114),
    .A1(_1532_));
 sg13g2_buf_1 _6475_ (.A(\i_music.i_sample.t1.genblk1[1].state.Q ),
    .X(_1536_));
 sg13g2_inv_2 _6476_ (.Y(_1537_),
    .A(net79));
 sg13g2_o21ai_1 _6477_ (.B1(net146),
    .Y(_1538_),
    .A1(net145),
    .A2(\i_music.i_sample.t3.genblk1[1].state.Q ));
 sg13g2_a22oi_1 _6478_ (.Y(_1539_),
    .B1(\i_music.i_sample.t4.genblk1[1].state.Q ),
    .B2(net112),
    .A2(\i_music.i_sample.t2.genblk1[1].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6479_ (.Y(_0242_),
    .B1(_1538_),
    .B2(_1539_),
    .A2(net114),
    .A1(_1537_));
 sg13g2_buf_1 _6480_ (.A(\i_music.i_sample.t1.genblk1[2].state.Q ),
    .X(_1540_));
 sg13g2_buf_1 _6481_ (.A(_1540_),
    .X(_1541_));
 sg13g2_inv_1 _6482_ (.Y(_1542_),
    .A(net76));
 sg13g2_buf_1 _6483_ (.A(_1542_),
    .X(_1543_));
 sg13g2_o21ai_1 _6484_ (.B1(net145),
    .Y(_1544_),
    .A1(net146),
    .A2(\i_music.i_sample.t4.genblk1[2].state.Q ));
 sg13g2_a22oi_1 _6485_ (.Y(_1545_),
    .B1(\i_music.i_sample.t3.genblk1[2].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t2.genblk1[2].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6486_ (.Y(_0243_),
    .B1(_1544_),
    .B2(_1545_),
    .A2(net114),
    .A1(_1543_));
 sg13g2_buf_1 _6487_ (.A(\i_music.i_sample.t1.genblk1[3].state.Q ),
    .X(_1546_));
 sg13g2_inv_1 _6488_ (.Y(_1547_),
    .A(net78));
 sg13g2_buf_1 _6489_ (.A(_1547_),
    .X(_1548_));
 sg13g2_buf_1 _6490_ (.A(net70),
    .X(_1549_));
 sg13g2_o21ai_1 _6491_ (.B1(net145),
    .Y(_1550_),
    .A1(net146),
    .A2(\i_music.i_sample.t4.genblk1[3].state.Q ));
 sg13g2_a22oi_1 _6492_ (.Y(_1551_),
    .B1(\i_music.i_sample.t3.genblk1[3].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t2.genblk1[3].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6493_ (.Y(_0244_),
    .B1(_1550_),
    .B2(_1551_),
    .A2(net114),
    .A1(net59));
 sg13g2_buf_1 _6494_ (.A(\i_music.i_sample.t1.genblk1[4].state.Q ),
    .X(_1552_));
 sg13g2_inv_1 _6495_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_buf_1 _6496_ (.A(net75),
    .X(_1554_));
 sg13g2_o21ai_1 _6497_ (.B1(net145),
    .Y(_1555_),
    .A1(net146),
    .A2(\i_music.i_sample.t4.genblk1[4].state.Q ));
 sg13g2_a22oi_1 _6498_ (.Y(_1556_),
    .B1(\i_music.i_sample.t3.genblk1[4].state.Q ),
    .B2(net123),
    .A2(\i_music.i_sample.t2.genblk1[4].state.Q ),
    .A1(_1534_));
 sg13g2_a22oi_1 _6499_ (.Y(_0245_),
    .B1(_1555_),
    .B2(_1556_),
    .A2(net114),
    .A1(_1554_));
 sg13g2_buf_1 _6500_ (.A(\i_music.i_sample.t1.genblk1[5].state.Q ),
    .X(_1557_));
 sg13g2_buf_1 _6501_ (.A(_1557_),
    .X(_1558_));
 sg13g2_inv_1 _6502_ (.Y(_1559_),
    .A(net74));
 sg13g2_buf_1 _6503_ (.A(net68),
    .X(_1560_));
 sg13g2_o21ai_1 _6504_ (.B1(net146),
    .Y(_1561_),
    .A1(net145),
    .A2(\i_music.i_sample.t3.genblk1[5].state.Q ));
 sg13g2_a22oi_1 _6505_ (.Y(_1562_),
    .B1(\i_music.i_sample.t4.genblk1[5].state.Q ),
    .B2(_1483_),
    .A2(\i_music.i_sample.t2.genblk1[5].state.Q ),
    .A1(_1534_));
 sg13g2_a22oi_1 _6506_ (.Y(_0246_),
    .B1(_1561_),
    .B2(_1562_),
    .A2(net114),
    .A1(_1560_));
 sg13g2_buf_1 _6507_ (.A(\i_music.i_sample.t1.genblk1[6].state.Q ),
    .X(_1563_));
 sg13g2_inv_1 _6508_ (.Y(_1564_),
    .A(_1563_));
 sg13g2_buf_1 _6509_ (.A(_1564_),
    .X(_1565_));
 sg13g2_o21ai_1 _6510_ (.B1(net146),
    .Y(_1566_),
    .A1(net145),
    .A2(\i_music.i_sample.t3.genblk1[6].state.Q ));
 sg13g2_a22oi_1 _6511_ (.Y(_1567_),
    .B1(\i_music.i_sample.t4.genblk1[6].state.Q ),
    .B2(net112),
    .A2(\i_music.i_sample.t2.genblk1[6].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6512_ (.Y(_0247_),
    .B1(_1566_),
    .B2(_1567_),
    .A2(net114),
    .A1(net67));
 sg13g2_buf_1 _6513_ (.A(\i_music.i_sample.t1.genblk1[7].state.Q ),
    .X(_1568_));
 sg13g2_inv_2 _6514_ (.Y(_1569_),
    .A(net77));
 sg13g2_o21ai_1 _6515_ (.B1(net146),
    .Y(_1570_),
    .A1(net145),
    .A2(\i_music.i_sample.t3.genblk1[7].state.Q ));
 sg13g2_a22oi_1 _6516_ (.Y(_1571_),
    .B1(\i_music.i_sample.t4.genblk1[7].state.Q ),
    .B2(net112),
    .A2(\i_music.i_sample.t2.genblk1[7].state.Q ),
    .A1(net100));
 sg13g2_a22oi_1 _6517_ (.Y(_0248_),
    .B1(_1570_),
    .B2(_1571_),
    .A2(net114),
    .A1(_1569_));
 sg13g2_inv_1 _6518_ (.Y(_1572_),
    .A(\i_music.count[24] ));
 sg13g2_inv_1 _6519_ (.Y(_1573_),
    .A(_1186_));
 sg13g2_inv_1 _6520_ (.Y(_1574_),
    .A(_1185_));
 sg13g2_inv_1 _6521_ (.Y(_1575_),
    .A(\i_music.count[23] ));
 sg13g2_buf_1 _6522_ (.A(\i_music.count[21] ),
    .X(_1576_));
 sg13g2_nand2_1 _6523_ (.Y(_1577_),
    .A(_1576_),
    .B(\i_music.count[20] ));
 sg13g2_inv_1 _6524_ (.Y(_1578_),
    .A(\i_music.count[19] ));
 sg13g2_inv_1 _6525_ (.Y(_1579_),
    .A(\i_music.count[17] ));
 sg13g2_inv_1 _6526_ (.Y(_1580_),
    .A(\i_music.count[15] ));
 sg13g2_inv_1 _6527_ (.Y(_1581_),
    .A(\i_music.count[13] ));
 sg13g2_nor2_1 _6528_ (.A(_1020_),
    .B(_1236_),
    .Y(_1582_));
 sg13g2_nand2_1 _6529_ (.Y(_1583_),
    .A(_1582_),
    .B(_4225_));
 sg13g2_nor2_1 _6530_ (.A(_1001_),
    .B(_1583_),
    .Y(_1584_));
 sg13g2_nand2_1 _6531_ (.Y(_1585_),
    .A(_1584_),
    .B(_4236_));
 sg13g2_nor2_1 _6532_ (.A(_1155_),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_buf_1 _6533_ (.A(\i_music.count[10] ),
    .X(_1587_));
 sg13g2_nand2_1 _6534_ (.Y(_1588_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_nor2b_1 _6535_ (.A(_1588_),
    .B_N(\i_music.count[11] ),
    .Y(_1589_));
 sg13g2_nand2_1 _6536_ (.Y(_1590_),
    .A(_1589_),
    .B(\i_music.count[12] ));
 sg13g2_nor2_1 _6537_ (.A(_1581_),
    .B(_1590_),
    .Y(_1591_));
 sg13g2_nand2_1 _6538_ (.Y(_1592_),
    .A(_1591_),
    .B(\i_music.count[14] ));
 sg13g2_nor2_1 _6539_ (.A(_1580_),
    .B(_1592_),
    .Y(_1593_));
 sg13g2_nand2_1 _6540_ (.Y(_1594_),
    .A(_1593_),
    .B(\i_music.count[16] ));
 sg13g2_nor2_1 _6541_ (.A(_1579_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_nand2_1 _6542_ (.Y(_1596_),
    .A(_1595_),
    .B(\i_music.count[18] ));
 sg13g2_nor2_1 _6543_ (.A(_1578_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_inv_1 _6544_ (.Y(_1598_),
    .A(_1597_));
 sg13g2_nor2_1 _6545_ (.A(_1577_),
    .B(_1598_),
    .Y(_1599_));
 sg13g2_buf_2 _6546_ (.A(\i_music.count[22] ),
    .X(_1600_));
 sg13g2_nand2_1 _6547_ (.Y(_1601_),
    .A(_1599_),
    .B(_1600_));
 sg13g2_nor2_1 _6548_ (.A(_1575_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_inv_1 _6549_ (.Y(_1603_),
    .A(_1602_));
 sg13g2_nor4_2 _6550_ (.A(_1572_),
    .B(_1573_),
    .C(_1574_),
    .Y(_1604_),
    .D(_1603_));
 sg13g2_nor2_1 _6551_ (.A(_1195_),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_and2_1 _6552_ (.A(_1604_),
    .B(_1195_),
    .X(_1606_));
 sg13g2_buf_1 _6553_ (.A(_1606_),
    .X(_1607_));
 sg13g2_nor3_1 _6554_ (.A(net147),
    .B(_1605_),
    .C(_1607_),
    .Y(_1608_));
 sg13g2_buf_2 _6555_ (.A(_1608_),
    .X(_0175_));
 sg13g2_inv_1 _6556_ (.Y(_1609_),
    .A(_0175_));
 sg13g2_inv_1 _6557_ (.Y(_1610_),
    .A(_1600_));
 sg13g2_nor4_1 _6558_ (.A(_1575_),
    .B(_1572_),
    .C(_1574_),
    .D(_1610_),
    .Y(_1611_));
 sg13g2_a21oi_1 _6559_ (.A1(_1599_),
    .A2(_1611_),
    .Y(_1612_),
    .B1(_1186_));
 sg13g2_nand2b_1 _6560_ (.Y(_1613_),
    .B(_4140_),
    .A_N(_1612_));
 sg13g2_nor2_1 _6561_ (.A(_1613_),
    .B(_1604_),
    .Y(_0174_));
 sg13g2_inv_1 _6562_ (.Y(_1614_),
    .A(_0174_));
 sg13g2_nor2_1 _6563_ (.A(_1572_),
    .B(_1603_),
    .Y(_1615_));
 sg13g2_xnor2_1 _6564_ (.Y(_1616_),
    .A(_1316_),
    .B(_1615_));
 sg13g2_nor2_1 _6565_ (.A(net147),
    .B(_1616_),
    .Y(_0173_));
 sg13g2_nand2_1 _6566_ (.Y(_1617_),
    .A(_1614_),
    .B(_0173_));
 sg13g2_inv_1 _6567_ (.Y(_1618_),
    .A(_0173_));
 sg13g2_nand3_1 _6568_ (.B(_1618_),
    .C(_1614_),
    .A(_1609_),
    .Y(_0151_));
 sg13g2_o21ai_1 _6569_ (.B1(_0151_),
    .Y(_0019_),
    .A1(_1609_),
    .A2(_1617_));
 sg13g2_nand2_1 _6570_ (.Y(_1619_),
    .A(_0173_),
    .B(_0174_));
 sg13g2_nor2_1 _6571_ (.A(_1614_),
    .B(_0175_),
    .Y(_0153_));
 sg13g2_a21oi_1 _6572_ (.A1(_0175_),
    .A2(_1619_),
    .Y(_0020_),
    .B1(_0153_));
 sg13g2_inv_1 _6573_ (.Y(_0154_),
    .A(_0153_));
 sg13g2_nand2_1 _6574_ (.Y(_0021_),
    .A(_0154_),
    .B(_1618_));
 sg13g2_nand2_1 _6575_ (.Y(_1620_),
    .A(_1618_),
    .B(_0174_));
 sg13g2_mux2_1 _6576_ (.A0(_1620_),
    .A1(_1617_),
    .S(_0175_),
    .X(_0022_));
 sg13g2_nand3_1 _6577_ (.B(_1620_),
    .C(_1617_),
    .A(_1609_),
    .Y(_0152_));
 sg13g2_nand2_1 _6578_ (.Y(_1621_),
    .A(_0175_),
    .B(_1619_));
 sg13g2_nand2_1 _6579_ (.Y(_0023_),
    .A(_0152_),
    .B(_1621_));
 sg13g2_nand2_1 _6580_ (.Y(_1622_),
    .A(_1258_),
    .B(net157));
 sg13g2_buf_1 _6581_ (.A(_1622_),
    .X(_1623_));
 sg13g2_nand2_1 _6582_ (.Y(_1624_),
    .A(net89),
    .B(\i_display.frame_crotchet[0] ));
 sg13g2_o21ai_1 _6583_ (.B1(_1624_),
    .Y(_0122_),
    .A1(_1574_),
    .A2(net89));
 sg13g2_nand2_1 _6584_ (.Y(_1625_),
    .A(net89),
    .B(\i_display.frame_crotchet[1] ));
 sg13g2_o21ai_1 _6585_ (.B1(_1625_),
    .Y(_0123_),
    .A1(_1187_),
    .A2(net89));
 sg13g2_buf_1 _6586_ (.A(\i_display.frame_crotchet[2] ),
    .X(_1626_));
 sg13g2_buf_1 _6587_ (.A(_1626_),
    .X(_1627_));
 sg13g2_nand2_1 _6588_ (.Y(_1628_),
    .A(net89),
    .B(net144));
 sg13g2_o21ai_1 _6589_ (.B1(_1628_),
    .Y(_0124_),
    .A1(_1197_),
    .A2(net89));
 sg13g2_buf_1 _6590_ (.A(\i_display.frame_crotchet[3] ),
    .X(_1629_));
 sg13g2_nand2_1 _6591_ (.Y(_1630_),
    .A(_1622_),
    .B(net156));
 sg13g2_o21ai_1 _6592_ (.B1(_1630_),
    .Y(_0125_),
    .A1(_1193_),
    .A2(net89));
 sg13g2_buf_2 _6593_ (.A(\i_display.frame_crotchet[4] ),
    .X(_1631_));
 sg13g2_a21o_1 _6594_ (.A2(net89),
    .A1(_1631_),
    .B1(_1479_),
    .X(_0126_));
 sg13g2_buf_2 _6595_ (.A(\i_display.frame_crotchet[5] ),
    .X(_1632_));
 sg13g2_nand2_1 _6596_ (.Y(_1633_),
    .A(_1622_),
    .B(_1632_));
 sg13g2_o21ai_1 _6597_ (.B1(_1633_),
    .Y(_0127_),
    .A1(net148),
    .A2(_1623_));
 sg13g2_buf_2 _6598_ (.A(\i_display.frame_crotchet[6] ),
    .X(_1634_));
 sg13g2_nand2_1 _6599_ (.Y(_1635_),
    .A(_1622_),
    .B(_1634_));
 sg13g2_o21ai_1 _6600_ (.B1(_1635_),
    .Y(_0128_),
    .A1(_1176_),
    .A2(_1623_));
 sg13g2_inv_1 _6601_ (.Y(_1636_),
    .A(\i_music.i_pwm.count[7] ));
 sg13g2_buf_1 _6602_ (.A(_1380_),
    .X(_1637_));
 sg13g2_o21ai_1 _6603_ (.B1(net143),
    .Y(_1638_),
    .A1(\i_music.i_pwm.sample[7] ),
    .A2(_1636_));
 sg13g2_nand2b_1 _6604_ (.Y(_1639_),
    .B(\i_music.i_pwm.count[6] ),
    .A_N(\i_music.i_pwm.sample[6] ));
 sg13g2_inv_1 _6605_ (.Y(_1640_),
    .A(\i_music.i_pwm.count[5] ));
 sg13g2_nor2_1 _6606_ (.A(\i_music.i_pwm.sample[5] ),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_inv_1 _6607_ (.Y(_1642_),
    .A(\i_music.i_pwm.count[4] ));
 sg13g2_nor2_1 _6608_ (.A(\i_music.i_pwm.sample[4] ),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_inv_1 _6609_ (.Y(_1644_),
    .A(\i_music.i_pwm.count[3] ));
 sg13g2_nor2_1 _6610_ (.A(\i_music.i_pwm.sample[3] ),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_nor2_1 _6611_ (.A(_1643_),
    .B(_1645_),
    .Y(_1646_));
 sg13g2_nor2b_1 _6612_ (.A(\i_music.i_pwm.count[0] ),
    .B_N(\i_music.i_pwm.sample[0] ),
    .Y(_1647_));
 sg13g2_inv_1 _6613_ (.Y(_1648_),
    .A(\i_music.i_pwm.sample[1] ));
 sg13g2_buf_1 _6614_ (.A(\i_music.i_pwm.count[1] ),
    .X(_1649_));
 sg13g2_nand2_1 _6615_ (.Y(_1650_),
    .A(_1648_),
    .B(_1649_));
 sg13g2_nor2_1 _6616_ (.A(_1649_),
    .B(_1648_),
    .Y(_1651_));
 sg13g2_a21oi_1 _6617_ (.A1(_1647_),
    .A2(_1650_),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_inv_1 _6618_ (.Y(_1653_),
    .A(\i_music.i_pwm.count[2] ));
 sg13g2_nor2_1 _6619_ (.A(\i_music.i_pwm.sample[2] ),
    .B(_1653_),
    .Y(_1654_));
 sg13g2_inv_1 _6620_ (.Y(_1655_),
    .A(_1654_));
 sg13g2_nand2b_1 _6621_ (.Y(_1656_),
    .B(_1655_),
    .A_N(_1652_));
 sg13g2_nand2_1 _6622_ (.Y(_1657_),
    .A(_1644_),
    .B(\i_music.i_pwm.sample[3] ));
 sg13g2_nand2_1 _6623_ (.Y(_1658_),
    .A(_1653_),
    .B(\i_music.i_pwm.sample[2] ));
 sg13g2_nand3_1 _6624_ (.B(_1657_),
    .C(_1658_),
    .A(_1656_),
    .Y(_1659_));
 sg13g2_a22oi_1 _6625_ (.Y(_1660_),
    .B1(_1646_),
    .B2(_1659_),
    .A2(\i_music.i_pwm.sample[4] ),
    .A1(_1642_));
 sg13g2_inv_1 _6626_ (.Y(_1661_),
    .A(\i_music.i_pwm.count[6] ));
 sg13g2_a22oi_1 _6627_ (.Y(_1662_),
    .B1(_1661_),
    .B2(\i_music.i_pwm.sample[6] ),
    .A2(\i_music.i_pwm.sample[5] ),
    .A1(_1640_));
 sg13g2_o21ai_1 _6628_ (.B1(_1662_),
    .Y(_1663_),
    .A1(_1641_),
    .A2(_1660_));
 sg13g2_a22oi_1 _6629_ (.Y(_1664_),
    .B1(_1639_),
    .B2(_1663_),
    .A2(\i_music.i_pwm.sample[7] ),
    .A1(_1636_));
 sg13g2_buf_1 _6630_ (.A(net147),
    .X(_1665_));
 sg13g2_buf_1 _6631_ (.A(net135),
    .X(_1666_));
 sg13g2_nand2_1 _6632_ (.Y(_1667_),
    .A(net128),
    .B(\i_music.i_pwm.pwm ));
 sg13g2_o21ai_1 _6633_ (.B1(_1667_),
    .Y(_0196_),
    .A1(_1638_),
    .A2(_1664_));
 sg13g2_inv_1 _6634_ (.Y(_1668_),
    .A(\i_music.i_sample.sample_acc[0] ));
 sg13g2_inv_1 _6635_ (.Y(_1669_),
    .A(\i_music.violin_note_idx[2][8] ));
 sg13g2_inv_1 _6636_ (.Y(_1670_),
    .A(\i_music.violin_note_idx[3][8] ));
 sg13g2_nor2b_1 _6637_ (.A(_4233_),
    .B_N(_0086_),
    .Y(_1671_));
 sg13g2_a221oi_1 _6638_ (.B2(net129),
    .C1(_1671_),
    .B1(_1670_),
    .A1(net124),
    .Y(_1672_),
    .A2(_1669_));
 sg13g2_buf_1 _6639_ (.A(_1672_),
    .X(_1673_));
 sg13g2_inv_1 _6640_ (.Y(_1674_),
    .A(\i_music.violin_note_idx[2][3] ));
 sg13g2_inv_1 _6641_ (.Y(_1675_),
    .A(\i_music.violin_note_idx[3][3] ));
 sg13g2_nand2_1 _6642_ (.Y(_1676_),
    .A(net138),
    .B(_0079_));
 sg13g2_inv_1 _6643_ (.Y(_1677_),
    .A(_1676_));
 sg13g2_a221oi_1 _6644_ (.B2(_1498_),
    .C1(_1677_),
    .B1(_1675_),
    .A1(_1481_),
    .Y(_1678_),
    .A2(_1674_));
 sg13g2_buf_2 _6645_ (.A(_1678_),
    .X(_1679_));
 sg13g2_buf_8 _6646_ (.A(_1679_),
    .X(_1680_));
 sg13g2_buf_1 _6647_ (.A(net107),
    .X(_1681_));
 sg13g2_buf_1 _6648_ (.A(\i_music.violin_note_idx[3][1] ),
    .X(_1682_));
 sg13g2_inv_1 _6649_ (.Y(_1683_),
    .A(\i_music.violin_note_idx[2][1] ));
 sg13g2_nand2_1 _6650_ (.Y(_1684_),
    .A(net138),
    .B(_0082_));
 sg13g2_inv_1 _6651_ (.Y(_1685_),
    .A(_1684_));
 sg13g2_a21oi_1 _6652_ (.A1(_1480_),
    .A2(_1683_),
    .Y(_1686_),
    .B1(_1685_));
 sg13g2_o21ai_1 _6653_ (.B1(_1686_),
    .Y(_1687_),
    .A1(_1682_),
    .A2(_4234_));
 sg13g2_buf_2 _6654_ (.A(_1687_),
    .X(_1688_));
 sg13g2_inv_1 _6655_ (.Y(_1689_),
    .A(\i_music.violin_note_idx[2][2] ));
 sg13g2_a22oi_1 _6656_ (.Y(_1690_),
    .B1(_1689_),
    .B2(net124),
    .A2(_0083_),
    .A1(_1157_));
 sg13g2_o21ai_1 _6657_ (.B1(_1690_),
    .Y(_1691_),
    .A1(\i_music.violin_note_idx[3][2] ),
    .A2(net136));
 sg13g2_buf_1 _6658_ (.A(_1691_),
    .X(_1692_));
 sg13g2_inv_2 _6659_ (.Y(_1693_),
    .A(net106));
 sg13g2_nor2_1 _6660_ (.A(_1688_),
    .B(net98),
    .Y(_1694_));
 sg13g2_inv_1 _6661_ (.Y(_1695_),
    .A(_1694_));
 sg13g2_inv_1 _6662_ (.Y(_1696_),
    .A(\i_music.violin_note_idx[2][5] ));
 sg13g2_inv_1 _6663_ (.Y(_1697_),
    .A(\i_music.violin_note_idx[3][5] ));
 sg13g2_nand2_1 _6664_ (.Y(_1698_),
    .A(net138),
    .B(_0078_));
 sg13g2_inv_1 _6665_ (.Y(_1699_),
    .A(_1698_));
 sg13g2_a221oi_1 _6666_ (.B2(net129),
    .C1(_1699_),
    .B1(_1697_),
    .A1(net124),
    .Y(_1700_),
    .A2(_1696_));
 sg13g2_buf_1 _6667_ (.A(_1700_),
    .X(_1701_));
 sg13g2_inv_1 _6668_ (.Y(_1702_),
    .A(\i_music.violin_note_idx[2][4] ));
 sg13g2_inv_1 _6669_ (.Y(_1703_),
    .A(\i_music.violin_note_idx[3][4] ));
 sg13g2_nand2_1 _6670_ (.Y(_1704_),
    .A(net138),
    .B(_0080_));
 sg13g2_inv_1 _6671_ (.Y(_1705_),
    .A(_1704_));
 sg13g2_a221oi_1 _6672_ (.B2(_1498_),
    .C1(_1705_),
    .B1(_1703_),
    .A1(net124),
    .Y(_1706_),
    .A2(_1702_));
 sg13g2_buf_1 _6673_ (.A(_1706_),
    .X(_1707_));
 sg13g2_nor2_2 _6674_ (.A(_1701_),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_inv_1 _6675_ (.Y(_1709_),
    .A(_1708_));
 sg13g2_inv_1 _6676_ (.Y(_1710_),
    .A(\i_music.violin_note_idx[2][6] ));
 sg13g2_inv_1 _6677_ (.Y(_1711_),
    .A(\i_music.violin_note_idx[3][6] ));
 sg13g2_nand2_1 _6678_ (.Y(_1712_),
    .A(net138),
    .B(_0081_));
 sg13g2_inv_1 _6679_ (.Y(_1713_),
    .A(_1712_));
 sg13g2_a221oi_1 _6680_ (.B2(_1499_),
    .C1(_1713_),
    .B1(_1711_),
    .A1(net124),
    .Y(_1714_),
    .A2(_1710_));
 sg13g2_buf_1 _6681_ (.A(_1714_),
    .X(_1715_));
 sg13g2_inv_1 _6682_ (.Y(_1716_),
    .A(\i_music.violin_note_idx[2][7] ));
 sg13g2_nand2_1 _6683_ (.Y(_1717_),
    .A(_1157_),
    .B(_0084_));
 sg13g2_inv_1 _6684_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_a221oi_1 _6685_ (.B2(_1499_),
    .C1(_1718_),
    .B1(_0085_),
    .A1(_1481_),
    .Y(_1719_),
    .A2(_1716_));
 sg13g2_buf_1 _6686_ (.A(_1719_),
    .X(_1720_));
 sg13g2_inv_1 _6687_ (.Y(_1721_),
    .A(_1720_));
 sg13g2_nor2_1 _6688_ (.A(_1715_),
    .B(_1721_),
    .Y(_1722_));
 sg13g2_inv_1 _6689_ (.Y(_1723_),
    .A(_1722_));
 sg13g2_nor2_1 _6690_ (.A(_1709_),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_inv_1 _6691_ (.Y(_1725_),
    .A(_1724_));
 sg13g2_nor4_1 _6692_ (.A(_1673_),
    .B(net99),
    .C(_1695_),
    .D(_1725_),
    .Y(_1726_));
 sg13g2_buf_1 _6693_ (.A(_1726_),
    .X(_1727_));
 sg13g2_buf_1 _6694_ (.A(net106),
    .X(_1728_));
 sg13g2_buf_2 _6695_ (.A(\i_music.violin_note_idx[3][0] ),
    .X(_1729_));
 sg13g2_inv_1 _6696_ (.Y(_1730_),
    .A(\i_music.violin_note_idx[2][0] ));
 sg13g2_nand2_1 _6697_ (.Y(_1731_),
    .A(net138),
    .B(_0103_));
 sg13g2_inv_1 _6698_ (.Y(_1732_),
    .A(_1731_));
 sg13g2_a21oi_1 _6699_ (.A1(_1480_),
    .A2(_1730_),
    .Y(_1733_),
    .B1(_1732_));
 sg13g2_o21ai_1 _6700_ (.B1(_1733_),
    .Y(_1734_),
    .A1(_1729_),
    .A2(net136));
 sg13g2_buf_1 _6701_ (.A(_1734_),
    .X(_1735_));
 sg13g2_inv_1 _6702_ (.Y(_1736_),
    .A(net105));
 sg13g2_inv_2 _6703_ (.Y(_1737_),
    .A(_1688_));
 sg13g2_nand2_1 _6704_ (.Y(_1738_),
    .A(_1736_),
    .B(_1737_));
 sg13g2_buf_2 _6705_ (.A(_1738_),
    .X(_1739_));
 sg13g2_nor2_1 _6706_ (.A(net97),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_buf_1 _6707_ (.A(_1701_),
    .X(_1741_));
 sg13g2_nor2_1 _6708_ (.A(_1741_),
    .B(_1723_),
    .Y(_1742_));
 sg13g2_inv_1 _6709_ (.Y(_1743_),
    .A(_1742_));
 sg13g2_inv_1 _6710_ (.Y(_1744_),
    .A(net110));
 sg13g2_buf_1 _6711_ (.A(_1744_),
    .X(_1745_));
 sg13g2_nor2_1 _6712_ (.A(net107),
    .B(net96),
    .Y(_1746_));
 sg13g2_nor2b_1 _6713_ (.A(_1743_),
    .B_N(_1746_),
    .Y(_1747_));
 sg13g2_buf_1 _6714_ (.A(_1741_),
    .X(_1748_));
 sg13g2_inv_2 _6715_ (.Y(_1749_),
    .A(_1679_));
 sg13g2_nor2_2 _6716_ (.A(_1749_),
    .B(_1744_),
    .Y(_1750_));
 sg13g2_nor2_2 _6717_ (.A(_1737_),
    .B(net98),
    .Y(_1751_));
 sg13g2_inv_1 _6718_ (.Y(_1752_),
    .A(_1751_));
 sg13g2_nor2_2 _6719_ (.A(_1679_),
    .B(net110),
    .Y(_1753_));
 sg13g2_nand2_2 _6720_ (.Y(_1754_),
    .A(_1751_),
    .B(_1735_));
 sg13g2_inv_1 _6721_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_a22oi_1 _6722_ (.Y(_1756_),
    .B1(_1753_),
    .B2(_1755_),
    .A2(_1752_),
    .A1(_1750_));
 sg13g2_buf_1 _6723_ (.A(_1749_),
    .X(_1757_));
 sg13g2_nand2_1 _6724_ (.Y(_1758_),
    .A(_1754_),
    .B(_1757_));
 sg13g2_nor2_1 _6725_ (.A(net105),
    .B(_1749_),
    .Y(_1759_));
 sg13g2_buf_2 _6726_ (.A(_1759_),
    .X(_1760_));
 sg13g2_nor2_1 _6727_ (.A(_1688_),
    .B(_1692_),
    .Y(_1761_));
 sg13g2_buf_2 _6728_ (.A(_1761_),
    .X(_1762_));
 sg13g2_nand2_1 _6729_ (.Y(_1763_),
    .A(_1760_),
    .B(_1762_));
 sg13g2_inv_1 _6730_ (.Y(_1764_),
    .A(_1701_));
 sg13g2_nor2_1 _6731_ (.A(net110),
    .B(_1764_),
    .Y(_1765_));
 sg13g2_buf_2 _6732_ (.A(_1765_),
    .X(_1766_));
 sg13g2_nand3_1 _6733_ (.B(_1763_),
    .C(_1766_),
    .A(_1758_),
    .Y(_1767_));
 sg13g2_o21ai_1 _6734_ (.B1(_1767_),
    .Y(_1768_),
    .A1(net95),
    .A2(_1756_));
 sg13g2_inv_2 _6735_ (.Y(_1769_),
    .A(_1715_));
 sg13g2_nor2_2 _6736_ (.A(_1769_),
    .B(_1721_),
    .Y(_1770_));
 sg13g2_a221oi_1 _6737_ (.B2(_1770_),
    .C1(_1673_),
    .B1(_1768_),
    .A1(_1740_),
    .Y(_1771_),
    .A2(_1747_));
 sg13g2_inv_1 _6738_ (.Y(_1772_),
    .A(_1771_));
 sg13g2_buf_1 _6739_ (.A(_1707_),
    .X(_1773_));
 sg13g2_nor2_2 _6740_ (.A(net105),
    .B(_1737_),
    .Y(_1774_));
 sg13g2_inv_1 _6741_ (.Y(_1775_),
    .A(_1774_));
 sg13g2_nor2_1 _6742_ (.A(net97),
    .B(_1775_),
    .Y(_1776_));
 sg13g2_nor2_1 _6743_ (.A(net103),
    .B(_1776_),
    .Y(_1777_));
 sg13g2_nor2_1 _6744_ (.A(net107),
    .B(_1752_),
    .Y(_1778_));
 sg13g2_inv_1 _6745_ (.Y(_1779_),
    .A(_1778_));
 sg13g2_nor2_1 _6746_ (.A(_1688_),
    .B(_1749_),
    .Y(_1780_));
 sg13g2_a21oi_1 _6747_ (.A1(_1780_),
    .A2(net98),
    .Y(_1781_),
    .B1(_1760_));
 sg13g2_a22oi_1 _6748_ (.Y(_1782_),
    .B1(net103),
    .B2(_1781_),
    .A2(_1779_),
    .A1(_1777_));
 sg13g2_nand2b_1 _6749_ (.Y(_1783_),
    .B(net95),
    .A_N(_1782_));
 sg13g2_nand2_1 _6750_ (.Y(_1784_),
    .A(_1737_),
    .B(net105));
 sg13g2_buf_1 _6751_ (.A(_1784_),
    .X(_1785_));
 sg13g2_o21ai_1 _6752_ (.B1(_1749_),
    .Y(_1786_),
    .A1(net106),
    .A2(_1785_));
 sg13g2_buf_1 _6753_ (.A(_1786_),
    .X(_1787_));
 sg13g2_nor2_1 _6754_ (.A(_1694_),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_nor2_1 _6755_ (.A(net98),
    .B(_1785_),
    .Y(_1789_));
 sg13g2_inv_2 _6756_ (.Y(_1790_),
    .A(_1789_));
 sg13g2_o21ai_1 _6757_ (.B1(_1790_),
    .Y(_1791_),
    .A1(net99),
    .A2(_1788_));
 sg13g2_nand2_1 _6758_ (.Y(_1792_),
    .A(_1791_),
    .B(_1708_));
 sg13g2_a21oi_1 _6759_ (.A1(_1783_),
    .A2(_1792_),
    .Y(_1793_),
    .B1(_1723_));
 sg13g2_nor2_1 _6760_ (.A(_1762_),
    .B(_1758_),
    .Y(_1794_));
 sg13g2_nor2_1 _6761_ (.A(net105),
    .B(net106),
    .Y(_1795_));
 sg13g2_inv_1 _6762_ (.Y(_1796_),
    .A(_1795_));
 sg13g2_nand2_1 _6763_ (.Y(_1797_),
    .A(_1794_),
    .B(_1796_));
 sg13g2_buf_1 _6764_ (.A(_1764_),
    .X(_1798_));
 sg13g2_nor2_2 _6765_ (.A(net93),
    .B(net96),
    .Y(_1799_));
 sg13g2_nand2_1 _6766_ (.Y(_1800_),
    .A(net99),
    .B(net98));
 sg13g2_nand3_1 _6767_ (.B(_1799_),
    .C(_1800_),
    .A(_1797_),
    .Y(_1801_));
 sg13g2_nand2_1 _6768_ (.Y(_1802_),
    .A(_1739_),
    .B(net97));
 sg13g2_nor2_1 _6769_ (.A(_1680_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_nor2_1 _6770_ (.A(net95),
    .B(_1753_),
    .Y(_1804_));
 sg13g2_o21ai_1 _6771_ (.B1(_1804_),
    .Y(_1805_),
    .A1(_1803_),
    .A2(_1777_));
 sg13g2_inv_1 _6772_ (.Y(_1806_),
    .A(_1776_));
 sg13g2_nor2_2 _6773_ (.A(_1795_),
    .B(_1749_),
    .Y(_1807_));
 sg13g2_inv_1 _6774_ (.Y(_1808_),
    .A(_1807_));
 sg13g2_nand2_1 _6775_ (.Y(_1809_),
    .A(_1806_),
    .B(_1808_));
 sg13g2_nand3_1 _6776_ (.B(net97),
    .C(net107),
    .A(_1739_),
    .Y(_1810_));
 sg13g2_nand3_1 _6777_ (.B(_1766_),
    .C(_1810_),
    .A(_1809_),
    .Y(_1811_));
 sg13g2_nand3_1 _6778_ (.B(_1805_),
    .C(_1811_),
    .A(_1801_),
    .Y(_1812_));
 sg13g2_inv_1 _6779_ (.Y(_1813_),
    .A(_1799_));
 sg13g2_buf_1 _6780_ (.A(net94),
    .X(_1814_));
 sg13g2_nor2_1 _6781_ (.A(net106),
    .B(_1736_),
    .Y(_1815_));
 sg13g2_inv_1 _6782_ (.Y(_1816_),
    .A(_1815_));
 sg13g2_a22oi_1 _6783_ (.Y(_1817_),
    .B1(_1688_),
    .B2(_1807_),
    .A2(_1816_),
    .A1(net88));
 sg13g2_nor2_1 _6784_ (.A(_1813_),
    .B(_1817_),
    .Y(_1818_));
 sg13g2_nor2_2 _6785_ (.A(net104),
    .B(net96),
    .Y(_1819_));
 sg13g2_nand2_1 _6786_ (.Y(_1820_),
    .A(_1778_),
    .B(_1709_));
 sg13g2_o21ai_1 _6787_ (.B1(_1820_),
    .Y(_1821_),
    .A1(_1819_),
    .A2(_1778_));
 sg13g2_nand2_1 _6788_ (.Y(_1822_),
    .A(_1790_),
    .B(net94));
 sg13g2_nand2_1 _6789_ (.Y(_1823_),
    .A(_1822_),
    .B(_1810_));
 sg13g2_nand2_1 _6790_ (.Y(_1824_),
    .A(_1823_),
    .B(_1766_));
 sg13g2_nand3_1 _6791_ (.B(_1824_),
    .C(_1715_),
    .A(_1821_),
    .Y(_1825_));
 sg13g2_o21ai_1 _6792_ (.B1(_1721_),
    .Y(_1826_),
    .A1(_1818_),
    .A2(_1825_));
 sg13g2_a21oi_1 _6793_ (.A1(_1812_),
    .A2(_1769_),
    .Y(_1827_),
    .B1(_1826_));
 sg13g2_nor3_1 _6794_ (.A(_1772_),
    .B(_1793_),
    .C(_1827_),
    .Y(_1828_));
 sg13g2_inv_1 _6795_ (.Y(_1829_),
    .A(_1753_));
 sg13g2_nor2b_1 _6796_ (.A(_1774_),
    .B_N(_1785_),
    .Y(_1830_));
 sg13g2_nor3_1 _6797_ (.A(net98),
    .B(_1829_),
    .C(_1830_),
    .Y(_1831_));
 sg13g2_nor2_1 _6798_ (.A(_1736_),
    .B(_1679_),
    .Y(_1832_));
 sg13g2_inv_2 _6799_ (.Y(_1833_),
    .A(_1673_));
 sg13g2_nor2_1 _6800_ (.A(_1715_),
    .B(_1720_),
    .Y(_1834_));
 sg13g2_inv_1 _6801_ (.Y(_1835_),
    .A(_1834_));
 sg13g2_nor2_1 _6802_ (.A(_1833_),
    .B(_1835_),
    .Y(_1836_));
 sg13g2_o21ai_1 _6803_ (.B1(_1836_),
    .Y(_1837_),
    .A1(_1709_),
    .A2(_1832_));
 sg13g2_a21oi_1 _6804_ (.A1(_1819_),
    .A2(_1763_),
    .Y(_1838_),
    .B1(_1837_));
 sg13g2_o21ai_1 _6805_ (.B1(_1838_),
    .Y(_1839_),
    .A1(net93),
    .A2(_1831_));
 sg13g2_nor2b_1 _6806_ (.A(_1828_),
    .B_N(_1839_),
    .Y(_1840_));
 sg13g2_buf_1 _6807_ (.A(_1840_),
    .X(_1841_));
 sg13g2_inv_2 _6808_ (.Y(_1842_),
    .A(_1841_));
 sg13g2_nor2_1 _6809_ (.A(_1727_),
    .B(_1842_),
    .Y(_1843_));
 sg13g2_nor2_1 _6810_ (.A(net106),
    .B(_1737_),
    .Y(_1844_));
 sg13g2_inv_1 _6811_ (.Y(_1845_),
    .A(_1844_));
 sg13g2_nor2_1 _6812_ (.A(_1736_),
    .B(net98),
    .Y(_1846_));
 sg13g2_inv_1 _6813_ (.Y(_1847_),
    .A(_1846_));
 sg13g2_nand2_1 _6814_ (.Y(_1848_),
    .A(_1847_),
    .B(_1796_));
 sg13g2_a221oi_1 _6815_ (.B2(net94),
    .C1(net96),
    .B1(_1848_),
    .A1(_1760_),
    .Y(_1849_),
    .A2(_1845_));
 sg13g2_nand2_1 _6816_ (.Y(_1850_),
    .A(_1830_),
    .B(net106));
 sg13g2_nor2_1 _6817_ (.A(net105),
    .B(_1679_),
    .Y(_1851_));
 sg13g2_a21oi_1 _6818_ (.A1(_1850_),
    .A2(_1807_),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_inv_1 _6819_ (.Y(_1853_),
    .A(_1760_));
 sg13g2_nand2_1 _6820_ (.Y(_1854_),
    .A(_1775_),
    .B(_1749_));
 sg13g2_a21oi_1 _6821_ (.A1(_1853_),
    .A2(_1854_),
    .Y(_1855_),
    .B1(net97));
 sg13g2_o21ai_1 _6822_ (.B1(net96),
    .Y(_1856_),
    .A1(_1789_),
    .A2(_1855_));
 sg13g2_nor2_1 _6823_ (.A(net105),
    .B(_1762_),
    .Y(_1857_));
 sg13g2_a21oi_1 _6824_ (.A1(_1737_),
    .A2(_1815_),
    .Y(_1858_),
    .B1(_1857_));
 sg13g2_nand2_1 _6825_ (.Y(_1859_),
    .A(_1858_),
    .B(net94));
 sg13g2_nand3_1 _6826_ (.B(net110),
    .C(_1853_),
    .A(_1859_),
    .Y(_1860_));
 sg13g2_a21oi_1 _6827_ (.A1(_1856_),
    .A2(_1860_),
    .Y(_1861_),
    .B1(net104));
 sg13g2_a221oi_1 _6828_ (.B2(_1852_),
    .C1(_1861_),
    .B1(_1766_),
    .A1(net104),
    .Y(_1862_),
    .A2(_1849_));
 sg13g2_nand2_1 _6829_ (.Y(_1863_),
    .A(_1862_),
    .B(_1715_));
 sg13g2_nor2_1 _6830_ (.A(_1679_),
    .B(_1857_),
    .Y(_1864_));
 sg13g2_inv_1 _6831_ (.Y(_1865_),
    .A(_1864_));
 sg13g2_o21ai_1 _6832_ (.B1(_1865_),
    .Y(_1866_),
    .A1(net94),
    .A2(_1739_));
 sg13g2_nor2_1 _6833_ (.A(net110),
    .B(_1760_),
    .Y(_1867_));
 sg13g2_a21o_1 _6834_ (.A2(net110),
    .A1(_1866_),
    .B1(_1867_),
    .X(_1868_));
 sg13g2_nand2_1 _6835_ (.Y(_1869_),
    .A(_1785_),
    .B(net98));
 sg13g2_nor2_1 _6836_ (.A(_1679_),
    .B(_1869_),
    .Y(_1870_));
 sg13g2_a21oi_1 _6837_ (.A1(_1845_),
    .A2(_1785_),
    .Y(_1871_),
    .B1(net94));
 sg13g2_o21ai_1 _6838_ (.B1(net96),
    .Y(_1872_),
    .A1(_1870_),
    .A2(_1871_));
 sg13g2_nor2_1 _6839_ (.A(net107),
    .B(_1694_),
    .Y(_1873_));
 sg13g2_a21oi_1 _6840_ (.A1(_1832_),
    .A2(_1844_),
    .Y(_1874_),
    .B1(_1744_));
 sg13g2_o21ai_1 _6841_ (.B1(_1874_),
    .Y(_1875_),
    .A1(_1760_),
    .A2(_1873_));
 sg13g2_a21oi_1 _6842_ (.A1(_1872_),
    .A2(_1875_),
    .Y(_1876_),
    .B1(net93));
 sg13g2_a21oi_1 _6843_ (.A1(_1868_),
    .A2(net93),
    .Y(_1877_),
    .B1(_1876_));
 sg13g2_a21oi_1 _6844_ (.A1(_1877_),
    .A2(_1769_),
    .Y(_1878_),
    .B1(_1720_));
 sg13g2_nand2_1 _6845_ (.Y(_1879_),
    .A(_1863_),
    .B(_1878_));
 sg13g2_inv_1 _6846_ (.Y(_1880_),
    .A(_1762_));
 sg13g2_a21oi_1 _6847_ (.A1(_1807_),
    .A2(_1880_),
    .Y(_1881_),
    .B1(_1866_));
 sg13g2_buf_1 _6848_ (.A(_1745_),
    .X(_1882_));
 sg13g2_a21oi_1 _6849_ (.A1(_1881_),
    .A2(net87),
    .Y(_1883_),
    .B1(_1743_));
 sg13g2_inv_1 _6850_ (.Y(_1884_),
    .A(_1822_));
 sg13g2_a21oi_1 _6851_ (.A1(_1884_),
    .A2(_1796_),
    .Y(_1885_),
    .B1(net87));
 sg13g2_o21ai_1 _6852_ (.B1(_1885_),
    .Y(_1886_),
    .A1(net88),
    .A2(_1857_));
 sg13g2_nor2_2 _6853_ (.A(_1774_),
    .B(net94),
    .Y(_1887_));
 sg13g2_nand2_1 _6854_ (.Y(_1888_),
    .A(_1785_),
    .B(net97));
 sg13g2_nand2_1 _6855_ (.Y(_1889_),
    .A(_1887_),
    .B(_1888_));
 sg13g2_nor2_1 _6856_ (.A(net110),
    .B(_1832_),
    .Y(_1890_));
 sg13g2_nand2_1 _6857_ (.Y(_1891_),
    .A(_1865_),
    .B(_1853_));
 sg13g2_a22oi_1 _6858_ (.Y(_1892_),
    .B1(net110),
    .B2(_1891_),
    .A2(_1890_),
    .A1(_1889_));
 sg13g2_o21ai_1 _6859_ (.B1(_1867_),
    .Y(_1893_),
    .A1(_1846_),
    .A2(_1787_));
 sg13g2_nor2_1 _6860_ (.A(_1736_),
    .B(_1694_),
    .Y(_1894_));
 sg13g2_a21oi_1 _6861_ (.A1(_1894_),
    .A2(_1746_),
    .Y(_1895_),
    .B1(net93));
 sg13g2_nand2_1 _6862_ (.Y(_1896_),
    .A(_1858_),
    .B(_1750_));
 sg13g2_nand3_1 _6863_ (.B(_1895_),
    .C(_1896_),
    .A(_1893_),
    .Y(_1897_));
 sg13g2_o21ai_1 _6864_ (.B1(_1897_),
    .Y(_1898_),
    .A1(net104),
    .A2(_1892_));
 sg13g2_nor2_2 _6865_ (.A(_1762_),
    .B(_1749_),
    .Y(_1899_));
 sg13g2_nor2_1 _6866_ (.A(_1760_),
    .B(_1899_),
    .Y(_1900_));
 sg13g2_nor2b_1 _6867_ (.A(_1900_),
    .B_N(_1888_),
    .Y(_1901_));
 sg13g2_inv_1 _6868_ (.Y(_1902_),
    .A(_1750_));
 sg13g2_inv_1 _6869_ (.Y(_1903_),
    .A(_1851_));
 sg13g2_o21ai_1 _6870_ (.B1(_1903_),
    .Y(_1904_),
    .A1(_1894_),
    .A2(_1902_));
 sg13g2_a22oi_1 _6871_ (.Y(_1905_),
    .B1(net104),
    .B2(_1904_),
    .A2(_1766_),
    .A1(_1901_));
 sg13g2_nor2_1 _6872_ (.A(_1723_),
    .B(_1905_),
    .Y(_1906_));
 sg13g2_a221oi_1 _6873_ (.B2(_1770_),
    .C1(_1906_),
    .B1(_1898_),
    .A1(_1883_),
    .Y(_1907_),
    .A2(_1886_));
 sg13g2_nand2_1 _6874_ (.Y(_1908_),
    .A(_1879_),
    .B(_1907_));
 sg13g2_a21oi_1 _6875_ (.A1(_1903_),
    .A2(_1739_),
    .Y(_1909_),
    .B1(net87));
 sg13g2_a21o_1 _6876_ (.A2(_1822_),
    .A1(_1867_),
    .B1(_1909_),
    .X(_1910_));
 sg13g2_nor2_1 _6877_ (.A(net95),
    .B(_1835_),
    .Y(_1911_));
 sg13g2_a21oi_1 _6878_ (.A1(_1910_),
    .A2(_1911_),
    .Y(_1912_),
    .B1(_1833_));
 sg13g2_a21oi_1 _6879_ (.A1(_1908_),
    .A2(_1833_),
    .Y(_1913_),
    .B1(_1912_));
 sg13g2_buf_2 _6880_ (.A(_1913_),
    .X(_1914_));
 sg13g2_inv_1 _6881_ (.Y(_1915_),
    .A(_1914_));
 sg13g2_nand2_1 _6882_ (.Y(_1916_),
    .A(_1774_),
    .B(net97));
 sg13g2_nor2_1 _6883_ (.A(_1681_),
    .B(_1916_),
    .Y(_1917_));
 sg13g2_nor2_1 _6884_ (.A(_1851_),
    .B(_1857_),
    .Y(_1918_));
 sg13g2_inv_1 _6885_ (.Y(_1919_),
    .A(_1918_));
 sg13g2_a22oi_1 _6886_ (.Y(_1920_),
    .B1(_1798_),
    .B2(_1919_),
    .A2(net87),
    .A1(_1917_));
 sg13g2_nor3_1 _6887_ (.A(_1708_),
    .B(_1835_),
    .C(_1920_),
    .Y(_1921_));
 sg13g2_nand2_1 _6888_ (.Y(_1922_),
    .A(_1739_),
    .B(_1693_));
 sg13g2_o21ai_1 _6889_ (.B1(_1808_),
    .Y(_1923_),
    .A1(net99),
    .A2(_1751_));
 sg13g2_a22oi_1 _6890_ (.Y(_1924_),
    .B1(net87),
    .B2(_1923_),
    .A2(_1750_),
    .A1(_1922_));
 sg13g2_o21ai_1 _6891_ (.B1(_1777_),
    .Y(_1925_),
    .A1(net99),
    .A2(_1754_));
 sg13g2_nand2_1 _6892_ (.Y(_1926_),
    .A(_1781_),
    .B(_1874_));
 sg13g2_nand3_1 _6893_ (.B(_1926_),
    .C(net95),
    .A(_1925_),
    .Y(_1927_));
 sg13g2_o21ai_1 _6894_ (.B1(_1927_),
    .Y(_1928_),
    .A1(_1748_),
    .A2(_1924_));
 sg13g2_nand2_1 _6895_ (.Y(_1929_),
    .A(_1850_),
    .B(net99));
 sg13g2_nand3_1 _6896_ (.B(_1929_),
    .C(_1708_),
    .A(_1797_),
    .Y(_1930_));
 sg13g2_nand3_1 _6897_ (.B(_1819_),
    .C(_1810_),
    .A(_1822_),
    .Y(_1931_));
 sg13g2_nand4_1 _6898_ (.B(_1770_),
    .C(_1767_),
    .A(_1930_),
    .Y(_1932_),
    .D(_1931_));
 sg13g2_nand2_1 _6899_ (.Y(_1933_),
    .A(_1932_),
    .B(_1833_));
 sg13g2_a21oi_1 _6900_ (.A1(_1722_),
    .A2(_1928_),
    .Y(_1934_),
    .B1(_1933_));
 sg13g2_nand2_1 _6901_ (.Y(_1935_),
    .A(_1780_),
    .B(_1847_));
 sg13g2_inv_1 _6902_ (.Y(_1936_),
    .A(_1935_));
 sg13g2_nor3_1 _6903_ (.A(net103),
    .B(_1936_),
    .C(_1794_),
    .Y(_1937_));
 sg13g2_o21ai_1 _6904_ (.B1(_1779_),
    .Y(_1938_),
    .A1(net88),
    .A2(_1916_));
 sg13g2_o21ai_1 _6905_ (.B1(net93),
    .Y(_1939_),
    .A1(net87),
    .A2(_1938_));
 sg13g2_a22oi_1 _6906_ (.Y(_1940_),
    .B1(_1802_),
    .B2(_1899_),
    .A2(_1815_),
    .A1(_1814_));
 sg13g2_nand2_1 _6907_ (.Y(_1941_),
    .A(_1847_),
    .B(_1814_));
 sg13g2_nand3_1 _6908_ (.B(_1754_),
    .C(net87),
    .A(_1941_),
    .Y(_1942_));
 sg13g2_o21ai_1 _6909_ (.B1(_1942_),
    .Y(_1943_),
    .A1(_1882_),
    .A2(_1940_));
 sg13g2_nand2_1 _6910_ (.Y(_1944_),
    .A(_1943_),
    .B(_1748_));
 sg13g2_o21ai_1 _6911_ (.B1(_1944_),
    .Y(_1945_),
    .A1(_1937_),
    .A2(_1939_));
 sg13g2_a21oi_1 _6912_ (.A1(_1806_),
    .A2(_1754_),
    .Y(_1946_),
    .B1(net88));
 sg13g2_o21ai_1 _6913_ (.B1(_1773_),
    .Y(_1947_),
    .A1(_1803_),
    .A2(_1946_));
 sg13g2_o21ai_1 _6914_ (.B1(_1947_),
    .Y(_1948_),
    .A1(_1773_),
    .A2(_1946_));
 sg13g2_a21oi_1 _6915_ (.A1(_1847_),
    .A2(_1775_),
    .Y(_1949_),
    .B1(_1680_));
 sg13g2_nor2b_1 _6916_ (.A(_1848_),
    .B_N(_1899_),
    .Y(_1950_));
 sg13g2_o21ai_1 _6917_ (.B1(_1766_),
    .Y(_1951_),
    .A1(_1949_),
    .A2(_1950_));
 sg13g2_nand2_1 _6918_ (.Y(_1952_),
    .A(_1735_),
    .B(_1688_));
 sg13g2_a21oi_1 _6919_ (.A1(_1952_),
    .A2(_1728_),
    .Y(_1953_),
    .B1(_1681_));
 sg13g2_o21ai_1 _6920_ (.B1(_1799_),
    .Y(_1954_),
    .A1(_1899_),
    .A2(_1953_));
 sg13g2_nand2_1 _6921_ (.Y(_1955_),
    .A(_1951_),
    .B(_1954_));
 sg13g2_a21oi_1 _6922_ (.A1(_1948_),
    .A2(_1798_),
    .Y(_1956_),
    .B1(_1955_));
 sg13g2_a21oi_1 _6923_ (.A1(_1956_),
    .A2(_1769_),
    .Y(_1957_),
    .B1(_1720_));
 sg13g2_o21ai_1 _6924_ (.B1(_1957_),
    .Y(_1958_),
    .A1(_1769_),
    .A2(_1945_));
 sg13g2_a22oi_1 _6925_ (.Y(_1959_),
    .B1(_1934_),
    .B2(_1958_),
    .A2(_1921_),
    .A1(_1673_));
 sg13g2_buf_2 _6926_ (.A(_1959_),
    .X(_1960_));
 sg13g2_nand2_1 _6927_ (.Y(_1961_),
    .A(_1915_),
    .B(_1960_));
 sg13g2_inv_2 _6928_ (.Y(_1962_),
    .A(_1960_));
 sg13g2_nand2_1 _6929_ (.Y(_1963_),
    .A(_1962_),
    .B(_1914_));
 sg13g2_inv_1 _6930_ (.Y(_1964_),
    .A(_1850_));
 sg13g2_nor2_1 _6931_ (.A(_1762_),
    .B(_1964_),
    .Y(_1965_));
 sg13g2_inv_1 _6932_ (.Y(_1966_),
    .A(_1965_));
 sg13g2_nand2_1 _6933_ (.Y(_1967_),
    .A(_1850_),
    .B(_1757_));
 sg13g2_nor2b_1 _6934_ (.A(_1967_),
    .B_N(_1922_),
    .Y(_1968_));
 sg13g2_a21oi_1 _6935_ (.A1(_1966_),
    .A2(net107),
    .Y(_1969_),
    .B1(_1968_));
 sg13g2_a21oi_1 _6936_ (.A1(_1869_),
    .A2(_1887_),
    .Y(_1970_),
    .B1(_1788_));
 sg13g2_a21oi_1 _6937_ (.A1(_1970_),
    .A2(net103),
    .Y(_1971_),
    .B1(net104));
 sg13g2_o21ai_1 _6938_ (.B1(_1971_),
    .Y(_1972_),
    .A1(net103),
    .A2(_1969_));
 sg13g2_o21ai_1 _6939_ (.B1(_1766_),
    .Y(_1973_),
    .A1(_1887_),
    .A2(_1968_));
 sg13g2_nand2_1 _6940_ (.Y(_1974_),
    .A(_1964_),
    .B(net107));
 sg13g2_nand4_1 _6941_ (.B(_1796_),
    .C(_1799_),
    .A(_1974_),
    .Y(_1975_),
    .D(_1779_));
 sg13g2_nand3_1 _6942_ (.B(_1973_),
    .C(_1975_),
    .A(_1972_),
    .Y(_1976_));
 sg13g2_a22oi_1 _6943_ (.Y(_1977_),
    .B1(net94),
    .B2(_1964_),
    .A2(_1887_),
    .A1(_1848_));
 sg13g2_inv_1 _6944_ (.Y(_1978_),
    .A(_1780_));
 sg13g2_a22oi_1 _6945_ (.Y(_1979_),
    .B1(_1808_),
    .B2(_1978_),
    .A2(_1775_),
    .A1(net97));
 sg13g2_nand3b_1 _6946_ (.B(_1745_),
    .C(_1854_),
    .Y(_1980_),
    .A_N(_1979_));
 sg13g2_o21ai_1 _6947_ (.B1(_1980_),
    .Y(_1981_),
    .A1(net87),
    .A2(_1977_));
 sg13g2_inv_1 _6948_ (.Y(_1982_),
    .A(_1967_));
 sg13g2_a21oi_1 _6949_ (.A1(_1982_),
    .A2(_1816_),
    .Y(_1983_),
    .B1(_1979_));
 sg13g2_inv_1 _6950_ (.Y(_1984_),
    .A(_1830_));
 sg13g2_a21oi_1 _6951_ (.A1(_1984_),
    .A2(_1899_),
    .Y(_1985_),
    .B1(net104));
 sg13g2_nor2_1 _6952_ (.A(_1819_),
    .B(_1985_),
    .Y(_1986_));
 sg13g2_a21oi_1 _6953_ (.A1(_1983_),
    .A2(net103),
    .Y(_1987_),
    .B1(_1986_));
 sg13g2_a21oi_1 _6954_ (.A1(_1981_),
    .A2(net95),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_a21oi_1 _6955_ (.A1(_1988_),
    .A2(_1769_),
    .Y(_1989_),
    .B1(_1720_));
 sg13g2_o21ai_1 _6956_ (.B1(_1989_),
    .Y(_1990_),
    .A1(_1769_),
    .A2(_1976_));
 sg13g2_nor2_1 _6957_ (.A(net107),
    .B(_1965_),
    .Y(_1991_));
 sg13g2_o21ai_1 _6958_ (.B1(_1819_),
    .Y(_1992_),
    .A1(_1815_),
    .A2(_1978_));
 sg13g2_nor2_1 _6959_ (.A(net106),
    .B(_1984_),
    .Y(_1993_));
 sg13g2_nor2b_1 _6960_ (.A(_1993_),
    .B_N(_1746_),
    .Y(_1994_));
 sg13g2_a22oi_1 _6961_ (.Y(_1995_),
    .B1(_1753_),
    .B2(_1789_),
    .A2(net96),
    .A1(_1774_));
 sg13g2_o21ai_1 _6962_ (.B1(_1995_),
    .Y(_1996_),
    .A1(_1858_),
    .A2(_1902_));
 sg13g2_o21ai_1 _6963_ (.B1(net104),
    .Y(_1997_),
    .A1(_1994_),
    .A2(_1996_));
 sg13g2_o21ai_1 _6964_ (.B1(_1997_),
    .Y(_1998_),
    .A1(_1991_),
    .A2(_1992_));
 sg13g2_nand2_1 _6965_ (.Y(_1999_),
    .A(_1974_),
    .B(_1763_));
 sg13g2_a21oi_1 _6966_ (.A1(net88),
    .A2(_1984_),
    .Y(_2000_),
    .B1(_1999_));
 sg13g2_a21oi_1 _6967_ (.A1(_1887_),
    .A2(_1695_),
    .Y(_2001_),
    .B1(net96));
 sg13g2_nand2_1 _6968_ (.Y(_2002_),
    .A(_2001_),
    .B(_1865_));
 sg13g2_inv_1 _6969_ (.Y(_2003_),
    .A(_1993_));
 sg13g2_a21oi_1 _6970_ (.A1(_2003_),
    .A2(_1890_),
    .Y(_2004_),
    .B1(net93));
 sg13g2_a22oi_1 _6971_ (.Y(_2005_),
    .B1(_2002_),
    .B2(_2004_),
    .A2(_1985_),
    .A1(_1885_));
 sg13g2_o21ai_1 _6972_ (.B1(_2005_),
    .Y(_2006_),
    .A1(_1709_),
    .A2(_2000_));
 sg13g2_o21ai_1 _6973_ (.B1(_1935_),
    .Y(_2007_),
    .A1(_1795_),
    .A2(_1737_));
 sg13g2_o21ai_1 _6974_ (.B1(_1833_),
    .Y(_2008_),
    .A1(_1725_),
    .A2(_2007_));
 sg13g2_a221oi_1 _6975_ (.B2(_1770_),
    .C1(_2008_),
    .B1(_2006_),
    .A1(_1998_),
    .Y(_2009_),
    .A2(_1722_));
 sg13g2_nand2_1 _6976_ (.Y(_2010_),
    .A(_1990_),
    .B(_2009_));
 sg13g2_o21ai_1 _6977_ (.B1(_1867_),
    .Y(_2011_),
    .A1(_1755_),
    .A2(_1787_));
 sg13g2_o21ai_1 _6978_ (.B1(net88),
    .Y(_2012_),
    .A1(net105),
    .A2(_1844_));
 sg13g2_nand2_1 _6979_ (.Y(_2013_),
    .A(_1807_),
    .B(_1916_));
 sg13g2_nand3_1 _6980_ (.B(net103),
    .C(_2013_),
    .A(_2012_),
    .Y(_2014_));
 sg13g2_nand3_1 _6981_ (.B(net93),
    .C(_2014_),
    .A(_2011_),
    .Y(_2015_));
 sg13g2_o21ai_1 _6982_ (.B1(net95),
    .Y(_2016_),
    .A1(_1829_),
    .A2(_1790_));
 sg13g2_nand3_1 _6983_ (.B(_1836_),
    .C(_2016_),
    .A(_2015_),
    .Y(_2017_));
 sg13g2_nand2_1 _6984_ (.Y(_2018_),
    .A(_2010_),
    .B(_2017_));
 sg13g2_buf_2 _6985_ (.A(_2018_),
    .X(_2019_));
 sg13g2_inv_1 _6986_ (.Y(_2020_),
    .A(_2019_));
 sg13g2_a21oi_1 _6987_ (.A1(_1961_),
    .A2(_1963_),
    .Y(_2021_),
    .B1(_2020_));
 sg13g2_nor2_1 _6988_ (.A(_1962_),
    .B(_2020_),
    .Y(_2022_));
 sg13g2_o21ai_1 _6989_ (.B1(_1841_),
    .Y(_2023_),
    .A1(_1914_),
    .A2(_2022_));
 sg13g2_o21ai_1 _6990_ (.B1(_2023_),
    .Y(_2024_),
    .A1(_1843_),
    .A2(_2021_));
 sg13g2_inv_1 _6991_ (.Y(_2025_),
    .A(_1491_));
 sg13g2_nand2_1 _6992_ (.Y(_2026_),
    .A(_2024_),
    .B(_2025_));
 sg13g2_xnor2_1 _6993_ (.Y(_2027_),
    .A(_1600_),
    .B(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3] ));
 sg13g2_inv_1 _6994_ (.Y(_2028_),
    .A(_2027_));
 sg13g2_inv_1 _6995_ (.Y(_2029_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[2] ));
 sg13g2_nor2_1 _6996_ (.A(_1576_),
    .B(\i_music.count[20] ),
    .Y(_2030_));
 sg13g2_inv_1 _6997_ (.Y(_2031_),
    .A(_1577_));
 sg13g2_nor2_1 _6998_ (.A(_2030_),
    .B(_2031_),
    .Y(_2032_));
 sg13g2_xor2_1 _6999_ (.B(_2032_),
    .A(_0077_),
    .X(_2033_));
 sg13g2_nor2_1 _7000_ (.A(_2029_),
    .B(_2033_),
    .Y(_2034_));
 sg13g2_xnor2_1 _7001_ (.Y(_2035_),
    .A(\i_music.count[19] ),
    .B(_1576_));
 sg13g2_o21ai_1 _7002_ (.B1(_2035_),
    .Y(_2036_),
    .A1(_2031_),
    .A2(_2030_));
 sg13g2_xnor2_1 _7003_ (.Y(_2037_),
    .A(_1600_),
    .B(_2036_));
 sg13g2_nor2b_1 _7004_ (.A(_2037_),
    .B_N(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1] ),
    .Y(_2038_));
 sg13g2_inv_1 _7005_ (.Y(_2039_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0] ));
 sg13g2_nand2_1 _7006_ (.Y(_2040_),
    .A(_2032_),
    .B(_2035_));
 sg13g2_xnor2_1 _7007_ (.Y(_2041_),
    .A(_1600_),
    .B(_2040_));
 sg13g2_nor2_1 _7008_ (.A(_2039_),
    .B(_2041_),
    .Y(_2042_));
 sg13g2_inv_1 _7009_ (.Y(_2043_),
    .A(_2042_));
 sg13g2_xnor2_1 _7010_ (.Y(_2044_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1] ),
    .B(_2037_));
 sg13g2_inv_1 _7011_ (.Y(_2045_),
    .A(_2044_));
 sg13g2_nor2_1 _7012_ (.A(_2043_),
    .B(_2045_),
    .Y(_2046_));
 sg13g2_nor2_1 _7013_ (.A(_2038_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_inv_1 _7014_ (.Y(_2048_),
    .A(_2047_));
 sg13g2_nand2_1 _7015_ (.Y(_2049_),
    .A(_2033_),
    .B(_2029_));
 sg13g2_o21ai_1 _7016_ (.B1(_2049_),
    .Y(_2050_),
    .A1(_2034_),
    .A2(_2048_));
 sg13g2_nor2_1 _7017_ (.A(_2028_),
    .B(_2050_),
    .Y(_2051_));
 sg13g2_a21oi_2 _7018_ (.B1(_2051_),
    .Y(_2052_),
    .A2(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3] ),
    .A1(_1610_));
 sg13g2_nand2b_1 _7019_ (.Y(_2053_),
    .B(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4] ),
    .A_N(_2052_));
 sg13g2_buf_1 _7020_ (.A(\i_music.violin_note_idx[1][7] ),
    .X(_2054_));
 sg13g2_nand2_1 _7021_ (.Y(_2055_),
    .A(_2054_),
    .B(\i_music.violin_note_idx[1][8] ));
 sg13g2_nand2_1 _7022_ (.Y(_2056_),
    .A(_1491_),
    .B(_2055_));
 sg13g2_inv_1 _7023_ (.Y(_2057_),
    .A(_2056_));
 sg13g2_nand2b_1 _7024_ (.Y(_2058_),
    .B(_2052_),
    .A_N(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4] ));
 sg13g2_nand3_1 _7025_ (.B(_2057_),
    .C(_2058_),
    .A(_2053_),
    .Y(_2059_));
 sg13g2_nand2_1 _7026_ (.Y(_2060_),
    .A(_2026_),
    .B(_2059_));
 sg13g2_nor2_1 _7027_ (.A(_2019_),
    .B(_1914_),
    .Y(_2061_));
 sg13g2_nor3_1 _7028_ (.A(_1842_),
    .B(_2061_),
    .C(_2022_),
    .Y(_2062_));
 sg13g2_nor2_1 _7029_ (.A(_1492_),
    .B(_1727_),
    .Y(_2063_));
 sg13g2_nand2_1 _7030_ (.Y(_2064_),
    .A(_2061_),
    .B(_1960_));
 sg13g2_nand3b_1 _7031_ (.B(_2063_),
    .C(_2064_),
    .Y(_2065_),
    .A_N(_2062_));
 sg13g2_inv_1 _7032_ (.Y(_2066_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[6] ));
 sg13g2_inv_1 _7033_ (.Y(_2067_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[5] ));
 sg13g2_nor3_1 _7034_ (.A(_0055_),
    .B(_2067_),
    .C(_2052_),
    .Y(_2068_));
 sg13g2_inv_1 _7035_ (.Y(_2069_),
    .A(_2068_));
 sg13g2_nor2_1 _7036_ (.A(_2066_),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_inv_1 _7037_ (.Y(_2071_),
    .A(_2070_));
 sg13g2_inv_1 _7038_ (.Y(_2072_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7] ));
 sg13g2_a21oi_1 _7039_ (.A1(_2071_),
    .A2(_2072_),
    .Y(_2073_),
    .B1(_2056_));
 sg13g2_nor2_1 _7040_ (.A(_2072_),
    .B(_2071_),
    .Y(_2074_));
 sg13g2_inv_1 _7041_ (.Y(_2075_),
    .A(_2074_));
 sg13g2_nand2_1 _7042_ (.Y(_2076_),
    .A(_2073_),
    .B(_2075_));
 sg13g2_nand2_1 _7043_ (.Y(_2077_),
    .A(_2065_),
    .B(_2076_));
 sg13g2_nand2_1 _7044_ (.Y(_2078_),
    .A(_2019_),
    .B(_1842_));
 sg13g2_nor2_1 _7045_ (.A(_1962_),
    .B(_2061_),
    .Y(_2079_));
 sg13g2_nor2_1 _7046_ (.A(_2020_),
    .B(_1915_),
    .Y(_2080_));
 sg13g2_inv_1 _7047_ (.Y(_2081_),
    .A(_2080_));
 sg13g2_a221oi_1 _7048_ (.B2(_2081_),
    .C1(_1727_),
    .B1(_2079_),
    .A1(_1962_),
    .Y(_2082_),
    .A2(_2078_));
 sg13g2_o21ai_1 _7049_ (.B1(_2067_),
    .Y(_2083_),
    .A1(_0055_),
    .A2(_2052_));
 sg13g2_nand3_1 _7050_ (.B(_2069_),
    .C(_2057_),
    .A(_2083_),
    .Y(_2084_));
 sg13g2_o21ai_1 _7051_ (.B1(_2084_),
    .Y(_2085_),
    .A1(net122),
    .A2(_2082_));
 sg13g2_nand2_1 _7052_ (.Y(_2086_),
    .A(_2081_),
    .B(_1962_));
 sg13g2_nor2_1 _7053_ (.A(_2061_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_o21ai_1 _7054_ (.B1(_1841_),
    .Y(_2088_),
    .A1(_2022_),
    .A2(_2087_));
 sg13g2_a21oi_1 _7055_ (.A1(_2079_),
    .A2(_1842_),
    .Y(_2089_),
    .B1(_1727_));
 sg13g2_a21oi_1 _7056_ (.A1(_2088_),
    .A2(_2089_),
    .Y(_2090_),
    .B1(net122));
 sg13g2_o21ai_1 _7057_ (.B1(_2066_),
    .Y(_2091_),
    .A1(_2067_),
    .A2(_2053_));
 sg13g2_nor3_1 _7058_ (.A(_2067_),
    .B(_2066_),
    .C(_2053_),
    .Y(_2092_));
 sg13g2_inv_1 _7059_ (.Y(_2093_),
    .A(_2092_));
 sg13g2_nand3_1 _7060_ (.B(_2093_),
    .C(_2057_),
    .A(_2091_),
    .Y(_2094_));
 sg13g2_nand2b_1 _7061_ (.Y(_2095_),
    .B(_2094_),
    .A_N(_2090_));
 sg13g2_nor4_1 _7062_ (.A(_2060_),
    .B(_2077_),
    .C(_2085_),
    .D(_2095_),
    .Y(_2096_));
 sg13g2_nand3_1 _7063_ (.B(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7] ),
    .C(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8] ),
    .A(_2092_),
    .Y(_2097_));
 sg13g2_nand3b_1 _7064_ (.B(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0] ),
    .C(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10] ),
    .Y(_2098_),
    .A_N(_2097_));
 sg13g2_inv_1 _7065_ (.Y(_2099_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10] ));
 sg13g2_o21ai_1 _7066_ (.B1(_2099_),
    .Y(_2100_),
    .A1(_2039_),
    .A2(_2097_));
 sg13g2_nand3_1 _7067_ (.B(_2100_),
    .C(_2057_),
    .A(_2098_),
    .Y(_2101_));
 sg13g2_nor2_1 _7068_ (.A(_1842_),
    .B(_2019_),
    .Y(_2102_));
 sg13g2_nand4_1 _7069_ (.B(_1914_),
    .C(_1960_),
    .A(_2102_),
    .Y(_2103_),
    .D(_2063_));
 sg13g2_inv_1 _7070_ (.Y(_2104_),
    .A(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8] ));
 sg13g2_o21ai_1 _7071_ (.B1(_2039_),
    .Y(_2105_),
    .A1(_2104_),
    .A2(_2075_));
 sg13g2_nand3_1 _7072_ (.B(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0] ),
    .C(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8] ),
    .A(_2074_),
    .Y(_2106_));
 sg13g2_nand3_1 _7073_ (.B(_2057_),
    .C(_2106_),
    .A(_2105_),
    .Y(_2107_));
 sg13g2_nand2_1 _7074_ (.Y(_2108_),
    .A(_2103_),
    .B(_2107_));
 sg13g2_a22oi_1 _7075_ (.Y(_2109_),
    .B1(_1842_),
    .B2(_2064_),
    .A2(_1960_),
    .A1(_2102_));
 sg13g2_nand2_1 _7076_ (.Y(_2110_),
    .A(_2109_),
    .B(_2025_));
 sg13g2_o21ai_1 _7077_ (.B1(_2104_),
    .Y(_2111_),
    .A1(_2072_),
    .A2(_2093_));
 sg13g2_nand3_1 _7078_ (.B(_2057_),
    .C(_2097_),
    .A(_2111_),
    .Y(_2112_));
 sg13g2_nand2_1 _7079_ (.Y(_2113_),
    .A(_2110_),
    .B(_2112_));
 sg13g2_nor2_1 _7080_ (.A(_2108_),
    .B(_2113_),
    .Y(_2114_));
 sg13g2_nand2_1 _7081_ (.Y(_2115_),
    .A(_2078_),
    .B(_1962_));
 sg13g2_inv_1 _7082_ (.Y(_2116_),
    .A(_2115_));
 sg13g2_o21ai_1 _7083_ (.B1(_1915_),
    .Y(_2117_),
    .A1(_2102_),
    .A2(_2116_));
 sg13g2_nor2_1 _7084_ (.A(_1727_),
    .B(_1915_),
    .Y(_2118_));
 sg13g2_a21oi_1 _7085_ (.A1(_2115_),
    .A2(_2118_),
    .Y(_2119_),
    .B1(net122));
 sg13g2_nand2_1 _7086_ (.Y(_2120_),
    .A(_2117_),
    .B(_2119_));
 sg13g2_nor2_1 _7087_ (.A(_2056_),
    .B(_2046_),
    .Y(_2121_));
 sg13g2_o21ai_1 _7088_ (.B1(_2121_),
    .Y(_2122_),
    .A1(_2042_),
    .A2(_2044_));
 sg13g2_nand2_1 _7089_ (.Y(_2123_),
    .A(_2120_),
    .B(_2122_));
 sg13g2_o21ai_1 _7090_ (.B1(_1842_),
    .Y(_2124_),
    .A1(_2079_),
    .A2(_2087_));
 sg13g2_nand2_1 _7091_ (.Y(_2125_),
    .A(_2022_),
    .B(_1914_));
 sg13g2_nand3_1 _7092_ (.B(_1841_),
    .C(_2125_),
    .A(_2086_),
    .Y(_2126_));
 sg13g2_nand2_1 _7093_ (.Y(_2127_),
    .A(_2124_),
    .B(_2126_));
 sg13g2_nand2_1 _7094_ (.Y(_2128_),
    .A(_2127_),
    .B(_2063_));
 sg13g2_nand2_1 _7095_ (.Y(_2129_),
    .A(_2041_),
    .B(_2039_));
 sg13g2_nand3_1 _7096_ (.B(_2129_),
    .C(_2055_),
    .A(_2043_),
    .Y(_2130_));
 sg13g2_inv_1 _7097_ (.Y(_2131_),
    .A(_1727_));
 sg13g2_nor2_1 _7098_ (.A(net122),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_a22oi_1 _7099_ (.Y(_2133_),
    .B1(_2132_),
    .B2(_1914_),
    .A2(_2130_),
    .A1(net122));
 sg13g2_nand2_1 _7100_ (.Y(_2134_),
    .A(_2128_),
    .B(_2133_));
 sg13g2_nand2b_1 _7101_ (.Y(_2135_),
    .B(_2134_),
    .A_N(_2123_));
 sg13g2_xnor2_1 _7102_ (.Y(_2136_),
    .A(_1960_),
    .B(_2019_));
 sg13g2_nand2b_1 _7103_ (.Y(_2137_),
    .B(_2118_),
    .A_N(_2136_));
 sg13g2_nand2b_1 _7104_ (.Y(_2138_),
    .B(_1915_),
    .A_N(_1843_));
 sg13g2_nand2_1 _7105_ (.Y(_2139_),
    .A(_2137_),
    .B(_2138_));
 sg13g2_a21oi_1 _7106_ (.A1(_2136_),
    .A2(_1843_),
    .Y(_2140_),
    .B1(_2139_));
 sg13g2_a21oi_1 _7107_ (.A1(_2050_),
    .A2(_2028_),
    .Y(_2141_),
    .B1(_2056_));
 sg13g2_nand2b_1 _7108_ (.Y(_2142_),
    .B(_2141_),
    .A_N(_2051_));
 sg13g2_o21ai_1 _7109_ (.B1(_2142_),
    .Y(_2143_),
    .A1(net122),
    .A2(_2140_));
 sg13g2_nand2_1 _7110_ (.Y(_2144_),
    .A(_2078_),
    .B(_2063_));
 sg13g2_nand2_1 _7111_ (.Y(_2145_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_a21oi_1 _7112_ (.A1(_2145_),
    .A2(_2081_),
    .Y(_2146_),
    .B1(_2102_));
 sg13g2_nor2b_1 _7113_ (.A(_2034_),
    .B_N(_2049_),
    .Y(_2147_));
 sg13g2_nor2b_1 _7114_ (.A(_2047_),
    .B_N(_2147_),
    .Y(_2148_));
 sg13g2_o21ai_1 _7115_ (.B1(_2055_),
    .Y(_2149_),
    .A1(_2147_),
    .A2(_2048_));
 sg13g2_o21ai_1 _7116_ (.B1(_1492_),
    .Y(_2150_),
    .A1(_2148_),
    .A2(_2149_));
 sg13g2_o21ai_1 _7117_ (.B1(_2150_),
    .Y(_2151_),
    .A1(_2144_),
    .A2(_2146_));
 sg13g2_nand2b_1 _7118_ (.Y(_2152_),
    .B(_2151_),
    .A_N(_2143_));
 sg13g2_nor2_1 _7119_ (.A(_2135_),
    .B(_2152_),
    .Y(_2153_));
 sg13g2_nand4_1 _7120_ (.B(_2101_),
    .C(_2114_),
    .A(_2096_),
    .Y(_2154_),
    .D(_2153_));
 sg13g2_buf_2 _7121_ (.A(_2154_),
    .X(_2155_));
 sg13g2_inv_1 _7122_ (.Y(_2156_),
    .A(net124));
 sg13g2_nor2_1 _7123_ (.A(\i_music.i_sample.t3.genblk1[5].state.Q ),
    .B(_2156_),
    .Y(_2157_));
 sg13g2_inv_1 _7124_ (.Y(_2158_),
    .A(\i_music.i_sample.t2.genblk1[5].state.Q ));
 sg13g2_inv_1 _7125_ (.Y(_2159_),
    .A(\i_music.i_sample.t4.genblk1[5].state.Q ));
 sg13g2_a22oi_1 _7126_ (.Y(_2160_),
    .B1(_2159_),
    .B2(net129),
    .A2(_2158_),
    .A1(net130));
 sg13g2_nor2b_1 _7127_ (.A(_2157_),
    .B_N(_2160_),
    .Y(_2161_));
 sg13g2_buf_1 _7128_ (.A(_2161_),
    .X(_2162_));
 sg13g2_inv_1 _7129_ (.Y(_2163_),
    .A(_2162_));
 sg13g2_buf_1 _7130_ (.A(_2163_),
    .X(_2164_));
 sg13g2_nor2_1 _7131_ (.A(\i_music.i_sample.t4.genblk1[4].state.Q ),
    .B(net136),
    .Y(_2165_));
 sg13g2_inv_1 _7132_ (.Y(_2166_),
    .A(\i_music.i_sample.t2.genblk1[4].state.Q ));
 sg13g2_inv_1 _7133_ (.Y(_2167_),
    .A(\i_music.i_sample.t3.genblk1[4].state.Q ));
 sg13g2_a22oi_1 _7134_ (.Y(_2168_),
    .B1(_2167_),
    .B2(_1482_),
    .A2(_2166_),
    .A1(net130));
 sg13g2_nor2b_1 _7135_ (.A(_2165_),
    .B_N(_2168_),
    .Y(_2169_));
 sg13g2_buf_1 _7136_ (.A(_2169_),
    .X(_2170_));
 sg13g2_buf_1 _7137_ (.A(net57),
    .X(_2171_));
 sg13g2_buf_1 _7138_ (.A(net49),
    .X(_2172_));
 sg13g2_nor2_1 _7139_ (.A(\i_music.i_sample.t4.genblk1[2].state.Q ),
    .B(net136),
    .Y(_2173_));
 sg13g2_inv_1 _7140_ (.Y(_2174_),
    .A(\i_music.i_sample.t2.genblk1[2].state.Q ));
 sg13g2_inv_1 _7141_ (.Y(_2175_),
    .A(\i_music.i_sample.t3.genblk1[2].state.Q ));
 sg13g2_a22oi_1 _7142_ (.Y(_2176_),
    .B1(_2175_),
    .B2(net116),
    .A2(_2174_),
    .A1(net130));
 sg13g2_nor2b_1 _7143_ (.A(_2173_),
    .B_N(_2176_),
    .Y(_2177_));
 sg13g2_buf_1 _7144_ (.A(_2177_),
    .X(_2178_));
 sg13g2_inv_2 _7145_ (.Y(_2179_),
    .A(_2178_));
 sg13g2_a22oi_1 _7146_ (.Y(_2180_),
    .B1(\i_music.i_sample.t4.genblk1[1].state.Q ),
    .B2(net129),
    .A2(\i_music.i_sample.t3.genblk1[1].state.Q ),
    .A1(net116));
 sg13g2_inv_1 _7147_ (.Y(_2181_),
    .A(_2180_));
 sg13g2_a21oi_1 _7148_ (.A1(net130),
    .A2(\i_music.i_sample.t2.genblk1[1].state.Q ),
    .Y(_2182_),
    .B1(_2181_));
 sg13g2_buf_1 _7149_ (.A(_2182_),
    .X(_2183_));
 sg13g2_nor2_2 _7150_ (.A(_2179_),
    .B(net56),
    .Y(_2184_));
 sg13g2_nor2_1 _7151_ (.A(\i_music.i_sample.t4.genblk1[3].state.Q ),
    .B(net136),
    .Y(_2185_));
 sg13g2_inv_1 _7152_ (.Y(_2186_),
    .A(\i_music.i_sample.t2.genblk1[3].state.Q ));
 sg13g2_inv_1 _7153_ (.Y(_2187_),
    .A(\i_music.i_sample.t3.genblk1[3].state.Q ));
 sg13g2_a22oi_1 _7154_ (.Y(_2188_),
    .B1(_2187_),
    .B2(net116),
    .A2(_2186_),
    .A1(net130));
 sg13g2_nor2b_1 _7155_ (.A(_2185_),
    .B_N(_2188_),
    .Y(_2189_));
 sg13g2_buf_1 _7156_ (.A(_2189_),
    .X(_2190_));
 sg13g2_inv_1 _7157_ (.Y(_2191_),
    .A(net55));
 sg13g2_buf_1 _7158_ (.A(_2191_),
    .X(_2192_));
 sg13g2_nor2_1 _7159_ (.A(\i_music.i_sample.t3.genblk1[0].state.Q ),
    .B(_2156_),
    .Y(_2193_));
 sg13g2_inv_1 _7160_ (.Y(_2194_),
    .A(\i_music.i_sample.t2.genblk1[0].state.Q ));
 sg13g2_inv_1 _7161_ (.Y(_2195_),
    .A(\i_music.i_sample.t4.genblk1[0].state.Q ));
 sg13g2_a22oi_1 _7162_ (.Y(_2196_),
    .B1(_2195_),
    .B2(net129),
    .A2(_2194_),
    .A1(net130));
 sg13g2_nor2b_1 _7163_ (.A(_2193_),
    .B_N(_2196_),
    .Y(_2197_));
 sg13g2_buf_1 _7164_ (.A(_2197_),
    .X(_2198_));
 sg13g2_inv_2 _7165_ (.Y(_2199_),
    .A(net54));
 sg13g2_inv_1 _7166_ (.Y(_2200_),
    .A(net56));
 sg13g2_buf_1 _7167_ (.A(_2200_),
    .X(_2201_));
 sg13g2_nor2_1 _7168_ (.A(_2199_),
    .B(net37),
    .Y(_2202_));
 sg13g2_nor2_1 _7169_ (.A(_2192_),
    .B(_2202_),
    .Y(_2203_));
 sg13g2_inv_1 _7170_ (.Y(_2204_),
    .A(_2203_));
 sg13g2_nor2_1 _7171_ (.A(_2178_),
    .B(net54),
    .Y(_2205_));
 sg13g2_buf_1 _7172_ (.A(_2205_),
    .X(_2206_));
 sg13g2_nor2_1 _7173_ (.A(_2190_),
    .B(_2206_),
    .Y(_2207_));
 sg13g2_inv_1 _7174_ (.Y(_2208_),
    .A(_2207_));
 sg13g2_o21ai_1 _7175_ (.B1(_2208_),
    .Y(_2209_),
    .A1(_2184_),
    .A2(_2204_));
 sg13g2_buf_1 _7176_ (.A(_2178_),
    .X(_2210_));
 sg13g2_nor2_1 _7177_ (.A(net54),
    .B(_2200_),
    .Y(_2211_));
 sg13g2_inv_1 _7178_ (.Y(_2212_),
    .A(_2211_));
 sg13g2_nor2_2 _7179_ (.A(_2199_),
    .B(net56),
    .Y(_2213_));
 sg13g2_inv_1 _7180_ (.Y(_2214_),
    .A(_2213_));
 sg13g2_nand2_2 _7181_ (.Y(_2215_),
    .A(_2212_),
    .B(_2214_));
 sg13g2_nor2_1 _7182_ (.A(_2210_),
    .B(_2215_),
    .Y(_2216_));
 sg13g2_inv_1 _7183_ (.Y(_2217_),
    .A(_2215_));
 sg13g2_nor2_1 _7184_ (.A(_2179_),
    .B(_2217_),
    .Y(_2218_));
 sg13g2_inv_1 _7185_ (.Y(_2219_),
    .A(_2218_));
 sg13g2_buf_1 _7186_ (.A(net55),
    .X(_2220_));
 sg13g2_nand3b_1 _7187_ (.B(_2219_),
    .C(net47),
    .Y(_2221_),
    .A_N(_2216_));
 sg13g2_nor2_2 _7188_ (.A(net55),
    .B(net37),
    .Y(_2222_));
 sg13g2_inv_1 _7189_ (.Y(_2223_),
    .A(_2169_));
 sg13g2_buf_1 _7190_ (.A(_2223_),
    .X(_2224_));
 sg13g2_a21oi_1 _7191_ (.A1(_2222_),
    .A2(_2206_),
    .Y(_2225_),
    .B1(net46));
 sg13g2_nand2_1 _7192_ (.Y(_2226_),
    .A(_2221_),
    .B(_2225_));
 sg13g2_o21ai_1 _7193_ (.B1(_2226_),
    .Y(_2227_),
    .A1(_2172_),
    .A2(_2209_));
 sg13g2_nor2_1 _7194_ (.A(net48),
    .B(_2199_),
    .Y(_2228_));
 sg13g2_nand2_1 _7195_ (.Y(_2229_),
    .A(_2228_),
    .B(net56));
 sg13g2_nand2_1 _7196_ (.Y(_2230_),
    .A(_2229_),
    .B(net47));
 sg13g2_a21oi_1 _7197_ (.A1(_2219_),
    .A2(_2230_),
    .Y(_2231_),
    .B1(net49));
 sg13g2_nand2_1 _7198_ (.Y(_2232_),
    .A(_2217_),
    .B(net48));
 sg13g2_buf_1 _7199_ (.A(_2220_),
    .X(_2233_));
 sg13g2_inv_1 _7200_ (.Y(_2234_),
    .A(_2228_));
 sg13g2_nand4_1 _7201_ (.B(net57),
    .C(_2233_),
    .A(_2232_),
    .Y(_2235_),
    .D(_2234_));
 sg13g2_buf_1 _7202_ (.A(_2162_),
    .X(_2236_));
 sg13g2_nor2_2 _7203_ (.A(net48),
    .B(net37),
    .Y(_2237_));
 sg13g2_inv_1 _7204_ (.Y(_2238_),
    .A(_2237_));
 sg13g2_nor2_1 _7205_ (.A(net47),
    .B(_2238_),
    .Y(_2239_));
 sg13g2_nand3_1 _7206_ (.B(net57),
    .C(net54),
    .A(_2239_),
    .Y(_2240_));
 sg13g2_nand3_1 _7207_ (.B(net45),
    .C(_2240_),
    .A(_2235_),
    .Y(_2241_));
 sg13g2_nor2_1 _7208_ (.A(\i_music.i_sample.t3.genblk1[6].state.Q ),
    .B(_2156_),
    .Y(_2242_));
 sg13g2_inv_1 _7209_ (.Y(_2243_),
    .A(\i_music.i_sample.t2.genblk1[6].state.Q ));
 sg13g2_inv_1 _7210_ (.Y(_2244_),
    .A(\i_music.i_sample.t4.genblk1[6].state.Q ));
 sg13g2_a22oi_1 _7211_ (.Y(_2245_),
    .B1(_2244_),
    .B2(net129),
    .A2(_2243_),
    .A1(net130));
 sg13g2_nor2b_1 _7212_ (.A(_2242_),
    .B_N(_2245_),
    .Y(_2246_));
 sg13g2_buf_1 _7213_ (.A(_2246_),
    .X(_2247_));
 sg13g2_nor2_1 _7214_ (.A(\i_music.i_sample.t3.genblk1[7].state.Q ),
    .B(_2156_),
    .Y(_2248_));
 sg13g2_inv_1 _7215_ (.Y(_2249_),
    .A(\i_music.i_sample.t2.genblk1[7].state.Q ));
 sg13g2_inv_1 _7216_ (.Y(_2250_),
    .A(\i_music.i_sample.t4.genblk1[7].state.Q ));
 sg13g2_a22oi_1 _7217_ (.Y(_2251_),
    .B1(_2250_),
    .B2(net129),
    .A2(_2249_),
    .A1(net130));
 sg13g2_nor2b_1 _7218_ (.A(_2248_),
    .B_N(_2251_),
    .Y(_2252_));
 sg13g2_buf_2 _7219_ (.A(_2252_),
    .X(_2253_));
 sg13g2_inv_2 _7220_ (.Y(_2254_),
    .A(_2253_));
 sg13g2_nor2_1 _7221_ (.A(net53),
    .B(_2254_),
    .Y(_2255_));
 sg13g2_o21ai_1 _7222_ (.B1(_2255_),
    .Y(_2256_),
    .A1(_2231_),
    .A2(_2241_));
 sg13g2_a21oi_1 _7223_ (.A1(_2164_),
    .A2(_2227_),
    .Y(_2257_),
    .B1(_2256_));
 sg13g2_buf_1 _7224_ (.A(_2224_),
    .X(_2258_));
 sg13g2_nor2_1 _7225_ (.A(net38),
    .B(_2183_),
    .Y(_2259_));
 sg13g2_nor2_1 _7226_ (.A(_2259_),
    .B(_2222_),
    .Y(_2260_));
 sg13g2_nand2_1 _7227_ (.Y(_2261_),
    .A(_2201_),
    .B(_2199_));
 sg13g2_buf_1 _7228_ (.A(net38),
    .X(_2262_));
 sg13g2_nand3_1 _7229_ (.B(_2261_),
    .C(_2262_),
    .A(_2238_),
    .Y(_2263_));
 sg13g2_o21ai_1 _7230_ (.B1(_2263_),
    .Y(_2264_),
    .A1(net54),
    .A2(_2260_));
 sg13g2_nor2_1 _7231_ (.A(_2179_),
    .B(_2200_),
    .Y(_2265_));
 sg13g2_buf_2 _7232_ (.A(_2265_),
    .X(_2266_));
 sg13g2_nor2_2 _7233_ (.A(_2210_),
    .B(net56),
    .Y(_2267_));
 sg13g2_nor2_2 _7234_ (.A(_2267_),
    .B(_2266_),
    .Y(_2268_));
 sg13g2_a22oi_1 _7235_ (.Y(_2269_),
    .B1(net54),
    .B2(_2268_),
    .A2(_2266_),
    .A1(_2262_));
 sg13g2_nor2_1 _7236_ (.A(net46),
    .B(_2269_),
    .Y(_2270_));
 sg13g2_a21oi_1 _7237_ (.A1(net35),
    .A2(_2264_),
    .Y(_2271_),
    .B1(_2270_));
 sg13g2_inv_1 _7238_ (.Y(_2272_),
    .A(_2247_));
 sg13g2_nor2_1 _7239_ (.A(_2254_),
    .B(net44),
    .Y(_2273_));
 sg13g2_o21ai_1 _7240_ (.B1(_2273_),
    .Y(_2274_),
    .A1(_2236_),
    .A2(_2271_));
 sg13g2_nor2_1 _7241_ (.A(net54),
    .B(_2179_),
    .Y(_2275_));
 sg13g2_nor2_1 _7242_ (.A(net48),
    .B(_2217_),
    .Y(_2276_));
 sg13g2_nor3_1 _7243_ (.A(_2220_),
    .B(_2275_),
    .C(_2276_),
    .Y(_2277_));
 sg13g2_nor2_1 _7244_ (.A(net38),
    .B(net37),
    .Y(_2278_));
 sg13g2_nor2_1 _7245_ (.A(net38),
    .B(_2179_),
    .Y(_2279_));
 sg13g2_inv_1 _7246_ (.Y(_2280_),
    .A(_2279_));
 sg13g2_nand2_1 _7247_ (.Y(_2281_),
    .A(_2280_),
    .B(_2223_));
 sg13g2_nor2_1 _7248_ (.A(_2278_),
    .B(_2281_),
    .Y(_2282_));
 sg13g2_nor2b_1 _7249_ (.A(_2277_),
    .B_N(_2282_),
    .Y(_2283_));
 sg13g2_nor4_1 _7250_ (.A(net33),
    .B(_2206_),
    .C(_2213_),
    .D(_2266_),
    .Y(_2284_));
 sg13g2_nor3_1 _7251_ (.A(net36),
    .B(_2216_),
    .C(_2218_),
    .Y(_2285_));
 sg13g2_nor3_1 _7252_ (.A(net35),
    .B(_2284_),
    .C(_2285_),
    .Y(_2286_));
 sg13g2_nor3_1 _7253_ (.A(net40),
    .B(_2283_),
    .C(_2286_),
    .Y(_2287_));
 sg13g2_nor2_1 _7254_ (.A(_2274_),
    .B(_2287_),
    .Y(_2288_));
 sg13g2_nor2_1 _7255_ (.A(_2179_),
    .B(_2199_),
    .Y(_2289_));
 sg13g2_buf_1 _7256_ (.A(_2289_),
    .X(_2290_));
 sg13g2_nor2_1 _7257_ (.A(_2206_),
    .B(_2290_),
    .Y(_2291_));
 sg13g2_inv_1 _7258_ (.Y(_2292_),
    .A(_2291_));
 sg13g2_nor2_1 _7259_ (.A(net55),
    .B(_2213_),
    .Y(_2293_));
 sg13g2_inv_1 _7260_ (.Y(_2294_),
    .A(_2293_));
 sg13g2_inv_1 _7261_ (.Y(_2295_),
    .A(_2268_));
 sg13g2_nor2_1 _7262_ (.A(_2294_),
    .B(_2295_),
    .Y(_2296_));
 sg13g2_a21oi_1 _7263_ (.A1(_2203_),
    .A2(_2292_),
    .Y(_2297_),
    .B1(_2296_));
 sg13g2_a21oi_1 _7264_ (.A1(_2297_),
    .A2(_2224_),
    .Y(_2298_),
    .B1(_2162_));
 sg13g2_inv_1 _7265_ (.Y(_2299_),
    .A(_2184_));
 sg13g2_nand2_1 _7266_ (.Y(_2300_),
    .A(_2299_),
    .B(net55));
 sg13g2_inv_1 _7267_ (.Y(_2301_),
    .A(_2300_));
 sg13g2_inv_1 _7268_ (.Y(_2302_),
    .A(_2275_));
 sg13g2_nor2_1 _7269_ (.A(net55),
    .B(_2199_),
    .Y(_2303_));
 sg13g2_a21oi_1 _7270_ (.A1(_2301_),
    .A2(_2302_),
    .Y(_2304_),
    .B1(_2303_));
 sg13g2_nor2_2 _7271_ (.A(net55),
    .B(_2184_),
    .Y(_2305_));
 sg13g2_nand2_1 _7272_ (.Y(_2306_),
    .A(_2305_),
    .B(_2238_));
 sg13g2_nand3_1 _7273_ (.B(net57),
    .C(_2306_),
    .A(_2304_),
    .Y(_2307_));
 sg13g2_nand2_1 _7274_ (.Y(_2308_),
    .A(_2212_),
    .B(_2234_));
 sg13g2_o21ai_1 _7275_ (.B1(_2308_),
    .Y(_2309_),
    .A1(net37),
    .A2(_2208_));
 sg13g2_nand2_1 _7276_ (.Y(_2310_),
    .A(_2305_),
    .B(_2302_));
 sg13g2_nor2_1 _7277_ (.A(net38),
    .B(_2213_),
    .Y(_2311_));
 sg13g2_a21oi_1 _7278_ (.A1(_2268_),
    .A2(_2311_),
    .Y(_2312_),
    .B1(net46));
 sg13g2_o21ai_1 _7279_ (.B1(_2312_),
    .Y(_2313_),
    .A1(_2310_),
    .A2(_2216_));
 sg13g2_o21ai_1 _7280_ (.B1(_2313_),
    .Y(_2314_),
    .A1(net49),
    .A2(_2309_));
 sg13g2_a221oi_1 _7281_ (.B2(net45),
    .C1(net44),
    .B1(_2314_),
    .A1(_2298_),
    .Y(_2315_),
    .A2(_2307_));
 sg13g2_nand2_1 _7282_ (.Y(_2316_),
    .A(_2223_),
    .B(_2179_));
 sg13g2_nand2_1 _7283_ (.Y(_2317_),
    .A(net46),
    .B(net38));
 sg13g2_o21ai_1 _7284_ (.B1(_2317_),
    .Y(_2318_),
    .A1(_2316_),
    .A2(_2212_));
 sg13g2_nor3_1 _7285_ (.A(net57),
    .B(_2199_),
    .C(_2237_),
    .Y(_2319_));
 sg13g2_o21ai_1 _7286_ (.B1(net33),
    .Y(_2320_),
    .A1(_2275_),
    .A2(_2215_));
 sg13g2_o21ai_1 _7287_ (.B1(_2320_),
    .Y(_2321_),
    .A1(_2318_),
    .A2(_2319_));
 sg13g2_nor2b_1 _7288_ (.A(_2299_),
    .B_N(_2303_),
    .Y(_2322_));
 sg13g2_a21oi_1 _7289_ (.A1(_2301_),
    .A2(_2261_),
    .Y(_2323_),
    .B1(_2322_));
 sg13g2_a21oi_1 _7290_ (.A1(_2323_),
    .A2(_2171_),
    .Y(_2324_),
    .B1(net45));
 sg13g2_a21oi_1 _7291_ (.A1(net47),
    .A2(_2211_),
    .Y(_2325_),
    .B1(_2277_));
 sg13g2_o21ai_1 _7292_ (.B1(_2306_),
    .Y(_2326_),
    .A1(net54),
    .A2(_2266_));
 sg13g2_nand2_1 _7293_ (.Y(_2327_),
    .A(_2326_),
    .B(_2170_));
 sg13g2_o21ai_1 _7294_ (.B1(_2327_),
    .Y(_2328_),
    .A1(net49),
    .A2(_2325_));
 sg13g2_a221oi_1 _7295_ (.B2(net45),
    .C1(net53),
    .B1(_2328_),
    .A1(_2321_),
    .Y(_2329_),
    .A2(_2324_));
 sg13g2_nor3_1 _7296_ (.A(_2253_),
    .B(_2315_),
    .C(_2329_),
    .Y(_2330_));
 sg13g2_nor3_1 _7297_ (.A(_2257_),
    .B(_2288_),
    .C(_2330_),
    .Y(_2331_));
 sg13g2_nand2_1 _7298_ (.Y(_2332_),
    .A(_2155_),
    .B(_2331_));
 sg13g2_nor2_1 _7299_ (.A(_1668_),
    .B(_2332_),
    .Y(_2333_));
 sg13g2_inv_1 _7300_ (.Y(_2334_),
    .A(_2333_));
 sg13g2_nor2_1 _7301_ (.A(_2294_),
    .B(_2308_),
    .Y(_2335_));
 sg13g2_inv_1 _7302_ (.Y(_2336_),
    .A(_2335_));
 sg13g2_a21oi_1 _7303_ (.A1(_2292_),
    .A2(_2278_),
    .Y(_2337_),
    .B1(net46));
 sg13g2_a21oi_1 _7304_ (.A1(_2311_),
    .A2(_2302_),
    .Y(_2338_),
    .B1(_2171_));
 sg13g2_a22oi_1 _7305_ (.Y(_2339_),
    .B1(_2338_),
    .B2(_2320_),
    .A2(_2337_),
    .A1(_2336_));
 sg13g2_inv_1 _7306_ (.Y(_2340_),
    .A(_2266_));
 sg13g2_inv_1 _7307_ (.Y(_2341_),
    .A(_2290_));
 sg13g2_nand2_1 _7308_ (.Y(_2342_),
    .A(_2340_),
    .B(_2341_));
 sg13g2_o21ai_1 _7309_ (.B1(net36),
    .Y(_2343_),
    .A1(_2342_),
    .A2(_2216_));
 sg13g2_inv_1 _7310_ (.Y(_2344_),
    .A(_2267_));
 sg13g2_nand3_1 _7311_ (.B(net33),
    .C(_2302_),
    .A(_2344_),
    .Y(_2345_));
 sg13g2_nand3_1 _7312_ (.B(net49),
    .C(_2345_),
    .A(_2343_),
    .Y(_2346_));
 sg13g2_nor2_1 _7313_ (.A(net48),
    .B(_2213_),
    .Y(_2347_));
 sg13g2_inv_1 _7314_ (.Y(_2348_),
    .A(_2347_));
 sg13g2_a21oi_1 _7315_ (.A1(_2348_),
    .A2(_2299_),
    .Y(_2349_),
    .B1(net47));
 sg13g2_nor2_1 _7316_ (.A(net49),
    .B(_2349_),
    .Y(_2350_));
 sg13g2_o21ai_1 _7317_ (.B1(net36),
    .Y(_2351_),
    .A1(_2275_),
    .A2(_2215_));
 sg13g2_a21oi_1 _7318_ (.A1(_2350_),
    .A2(_2351_),
    .Y(_2352_),
    .B1(net40));
 sg13g2_a221oi_1 _7319_ (.B2(_2352_),
    .C1(_2254_),
    .B1(_2346_),
    .A1(_2339_),
    .Y(_2353_),
    .A2(net40));
 sg13g2_a221oi_1 _7320_ (.B2(_2233_),
    .C1(_2162_),
    .B1(_2291_),
    .A1(_2207_),
    .Y(_2354_),
    .A2(net56));
 sg13g2_inv_1 _7321_ (.Y(_2355_),
    .A(_2222_));
 sg13g2_o21ai_1 _7322_ (.B1(_2162_),
    .Y(_2356_),
    .A1(_2290_),
    .A2(_2260_));
 sg13g2_a21oi_1 _7323_ (.A1(_2292_),
    .A2(_2355_),
    .Y(_2357_),
    .B1(_2356_));
 sg13g2_nor3_1 _7324_ (.A(net49),
    .B(_2354_),
    .C(_2357_),
    .Y(_2358_));
 sg13g2_nor2_1 _7325_ (.A(net33),
    .B(_2302_),
    .Y(_2359_));
 sg13g2_a21o_1 _7326_ (.A2(_2163_),
    .A1(_2301_),
    .B1(_2222_),
    .X(_2360_));
 sg13g2_a22oi_1 _7327_ (.Y(_2361_),
    .B1(_2234_),
    .B2(_2360_),
    .A2(_2359_),
    .A1(_2162_));
 sg13g2_o21ai_1 _7328_ (.B1(_2254_),
    .Y(_2362_),
    .A1(net35),
    .A2(_2361_));
 sg13g2_o21ai_1 _7329_ (.B1(_2247_),
    .Y(_2363_),
    .A1(_2358_),
    .A2(_2362_));
 sg13g2_nor2_1 _7330_ (.A(net56),
    .B(_2290_),
    .Y(_2364_));
 sg13g2_inv_1 _7331_ (.Y(_2365_),
    .A(_2364_));
 sg13g2_a21oi_1 _7332_ (.A1(_2203_),
    .A2(_2365_),
    .Y(_2366_),
    .B1(_2349_));
 sg13g2_nand2_1 _7333_ (.Y(_2367_),
    .A(_2366_),
    .B(_2170_));
 sg13g2_o21ai_1 _7334_ (.B1(_2282_),
    .Y(_2368_),
    .A1(_2208_),
    .A2(_2365_));
 sg13g2_nand3_1 _7335_ (.B(net45),
    .C(_2368_),
    .A(_2367_),
    .Y(_2369_));
 sg13g2_nor2_1 _7336_ (.A(net55),
    .B(net48),
    .Y(_2370_));
 sg13g2_nor2_1 _7337_ (.A(_2370_),
    .B(_2293_),
    .Y(_2371_));
 sg13g2_o21ai_1 _7338_ (.B1(net47),
    .Y(_2372_),
    .A1(net56),
    .A2(_2292_));
 sg13g2_o21ai_1 _7339_ (.B1(_2372_),
    .Y(_2373_),
    .A1(_2267_),
    .A2(_2371_));
 sg13g2_o21ai_1 _7340_ (.B1(_2223_),
    .Y(_2374_),
    .A1(net38),
    .A2(net37));
 sg13g2_nor3_1 _7341_ (.A(_2267_),
    .B(_2303_),
    .C(_2374_),
    .Y(_2375_));
 sg13g2_nor2_1 _7342_ (.A(_2162_),
    .B(_2375_),
    .Y(_2376_));
 sg13g2_o21ai_1 _7343_ (.B1(_2376_),
    .Y(_2377_),
    .A1(net46),
    .A2(_2373_));
 sg13g2_a21oi_1 _7344_ (.A1(_2369_),
    .A2(_2377_),
    .Y(_2378_),
    .B1(_2253_));
 sg13g2_nor2_1 _7345_ (.A(net47),
    .B(_2211_),
    .Y(_2379_));
 sg13g2_nor2_1 _7346_ (.A(_2192_),
    .B(_2341_),
    .Y(_2380_));
 sg13g2_o21ai_1 _7347_ (.B1(net38),
    .Y(_2381_),
    .A1(net37),
    .A2(_2341_));
 sg13g2_nand3b_1 _7348_ (.B(_2381_),
    .C(net57),
    .Y(_2382_),
    .A_N(_2380_));
 sg13g2_o21ai_1 _7349_ (.B1(_2382_),
    .Y(_2383_),
    .A1(_2379_),
    .A2(_2374_));
 sg13g2_a22oi_1 _7350_ (.Y(_2384_),
    .B1(_2341_),
    .B2(_2379_),
    .A2(_2344_),
    .A1(_2203_));
 sg13g2_nand2b_1 _7351_ (.Y(_2385_),
    .B(net35),
    .A_N(_2384_));
 sg13g2_nor2_1 _7352_ (.A(net46),
    .B(_2207_),
    .Y(_2386_));
 sg13g2_a21oi_1 _7353_ (.A1(_2386_),
    .A2(_2365_),
    .Y(_2387_),
    .B1(_2163_));
 sg13g2_a221oi_1 _7354_ (.B2(_2387_),
    .C1(_2254_),
    .B1(_2385_),
    .A1(_2383_),
    .Y(_2388_),
    .A2(_2163_));
 sg13g2_o21ai_1 _7355_ (.B1(net44),
    .Y(_2389_),
    .A1(_2378_),
    .A2(_2388_));
 sg13g2_o21ai_1 _7356_ (.B1(_2389_),
    .Y(_2390_),
    .A1(_2353_),
    .A2(_2363_));
 sg13g2_nand2b_1 _7357_ (.Y(_2391_),
    .B(_2155_),
    .A_N(_2390_));
 sg13g2_xor2_1 _7358_ (.B(_2391_),
    .A(\i_music.i_sample.sample_acc[1] ),
    .X(_2392_));
 sg13g2_xnor2_1 _7359_ (.Y(_2393_),
    .A(_2334_),
    .B(_2392_));
 sg13g2_nor2_1 _7360_ (.A(net147),
    .B(net136),
    .Y(_2394_));
 sg13g2_buf_1 _7361_ (.A(_2394_),
    .X(_2395_));
 sg13g2_buf_1 _7362_ (.A(_2395_),
    .X(_2396_));
 sg13g2_nor2_1 _7363_ (.A(\i_music.i_pwm.sample[0] ),
    .B(net113),
    .Y(_2397_));
 sg13g2_a21oi_1 _7364_ (.A1(_2393_),
    .A2(net113),
    .Y(_0197_),
    .B1(_2397_));
 sg13g2_inv_1 _7365_ (.Y(_2398_),
    .A(\i_music.i_sample.sample_acc[2] ));
 sg13g2_inv_1 _7366_ (.Y(_2399_),
    .A(_2305_));
 sg13g2_nor2_1 _7367_ (.A(_2290_),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_nor2_1 _7368_ (.A(_2266_),
    .B(_2230_),
    .Y(_2401_));
 sg13g2_o21ai_1 _7369_ (.B1(net39),
    .Y(_2402_),
    .A1(_2400_),
    .A2(_2401_));
 sg13g2_inv_1 _7370_ (.Y(_2403_),
    .A(_2281_));
 sg13g2_o21ai_1 _7371_ (.B1(_2403_),
    .Y(_2404_),
    .A1(net36),
    .A2(_2344_));
 sg13g2_nand3_1 _7372_ (.B(net40),
    .C(_2404_),
    .A(_2402_),
    .Y(_2405_));
 sg13g2_nor2_1 _7373_ (.A(net57),
    .B(_2370_),
    .Y(_2406_));
 sg13g2_nand2_1 _7374_ (.Y(_2407_),
    .A(_2179_),
    .B(net47));
 sg13g2_nand2_1 _7375_ (.Y(_2408_),
    .A(_2407_),
    .B(net57));
 sg13g2_nor2_1 _7376_ (.A(net33),
    .B(_2214_),
    .Y(_2409_));
 sg13g2_o21ai_1 _7377_ (.B1(net45),
    .Y(_2410_),
    .A1(_2408_),
    .A2(_2409_));
 sg13g2_a21o_1 _7378_ (.A2(_2406_),
    .A1(net37),
    .B1(_2410_),
    .X(_2411_));
 sg13g2_and3_1 _7379_ (.X(_2412_),
    .A(_2405_),
    .B(net44),
    .C(_2411_));
 sg13g2_nor2_1 _7380_ (.A(_2407_),
    .B(_2213_),
    .Y(_2413_));
 sg13g2_inv_1 _7381_ (.Y(_2414_),
    .A(_2413_));
 sg13g2_nand2_1 _7382_ (.Y(_2415_),
    .A(_2336_),
    .B(_2414_));
 sg13g2_nand2_1 _7383_ (.Y(_2416_),
    .A(_2415_),
    .B(net39));
 sg13g2_inv_1 _7384_ (.Y(_2417_),
    .A(_2406_));
 sg13g2_nor2_1 _7385_ (.A(_2222_),
    .B(_2417_),
    .Y(_2418_));
 sg13g2_inv_1 _7386_ (.Y(_2419_),
    .A(_2259_));
 sg13g2_nor2_1 _7387_ (.A(_2228_),
    .B(_2419_),
    .Y(_2420_));
 sg13g2_inv_1 _7388_ (.Y(_2421_),
    .A(_2420_));
 sg13g2_a21oi_1 _7389_ (.A1(_2418_),
    .A2(_2421_),
    .Y(_2422_),
    .B1(net40));
 sg13g2_nor2_1 _7390_ (.A(_2317_),
    .B(_2232_),
    .Y(_2423_));
 sg13g2_nor3_1 _7391_ (.A(net39),
    .B(_2206_),
    .C(_2300_),
    .Y(_2424_));
 sg13g2_nand3_1 _7392_ (.B(net36),
    .C(_2234_),
    .A(_2212_),
    .Y(_2425_));
 sg13g2_nor2_1 _7393_ (.A(net46),
    .B(_2239_),
    .Y(_2426_));
 sg13g2_inv_1 _7394_ (.Y(_2427_),
    .A(_2426_));
 sg13g2_a21oi_1 _7395_ (.A1(_2425_),
    .A2(_2381_),
    .Y(_2428_),
    .B1(_2427_));
 sg13g2_nor3_1 _7396_ (.A(_2423_),
    .B(_2424_),
    .C(_2428_),
    .Y(_2429_));
 sg13g2_a221oi_1 _7397_ (.B2(net40),
    .C1(net44),
    .B1(_2429_),
    .A1(_2416_),
    .Y(_2430_),
    .A2(_2422_));
 sg13g2_o21ai_1 _7398_ (.B1(_2253_),
    .Y(_2431_),
    .A1(_2412_),
    .A2(_2430_));
 sg13g2_nor3_1 _7399_ (.A(_2258_),
    .B(_2420_),
    .C(_2296_),
    .Y(_2432_));
 sg13g2_nor3_1 _7400_ (.A(_2290_),
    .B(_2237_),
    .C(_2208_),
    .Y(_2433_));
 sg13g2_nor3_1 _7401_ (.A(_2172_),
    .B(_2433_),
    .C(_2284_),
    .Y(_2434_));
 sg13g2_nor3_1 _7402_ (.A(net45),
    .B(_2432_),
    .C(_2434_),
    .Y(_2435_));
 sg13g2_a21oi_1 _7403_ (.A1(_2311_),
    .A2(_2340_),
    .Y(_2436_),
    .B1(_2417_));
 sg13g2_nor2_1 _7404_ (.A(_2237_),
    .B(_2371_),
    .Y(_2437_));
 sg13g2_inv_1 _7405_ (.Y(_2438_),
    .A(_2437_));
 sg13g2_nand3_1 _7406_ (.B(net36),
    .C(_2302_),
    .A(_2229_),
    .Y(_2439_));
 sg13g2_a21oi_1 _7407_ (.A1(_2438_),
    .A2(_2439_),
    .Y(_2440_),
    .B1(net35));
 sg13g2_o21ai_1 _7408_ (.B1(net45),
    .Y(_2441_),
    .A1(_2436_),
    .A2(_2440_));
 sg13g2_nand2b_1 _7409_ (.Y(_2442_),
    .B(_2441_),
    .A_N(_2435_));
 sg13g2_nand2_1 _7410_ (.Y(_2443_),
    .A(_2303_),
    .B(net48));
 sg13g2_nor2_1 _7411_ (.A(net35),
    .B(_2359_),
    .Y(_2444_));
 sg13g2_o21ai_1 _7412_ (.B1(_2212_),
    .Y(_2445_),
    .A1(_2380_),
    .A2(_2437_));
 sg13g2_a22oi_1 _7413_ (.Y(_2446_),
    .B1(net35),
    .B2(_2445_),
    .A2(_2444_),
    .A1(_2443_));
 sg13g2_nor2_1 _7414_ (.A(_2407_),
    .B(_2211_),
    .Y(_2447_));
 sg13g2_nor2_1 _7415_ (.A(_2399_),
    .B(_2217_),
    .Y(_2448_));
 sg13g2_nor3_1 _7416_ (.A(net49),
    .B(_2447_),
    .C(_2448_),
    .Y(_2449_));
 sg13g2_nor2_1 _7417_ (.A(net33),
    .B(_2215_),
    .Y(_2450_));
 sg13g2_inv_1 _7418_ (.Y(_2451_),
    .A(_2450_));
 sg13g2_a21oi_1 _7419_ (.A1(_2451_),
    .A2(net48),
    .Y(_2452_),
    .B1(_2408_));
 sg13g2_nor2_1 _7420_ (.A(_2449_),
    .B(_2452_),
    .Y(_2453_));
 sg13g2_nor2_1 _7421_ (.A(net40),
    .B(_2453_),
    .Y(_2454_));
 sg13g2_a21oi_1 _7422_ (.A1(_2446_),
    .A2(net40),
    .Y(_2455_),
    .B1(_2454_));
 sg13g2_a21oi_1 _7423_ (.A1(_2455_),
    .A2(net53),
    .Y(_2456_),
    .B1(_2253_));
 sg13g2_o21ai_1 _7424_ (.B1(_2456_),
    .Y(_2457_),
    .A1(net53),
    .A2(_2442_));
 sg13g2_nand3_1 _7425_ (.B(_2431_),
    .C(_2457_),
    .A(_2155_),
    .Y(_2458_));
 sg13g2_xnor2_1 _7426_ (.Y(_2459_),
    .A(_2398_),
    .B(_2458_));
 sg13g2_nand2b_1 _7427_ (.Y(_2460_),
    .B(\i_music.i_sample.sample_acc[1] ),
    .A_N(_2391_));
 sg13g2_o21ai_1 _7428_ (.B1(_2460_),
    .Y(_2461_),
    .A1(_2334_),
    .A2(_2392_));
 sg13g2_xor2_1 _7429_ (.B(_2461_),
    .A(_2459_),
    .X(_2462_));
 sg13g2_nor2_1 _7430_ (.A(\i_music.i_pwm.sample[1] ),
    .B(net113),
    .Y(_2463_));
 sg13g2_a21oi_1 _7431_ (.A1(_2462_),
    .A2(net113),
    .Y(_0198_),
    .B1(_2463_));
 sg13g2_buf_1 _7432_ (.A(net39),
    .X(_2464_));
 sg13g2_nand2_1 _7433_ (.Y(_2465_),
    .A(_2348_),
    .B(net36));
 sg13g2_inv_1 _7434_ (.Y(_2466_),
    .A(_2465_));
 sg13g2_nor2_1 _7435_ (.A(_2464_),
    .B(_2466_),
    .Y(_2467_));
 sg13g2_buf_1 _7436_ (.A(net35),
    .X(_2468_));
 sg13g2_a21oi_1 _7437_ (.A1(_2263_),
    .A2(_2204_),
    .Y(_2469_),
    .B1(_2468_));
 sg13g2_buf_1 _7438_ (.A(_2164_),
    .X(_2470_));
 sg13g2_a21oi_2 _7439_ (.B1(net30),
    .Y(_2471_),
    .A2(_2468_),
    .A1(_2305_));
 sg13g2_o21ai_1 _7440_ (.B1(_2471_),
    .Y(_2472_),
    .A1(_2467_),
    .A2(_2469_));
 sg13g2_nand2_1 _7441_ (.Y(_2473_),
    .A(_2278_),
    .B(_2198_));
 sg13g2_nand2_1 _7442_ (.Y(_2474_),
    .A(_2295_),
    .B(_2473_));
 sg13g2_buf_1 _7443_ (.A(_2236_),
    .X(_2475_));
 sg13g2_a221oi_1 _7444_ (.B2(net32),
    .C1(net34),
    .B1(_2474_),
    .A1(_2268_),
    .Y(_2476_),
    .A2(_2294_));
 sg13g2_nor2_1 _7445_ (.A(net44),
    .B(_2476_),
    .Y(_2477_));
 sg13g2_nand2_1 _7446_ (.Y(_2478_),
    .A(_2280_),
    .B(net32));
 sg13g2_a21oi_1 _7447_ (.A1(_2268_),
    .A2(_2406_),
    .Y(_2479_),
    .B1(net30));
 sg13g2_inv_1 _7448_ (.Y(_2480_),
    .A(_2239_));
 sg13g2_o21ai_1 _7449_ (.B1(net39),
    .Y(_2481_),
    .A1(_2447_),
    .A2(_2400_));
 sg13g2_o21ai_1 _7450_ (.B1(_2481_),
    .Y(_2482_),
    .A1(net32),
    .A2(_2480_));
 sg13g2_a22oi_1 _7451_ (.Y(_2483_),
    .B1(net30),
    .B2(_2482_),
    .A2(_2479_),
    .A1(_2478_));
 sg13g2_a221oi_1 _7452_ (.B2(net44),
    .C1(_2254_),
    .B1(_2483_),
    .A1(_2472_),
    .Y(_2484_),
    .A2(_2477_));
 sg13g2_nand3_1 _7453_ (.B(_2340_),
    .C(net33),
    .A(_2365_),
    .Y(_2485_));
 sg13g2_a21oi_1 _7454_ (.A1(_2485_),
    .A2(_2414_),
    .Y(_2486_),
    .B1(_2258_));
 sg13g2_a221oi_1 _7455_ (.B2(_2403_),
    .C1(_2486_),
    .B1(_2199_),
    .A1(net31),
    .Y(_2487_),
    .A2(_2266_));
 sg13g2_nand2b_1 _7456_ (.Y(_2488_),
    .B(net30),
    .A_N(_2487_));
 sg13g2_o21ai_1 _7457_ (.B1(_2438_),
    .Y(_2489_),
    .A1(_2300_),
    .A2(_2276_));
 sg13g2_nand2_1 _7458_ (.Y(_2490_),
    .A(_2489_),
    .B(net39));
 sg13g2_o21ai_1 _7459_ (.B1(_2490_),
    .Y(_2491_),
    .A1(net32),
    .A2(_2409_));
 sg13g2_a21oi_1 _7460_ (.A1(_2491_),
    .A2(net34),
    .Y(_2492_),
    .B1(net53));
 sg13g2_a22oi_1 _7461_ (.Y(_2493_),
    .B1(_2207_),
    .B2(_2238_),
    .A2(_2206_),
    .A1(_2278_));
 sg13g2_nor2_1 _7462_ (.A(_2341_),
    .B(_2419_),
    .Y(_2494_));
 sg13g2_nand2_1 _7463_ (.Y(_2495_),
    .A(_2494_),
    .B(net39));
 sg13g2_o21ai_1 _7464_ (.B1(_2495_),
    .Y(_2496_),
    .A1(_2464_),
    .A2(_2493_));
 sg13g2_a21oi_1 _7465_ (.A1(net33),
    .A2(_2184_),
    .Y(_2497_),
    .B1(_2450_));
 sg13g2_nor2_1 _7466_ (.A(net39),
    .B(_2400_),
    .Y(_2498_));
 sg13g2_a221oi_1 _7467_ (.B2(_2498_),
    .C1(net34),
    .B1(_2221_),
    .A1(net32),
    .Y(_2499_),
    .A2(_2497_));
 sg13g2_a21oi_1 _7468_ (.A1(net34),
    .A2(_2496_),
    .Y(_2500_),
    .B1(_2499_));
 sg13g2_a221oi_1 _7469_ (.B2(net53),
    .C1(_2253_),
    .B1(_2500_),
    .A1(_2488_),
    .Y(_2501_),
    .A2(_2492_));
 sg13g2_nor2_1 _7470_ (.A(_2484_),
    .B(_2501_),
    .Y(_2502_));
 sg13g2_nand2_1 _7471_ (.Y(_2503_),
    .A(_2155_),
    .B(_2502_));
 sg13g2_xnor2_1 _7472_ (.Y(_2504_),
    .A(\i_music.i_sample.sample_acc[3] ),
    .B(_2503_));
 sg13g2_nand2b_1 _7473_ (.Y(_2505_),
    .B(_2461_),
    .A_N(_2459_));
 sg13g2_o21ai_1 _7474_ (.B1(_2505_),
    .Y(_2506_),
    .A1(_2398_),
    .A2(_2458_));
 sg13g2_xnor2_1 _7475_ (.Y(_2507_),
    .A(_2504_),
    .B(_2506_));
 sg13g2_nor2_1 _7476_ (.A(\i_music.i_pwm.sample[2] ),
    .B(_2395_),
    .Y(_2508_));
 sg13g2_a21oi_1 _7477_ (.A1(_2507_),
    .A2(net113),
    .Y(_0199_),
    .B1(_2508_));
 sg13g2_nor2_1 _7478_ (.A(net31),
    .B(_2305_),
    .Y(_2509_));
 sg13g2_nand3_1 _7479_ (.B(_2421_),
    .C(_2473_),
    .A(_2509_),
    .Y(_2510_));
 sg13g2_o21ai_1 _7480_ (.B1(net31),
    .Y(_2511_),
    .A1(_2322_),
    .A2(_2301_));
 sg13g2_nand2_1 _7481_ (.Y(_2512_),
    .A(_2419_),
    .B(_2280_));
 sg13g2_nand2b_1 _7482_ (.Y(_2513_),
    .B(_2426_),
    .A_N(_2512_));
 sg13g2_a21oi_1 _7483_ (.A1(_2511_),
    .A2(_2513_),
    .Y(_2514_),
    .B1(net34));
 sg13g2_a21o_1 _7484_ (.A2(_2510_),
    .A1(_2471_),
    .B1(_2514_),
    .X(_2515_));
 sg13g2_o21ai_1 _7485_ (.B1(net53),
    .Y(_2516_),
    .A1(_2470_),
    .A2(_2318_));
 sg13g2_nand2_1 _7486_ (.Y(_2517_),
    .A(_2237_),
    .B(net36));
 sg13g2_nand3_1 _7487_ (.B(net31),
    .C(_2517_),
    .A(_2425_),
    .Y(_2518_));
 sg13g2_o21ai_1 _7488_ (.B1(net32),
    .Y(_2519_),
    .A1(_2413_),
    .A2(_2494_));
 sg13g2_and3_1 _7489_ (.X(_2520_),
    .A(_2518_),
    .B(net30),
    .C(_2519_));
 sg13g2_nand3_1 _7490_ (.B(_2421_),
    .C(_2517_),
    .A(_2485_),
    .Y(_2521_));
 sg13g2_nor2_1 _7491_ (.A(net30),
    .B(_2403_),
    .Y(_2522_));
 sg13g2_o21ai_1 _7492_ (.B1(_2522_),
    .Y(_2523_),
    .A1(net31),
    .A2(_2521_));
 sg13g2_a21oi_1 _7493_ (.A1(_2280_),
    .A2(_2201_),
    .Y(_2524_),
    .B1(net32));
 sg13g2_nor2_1 _7494_ (.A(net31),
    .B(_2465_),
    .Y(_2525_));
 sg13g2_nor2_1 _7495_ (.A(net34),
    .B(_2525_),
    .Y(_2526_));
 sg13g2_o21ai_1 _7496_ (.B1(_2526_),
    .Y(_2527_),
    .A1(_2426_),
    .A2(_2524_));
 sg13g2_a21o_1 _7497_ (.A2(_2527_),
    .A1(_2523_),
    .B1(net53),
    .X(_2528_));
 sg13g2_o21ai_1 _7498_ (.B1(_2528_),
    .Y(_2529_),
    .A1(_2516_),
    .A2(_2520_));
 sg13g2_inv_1 _7499_ (.Y(_2530_),
    .A(_2255_));
 sg13g2_nor2_1 _7500_ (.A(net31),
    .B(_2280_),
    .Y(_2531_));
 sg13g2_o21ai_1 _7501_ (.B1(net34),
    .Y(_2532_),
    .A1(_2259_),
    .A2(_2281_));
 sg13g2_nor2_1 _7502_ (.A(net32),
    .B(_2239_),
    .Y(_2533_));
 sg13g2_nor2_1 _7503_ (.A(_2478_),
    .B(_2400_),
    .Y(_2534_));
 sg13g2_o21ai_1 _7504_ (.B1(net30),
    .Y(_2535_),
    .A1(_2533_),
    .A2(_2534_));
 sg13g2_o21ai_1 _7505_ (.B1(_2535_),
    .Y(_2536_),
    .A1(_2531_),
    .A2(_2532_));
 sg13g2_nor2b_1 _7506_ (.A(_2530_),
    .B_N(_2536_),
    .Y(_2537_));
 sg13g2_a221oi_1 _7507_ (.B2(_2254_),
    .C1(_2537_),
    .B1(_2529_),
    .A1(_2515_),
    .Y(_2538_),
    .A2(_2273_));
 sg13g2_nand2_1 _7508_ (.Y(_2539_),
    .A(_2155_),
    .B(_2538_));
 sg13g2_xnor2_1 _7509_ (.Y(_2540_),
    .A(\i_music.i_sample.sample_acc[4] ),
    .B(_2539_));
 sg13g2_inv_1 _7510_ (.Y(_2541_),
    .A(\i_music.i_sample.sample_acc[3] ));
 sg13g2_nand2_1 _7511_ (.Y(_2542_),
    .A(_2506_),
    .B(_2504_));
 sg13g2_o21ai_1 _7512_ (.B1(_2542_),
    .Y(_2543_),
    .A1(_2541_),
    .A2(_2503_));
 sg13g2_xnor2_1 _7513_ (.Y(_2544_),
    .A(_2540_),
    .B(_2543_));
 sg13g2_nor2_1 _7514_ (.A(\i_music.i_pwm.sample[3] ),
    .B(_2395_),
    .Y(_2545_));
 sg13g2_a21oi_1 _7515_ (.A1(_2544_),
    .A2(net113),
    .Y(_0200_),
    .B1(_2545_));
 sg13g2_buf_1 _7516_ (.A(_2155_),
    .X(_2546_));
 sg13g2_inv_1 _7517_ (.Y(_2547_),
    .A(_2509_));
 sg13g2_o21ai_1 _7518_ (.B1(_2471_),
    .Y(_2548_),
    .A1(_2547_),
    .A2(_2466_));
 sg13g2_o21ai_1 _7519_ (.B1(net31),
    .Y(_2549_),
    .A1(_2183_),
    .A2(_2280_));
 sg13g2_nand3_1 _7520_ (.B(net30),
    .C(_2549_),
    .A(_2427_),
    .Y(_2550_));
 sg13g2_nand2_1 _7521_ (.Y(_2551_),
    .A(_2548_),
    .B(_2550_));
 sg13g2_nor3_1 _7522_ (.A(_2475_),
    .B(_2525_),
    .C(_2467_),
    .Y(_2552_));
 sg13g2_o21ai_1 _7523_ (.B1(_2316_),
    .Y(_2553_),
    .A1(_2470_),
    .A2(_2317_));
 sg13g2_o21ai_1 _7524_ (.B1(net44),
    .Y(_2554_),
    .A1(_2553_),
    .A2(_2525_));
 sg13g2_o21ai_1 _7525_ (.B1(_2554_),
    .Y(_2555_),
    .A1(_2516_),
    .A2(_2552_));
 sg13g2_o21ai_1 _7526_ (.B1(_2532_),
    .Y(_2556_),
    .A1(net34),
    .A2(_2531_));
 sg13g2_nor2_1 _7527_ (.A(_2530_),
    .B(_2556_),
    .Y(_2557_));
 sg13g2_a221oi_1 _7528_ (.B2(_2254_),
    .C1(_2557_),
    .B1(_2555_),
    .A1(_2273_),
    .Y(_2558_),
    .A2(_2551_));
 sg13g2_nand2_1 _7529_ (.Y(_2559_),
    .A(net29),
    .B(_2558_));
 sg13g2_xnor2_1 _7530_ (.Y(_2560_),
    .A(\i_music.i_sample.sample_acc[5] ),
    .B(_2559_));
 sg13g2_inv_1 _7531_ (.Y(_2561_),
    .A(\i_music.i_sample.sample_acc[4] ));
 sg13g2_nor2_1 _7532_ (.A(_2561_),
    .B(_2539_),
    .Y(_2562_));
 sg13g2_a21o_1 _7533_ (.A2(_2540_),
    .A1(_2543_),
    .B1(_2562_),
    .X(_2563_));
 sg13g2_xnor2_1 _7534_ (.Y(_2564_),
    .A(_2560_),
    .B(_2563_));
 sg13g2_nor2_1 _7535_ (.A(\i_music.i_pwm.sample[4] ),
    .B(_2395_),
    .Y(_2565_));
 sg13g2_a21oi_1 _7536_ (.A1(_2564_),
    .A2(_2396_),
    .Y(_0201_),
    .B1(_2565_));
 sg13g2_nand3_1 _7537_ (.B(_2273_),
    .C(_2547_),
    .A(_2471_),
    .Y(_2566_));
 sg13g2_o21ai_1 _7538_ (.B1(_2272_),
    .Y(_2567_),
    .A1(_2475_),
    .A2(_2317_));
 sg13g2_a21o_1 _7539_ (.A2(_2567_),
    .A1(_2516_),
    .B1(_2253_),
    .X(_2568_));
 sg13g2_nand3_1 _7540_ (.B(_2566_),
    .C(_2568_),
    .A(net29),
    .Y(_2569_));
 sg13g2_xor2_1 _7541_ (.B(_2569_),
    .A(\i_music.i_sample.sample_acc[6] ),
    .X(_2570_));
 sg13g2_nand2_1 _7542_ (.Y(_2571_),
    .A(_2563_),
    .B(_2560_));
 sg13g2_nand3_1 _7543_ (.B(\i_music.i_sample.sample_acc[5] ),
    .C(_2558_),
    .A(net29),
    .Y(_2572_));
 sg13g2_nand2_1 _7544_ (.Y(_2573_),
    .A(_2571_),
    .B(_2572_));
 sg13g2_xnor2_1 _7545_ (.Y(_2574_),
    .A(_2570_),
    .B(_2573_));
 sg13g2_nor2_1 _7546_ (.A(\i_music.i_pwm.sample[5] ),
    .B(_2395_),
    .Y(_2575_));
 sg13g2_a21oi_1 _7547_ (.A1(_2574_),
    .A2(net113),
    .Y(_0202_),
    .B1(_2575_));
 sg13g2_nor2b_1 _7548_ (.A(_0064_),
    .B_N(_2570_),
    .Y(_2576_));
 sg13g2_nand4_1 _7549_ (.B(_2540_),
    .C(_2560_),
    .A(_2543_),
    .Y(_2577_),
    .D(_2576_));
 sg13g2_nand2_1 _7550_ (.Y(_2578_),
    .A(_2560_),
    .B(_2562_));
 sg13g2_nand2_1 _7551_ (.Y(_2579_),
    .A(_2578_),
    .B(_2572_));
 sg13g2_nand2_1 _7552_ (.Y(_2580_),
    .A(_2569_),
    .B(\i_music.i_sample.sample_acc[6] ));
 sg13g2_nor2_1 _7553_ (.A(_0064_),
    .B(_2580_),
    .Y(_2581_));
 sg13g2_a21oi_1 _7554_ (.A1(_2576_),
    .A2(_2579_),
    .Y(_2582_),
    .B1(_2581_));
 sg13g2_nand2_1 _7555_ (.Y(_2583_),
    .A(_2577_),
    .B(_2582_));
 sg13g2_nand2_1 _7556_ (.Y(_2584_),
    .A(_2573_),
    .B(_2570_));
 sg13g2_nand3_1 _7557_ (.B(_0064_),
    .C(_2580_),
    .A(_2584_),
    .Y(_2585_));
 sg13g2_nand2b_1 _7558_ (.Y(_2586_),
    .B(_2585_),
    .A_N(_2583_));
 sg13g2_nor2_1 _7559_ (.A(\i_music.i_pwm.sample[6] ),
    .B(_2395_),
    .Y(_2587_));
 sg13g2_a21oi_1 _7560_ (.A1(_2586_),
    .A2(net113),
    .Y(_0203_),
    .B1(_2587_));
 sg13g2_xnor2_1 _7561_ (.Y(_2588_),
    .A(\i_music.i_sample.sample_acc[8] ),
    .B(_2583_));
 sg13g2_nor2_1 _7562_ (.A(\i_music.i_pwm.sample[7] ),
    .B(_2395_),
    .Y(_2589_));
 sg13g2_a21oi_1 _7563_ (.A1(_2588_),
    .A2(_2396_),
    .Y(_0204_),
    .B1(_2589_));
 sg13g2_nor2_1 _7564_ (.A(_4230_),
    .B(_4239_),
    .Y(_2590_));
 sg13g2_inv_1 _7565_ (.Y(_2591_),
    .A(_2590_));
 sg13g2_inv_1 _7566_ (.Y(_2592_),
    .A(_1746_));
 sg13g2_a21oi_1 _7567_ (.A1(_1806_),
    .A2(_1790_),
    .Y(_2593_),
    .B1(_2592_));
 sg13g2_o21ai_1 _7568_ (.B1(net95),
    .Y(_2594_),
    .A1(_1829_),
    .A2(_2003_));
 sg13g2_nand3b_1 _7569_ (.B(_1787_),
    .C(_1800_),
    .Y(_2595_),
    .A_N(_1887_));
 sg13g2_a22oi_1 _7570_ (.Y(_2596_),
    .B1(_1819_),
    .B2(_2595_),
    .A2(_1708_),
    .A1(_1974_));
 sg13g2_o21ai_1 _7571_ (.B1(_2596_),
    .Y(_2597_),
    .A1(_2593_),
    .A2(_2594_));
 sg13g2_nand2_1 _7572_ (.Y(_2598_),
    .A(_2597_),
    .B(_1770_));
 sg13g2_a21oi_1 _7573_ (.A1(_1806_),
    .A2(_1790_),
    .Y(_2599_),
    .B1(net88));
 sg13g2_nor2b_1 _7574_ (.A(_1917_),
    .B_N(_1766_),
    .Y(_2600_));
 sg13g2_o21ai_1 _7575_ (.B1(_2600_),
    .Y(_2601_),
    .A1(_1984_),
    .A2(_1800_));
 sg13g2_o21ai_1 _7576_ (.B1(_2601_),
    .Y(_2602_),
    .A1(_1813_),
    .A2(_2599_));
 sg13g2_nand2_1 _7577_ (.Y(_2603_),
    .A(_2602_),
    .B(_1722_));
 sg13g2_nor3_1 _7578_ (.A(_1769_),
    .B(_1720_),
    .C(_1813_),
    .Y(_2604_));
 sg13g2_a22oi_1 _7579_ (.Y(_2605_),
    .B1(_1936_),
    .B2(_2604_),
    .A2(_1911_),
    .A1(_1902_));
 sg13g2_nand3_1 _7580_ (.B(net103),
    .C(_1900_),
    .A(_1967_),
    .Y(_2606_));
 sg13g2_a21oi_1 _7581_ (.A1(net99),
    .A2(_1751_),
    .Y(_2607_),
    .B1(_1949_));
 sg13g2_nand2_1 _7582_ (.Y(_2608_),
    .A(_2607_),
    .B(_1882_));
 sg13g2_nand3_1 _7583_ (.B(_2608_),
    .C(_1742_),
    .A(_2606_),
    .Y(_2609_));
 sg13g2_nand4_1 _7584_ (.B(_2603_),
    .C(_2605_),
    .A(_2598_),
    .Y(_2610_),
    .D(_2609_));
 sg13g2_nand2_1 _7585_ (.Y(_2611_),
    .A(_2610_),
    .B(_1833_));
 sg13g2_o21ai_1 _7586_ (.B1(_2611_),
    .Y(_2612_),
    .A1(_1833_),
    .A2(_1911_));
 sg13g2_nand2_1 _7587_ (.Y(_2613_),
    .A(_2612_),
    .B(\i_music.count[24] ));
 sg13g2_nand3_1 _7588_ (.B(_0077_),
    .C(_1575_),
    .A(_2613_),
    .Y(_2614_));
 sg13g2_o21ai_1 _7589_ (.B1(net88),
    .Y(_2615_),
    .A1(_1728_),
    .A2(_1739_));
 sg13g2_a21oi_1 _7590_ (.A1(_2615_),
    .A2(_1799_),
    .Y(_2616_),
    .B1(_1835_));
 sg13g2_and3_1 _7591_ (.X(_2617_),
    .A(_2604_),
    .B(net99),
    .C(_1754_));
 sg13g2_nor4_1 _7592_ (.A(_1673_),
    .B(_1724_),
    .C(_2616_),
    .D(_2617_),
    .Y(_2618_));
 sg13g2_o21ai_1 _7593_ (.B1(_2618_),
    .Y(_2619_),
    .A1(_0077_),
    .A2(_2612_));
 sg13g2_nand2_1 _7594_ (.Y(_2620_),
    .A(_2614_),
    .B(_2619_));
 sg13g2_nor4_1 _7595_ (.A(_4238_),
    .B(\i_music.count[11] ),
    .C(_1587_),
    .D(\i_music.count[13] ),
    .Y(_2621_));
 sg13g2_nand2_1 _7596_ (.Y(_2622_),
    .A(_1160_),
    .B(_1155_));
 sg13g2_inv_1 _7597_ (.Y(_2623_),
    .A(_2030_));
 sg13g2_nor2_1 _7598_ (.A(_2622_),
    .B(_2623_),
    .Y(_2624_));
 sg13g2_nand2b_1 _7599_ (.Y(_2625_),
    .B(_1578_),
    .A_N(\i_music.count[16] ));
 sg13g2_inv_1 _7600_ (.Y(_2626_),
    .A(\i_music.count[12] ));
 sg13g2_inv_1 _7601_ (.Y(_2627_),
    .A(\i_music.count[14] ));
 sg13g2_nand4_1 _7602_ (.B(_1580_),
    .C(_2627_),
    .A(_2626_),
    .Y(_2628_),
    .D(_1579_));
 sg13g2_nor4_1 _7603_ (.A(\i_music.count[18] ),
    .B(_2625_),
    .C(_4229_),
    .D(_2628_),
    .Y(_2629_));
 sg13g2_nand4_1 _7604_ (.B(_2621_),
    .C(_2624_),
    .A(_2620_),
    .Y(_2630_),
    .D(_2629_));
 sg13g2_nor4_2 _7605_ (.A(_1050_),
    .B(_1489_),
    .C(_2591_),
    .Y(_2631_),
    .D(_2630_));
 sg13g2_nor2_1 _7606_ (.A(net147),
    .B(_2631_),
    .Y(_2632_));
 sg13g2_buf_1 _7607_ (.A(_2632_),
    .X(_2633_));
 sg13g2_buf_1 _7608_ (.A(_1665_),
    .X(_2634_));
 sg13g2_buf_1 _7609_ (.A(\i_music.violin_note_idx[1][3] ),
    .X(_2635_));
 sg13g2_inv_1 _7610_ (.Y(_2636_),
    .A(\i_music.violin_note_idx[1][8] ));
 sg13g2_nor4_1 _7611_ (.A(_2635_),
    .B(_2054_),
    .C(\i_music.violin_note_idx[1][6] ),
    .D(_2636_),
    .Y(_2637_));
 sg13g2_inv_1 _7612_ (.Y(_2638_),
    .A(\i_music.violin_note_idx[1][2] ));
 sg13g2_inv_1 _7613_ (.Y(_2639_),
    .A(\i_music.violin_note_idx[1][5] ));
 sg13g2_nor2_1 _7614_ (.A(\i_music.violin_note_idx[1][4] ),
    .B(_2639_),
    .Y(_2640_));
 sg13g2_nor2_1 _7615_ (.A(\i_music.violin_note_idx[1][1] ),
    .B(\i_music.violin_note_idx[1][0] ),
    .Y(_2641_));
 sg13g2_nand4_1 _7616_ (.B(_2638_),
    .C(_2640_),
    .A(_2637_),
    .Y(_2642_),
    .D(_2641_));
 sg13g2_buf_2 _7617_ (.A(_2642_),
    .X(_2643_));
 sg13g2_inv_1 _7618_ (.Y(_2644_),
    .A(_2643_));
 sg13g2_nor3_1 _7619_ (.A(net127),
    .B(_0103_),
    .C(net120),
    .Y(_2645_));
 sg13g2_nand2_1 _7620_ (.Y(_2646_),
    .A(net43),
    .B(\i_music.violin_note_idx[1][0] ));
 sg13g2_o21ai_1 _7621_ (.B1(_2646_),
    .Y(_0214_),
    .A1(net43),
    .A2(_2645_));
 sg13g2_inv_1 _7622_ (.Y(_2647_),
    .A(\i_music.violin_note_idx[1][1] ));
 sg13g2_inv_1 _7623_ (.Y(_2648_),
    .A(_2633_));
 sg13g2_nand2_1 _7624_ (.Y(_2649_),
    .A(\i_music.violin_note_idx[1][1] ),
    .B(\i_music.violin_note_idx[1][0] ));
 sg13g2_nor2b_1 _7625_ (.A(_2641_),
    .B_N(_2649_),
    .Y(_2650_));
 sg13g2_a21oi_1 _7626_ (.A1(_2631_),
    .A2(_2650_),
    .Y(_2651_),
    .B1(net128));
 sg13g2_o21ai_1 _7627_ (.B1(_2651_),
    .Y(_0215_),
    .A1(_2647_),
    .A2(_2648_));
 sg13g2_xnor2_1 _7628_ (.Y(_2652_),
    .A(_0083_),
    .B(_2649_));
 sg13g2_nor2_1 _7629_ (.A(_2652_),
    .B(net120),
    .Y(_2653_));
 sg13g2_a21oi_1 _7630_ (.A1(_2631_),
    .A2(_2653_),
    .Y(_2654_),
    .B1(net128));
 sg13g2_o21ai_1 _7631_ (.B1(_2654_),
    .Y(_0216_),
    .A1(_2638_),
    .A2(_2648_));
 sg13g2_inv_1 _7632_ (.Y(_2655_),
    .A(_2635_));
 sg13g2_nor2_1 _7633_ (.A(_2638_),
    .B(_2649_),
    .Y(_2656_));
 sg13g2_nand2_1 _7634_ (.Y(_2657_),
    .A(_2656_),
    .B(_2635_));
 sg13g2_inv_1 _7635_ (.Y(_2658_),
    .A(_2657_));
 sg13g2_nor2_1 _7636_ (.A(_2635_),
    .B(_2656_),
    .Y(_2659_));
 sg13g2_o21ai_1 _7637_ (.B1(_2643_),
    .Y(_2660_),
    .A1(_2658_),
    .A2(_2659_));
 sg13g2_nand3_1 _7638_ (.B(net143),
    .C(_2660_),
    .A(_2631_),
    .Y(_2661_));
 sg13g2_o21ai_1 _7639_ (.B1(_2661_),
    .Y(_0217_),
    .A1(_2655_),
    .A2(_2648_));
 sg13g2_inv_1 _7640_ (.Y(_2662_),
    .A(\i_music.violin_note_idx[1][4] ));
 sg13g2_xnor2_1 _7641_ (.Y(_2663_),
    .A(_0080_),
    .B(_2657_));
 sg13g2_o21ai_1 _7642_ (.B1(net143),
    .Y(_2664_),
    .A1(_2663_),
    .A2(net120));
 sg13g2_inv_1 _7643_ (.Y(_2665_),
    .A(net1));
 sg13g2_nor2_1 _7644_ (.A(net157),
    .B(_2665_),
    .Y(_2666_));
 sg13g2_inv_1 _7645_ (.Y(_2667_),
    .A(_2666_));
 sg13g2_nand3_1 _7646_ (.B(_2664_),
    .C(_2667_),
    .A(_2648_),
    .Y(_2668_));
 sg13g2_o21ai_1 _7647_ (.B1(_2668_),
    .Y(_0218_),
    .A1(_2662_),
    .A2(_2648_));
 sg13g2_nor2_1 _7648_ (.A(_2662_),
    .B(_2657_),
    .Y(_2669_));
 sg13g2_nor2_1 _7649_ (.A(\i_music.violin_note_idx[1][5] ),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_inv_1 _7650_ (.Y(_2671_),
    .A(_2669_));
 sg13g2_nor2_1 _7651_ (.A(_2639_),
    .B(_2671_),
    .Y(_2672_));
 sg13g2_nor3_1 _7652_ (.A(net135),
    .B(_2670_),
    .C(_2672_),
    .Y(_2673_));
 sg13g2_inv_1 _7653_ (.Y(_2674_),
    .A(net2));
 sg13g2_nor2_1 _7654_ (.A(net157),
    .B(net2),
    .Y(_2675_));
 sg13g2_nand2_1 _7655_ (.Y(_2676_),
    .A(_2675_),
    .B(_2665_));
 sg13g2_o21ai_1 _7656_ (.B1(_2676_),
    .Y(_2677_),
    .A1(_2674_),
    .A2(_2667_));
 sg13g2_nor3_1 _7657_ (.A(_2673_),
    .B(_2677_),
    .C(net43),
    .Y(_2678_));
 sg13g2_a21oi_1 _7658_ (.A1(_2639_),
    .A2(net43),
    .Y(_0219_),
    .B1(_2678_));
 sg13g2_inv_1 _7659_ (.Y(_2679_),
    .A(\i_music.violin_note_idx[1][6] ));
 sg13g2_xnor2_1 _7660_ (.Y(_2680_),
    .A(_2679_),
    .B(_2672_));
 sg13g2_o21ai_1 _7661_ (.B1(net143),
    .Y(_2681_),
    .A1(net120),
    .A2(_2680_));
 sg13g2_nor2b_1 _7662_ (.A(net43),
    .B_N(_2676_),
    .Y(_2682_));
 sg13g2_a22oi_1 _7663_ (.Y(_0220_),
    .B1(_2681_),
    .B2(_2682_),
    .A2(net43),
    .A1(_2679_));
 sg13g2_inv_1 _7664_ (.Y(_2683_),
    .A(_2054_));
 sg13g2_inv_1 _7665_ (.Y(_2684_),
    .A(_2672_));
 sg13g2_nor2_1 _7666_ (.A(_2679_),
    .B(_2684_),
    .Y(_2685_));
 sg13g2_nor2_1 _7667_ (.A(_2054_),
    .B(_2685_),
    .Y(_2686_));
 sg13g2_inv_1 _7668_ (.Y(_2687_),
    .A(_2685_));
 sg13g2_nor2_1 _7669_ (.A(_2683_),
    .B(_2687_),
    .Y(_2688_));
 sg13g2_o21ai_1 _7670_ (.B1(_2643_),
    .Y(_2689_),
    .A1(_2686_),
    .A2(_2688_));
 sg13g2_buf_1 _7671_ (.A(net143),
    .X(_2690_));
 sg13g2_nand2_1 _7672_ (.Y(_2691_),
    .A(_2689_),
    .B(net134));
 sg13g2_a22oi_1 _7673_ (.Y(_0221_),
    .B1(_2691_),
    .B2(_2682_),
    .A2(net43),
    .A1(_2683_));
 sg13g2_nor3_1 _7674_ (.A(_2683_),
    .B(\i_music.violin_note_idx[1][8] ),
    .C(_2687_),
    .Y(_2692_));
 sg13g2_nor2_1 _7675_ (.A(_2636_),
    .B(_2688_),
    .Y(_2693_));
 sg13g2_o21ai_1 _7676_ (.B1(net143),
    .Y(_2694_),
    .A1(_2692_),
    .A2(_2693_));
 sg13g2_a22oi_1 _7677_ (.Y(_0222_),
    .B1(_2694_),
    .B2(_2682_),
    .A2(net43),
    .A1(_2636_));
 sg13g2_nor4_1 _7678_ (.A(\i_music.count[17] ),
    .B(\i_music.count[18] ),
    .C(_2623_),
    .D(_2625_),
    .Y(_2695_));
 sg13g2_nand4_1 _7679_ (.B(_2626_),
    .C(_1580_),
    .A(_1581_),
    .Y(_2696_),
    .D(_2627_));
 sg13g2_nor4_1 _7680_ (.A(\i_music.count[11] ),
    .B(_1587_),
    .C(_2622_),
    .D(_2696_),
    .Y(_2697_));
 sg13g2_nor4_1 _7681_ (.A(_4238_),
    .B(_2156_),
    .C(_2591_),
    .D(_4229_),
    .Y(_2698_));
 sg13g2_nand4_1 _7682_ (.B(_2695_),
    .C(_2697_),
    .A(_2620_),
    .Y(_2699_),
    .D(_2698_));
 sg13g2_nand2_1 _7683_ (.Y(_2700_),
    .A(_2699_),
    .B(net157));
 sg13g2_buf_2 _7684_ (.A(_2700_),
    .X(_2701_));
 sg13g2_buf_1 _7685_ (.A(_2701_),
    .X(_2702_));
 sg13g2_nand4_1 _7686_ (.B(\i_music.violin_note_idx[1][0] ),
    .C(_2635_),
    .A(_2647_),
    .Y(_2703_),
    .D(\i_music.violin_note_idx[1][6] ));
 sg13g2_nor2_1 _7687_ (.A(_2055_),
    .B(_2703_),
    .Y(_2704_));
 sg13g2_and3_1 _7688_ (.X(_2705_),
    .A(_2704_),
    .B(_2638_),
    .C(_2640_));
 sg13g2_buf_1 _7689_ (.A(_2705_),
    .X(_2706_));
 sg13g2_inv_1 _7690_ (.Y(_2707_),
    .A(_2706_));
 sg13g2_nand2_2 _7691_ (.Y(_2708_),
    .A(_2707_),
    .B(_2643_));
 sg13g2_nor2_1 _7692_ (.A(net135),
    .B(_2708_),
    .Y(_2709_));
 sg13g2_inv_1 _7693_ (.Y(_2710_),
    .A(_2709_));
 sg13g2_o21ai_1 _7694_ (.B1(_2702_),
    .Y(_2711_),
    .A1(_0104_),
    .A2(_2710_));
 sg13g2_o21ai_1 _7695_ (.B1(_2711_),
    .Y(_0223_),
    .A1(_1730_),
    .A2(net42));
 sg13g2_nand2_1 _7696_ (.Y(_2712_),
    .A(\i_music.violin_note_idx[2][1] ),
    .B(\i_music.violin_note_idx[2][0] ));
 sg13g2_inv_1 _7697_ (.Y(_2713_),
    .A(_2712_));
 sg13g2_nor2_1 _7698_ (.A(\i_music.violin_note_idx[2][1] ),
    .B(\i_music.violin_note_idx[2][0] ),
    .Y(_2714_));
 sg13g2_nor3_1 _7699_ (.A(_2713_),
    .B(_2714_),
    .C(_2708_),
    .Y(_2715_));
 sg13g2_o21ai_1 _7700_ (.B1(_2701_),
    .Y(_2716_),
    .A1(net127),
    .A2(_2715_));
 sg13g2_o21ai_1 _7701_ (.B1(_2716_),
    .Y(_0224_),
    .A1(_1683_),
    .A2(net42));
 sg13g2_nor2_1 _7702_ (.A(_1689_),
    .B(_2712_),
    .Y(_2717_));
 sg13g2_nor2_1 _7703_ (.A(\i_music.violin_note_idx[2][2] ),
    .B(_2713_),
    .Y(_2718_));
 sg13g2_nor3_1 _7704_ (.A(_2717_),
    .B(_2718_),
    .C(_2708_),
    .Y(_2719_));
 sg13g2_o21ai_1 _7705_ (.B1(_2701_),
    .Y(_2720_),
    .A1(net127),
    .A2(_2719_));
 sg13g2_o21ai_1 _7706_ (.B1(_2720_),
    .Y(_0225_),
    .A1(_1689_),
    .A2(net42));
 sg13g2_nor2_1 _7707_ (.A(\i_music.violin_note_idx[2][3] ),
    .B(_2717_),
    .Y(_2721_));
 sg13g2_inv_1 _7708_ (.Y(_2722_),
    .A(_2717_));
 sg13g2_nor2_1 _7709_ (.A(_1674_),
    .B(_2722_),
    .Y(_2723_));
 sg13g2_nor3_1 _7710_ (.A(_2721_),
    .B(_2723_),
    .C(_2708_),
    .Y(_2724_));
 sg13g2_o21ai_1 _7711_ (.B1(_2701_),
    .Y(_2725_),
    .A1(net127),
    .A2(_2724_));
 sg13g2_o21ai_1 _7712_ (.B1(_2725_),
    .Y(_0226_),
    .A1(_1674_),
    .A2(_2702_));
 sg13g2_nand2_1 _7713_ (.Y(_2726_),
    .A(_2723_),
    .B(\i_music.violin_note_idx[2][4] ));
 sg13g2_o21ai_1 _7714_ (.B1(_1702_),
    .Y(_2727_),
    .A1(_1674_),
    .A2(_2722_));
 sg13g2_nand4_1 _7715_ (.B(_2709_),
    .C(_2726_),
    .A(_2701_),
    .Y(_2728_),
    .D(_2727_));
 sg13g2_nand3_1 _7716_ (.B(net143),
    .C(\i_music.violin_note_idx[2][4] ),
    .A(_2699_),
    .Y(_2729_));
 sg13g2_nand3_1 _7717_ (.B(_2729_),
    .C(_2667_),
    .A(_2728_),
    .Y(_0227_));
 sg13g2_nor2_1 _7718_ (.A(net157),
    .B(_2674_),
    .Y(_2730_));
 sg13g2_inv_1 _7719_ (.Y(_2731_),
    .A(_2730_));
 sg13g2_nor2_1 _7720_ (.A(_1696_),
    .B(_2726_),
    .Y(_2732_));
 sg13g2_a21oi_1 _7721_ (.A1(_2723_),
    .A2(\i_music.violin_note_idx[2][4] ),
    .Y(_2733_),
    .B1(\i_music.violin_note_idx[2][5] ));
 sg13g2_o21ai_1 _7722_ (.B1(_2709_),
    .Y(_2734_),
    .A1(_2732_),
    .A2(_2733_));
 sg13g2_nand3_1 _7723_ (.B(_2731_),
    .C(_2734_),
    .A(_2701_),
    .Y(_2735_));
 sg13g2_o21ai_1 _7724_ (.B1(_2735_),
    .Y(_0228_),
    .A1(_1696_),
    .A2(net42));
 sg13g2_inv_1 _7725_ (.Y(_2736_),
    .A(_2732_));
 sg13g2_a21oi_1 _7726_ (.A1(_1710_),
    .A2(_2736_),
    .Y(_2737_),
    .B1(net120));
 sg13g2_nor2_1 _7727_ (.A(_1710_),
    .B(_2736_),
    .Y(_2738_));
 sg13g2_inv_1 _7728_ (.Y(_2739_),
    .A(_2738_));
 sg13g2_nor2_2 _7729_ (.A(_1308_),
    .B(_2706_),
    .Y(_2740_));
 sg13g2_inv_1 _7730_ (.Y(_2741_),
    .A(_2740_));
 sg13g2_a21oi_1 _7731_ (.A1(_2737_),
    .A2(_2739_),
    .Y(_2742_),
    .B1(_2741_));
 sg13g2_o21ai_1 _7732_ (.B1(_2731_),
    .Y(_2743_),
    .A1(\i_music.violin_note_idx[2][6] ),
    .A2(_2701_));
 sg13g2_a21oi_1 _7733_ (.A1(net42),
    .A2(_2742_),
    .Y(_0229_),
    .B1(_2743_));
 sg13g2_nand2_1 _7734_ (.Y(_2744_),
    .A(_2739_),
    .B(_1716_));
 sg13g2_nand2_1 _7735_ (.Y(_2745_),
    .A(_2738_),
    .B(\i_music.violin_note_idx[2][7] ));
 sg13g2_nand3_1 _7736_ (.B(_2643_),
    .C(_2745_),
    .A(_2744_),
    .Y(_2746_));
 sg13g2_nand2_1 _7737_ (.Y(_2747_),
    .A(_2746_),
    .B(_2740_));
 sg13g2_nand3_1 _7738_ (.B(_2731_),
    .C(_2747_),
    .A(_2701_),
    .Y(_2748_));
 sg13g2_o21ai_1 _7739_ (.B1(_2748_),
    .Y(_0230_),
    .A1(_1716_),
    .A2(net42));
 sg13g2_xnor2_1 _7740_ (.Y(_2749_),
    .A(_1669_),
    .B(_2745_));
 sg13g2_a21oi_1 _7741_ (.A1(_2749_),
    .A2(_2709_),
    .Y(_2750_),
    .B1(_2730_));
 sg13g2_nand2_1 _7742_ (.Y(_2751_),
    .A(net42),
    .B(_2750_));
 sg13g2_o21ai_1 _7743_ (.B1(_2751_),
    .Y(_0231_),
    .A1(_1669_),
    .A2(net42));
 sg13g2_o21ai_1 _7744_ (.B1(_2740_),
    .Y(_2752_),
    .A1(_1729_),
    .A2(net120));
 sg13g2_nor3_2 _7745_ (.A(net136),
    .B(_2591_),
    .C(_2630_),
    .Y(_2753_));
 sg13g2_nor2_1 _7746_ (.A(_1308_),
    .B(_2753_),
    .Y(_2754_));
 sg13g2_inv_1 _7747_ (.Y(_2755_),
    .A(_2754_));
 sg13g2_mux2_1 _7748_ (.A0(_1729_),
    .A1(_2752_),
    .S(net41),
    .X(_0232_));
 sg13g2_inv_1 _7749_ (.Y(_2756_),
    .A(_1682_));
 sg13g2_xnor2_1 _7750_ (.Y(_2757_),
    .A(_1682_),
    .B(_1729_));
 sg13g2_a21oi_1 _7751_ (.A1(_2643_),
    .A2(_2757_),
    .Y(_2758_),
    .B1(_2706_));
 sg13g2_a21oi_1 _7752_ (.A1(_2753_),
    .A2(_2758_),
    .Y(_2759_),
    .B1(_1666_));
 sg13g2_o21ai_1 _7753_ (.B1(_2759_),
    .Y(_0233_),
    .A1(_2756_),
    .A2(net41));
 sg13g2_inv_1 _7754_ (.Y(_2760_),
    .A(\i_music.violin_note_idx[3][2] ));
 sg13g2_nand2_1 _7755_ (.Y(_2761_),
    .A(_1682_),
    .B(_1729_));
 sg13g2_nor2_1 _7756_ (.A(_2760_),
    .B(_2761_),
    .Y(_2762_));
 sg13g2_a21oi_1 _7757_ (.A1(_1682_),
    .A2(_1729_),
    .Y(_2763_),
    .B1(\i_music.violin_note_idx[3][2] ));
 sg13g2_nor3_1 _7758_ (.A(_2762_),
    .B(_2763_),
    .C(_2708_),
    .Y(_2764_));
 sg13g2_a21oi_1 _7759_ (.A1(_2753_),
    .A2(_2764_),
    .Y(_2765_),
    .B1(net128));
 sg13g2_o21ai_1 _7760_ (.B1(_2765_),
    .Y(_0234_),
    .A1(_2760_),
    .A2(net41));
 sg13g2_xnor2_1 _7761_ (.Y(_2766_),
    .A(\i_music.violin_note_idx[3][3] ),
    .B(_2762_));
 sg13g2_o21ai_1 _7762_ (.B1(_2707_),
    .Y(_2767_),
    .A1(_2766_),
    .A2(net120));
 sg13g2_nand3_1 _7763_ (.B(_1637_),
    .C(_2767_),
    .A(_2753_),
    .Y(_2768_));
 sg13g2_o21ai_1 _7764_ (.B1(_2768_),
    .Y(_0235_),
    .A1(_1675_),
    .A2(net41));
 sg13g2_nor3_1 _7765_ (.A(_1675_),
    .B(_2760_),
    .C(_2761_),
    .Y(_2769_));
 sg13g2_inv_1 _7766_ (.Y(_2770_),
    .A(_2769_));
 sg13g2_nor2_1 _7767_ (.A(_1703_),
    .B(_2770_),
    .Y(_2771_));
 sg13g2_inv_1 _7768_ (.Y(_2772_),
    .A(_2771_));
 sg13g2_nand2_1 _7769_ (.Y(_2773_),
    .A(_2770_),
    .B(_1703_));
 sg13g2_nand3_1 _7770_ (.B(_2772_),
    .C(_2773_),
    .A(_2643_),
    .Y(_2774_));
 sg13g2_a22oi_1 _7771_ (.Y(_2775_),
    .B1(_2740_),
    .B2(_2774_),
    .A2(_2665_),
    .A1(_1665_));
 sg13g2_nor2_1 _7772_ (.A(_2775_),
    .B(_2754_),
    .Y(_2776_));
 sg13g2_a21oi_1 _7773_ (.A1(_1703_),
    .A2(_2754_),
    .Y(_0236_),
    .B1(_2776_));
 sg13g2_nand2_1 _7774_ (.Y(_2777_),
    .A(_2772_),
    .B(_1697_));
 sg13g2_nand2_1 _7775_ (.Y(_2778_),
    .A(_2771_),
    .B(\i_music.violin_note_idx[3][5] ));
 sg13g2_a21oi_1 _7776_ (.A1(_2777_),
    .A2(_2778_),
    .Y(_2779_),
    .B1(net120));
 sg13g2_nor2_1 _7777_ (.A(_2741_),
    .B(_2779_),
    .Y(_2780_));
 sg13g2_o21ai_1 _7778_ (.B1(net41),
    .Y(_2781_),
    .A1(_2675_),
    .A2(_2780_));
 sg13g2_o21ai_1 _7779_ (.B1(_2781_),
    .Y(_0237_),
    .A1(_1697_),
    .A2(_2755_));
 sg13g2_a21oi_1 _7780_ (.A1(_1711_),
    .A2(_2778_),
    .Y(_2782_),
    .B1(_2644_));
 sg13g2_nor2_1 _7781_ (.A(_1711_),
    .B(_2778_),
    .Y(_2783_));
 sg13g2_inv_1 _7782_ (.Y(_2784_),
    .A(_2783_));
 sg13g2_a21oi_1 _7783_ (.A1(_2782_),
    .A2(_2784_),
    .Y(_2785_),
    .B1(_2741_));
 sg13g2_nor2_1 _7784_ (.A(_2730_),
    .B(_2754_),
    .Y(_2786_));
 sg13g2_nand2b_1 _7785_ (.Y(_2787_),
    .B(_2786_),
    .A_N(_2785_));
 sg13g2_o21ai_1 _7786_ (.B1(_2787_),
    .Y(_0238_),
    .A1(_1711_),
    .A2(net41));
 sg13g2_inv_1 _7787_ (.Y(_2788_),
    .A(\i_music.violin_note_idx[3][7] ));
 sg13g2_nor2b_1 _7788_ (.A(_2783_),
    .B_N(_0085_),
    .Y(_2789_));
 sg13g2_nor2_1 _7789_ (.A(_0085_),
    .B(_2784_),
    .Y(_2790_));
 sg13g2_nor3_1 _7790_ (.A(_2644_),
    .B(_2789_),
    .C(_2790_),
    .Y(_2791_));
 sg13g2_o21ai_1 _7791_ (.B1(_2786_),
    .Y(_2792_),
    .A1(_2741_),
    .A2(_2791_));
 sg13g2_o21ai_1 _7792_ (.B1(_2792_),
    .Y(_0239_),
    .A1(_2788_),
    .A2(net41));
 sg13g2_nand2_1 _7793_ (.Y(_2793_),
    .A(_2783_),
    .B(\i_music.violin_note_idx[3][7] ));
 sg13g2_xnor2_1 _7794_ (.Y(_2794_),
    .A(\i_music.violin_note_idx[3][8] ),
    .B(_2793_));
 sg13g2_o21ai_1 _7795_ (.B1(_2786_),
    .Y(_2795_),
    .A1(_2710_),
    .A2(_2794_));
 sg13g2_o21ai_1 _7796_ (.B1(_2795_),
    .Y(_0240_),
    .A1(_1670_),
    .A2(net41));
 sg13g2_inv_1 _7797_ (.Y(_2796_),
    .A(_0026_));
 sg13g2_nand3_1 _7798_ (.B(_1109_),
    .C(_1146_),
    .A(_1000_),
    .Y(_2797_));
 sg13g2_buf_1 _7799_ (.A(_2797_),
    .X(_2798_));
 sg13g2_inv_1 _7800_ (.Y(_2799_),
    .A(_2798_));
 sg13g2_nor2_1 _7801_ (.A(net135),
    .B(_0640_),
    .Y(_2800_));
 sg13g2_o21ai_1 _7802_ (.B1(_2800_),
    .Y(_2801_),
    .A1(\i_display.in_line ),
    .A2(_2799_));
 sg13g2_a21oi_1 _7803_ (.A1(_2796_),
    .A2(_2799_),
    .Y(_0140_),
    .B1(_2801_));
 sg13g2_o21ai_1 _7804_ (.B1(_2800_),
    .Y(_2802_),
    .A1(_0101_),
    .A2(_2798_));
 sg13g2_a21oi_1 _7805_ (.A1(_4174_),
    .A2(_2798_),
    .Y(_0141_),
    .B1(_2802_));
 sg13g2_nand2_1 _7806_ (.Y(_2803_),
    .A(_4273_),
    .B(_4196_));
 sg13g2_o21ai_1 _7807_ (.B1(_2800_),
    .Y(_2804_),
    .A1(_4294_),
    .A2(_2799_));
 sg13g2_a21oi_1 _7808_ (.A1(_2799_),
    .A2(_2803_),
    .Y(_0142_),
    .B1(_2804_));
 sg13g2_nor3_1 _7809_ (.A(_1271_),
    .B(_1431_),
    .C(_1365_),
    .Y(_0150_));
 sg13g2_nand4_1 _7810_ (.B(\i_music.i_pwm.count[2] ),
    .C(\i_music.i_pwm.count[4] ),
    .A(\i_music.i_pwm.count[3] ),
    .Y(_2805_),
    .D(\i_music.i_pwm.count[7] ));
 sg13g2_nor2b_1 _7811_ (.A(\i_music.i_pwm.count[0] ),
    .B_N(_1649_),
    .Y(_2806_));
 sg13g2_nand3_1 _7812_ (.B(\i_music.i_pwm.count[5] ),
    .C(\i_music.i_pwm.count[6] ),
    .A(_2806_),
    .Y(_2807_));
 sg13g2_o21ai_1 _7813_ (.B1(net157),
    .Y(_2808_),
    .A1(_2805_),
    .A2(_2807_));
 sg13g2_buf_2 _7814_ (.A(_2808_),
    .X(_2809_));
 sg13g2_nor2b_1 _7815_ (.A(_2809_),
    .B_N(_0105_),
    .Y(_0188_));
 sg13g2_nor2_1 _7816_ (.A(\i_music.i_pwm.count[0] ),
    .B(_1649_),
    .Y(_2810_));
 sg13g2_nand2_1 _7817_ (.Y(_2811_),
    .A(\i_music.i_pwm.count[0] ),
    .B(_1649_));
 sg13g2_inv_1 _7818_ (.Y(_2812_),
    .A(_2811_));
 sg13g2_nor3_1 _7819_ (.A(_2810_),
    .B(_2812_),
    .C(_2809_),
    .Y(_0189_));
 sg13g2_nor2_1 _7820_ (.A(\i_music.i_pwm.count[2] ),
    .B(_2812_),
    .Y(_2813_));
 sg13g2_nor2_1 _7821_ (.A(_1653_),
    .B(_2811_),
    .Y(_2814_));
 sg13g2_nor3_1 _7822_ (.A(_2813_),
    .B(_2814_),
    .C(_2809_),
    .Y(_0190_));
 sg13g2_nor2_1 _7823_ (.A(\i_music.i_pwm.count[3] ),
    .B(_2814_),
    .Y(_2815_));
 sg13g2_nand2_1 _7824_ (.Y(_2816_),
    .A(_2814_),
    .B(\i_music.i_pwm.count[3] ));
 sg13g2_inv_1 _7825_ (.Y(_2817_),
    .A(_2816_));
 sg13g2_nor3_1 _7826_ (.A(_2815_),
    .B(_2817_),
    .C(_2809_),
    .Y(_0191_));
 sg13g2_nor2_1 _7827_ (.A(\i_music.i_pwm.count[4] ),
    .B(_2817_),
    .Y(_2818_));
 sg13g2_nor2_1 _7828_ (.A(_1642_),
    .B(_2816_),
    .Y(_2819_));
 sg13g2_nor3_1 _7829_ (.A(_2818_),
    .B(_2819_),
    .C(_2809_),
    .Y(_0192_));
 sg13g2_nor2_1 _7830_ (.A(\i_music.i_pwm.count[5] ),
    .B(_2819_),
    .Y(_2820_));
 sg13g2_inv_1 _7831_ (.Y(_2821_),
    .A(_2819_));
 sg13g2_nor2_1 _7832_ (.A(_1640_),
    .B(_2821_),
    .Y(_2822_));
 sg13g2_nor3_1 _7833_ (.A(_2820_),
    .B(_2822_),
    .C(_2809_),
    .Y(_0193_));
 sg13g2_nor3_1 _7834_ (.A(_1640_),
    .B(_1661_),
    .C(_2821_),
    .Y(_2823_));
 sg13g2_nor2_1 _7835_ (.A(\i_music.i_pwm.count[6] ),
    .B(_2822_),
    .Y(_2824_));
 sg13g2_nor3_1 _7836_ (.A(_2809_),
    .B(_2823_),
    .C(_2824_),
    .Y(_0194_));
 sg13g2_xnor2_1 _7837_ (.Y(_2825_),
    .A(\i_music.i_pwm.count[7] ),
    .B(_2823_));
 sg13g2_nor2_1 _7838_ (.A(_2809_),
    .B(_2825_),
    .Y(_0195_));
 sg13g2_inv_4 _7839_ (.A(_1632_),
    .Y(_2826_));
 sg13g2_nor2_1 _7840_ (.A(_1631_),
    .B(_2826_),
    .Y(_2827_));
 sg13g2_inv_1 _7841_ (.Y(_2828_),
    .A(_2827_));
 sg13g2_nor2_1 _7842_ (.A(_1629_),
    .B(_2828_),
    .Y(_2829_));
 sg13g2_inv_1 _7843_ (.Y(_2830_),
    .A(_2829_));
 sg13g2_nand4_1 _7844_ (.B(_1631_),
    .C(_1626_),
    .A(_2826_),
    .Y(_2831_),
    .D(\i_display.frame_crotchet[3] ));
 sg13g2_buf_1 _7845_ (.A(_2831_),
    .X(_2832_));
 sg13g2_a21oi_1 _7846_ (.A1(_2830_),
    .A2(net126),
    .Y(_2833_),
    .B1(_4288_));
 sg13g2_inv_1 _7847_ (.Y(_2834_),
    .A(_2833_));
 sg13g2_buf_1 _7848_ (.A(_4556_),
    .X(_2835_));
 sg13g2_nand2_1 _7849_ (.Y(_2836_),
    .A(net126),
    .B(net142));
 sg13g2_xnor2_1 _7850_ (.Y(_2837_),
    .A(_1012_),
    .B(_2836_));
 sg13g2_nand2_1 _7851_ (.Y(_2838_),
    .A(net126),
    .B(_4431_));
 sg13g2_nor2_1 _7852_ (.A(_1040_),
    .B(_2838_),
    .Y(_2839_));
 sg13g2_inv_2 _7853_ (.Y(_2840_),
    .A(net126));
 sg13g2_nor3_1 _7854_ (.A(_4495_),
    .B(_1065_),
    .C(_2840_),
    .Y(_2841_));
 sg13g2_a21oi_1 _7855_ (.A1(net126),
    .A2(net160),
    .Y(_2842_),
    .B1(_1066_));
 sg13g2_nor2_1 _7856_ (.A(_2842_),
    .B(_2841_),
    .Y(_2843_));
 sg13g2_nand2_1 _7857_ (.Y(_2844_),
    .A(net126),
    .B(_4413_));
 sg13g2_nor2_1 _7858_ (.A(_1052_),
    .B(_2844_),
    .Y(_2845_));
 sg13g2_nand2_1 _7859_ (.Y(_2846_),
    .A(_2843_),
    .B(_2845_));
 sg13g2_nand2b_1 _7860_ (.Y(_2847_),
    .B(_2846_),
    .A_N(_2841_));
 sg13g2_xnor2_1 _7861_ (.Y(_2848_),
    .A(_1039_),
    .B(_2838_));
 sg13g2_nand2_1 _7862_ (.Y(_2849_),
    .A(_2847_),
    .B(_2848_));
 sg13g2_nand2b_1 _7863_ (.Y(_2850_),
    .B(_2849_),
    .A_N(_2839_));
 sg13g2_a21oi_1 _7864_ (.A1(net126),
    .A2(net152),
    .Y(_2851_),
    .B1(_1081_));
 sg13g2_nand3_1 _7865_ (.B(net152),
    .C(_1081_),
    .A(net126),
    .Y(_2852_));
 sg13g2_nor2b_1 _7866_ (.A(_2851_),
    .B_N(_2852_),
    .Y(_2853_));
 sg13g2_nand2_1 _7867_ (.Y(_2854_),
    .A(_2850_),
    .B(_2853_));
 sg13g2_nand2_1 _7868_ (.Y(_2855_),
    .A(_2854_),
    .B(_2852_));
 sg13g2_xnor2_1 _7869_ (.Y(_2856_),
    .A(_2837_),
    .B(_2855_));
 sg13g2_nor2_1 _7870_ (.A(_2834_),
    .B(_2856_),
    .Y(_2857_));
 sg13g2_inv_2 _7871_ (.Y(_2858_),
    .A(_2856_));
 sg13g2_xor2_1 _7872_ (.B(_2847_),
    .A(_2848_),
    .X(_2859_));
 sg13g2_xnor2_1 _7873_ (.Y(_2860_),
    .A(_2853_),
    .B(_2850_));
 sg13g2_buf_2 _7874_ (.A(_2860_),
    .X(_2861_));
 sg13g2_xor2_1 _7875_ (.B(_2861_),
    .A(_2859_),
    .X(_2862_));
 sg13g2_inv_1 _7876_ (.Y(_2863_),
    .A(_2862_));
 sg13g2_xnor2_1 _7877_ (.Y(_2864_),
    .A(_1051_),
    .B(_2844_));
 sg13g2_xnor2_1 _7878_ (.Y(_2865_),
    .A(_2864_),
    .B(_2861_));
 sg13g2_nand2_1 _7879_ (.Y(_2866_),
    .A(_2863_),
    .B(_2865_));
 sg13g2_xor2_1 _7880_ (.B(_2843_),
    .A(_2845_),
    .X(_2867_));
 sg13g2_xor2_1 _7881_ (.B(_2861_),
    .A(_2867_),
    .X(_2868_));
 sg13g2_nand2_1 _7882_ (.Y(_2869_),
    .A(_2868_),
    .B(_2865_));
 sg13g2_xor2_1 _7883_ (.B(_2861_),
    .A(_2864_),
    .X(_2870_));
 sg13g2_xnor2_1 _7884_ (.Y(_2871_),
    .A(_2867_),
    .B(_2861_));
 sg13g2_nand2_1 _7885_ (.Y(_2872_),
    .A(_2870_),
    .B(_2871_));
 sg13g2_nand3_1 _7886_ (.B(_2869_),
    .C(_2872_),
    .A(_2866_),
    .Y(_2873_));
 sg13g2_xnor2_1 _7887_ (.Y(_2874_),
    .A(_2858_),
    .B(_2873_));
 sg13g2_inv_2 _7888_ (.Y(_2875_),
    .A(_1626_));
 sg13g2_nand2_1 _7889_ (.Y(_2876_),
    .A(_2875_),
    .B(net152));
 sg13g2_xnor2_1 _7890_ (.Y(_2877_),
    .A(net142),
    .B(_2876_));
 sg13g2_a22oi_1 _7891_ (.Y(_2878_),
    .B1(_4350_),
    .B2(_2840_),
    .A2(_2829_),
    .A1(_2877_));
 sg13g2_buf_1 _7892_ (.A(_2878_),
    .X(_2879_));
 sg13g2_nor2_1 _7893_ (.A(_1626_),
    .B(_2830_),
    .Y(_2880_));
 sg13g2_nand2_1 _7894_ (.Y(_2881_),
    .A(_4463_),
    .B(net142));
 sg13g2_nor2_1 _7895_ (.A(_4571_),
    .B(_2881_),
    .Y(_2882_));
 sg13g2_a21o_1 _7896_ (.A2(_2881_),
    .A1(_2880_),
    .B1(_2840_),
    .X(_2883_));
 sg13g2_nor2_1 _7897_ (.A(_2835_),
    .B(net158),
    .Y(_2884_));
 sg13g2_inv_1 _7898_ (.Y(_2885_),
    .A(_2884_));
 sg13g2_nand2_1 _7899_ (.Y(_2886_),
    .A(_2835_),
    .B(net158));
 sg13g2_nor2_1 _7900_ (.A(_2875_),
    .B(_2830_),
    .Y(_2887_));
 sg13g2_inv_1 _7901_ (.Y(_2888_),
    .A(_2887_));
 sg13g2_a21oi_1 _7902_ (.A1(_2885_),
    .A2(_2886_),
    .Y(_2889_),
    .B1(_2888_));
 sg13g2_a221oi_1 _7903_ (.B2(_4571_),
    .C1(_2889_),
    .B1(_2883_),
    .A1(_2880_),
    .Y(_2890_),
    .A2(_2882_));
 sg13g2_buf_1 _7904_ (.A(_2890_),
    .X(_2891_));
 sg13g2_nand2_1 _7905_ (.Y(_2892_),
    .A(_2872_),
    .B(_2862_));
 sg13g2_nand2_1 _7906_ (.Y(_2893_),
    .A(_2892_),
    .B(_2869_));
 sg13g2_xnor2_1 _7907_ (.Y(_2894_),
    .A(_2858_),
    .B(_2893_));
 sg13g2_nor2_1 _7908_ (.A(_2891_),
    .B(_2894_),
    .Y(_2895_));
 sg13g2_a21oi_1 _7909_ (.A1(_2874_),
    .A2(_2879_),
    .Y(_2896_),
    .B1(_2895_));
 sg13g2_nand3_1 _7910_ (.B(_2874_),
    .C(_2879_),
    .A(_2895_),
    .Y(_2897_));
 sg13g2_buf_1 _7911_ (.A(_2897_),
    .X(_2898_));
 sg13g2_nand2b_1 _7912_ (.Y(_2899_),
    .B(_2898_),
    .A_N(_2896_));
 sg13g2_inv_1 _7913_ (.Y(_2900_),
    .A(_2894_));
 sg13g2_nand2_1 _7914_ (.Y(_2901_),
    .A(_2900_),
    .B(_2879_));
 sg13g2_inv_1 _7915_ (.Y(_2902_),
    .A(_2901_));
 sg13g2_inv_1 _7916_ (.Y(_2903_),
    .A(_2891_));
 sg13g2_mux2_1 _7917_ (.A0(_2872_),
    .A1(_2869_),
    .S(_2862_),
    .X(_2904_));
 sg13g2_xnor2_1 _7918_ (.Y(_2905_),
    .A(_2858_),
    .B(_2904_));
 sg13g2_nand3_1 _7919_ (.B(_2903_),
    .C(_2905_),
    .A(_2902_),
    .Y(_2906_));
 sg13g2_buf_1 _7920_ (.A(_2906_),
    .X(_2907_));
 sg13g2_nand2_1 _7921_ (.Y(_2908_),
    .A(_2899_),
    .B(_2907_));
 sg13g2_inv_1 _7922_ (.Y(_2909_),
    .A(_2905_));
 sg13g2_xnor2_1 _7923_ (.Y(_2910_),
    .A(_4342_),
    .B(_2884_));
 sg13g2_a21oi_1 _7924_ (.A1(_4393_),
    .A2(net142),
    .Y(_2911_),
    .B1(_0413_));
 sg13g2_xnor2_1 _7925_ (.Y(_2912_),
    .A(_0410_),
    .B(_2911_));
 sg13g2_nor2_1 _7926_ (.A(_4343_),
    .B(_2832_),
    .Y(_2913_));
 sg13g2_a221oi_1 _7927_ (.B2(_2880_),
    .C1(_2913_),
    .B1(_2912_),
    .A1(_2887_),
    .Y(_2914_),
    .A2(_2910_));
 sg13g2_buf_1 _7928_ (.A(_2914_),
    .X(_2915_));
 sg13g2_nor2b_1 _7929_ (.A(_2909_),
    .B_N(_2915_),
    .Y(_2916_));
 sg13g2_nor2_1 _7930_ (.A(_2907_),
    .B(_2899_),
    .Y(_2917_));
 sg13g2_a21oi_2 _7931_ (.B1(_2917_),
    .Y(_2918_),
    .A2(_2916_),
    .A1(_2908_));
 sg13g2_nor2b_1 _7932_ (.A(_2894_),
    .B_N(_2915_),
    .Y(_2919_));
 sg13g2_a21oi_1 _7933_ (.A1(_2865_),
    .A2(_2871_),
    .Y(_2920_),
    .B1(_2863_));
 sg13g2_xnor2_1 _7934_ (.Y(_2921_),
    .A(_2856_),
    .B(_2920_));
 sg13g2_inv_1 _7935_ (.Y(_2922_),
    .A(_2921_));
 sg13g2_nor2b_1 _7936_ (.A(_2922_),
    .B_N(_2879_),
    .Y(_2923_));
 sg13g2_nand2_1 _7937_ (.Y(_2924_),
    .A(_2874_),
    .B(_2903_));
 sg13g2_inv_1 _7938_ (.Y(_2925_),
    .A(_2880_));
 sg13g2_a21oi_1 _7939_ (.A1(_2881_),
    .A2(_0414_),
    .Y(_2926_),
    .B1(_0411_));
 sg13g2_xnor2_1 _7940_ (.Y(_2927_),
    .A(_0464_),
    .B(_2926_));
 sg13g2_a21oi_1 _7941_ (.A1(_0414_),
    .A2(_4350_),
    .Y(_2928_),
    .B1(_0411_));
 sg13g2_nand2b_1 _7942_ (.Y(_2929_),
    .B(_4576_),
    .A_N(_2928_));
 sg13g2_nand2_1 _7943_ (.Y(_2930_),
    .A(_2928_),
    .B(_4575_));
 sg13g2_nand3_1 _7944_ (.B(_2929_),
    .C(_2930_),
    .A(_2887_),
    .Y(_2931_));
 sg13g2_o21ai_1 _7945_ (.B1(_2931_),
    .Y(_2932_),
    .A1(_2925_),
    .A2(_2927_));
 sg13g2_a21oi_2 _7946_ (.B1(_2932_),
    .Y(_2933_),
    .A2(_2840_),
    .A1(_4575_));
 sg13g2_nand2_1 _7947_ (.Y(_2934_),
    .A(_2905_),
    .B(_2933_));
 sg13g2_xnor2_1 _7948_ (.Y(_2935_),
    .A(_2924_),
    .B(_2934_));
 sg13g2_xor2_1 _7949_ (.B(_2935_),
    .A(_2923_),
    .X(_2936_));
 sg13g2_xnor2_1 _7950_ (.Y(_2937_),
    .A(_2898_),
    .B(_2936_));
 sg13g2_xor2_1 _7951_ (.B(_2937_),
    .A(_2919_),
    .X(_2938_));
 sg13g2_xnor2_1 _7952_ (.Y(_2939_),
    .A(_2918_),
    .B(_2938_));
 sg13g2_xor2_1 _7953_ (.B(_2939_),
    .A(_2857_),
    .X(_2940_));
 sg13g2_nand2_1 _7954_ (.Y(_2941_),
    .A(_2905_),
    .B(_2891_));
 sg13g2_inv_1 _7955_ (.Y(_2942_),
    .A(_2874_));
 sg13g2_o21ai_1 _7956_ (.B1(_2942_),
    .Y(_2943_),
    .A1(_2901_),
    .A2(_2941_));
 sg13g2_o21ai_1 _7957_ (.B1(_2901_),
    .Y(_2944_),
    .A1(_2891_),
    .A2(_2909_));
 sg13g2_nand3_1 _7958_ (.B(_2833_),
    .C(_2944_),
    .A(_2943_),
    .Y(_2945_));
 sg13g2_nor2_1 _7959_ (.A(_2834_),
    .B(_2922_),
    .Y(_2946_));
 sg13g2_xnor2_1 _7960_ (.Y(_2947_),
    .A(_2907_),
    .B(_2899_));
 sg13g2_xor2_1 _7961_ (.B(_2947_),
    .A(_2916_),
    .X(_2948_));
 sg13g2_nor2b_1 _7962_ (.A(_2946_),
    .B_N(_2948_),
    .Y(_2949_));
 sg13g2_nand2b_1 _7963_ (.Y(_2950_),
    .B(_2946_),
    .A_N(_2948_));
 sg13g2_o21ai_1 _7964_ (.B1(_2950_),
    .Y(_2951_),
    .A1(_2945_),
    .A2(_2949_));
 sg13g2_nor2b_1 _7965_ (.A(_2940_),
    .B_N(_2951_),
    .Y(_2952_));
 sg13g2_nand2_1 _7966_ (.Y(_2953_),
    .A(_2936_),
    .B(_2898_));
 sg13g2_nor2_1 _7967_ (.A(_2898_),
    .B(_2936_),
    .Y(_2954_));
 sg13g2_a21oi_1 _7968_ (.A1(_2953_),
    .A2(_2919_),
    .Y(_2955_),
    .B1(_2954_));
 sg13g2_nor2b_1 _7969_ (.A(_2942_),
    .B_N(_2915_),
    .Y(_2956_));
 sg13g2_nand2_1 _7970_ (.Y(_2957_),
    .A(_2934_),
    .B(_2924_));
 sg13g2_nor2_1 _7971_ (.A(_2924_),
    .B(_2934_),
    .Y(_2958_));
 sg13g2_a21oi_1 _7972_ (.A1(_2957_),
    .A2(_2923_),
    .Y(_2959_),
    .B1(_2958_));
 sg13g2_nand2_1 _7973_ (.Y(_2960_),
    .A(_2900_),
    .B(_2933_));
 sg13g2_nand2_1 _7974_ (.Y(_2961_),
    .A(_2921_),
    .B(_2903_));
 sg13g2_nand2_1 _7975_ (.Y(_2962_),
    .A(_2960_),
    .B(_2961_));
 sg13g2_nand2_1 _7976_ (.Y(_2963_),
    .A(_2921_),
    .B(_2933_));
 sg13g2_nand2b_1 _7977_ (.Y(_2964_),
    .B(_2895_),
    .A_N(_2963_));
 sg13g2_nor2b_1 _7978_ (.A(_2856_),
    .B_N(_2879_),
    .Y(_2965_));
 sg13g2_a21oi_1 _7979_ (.A1(_2962_),
    .A2(_2964_),
    .Y(_2966_),
    .B1(_2965_));
 sg13g2_nand3_1 _7980_ (.B(_2964_),
    .C(_2965_),
    .A(_2962_),
    .Y(_2967_));
 sg13g2_nand2b_1 _7981_ (.Y(_2968_),
    .B(_2967_),
    .A_N(_2966_));
 sg13g2_nor2_1 _7982_ (.A(_2959_),
    .B(_2968_),
    .Y(_2969_));
 sg13g2_nand2_1 _7983_ (.Y(_2970_),
    .A(_2968_),
    .B(_2959_));
 sg13g2_nor2b_1 _7984_ (.A(_2969_),
    .B_N(_2970_),
    .Y(_2971_));
 sg13g2_xnor2_1 _7985_ (.Y(_2972_),
    .A(_2956_),
    .B(_2971_));
 sg13g2_xor2_1 _7986_ (.B(_2972_),
    .A(_2955_),
    .X(_2973_));
 sg13g2_nand2_1 _7987_ (.Y(_2974_),
    .A(_2938_),
    .B(_2918_));
 sg13g2_nor2_1 _7988_ (.A(_2918_),
    .B(_2938_),
    .Y(_2975_));
 sg13g2_a21oi_1 _7989_ (.A1(_2974_),
    .A2(_2857_),
    .Y(_2976_),
    .B1(_2975_));
 sg13g2_xnor2_1 _7990_ (.Y(_2977_),
    .A(_2973_),
    .B(_2976_));
 sg13g2_nor2_1 _7991_ (.A(_2955_),
    .B(_2972_),
    .Y(_2978_));
 sg13g2_a21oi_1 _7992_ (.A1(_2970_),
    .A2(_2956_),
    .Y(_2979_),
    .B1(_2969_));
 sg13g2_nor2b_1 _7993_ (.A(_2922_),
    .B_N(_2915_),
    .Y(_2980_));
 sg13g2_nand2_1 _7994_ (.Y(_2981_),
    .A(_2858_),
    .B(_2903_));
 sg13g2_nand2_1 _7995_ (.Y(_2982_),
    .A(_2874_),
    .B(_2933_));
 sg13g2_xnor2_1 _7996_ (.Y(_2983_),
    .A(_2981_),
    .B(_2982_));
 sg13g2_and2_1 _7997_ (.A(_2967_),
    .B(_2964_),
    .X(_2984_));
 sg13g2_nor2_1 _7998_ (.A(_2983_),
    .B(_2984_),
    .Y(_2985_));
 sg13g2_nand2_1 _7999_ (.Y(_2986_),
    .A(_2984_),
    .B(_2983_));
 sg13g2_nor2b_1 _8000_ (.A(_2985_),
    .B_N(_2986_),
    .Y(_2987_));
 sg13g2_xnor2_1 _8001_ (.Y(_2988_),
    .A(_2980_),
    .B(_2987_));
 sg13g2_xnor2_1 _8002_ (.Y(_2989_),
    .A(_2979_),
    .B(_2988_));
 sg13g2_xnor2_1 _8003_ (.Y(_2990_),
    .A(_2978_),
    .B(_2989_));
 sg13g2_nand2_1 _8004_ (.Y(_2991_),
    .A(_2858_),
    .B(_2915_));
 sg13g2_nor2_1 _8005_ (.A(_2981_),
    .B(_2982_),
    .Y(_2992_));
 sg13g2_xor2_1 _8006_ (.B(_2992_),
    .A(_2963_),
    .X(_2993_));
 sg13g2_xor2_1 _8007_ (.B(_2993_),
    .A(_2991_),
    .X(_2994_));
 sg13g2_a21oi_1 _8008_ (.A1(_2986_),
    .A2(_2980_),
    .Y(_2995_),
    .B1(_2985_));
 sg13g2_xnor2_1 _8009_ (.Y(_2996_),
    .A(_2994_),
    .B(_2995_));
 sg13g2_nor2_1 _8010_ (.A(_2979_),
    .B(_2988_),
    .Y(_2997_));
 sg13g2_xor2_1 _8011_ (.B(_2997_),
    .A(_2996_),
    .X(_2998_));
 sg13g2_inv_1 _8012_ (.Y(_2999_),
    .A(_2998_));
 sg13g2_nor2_1 _8013_ (.A(_2991_),
    .B(_2993_),
    .Y(_3000_));
 sg13g2_a21oi_1 _8014_ (.A1(_2921_),
    .A2(_2992_),
    .Y(_3001_),
    .B1(_3000_));
 sg13g2_nor2b_1 _8015_ (.A(_2856_),
    .B_N(_2933_),
    .Y(_3002_));
 sg13g2_nand2_1 _8016_ (.Y(_3003_),
    .A(_3001_),
    .B(_3002_));
 sg13g2_nor2b_1 _8017_ (.A(_2995_),
    .B_N(_2994_),
    .Y(_3004_));
 sg13g2_xnor2_1 _8018_ (.Y(_3005_),
    .A(_3003_),
    .B(_3004_));
 sg13g2_nor2b_1 _8019_ (.A(_2999_),
    .B_N(_3005_),
    .Y(_3006_));
 sg13g2_nand4_1 _8020_ (.B(_2977_),
    .C(_2990_),
    .A(_2952_),
    .Y(_3007_),
    .D(_3006_));
 sg13g2_inv_1 _8021_ (.Y(_3008_),
    .A(_2990_));
 sg13g2_nand2b_1 _8022_ (.Y(_3009_),
    .B(_2973_),
    .A_N(_2976_));
 sg13g2_nand2b_1 _8023_ (.Y(_3010_),
    .B(_2978_),
    .A_N(_2989_));
 sg13g2_o21ai_1 _8024_ (.B1(_3010_),
    .Y(_3011_),
    .A1(_3008_),
    .A2(_3009_));
 sg13g2_nand2_1 _8025_ (.Y(_3012_),
    .A(_3011_),
    .B(_3006_));
 sg13g2_inv_1 _8026_ (.Y(_3013_),
    .A(_3003_));
 sg13g2_and3_1 _8027_ (.X(_3014_),
    .A(_3005_),
    .B(_2997_),
    .C(_2996_));
 sg13g2_a21oi_1 _8028_ (.A1(_3004_),
    .A2(_3013_),
    .Y(_3015_),
    .B1(_3014_));
 sg13g2_nand4_1 _8029_ (.B(_3012_),
    .C(_3001_),
    .A(_3007_),
    .Y(_3016_),
    .D(_3015_));
 sg13g2_inv_1 _8030_ (.Y(_3017_),
    .A(_0068_));
 sg13g2_nor2_1 _8031_ (.A(_3017_),
    .B(_2840_),
    .Y(_3018_));
 sg13g2_inv_1 _8032_ (.Y(_3019_),
    .A(_3018_));
 sg13g2_inv_1 _8033_ (.Y(_3020_),
    .A(_1015_));
 sg13g2_a21oi_2 _8034_ (.B1(_2829_),
    .Y(_3021_),
    .A2(_2826_),
    .A1(_1476_));
 sg13g2_nor2_1 _8035_ (.A(_4432_),
    .B(_3021_),
    .Y(_3022_));
 sg13g2_xnor2_1 _8036_ (.Y(_3023_),
    .A(_3020_),
    .B(_3022_));
 sg13g2_a21oi_1 _8037_ (.A1(_3016_),
    .A2(_3019_),
    .Y(_3024_),
    .B1(_3023_));
 sg13g2_nand3_1 _8038_ (.B(_3019_),
    .C(_3023_),
    .A(_3016_),
    .Y(_3025_));
 sg13g2_nand2b_1 _8039_ (.Y(_3026_),
    .B(_3025_),
    .A_N(_3024_));
 sg13g2_nand2_1 _8040_ (.Y(_3027_),
    .A(_2952_),
    .B(_2977_));
 sg13g2_nand2_1 _8041_ (.Y(_3028_),
    .A(_3027_),
    .B(_3009_));
 sg13g2_nand2_1 _8042_ (.Y(_3029_),
    .A(_3028_),
    .B(_2990_));
 sg13g2_nand2_1 _8043_ (.Y(_3030_),
    .A(_3029_),
    .B(_3010_));
 sg13g2_nand2_1 _8044_ (.Y(_3031_),
    .A(_3030_),
    .B(_2998_));
 sg13g2_a21oi_1 _8045_ (.A1(_2997_),
    .A2(_2996_),
    .Y(_3032_),
    .B1(_3005_));
 sg13g2_nand2_1 _8046_ (.Y(_3033_),
    .A(_3031_),
    .B(_3032_));
 sg13g2_nand3_1 _8047_ (.B(_3005_),
    .C(_2998_),
    .A(_3030_),
    .Y(_3034_));
 sg13g2_nor2_1 _8048_ (.A(_3018_),
    .B(_3014_),
    .Y(_3035_));
 sg13g2_inv_1 _8049_ (.Y(_3036_),
    .A(_1085_));
 sg13g2_o21ai_1 _8050_ (.B1(_3036_),
    .Y(_3037_),
    .A1(_4495_),
    .A2(_3021_));
 sg13g2_inv_1 _8051_ (.Y(_3038_),
    .A(_3021_));
 sg13g2_nand3_1 _8052_ (.B(net160),
    .C(_1085_),
    .A(_3038_),
    .Y(_3039_));
 sg13g2_and2_1 _8053_ (.A(_3037_),
    .B(_3039_),
    .X(_3040_));
 sg13g2_nand4_1 _8054_ (.B(_3034_),
    .C(_3035_),
    .A(_3033_),
    .Y(_3041_),
    .D(_3040_));
 sg13g2_nand2_1 _8055_ (.Y(_3042_),
    .A(_3041_),
    .B(_3039_));
 sg13g2_nand2b_1 _8056_ (.Y(_3043_),
    .B(_3042_),
    .A_N(_3026_));
 sg13g2_inv_1 _8057_ (.Y(_3044_),
    .A(_3040_));
 sg13g2_nand3_1 _8058_ (.B(_3034_),
    .C(_3035_),
    .A(_3033_),
    .Y(_3045_));
 sg13g2_nor2_1 _8059_ (.A(_3044_),
    .B(_3045_),
    .Y(_3046_));
 sg13g2_nor2b_1 _8060_ (.A(_3046_),
    .B_N(_3039_),
    .Y(_3047_));
 sg13g2_nand2_1 _8061_ (.Y(_3048_),
    .A(_3047_),
    .B(_3026_));
 sg13g2_nand2_1 _8062_ (.Y(_3049_),
    .A(_3043_),
    .B(_3048_));
 sg13g2_nand3_1 _8063_ (.B(_2999_),
    .C(_3010_),
    .A(_3029_),
    .Y(_3050_));
 sg13g2_a21oi_1 _8064_ (.A1(_3038_),
    .A2(_4413_),
    .Y(_3051_),
    .B1(_1043_));
 sg13g2_nand3_1 _8065_ (.B(_4413_),
    .C(_1043_),
    .A(_3038_),
    .Y(_3052_));
 sg13g2_nor2b_1 _8066_ (.A(_3051_),
    .B_N(_3052_),
    .Y(_3053_));
 sg13g2_nand4_1 _8067_ (.B(_3050_),
    .C(_3019_),
    .A(_3031_),
    .Y(_3054_),
    .D(_3053_));
 sg13g2_and2_1 _8068_ (.A(_3054_),
    .B(_3052_),
    .X(_3055_));
 sg13g2_buf_1 _8069_ (.A(_3055_),
    .X(_3056_));
 sg13g2_nand2_1 _8070_ (.Y(_3057_),
    .A(_3045_),
    .B(_3044_));
 sg13g2_nand2_1 _8071_ (.Y(_3058_),
    .A(_3057_),
    .B(_3041_));
 sg13g2_xnor2_1 _8072_ (.Y(_3059_),
    .A(_3056_),
    .B(_3058_));
 sg13g2_nor2_1 _8073_ (.A(_3049_),
    .B(_3059_),
    .Y(_3060_));
 sg13g2_nand3_1 _8074_ (.B(_3050_),
    .C(_3019_),
    .A(_3031_),
    .Y(_3061_));
 sg13g2_nand2b_1 _8075_ (.Y(_3062_),
    .B(_3061_),
    .A_N(_3053_));
 sg13g2_inv_1 _8076_ (.Y(_3063_),
    .A(_1055_));
 sg13g2_xnor2_1 _8077_ (.Y(_3064_),
    .A(_2977_),
    .B(_2952_));
 sg13g2_nor2_1 _8078_ (.A(_3063_),
    .B(_3064_),
    .Y(_3065_));
 sg13g2_o21ai_1 _8079_ (.B1(_3019_),
    .Y(_3066_),
    .A1(_1069_),
    .A2(_3065_));
 sg13g2_xnor2_1 _8080_ (.Y(_3067_),
    .A(_3008_),
    .B(_3028_));
 sg13g2_a21oi_1 _8081_ (.A1(_1069_),
    .A2(_3065_),
    .Y(_3068_),
    .B1(_3067_));
 sg13g2_nor2_1 _8082_ (.A(_3066_),
    .B(_3068_),
    .Y(_3069_));
 sg13g2_and3_1 _8083_ (.X(_3070_),
    .A(_3062_),
    .B(_3054_),
    .C(_3069_));
 sg13g2_buf_1 _8084_ (.A(_3070_),
    .X(_3071_));
 sg13g2_nand2_1 _8085_ (.Y(_3072_),
    .A(_3060_),
    .B(_3071_));
 sg13g2_nor2_1 _8086_ (.A(_3056_),
    .B(_3058_),
    .Y(_3073_));
 sg13g2_inv_1 _8087_ (.Y(_3074_),
    .A(_3043_));
 sg13g2_a21oi_1 _8088_ (.A1(_3073_),
    .A2(_3048_),
    .Y(_3075_),
    .B1(_3074_));
 sg13g2_nand2_1 _8089_ (.Y(_3076_),
    .A(_3072_),
    .B(_3075_));
 sg13g2_a21oi_1 _8090_ (.A1(_3038_),
    .A2(net152),
    .Y(_3077_),
    .B1(_1025_));
 sg13g2_nand3_1 _8091_ (.B(net152),
    .C(_1025_),
    .A(_3038_),
    .Y(_3078_));
 sg13g2_nor2b_1 _8092_ (.A(_3077_),
    .B_N(_3078_),
    .Y(_3079_));
 sg13g2_nand2_1 _8093_ (.Y(_3080_),
    .A(_3022_),
    .B(_1015_));
 sg13g2_nand2_1 _8094_ (.Y(_3081_),
    .A(_3025_),
    .B(_3080_));
 sg13g2_xor2_1 _8095_ (.B(_3081_),
    .A(_3079_),
    .X(_3082_));
 sg13g2_nand2_1 _8096_ (.Y(_3083_),
    .A(_3076_),
    .B(_3082_));
 sg13g2_inv_1 _8097_ (.Y(_3084_),
    .A(_3082_));
 sg13g2_nand3_1 _8098_ (.B(_3084_),
    .C(_3075_),
    .A(_3072_),
    .Y(_3085_));
 sg13g2_buf_1 _8099_ (.A(_3085_),
    .X(_3086_));
 sg13g2_nand2_2 _8100_ (.Y(_3087_),
    .A(_3083_),
    .B(_3086_));
 sg13g2_xnor2_1 _8101_ (.Y(_3088_),
    .A(_3071_),
    .B(_3059_));
 sg13g2_inv_2 _8102_ (.Y(_3089_),
    .A(_3088_));
 sg13g2_nand2_1 _8103_ (.Y(_3090_),
    .A(_3058_),
    .B(_3056_));
 sg13g2_a21oi_1 _8104_ (.A1(_3090_),
    .A2(_3071_),
    .Y(_3091_),
    .B1(_3073_));
 sg13g2_xnor2_1 _8105_ (.Y(_3092_),
    .A(_3049_),
    .B(_3091_));
 sg13g2_nor2_1 _8106_ (.A(_3089_),
    .B(_3092_),
    .Y(_3093_));
 sg13g2_nor2b_1 _8107_ (.A(_3087_),
    .B_N(_3093_),
    .Y(_3094_));
 sg13g2_inv_1 _8108_ (.Y(_3095_),
    .A(_3094_));
 sg13g2_nor2_1 _8109_ (.A(_4557_),
    .B(_3021_),
    .Y(_3096_));
 sg13g2_xnor2_1 _8110_ (.Y(_3097_),
    .A(_1099_),
    .B(_3096_));
 sg13g2_xnor2_1 _8111_ (.Y(_3098_),
    .A(_3078_),
    .B(_3097_));
 sg13g2_nand2_1 _8112_ (.Y(_3099_),
    .A(_3062_),
    .B(_3054_));
 sg13g2_nand2_1 _8113_ (.Y(_3100_),
    .A(_3067_),
    .B(_3019_));
 sg13g2_nor2_1 _8114_ (.A(_1070_),
    .B(_3100_),
    .Y(_3101_));
 sg13g2_nor2b_1 _8115_ (.A(_3099_),
    .B_N(_3101_),
    .Y(_3102_));
 sg13g2_a21oi_1 _8116_ (.A1(_3090_),
    .A2(_3102_),
    .Y(_3103_),
    .B1(_3073_));
 sg13g2_inv_1 _8117_ (.Y(_3104_),
    .A(_3103_));
 sg13g2_nor2_1 _8118_ (.A(_3084_),
    .B(_3049_),
    .Y(_3105_));
 sg13g2_nand2_1 _8119_ (.Y(_3106_),
    .A(_3081_),
    .B(_3079_));
 sg13g2_o21ai_1 _8120_ (.B1(_3106_),
    .Y(_3107_),
    .A1(_3043_),
    .A2(_3084_));
 sg13g2_a21oi_1 _8121_ (.A1(_3104_),
    .A2(_3105_),
    .Y(_3108_),
    .B1(_3107_));
 sg13g2_xor2_1 _8122_ (.B(_3099_),
    .A(_3101_),
    .X(_3109_));
 sg13g2_nor2_1 _8123_ (.A(_3109_),
    .B(_3059_),
    .Y(_3110_));
 sg13g2_xnor2_1 _8124_ (.Y(_3111_),
    .A(_1070_),
    .B(_3100_));
 sg13g2_nor4_1 _8125_ (.A(_3063_),
    .B(_3018_),
    .C(_3064_),
    .D(_3111_),
    .Y(_3112_));
 sg13g2_nand3_1 _8126_ (.B(_3105_),
    .C(_3112_),
    .A(_3110_),
    .Y(_3113_));
 sg13g2_nand2_1 _8127_ (.Y(_3114_),
    .A(_3108_),
    .B(_3113_));
 sg13g2_xnor2_1 _8128_ (.Y(_3115_),
    .A(_3098_),
    .B(_3114_));
 sg13g2_nand2_1 _8129_ (.Y(_3116_),
    .A(_3095_),
    .B(_3115_));
 sg13g2_inv_1 _8130_ (.Y(_3117_),
    .A(_3098_));
 sg13g2_xnor2_1 _8131_ (.Y(_3118_),
    .A(_3117_),
    .B(_3114_));
 sg13g2_nand2_1 _8132_ (.Y(_3119_),
    .A(_3118_),
    .B(_3094_));
 sg13g2_nand2_1 _8133_ (.Y(_3120_),
    .A(_1632_),
    .B(_1631_));
 sg13g2_inv_1 _8134_ (.Y(_3121_),
    .A(_3120_));
 sg13g2_inv_1 _8135_ (.Y(_3122_),
    .A(\i_display.in_line ));
 sg13g2_nor4_1 _8136_ (.A(_1632_),
    .B(_1631_),
    .C(net144),
    .D(net156),
    .Y(_3123_));
 sg13g2_inv_1 _8137_ (.Y(_3124_),
    .A(_3123_));
 sg13g2_nor2_2 _8138_ (.A(_3122_),
    .B(_3124_),
    .Y(_3125_));
 sg13g2_nand2_1 _8139_ (.Y(_3126_),
    .A(_2827_),
    .B(net156));
 sg13g2_xnor2_1 _8140_ (.Y(_3127_),
    .A(_0026_),
    .B(_3126_));
 sg13g2_nor2_1 _8141_ (.A(_3123_),
    .B(_3127_),
    .Y(_3128_));
 sg13g2_nor3_1 _8142_ (.A(_3121_),
    .B(_3125_),
    .C(_3128_),
    .Y(_3129_));
 sg13g2_nand3_1 _8143_ (.B(_3119_),
    .C(_3129_),
    .A(_3116_),
    .Y(_3130_));
 sg13g2_nor2_1 _8144_ (.A(_1054_),
    .B(_1052_),
    .Y(_3131_));
 sg13g2_inv_1 _8145_ (.Y(_3132_),
    .A(_3131_));
 sg13g2_inv_1 _8146_ (.Y(_3133_),
    .A(_1025_));
 sg13g2_nand2_1 _8147_ (.Y(_3134_),
    .A(_1041_),
    .B(_1083_));
 sg13g2_inv_1 _8148_ (.Y(_3135_),
    .A(_3134_));
 sg13g2_nor2_1 _8149_ (.A(_1013_),
    .B(_3135_),
    .Y(_3136_));
 sg13g2_nor2_1 _8150_ (.A(_3133_),
    .B(_3136_),
    .Y(_3137_));
 sg13g2_nor2_1 _8151_ (.A(_1099_),
    .B(_3137_),
    .Y(_3138_));
 sg13g2_inv_1 _8152_ (.Y(_3139_),
    .A(_3138_));
 sg13g2_nor2_1 _8153_ (.A(_1005_),
    .B(_3139_),
    .Y(_3140_));
 sg13g2_inv_1 _8154_ (.Y(_3141_),
    .A(_3140_));
 sg13g2_nand2_1 _8155_ (.Y(_3142_),
    .A(_3141_),
    .B(_0982_));
 sg13g2_nand2_1 _8156_ (.Y(_3143_),
    .A(_3142_),
    .B(_0713_));
 sg13g2_nand3_1 _8157_ (.B(_0982_),
    .C(_0714_),
    .A(_3141_),
    .Y(_3144_));
 sg13g2_nand2_1 _8158_ (.Y(_3145_),
    .A(_3143_),
    .B(_3144_));
 sg13g2_buf_1 _8159_ (.A(_3145_),
    .X(_3146_));
 sg13g2_nor2_1 _8160_ (.A(_1053_),
    .B(_1068_),
    .Y(_3147_));
 sg13g2_nor2_1 _8161_ (.A(_1152_),
    .B(_3147_),
    .Y(_3148_));
 sg13g2_nor3_1 _8162_ (.A(net150),
    .B(_3148_),
    .C(net81),
    .Y(_3149_));
 sg13g2_a21oi_1 _8163_ (.A1(_1069_),
    .A2(net81),
    .Y(_3150_),
    .B1(_3149_));
 sg13g2_nor2_1 _8164_ (.A(_1011_),
    .B(_1021_),
    .Y(_3151_));
 sg13g2_nand2_1 _8165_ (.Y(_3152_),
    .A(_3151_),
    .B(_1097_));
 sg13g2_nand2_1 _8166_ (.Y(_3153_),
    .A(_3152_),
    .B(_1002_));
 sg13g2_nor2_1 _8167_ (.A(_1160_),
    .B(_3153_),
    .Y(_3154_));
 sg13g2_or2_1 _8168_ (.X(_3155_),
    .B(_3154_),
    .A(_0710_));
 sg13g2_nand2_1 _8169_ (.Y(_3156_),
    .A(_3154_),
    .B(_0710_));
 sg13g2_nand2_1 _8170_ (.Y(_3157_),
    .A(_3155_),
    .B(_3156_));
 sg13g2_inv_2 _8171_ (.Y(_3158_),
    .A(_3157_));
 sg13g2_nor2_1 _8172_ (.A(net124),
    .B(_1485_),
    .Y(_3159_));
 sg13g2_inv_1 _8173_ (.Y(_3160_),
    .A(_3159_));
 sg13g2_nor2_1 _8174_ (.A(net131),
    .B(_3158_),
    .Y(_3161_));
 sg13g2_a22oi_1 _8175_ (.Y(_3162_),
    .B1(_3160_),
    .B2(_3161_),
    .A2(_3158_),
    .A1(_1066_));
 sg13g2_xnor2_1 _8176_ (.Y(_3163_),
    .A(_3150_),
    .B(_3162_));
 sg13g2_nor2_1 _8177_ (.A(_3132_),
    .B(_3163_),
    .Y(_3164_));
 sg13g2_inv_1 _8178_ (.Y(_3165_),
    .A(_3164_));
 sg13g2_nand2_1 _8179_ (.Y(_3166_),
    .A(_3163_),
    .B(_3132_));
 sg13g2_nand2_2 _8180_ (.Y(_3167_),
    .A(_3165_),
    .B(_3166_));
 sg13g2_inv_1 _8181_ (.Y(_3168_),
    .A(_3167_));
 sg13g2_inv_2 _8182_ (.Y(_3169_),
    .A(_1634_));
 sg13g2_a21oi_1 _8183_ (.A1(_3168_),
    .A2(_3125_),
    .Y(_3170_),
    .B1(_3169_));
 sg13g2_nand2_1 _8184_ (.Y(_3171_),
    .A(_3130_),
    .B(_3170_));
 sg13g2_inv_1 _8185_ (.Y(_3172_),
    .A(_3092_));
 sg13g2_nand2_1 _8186_ (.Y(_3173_),
    .A(_3172_),
    .B(_3089_));
 sg13g2_nor2_1 _8187_ (.A(_3173_),
    .B(_3087_),
    .Y(_3174_));
 sg13g2_xnor2_1 _8188_ (.Y(_3175_),
    .A(_3174_),
    .B(_3115_));
 sg13g2_nor2_2 _8189_ (.A(_3122_),
    .B(_3120_),
    .Y(_3176_));
 sg13g2_a21oi_1 _8190_ (.A1(_3128_),
    .A2(_3120_),
    .Y(_3177_),
    .B1(_3176_));
 sg13g2_inv_1 _8191_ (.Y(_3178_),
    .A(_3177_));
 sg13g2_nand2_1 _8192_ (.Y(_3179_),
    .A(_3175_),
    .B(_3178_));
 sg13g2_nor2b_1 _8193_ (.A(_3171_),
    .B_N(_3179_),
    .Y(_3180_));
 sg13g2_nor2_1 _8194_ (.A(_3150_),
    .B(_3162_),
    .Y(_3181_));
 sg13g2_inv_1 _8195_ (.Y(_3182_),
    .A(_1043_));
 sg13g2_o21ai_1 _8196_ (.B1(_1042_),
    .Y(_3183_),
    .A1(_1069_),
    .A2(_1055_));
 sg13g2_nor2_1 _8197_ (.A(_1053_),
    .B(_1067_),
    .Y(_3184_));
 sg13g2_inv_1 _8198_ (.Y(_3185_),
    .A(_3184_));
 sg13g2_nor2_1 _8199_ (.A(_3185_),
    .B(_3182_),
    .Y(_3186_));
 sg13g2_nor2_1 _8200_ (.A(_3186_),
    .B(_3146_),
    .Y(_3187_));
 sg13g2_a22oi_1 _8201_ (.Y(_3188_),
    .B1(_3183_),
    .B2(_3187_),
    .A2(net81),
    .A1(_3182_));
 sg13g2_nand2_1 _8202_ (.Y(_3189_),
    .A(_1039_),
    .B(_2025_));
 sg13g2_o21ai_1 _8203_ (.B1(_0707_),
    .Y(_3190_),
    .A1(_4230_),
    .A2(_2025_));
 sg13g2_nor2_1 _8204_ (.A(_3190_),
    .B(_3158_),
    .Y(_3191_));
 sg13g2_a22oi_1 _8205_ (.Y(_3192_),
    .B1(_3189_),
    .B2(_3191_),
    .A2(_3158_),
    .A1(_1039_));
 sg13g2_xor2_1 _8206_ (.B(_3192_),
    .A(_3188_),
    .X(_3193_));
 sg13g2_o21ai_1 _8207_ (.B1(_3193_),
    .Y(_3194_),
    .A1(_3181_),
    .A2(_3164_));
 sg13g2_nor2_1 _8208_ (.A(_3181_),
    .B(_3164_),
    .Y(_3195_));
 sg13g2_nand2b_1 _8209_ (.Y(_3196_),
    .B(_3195_),
    .A_N(_3193_));
 sg13g2_nand2_1 _8210_ (.Y(_3197_),
    .A(_3194_),
    .B(_3196_));
 sg13g2_buf_2 _8211_ (.A(_3197_),
    .X(_3198_));
 sg13g2_inv_2 _8212_ (.Y(_3199_),
    .A(_3198_));
 sg13g2_xnor2_1 _8213_ (.Y(_3200_),
    .A(_1096_),
    .B(_3151_));
 sg13g2_and3_1 _8214_ (.X(_3201_),
    .A(_3190_),
    .B(_1011_),
    .C(_1082_));
 sg13g2_buf_1 _8215_ (.A(_3201_),
    .X(_3202_));
 sg13g2_xor2_1 _8216_ (.B(_1021_),
    .A(_1011_),
    .X(_3203_));
 sg13g2_a21oi_1 _8217_ (.A1(_3202_),
    .A2(_3203_),
    .Y(_3204_),
    .B1(_3158_));
 sg13g2_xor2_1 _8218_ (.B(_3204_),
    .A(_3200_),
    .X(_3205_));
 sg13g2_nor2_1 _8219_ (.A(net150),
    .B(_3136_),
    .Y(_3206_));
 sg13g2_a21oi_1 _8220_ (.A1(_1229_),
    .A2(_3206_),
    .Y(_3207_),
    .B1(_3138_));
 sg13g2_inv_1 _8221_ (.Y(_3208_),
    .A(_3206_));
 sg13g2_a21oi_1 _8222_ (.A1(_1013_),
    .A2(_3135_),
    .Y(_3209_),
    .B1(_3208_));
 sg13g2_xnor2_1 _8223_ (.Y(_3210_),
    .A(_1085_),
    .B(_1043_));
 sg13g2_nand3_1 _8224_ (.B(_3186_),
    .C(_3210_),
    .A(_3209_),
    .Y(_3211_));
 sg13g2_xnor2_1 _8225_ (.Y(_3212_),
    .A(_1025_),
    .B(_3206_));
 sg13g2_nand2b_1 _8226_ (.Y(_3213_),
    .B(_3212_),
    .A_N(_3211_));
 sg13g2_xnor2_1 _8227_ (.Y(_3214_),
    .A(_3207_),
    .B(_3213_));
 sg13g2_nor2_1 _8228_ (.A(net81),
    .B(_3214_),
    .Y(_3215_));
 sg13g2_a21oi_1 _8229_ (.A1(net81),
    .A2(_3207_),
    .Y(_3216_),
    .B1(_3215_));
 sg13g2_xnor2_1 _8230_ (.Y(_3217_),
    .A(_3205_),
    .B(_3216_));
 sg13g2_inv_1 _8231_ (.Y(_3218_),
    .A(net81));
 sg13g2_nand2_1 _8232_ (.Y(_3219_),
    .A(_3218_),
    .B(_3211_));
 sg13g2_xnor2_1 _8233_ (.Y(_3220_),
    .A(_3212_),
    .B(_3219_));
 sg13g2_nor2_1 _8234_ (.A(_3202_),
    .B(_3158_),
    .Y(_3221_));
 sg13g2_xor2_1 _8235_ (.B(_3221_),
    .A(_3203_),
    .X(_3222_));
 sg13g2_a21oi_1 _8236_ (.A1(_3186_),
    .A2(_3210_),
    .Y(_3223_),
    .B1(_3146_));
 sg13g2_xor2_1 _8237_ (.B(_3223_),
    .A(_3209_),
    .X(_3224_));
 sg13g2_a221oi_1 _8238_ (.B2(_3156_),
    .C1(net131),
    .B1(_3155_),
    .A1(_1491_),
    .Y(_3225_),
    .A2(_2590_));
 sg13g2_nor2_1 _8239_ (.A(_1012_),
    .B(_3225_),
    .Y(_3226_));
 sg13g2_a21oi_1 _8240_ (.A1(_1010_),
    .A2(_3225_),
    .Y(_3227_),
    .B1(_3226_));
 sg13g2_inv_1 _8241_ (.Y(_3228_),
    .A(_3227_));
 sg13g2_xnor2_1 _8242_ (.Y(_3229_),
    .A(_3210_),
    .B(_3187_));
 sg13g2_inv_1 _8243_ (.Y(_3230_),
    .A(_3229_));
 sg13g2_xnor2_1 _8244_ (.Y(_3231_),
    .A(_1082_),
    .B(_3191_));
 sg13g2_inv_1 _8245_ (.Y(_3232_),
    .A(_3231_));
 sg13g2_xnor2_1 _8246_ (.Y(_3233_),
    .A(_3229_),
    .B(_3231_));
 sg13g2_nor2_1 _8247_ (.A(_3188_),
    .B(_3192_),
    .Y(_3234_));
 sg13g2_nor2b_1 _8248_ (.A(_3234_),
    .B_N(_3194_),
    .Y(_3235_));
 sg13g2_or2_1 _8249_ (.X(_3236_),
    .B(_3235_),
    .A(_3233_));
 sg13g2_o21ai_1 _8250_ (.B1(_3236_),
    .Y(_3237_),
    .A1(_3230_),
    .A2(_3232_));
 sg13g2_xnor2_1 _8251_ (.Y(_3238_),
    .A(_3224_),
    .B(_3227_));
 sg13g2_nand2_1 _8252_ (.Y(_3239_),
    .A(_3237_),
    .B(_3238_));
 sg13g2_o21ai_1 _8253_ (.B1(_3239_),
    .Y(_3240_),
    .A1(_3224_),
    .A2(_3228_));
 sg13g2_xor2_1 _8254_ (.B(_3222_),
    .A(_3220_),
    .X(_3241_));
 sg13g2_nand2_1 _8255_ (.Y(_3242_),
    .A(_3240_),
    .B(_3241_));
 sg13g2_o21ai_1 _8256_ (.B1(_3242_),
    .Y(_3243_),
    .A1(_3220_),
    .A2(_3222_));
 sg13g2_or2_1 _8257_ (.X(_3244_),
    .B(_3243_),
    .A(_3217_));
 sg13g2_nand2_1 _8258_ (.Y(_3245_),
    .A(_3243_),
    .B(_3217_));
 sg13g2_nand2_1 _8259_ (.Y(_3246_),
    .A(_3244_),
    .B(_3245_));
 sg13g2_buf_2 _8260_ (.A(_3246_),
    .X(_3247_));
 sg13g2_inv_1 _8261_ (.Y(_3248_),
    .A(_3247_));
 sg13g2_xnor2_1 _8262_ (.Y(_3249_),
    .A(_1005_),
    .B(_3138_));
 sg13g2_nor2_1 _8263_ (.A(_1099_),
    .B(_3213_),
    .Y(_3250_));
 sg13g2_nor2_1 _8264_ (.A(net81),
    .B(_3250_),
    .Y(_3251_));
 sg13g2_xnor2_1 _8265_ (.Y(_3252_),
    .A(_3249_),
    .B(_3251_));
 sg13g2_xor2_1 _8266_ (.B(_3152_),
    .A(_1002_),
    .X(_3253_));
 sg13g2_nand3_1 _8267_ (.B(_3200_),
    .C(_3203_),
    .A(_3202_),
    .Y(_3254_));
 sg13g2_nor2_1 _8268_ (.A(_3253_),
    .B(_3254_),
    .Y(_3255_));
 sg13g2_inv_1 _8269_ (.Y(_3256_),
    .A(_3255_));
 sg13g2_a21oi_1 _8270_ (.A1(_3253_),
    .A2(_3254_),
    .Y(_3257_),
    .B1(_3158_));
 sg13g2_a22oi_1 _8271_ (.Y(_3258_),
    .B1(_3256_),
    .B2(_3257_),
    .A2(_3253_),
    .A1(_3158_));
 sg13g2_xnor2_1 _8272_ (.Y(_3259_),
    .A(_3252_),
    .B(_3258_));
 sg13g2_inv_1 _8273_ (.Y(_3260_),
    .A(_3216_));
 sg13g2_o21ai_1 _8274_ (.B1(_3245_),
    .Y(_3261_),
    .A1(_3205_),
    .A2(_3260_));
 sg13g2_xnor2_1 _8275_ (.Y(_3262_),
    .A(_3259_),
    .B(_3261_));
 sg13g2_xnor2_1 _8276_ (.Y(_3263_),
    .A(_0310_),
    .B(_3262_));
 sg13g2_a21oi_1 _8277_ (.A1(_4575_),
    .A2(_3248_),
    .Y(_3264_),
    .B1(_3263_));
 sg13g2_nor2_1 _8278_ (.A(_4393_),
    .B(_3198_),
    .Y(_3265_));
 sg13g2_nor2_1 _8279_ (.A(_4288_),
    .B(_3199_),
    .Y(_3266_));
 sg13g2_or2_1 _8280_ (.X(_3267_),
    .B(_3240_),
    .A(_3241_));
 sg13g2_nand2_1 _8281_ (.Y(_3268_),
    .A(_3267_),
    .B(_3242_));
 sg13g2_buf_1 _8282_ (.A(_3268_),
    .X(_3269_));
 sg13g2_nor2_1 _8283_ (.A(net159),
    .B(net66),
    .Y(_3270_));
 sg13g2_nand2_1 _8284_ (.Y(_3271_),
    .A(net66),
    .B(_0410_));
 sg13g2_or2_1 _8285_ (.X(_3272_),
    .B(_3237_),
    .A(_3238_));
 sg13g2_nand2_1 _8286_ (.Y(_3273_),
    .A(_3272_),
    .B(_3239_));
 sg13g2_buf_2 _8287_ (.A(_3273_),
    .X(_3274_));
 sg13g2_xnor2_1 _8288_ (.Y(_3275_),
    .A(net161),
    .B(_3274_));
 sg13g2_nand3b_1 _8289_ (.B(_3271_),
    .C(_3275_),
    .Y(_3276_),
    .A_N(_3270_));
 sg13g2_inv_1 _8290_ (.Y(_3277_),
    .A(_3276_));
 sg13g2_nand2_1 _8291_ (.Y(_3278_),
    .A(_3235_),
    .B(_3233_));
 sg13g2_nand2_1 _8292_ (.Y(_3279_),
    .A(_3236_),
    .B(_3278_));
 sg13g2_buf_2 _8293_ (.A(_3279_),
    .X(_3280_));
 sg13g2_xnor2_1 _8294_ (.Y(_3281_),
    .A(_4350_),
    .B(_3280_));
 sg13g2_nand2_1 _8295_ (.Y(_3282_),
    .A(_3277_),
    .B(_3281_));
 sg13g2_nor3_1 _8296_ (.A(_3265_),
    .B(_3266_),
    .C(_3282_),
    .Y(_3283_));
 sg13g2_nor2_1 _8297_ (.A(_4575_),
    .B(_3248_),
    .Y(_3284_));
 sg13g2_inv_1 _8298_ (.Y(_3285_),
    .A(_3284_));
 sg13g2_xnor2_1 _8299_ (.Y(_3286_),
    .A(_1055_),
    .B(_1051_));
 sg13g2_xnor2_1 _8300_ (.Y(_3287_),
    .A(_4283_),
    .B(_3286_));
 sg13g2_xnor2_1 _8301_ (.Y(_3288_),
    .A(_4266_),
    .B(_3167_));
 sg13g2_nor2_1 _8302_ (.A(_3287_),
    .B(_3288_),
    .Y(_3289_));
 sg13g2_and4_1 _8303_ (.A(_3264_),
    .B(_3283_),
    .C(_3285_),
    .D(_3289_),
    .X(_3290_));
 sg13g2_inv_1 _8304_ (.Y(_3291_),
    .A(_3288_));
 sg13g2_o21ai_1 _8305_ (.B1(_3291_),
    .Y(_3292_),
    .A1(net160),
    .A2(_3286_));
 sg13g2_o21ai_1 _8306_ (.B1(_3292_),
    .Y(_3293_),
    .A1(_4432_),
    .A2(_3168_));
 sg13g2_nand2_1 _8307_ (.Y(_3294_),
    .A(_3283_),
    .B(_3293_));
 sg13g2_a22oi_1 _8308_ (.Y(_3295_),
    .B1(_3266_),
    .B2(_3281_),
    .A2(_3280_),
    .A1(net142));
 sg13g2_nand2b_1 _8309_ (.Y(_3296_),
    .B(_3277_),
    .A_N(_3295_));
 sg13g2_nand2_1 _8310_ (.Y(_3297_),
    .A(_3274_),
    .B(net158));
 sg13g2_a21o_1 _8311_ (.A2(_3297_),
    .A1(_3271_),
    .B1(_3270_),
    .X(_3298_));
 sg13g2_nand4_1 _8312_ (.B(_3285_),
    .C(_3296_),
    .A(_3294_),
    .Y(_3299_),
    .D(_3298_));
 sg13g2_a22oi_1 _8313_ (.Y(_3300_),
    .B1(_3264_),
    .B2(_3299_),
    .A2(_3262_),
    .A1(_0440_));
 sg13g2_xnor2_1 _8314_ (.Y(_3301_),
    .A(_0980_),
    .B(_3153_));
 sg13g2_nand2_1 _8315_ (.Y(_3302_),
    .A(_3256_),
    .B(_3157_));
 sg13g2_xor2_1 _8316_ (.B(_3302_),
    .A(_3301_),
    .X(_3303_));
 sg13g2_xnor2_1 _8317_ (.Y(_3304_),
    .A(_0982_),
    .B(_3140_));
 sg13g2_inv_1 _8318_ (.Y(_3305_),
    .A(_3304_));
 sg13g2_a21oi_1 _8319_ (.A1(_3250_),
    .A2(_3249_),
    .Y(_3306_),
    .B1(net81));
 sg13g2_xnor2_1 _8320_ (.Y(_3307_),
    .A(_3305_),
    .B(_3306_));
 sg13g2_xor2_1 _8321_ (.B(_3307_),
    .A(_3303_),
    .X(_3308_));
 sg13g2_nor2b_1 _8322_ (.A(_3258_),
    .B_N(_3252_),
    .Y(_3309_));
 sg13g2_a21o_1 _8323_ (.A2(_3259_),
    .A1(_3261_),
    .B1(_3309_),
    .X(_3310_));
 sg13g2_xnor2_1 _8324_ (.Y(_3311_),
    .A(_3308_),
    .B(_3310_));
 sg13g2_nand2_1 _8325_ (.Y(_3312_),
    .A(_3311_),
    .B(_0367_));
 sg13g2_o21ai_1 _8326_ (.B1(_3312_),
    .Y(_3313_),
    .A1(_3290_),
    .A2(_3300_));
 sg13g2_nand2_1 _8327_ (.Y(_3314_),
    .A(_3310_),
    .B(_3308_));
 sg13g2_nand2_1 _8328_ (.Y(_3315_),
    .A(_3307_),
    .B(_3303_));
 sg13g2_nand3_1 _8329_ (.B(_3255_),
    .C(_3301_),
    .A(_3157_),
    .Y(_3316_));
 sg13g2_nand4_1 _8330_ (.B(_3218_),
    .C(_3305_),
    .A(_3250_),
    .Y(_3317_),
    .D(_3249_));
 sg13g2_xnor2_1 _8331_ (.Y(_3318_),
    .A(_3316_),
    .B(_3317_));
 sg13g2_nand3_1 _8332_ (.B(_3315_),
    .C(_3318_),
    .A(_3314_),
    .Y(_3319_));
 sg13g2_o21ai_1 _8333_ (.B1(_1631_),
    .Y(_3320_),
    .A1(_0367_),
    .A2(_3311_));
 sg13g2_nor2_1 _8334_ (.A(_3319_),
    .B(_3320_),
    .Y(_3321_));
 sg13g2_nand2_2 _8335_ (.Y(_3322_),
    .A(_3313_),
    .B(_3321_));
 sg13g2_a21oi_1 _8336_ (.A1(\i_display.frame_crotchet[1] ),
    .A2(_3199_),
    .Y(_3323_),
    .B1(_3322_));
 sg13g2_a21oi_1 _8337_ (.A1(_3122_),
    .A2(_0024_),
    .Y(_3324_),
    .B1(_1632_));
 sg13g2_nand2_1 _8338_ (.Y(_3325_),
    .A(_3322_),
    .B(_3324_));
 sg13g2_nor2_1 _8339_ (.A(_3262_),
    .B(_3311_),
    .Y(_3326_));
 sg13g2_nand2_1 _8340_ (.Y(_3327_),
    .A(_3247_),
    .B(net66));
 sg13g2_a21oi_1 _8341_ (.A1(_3326_),
    .A2(_3327_),
    .Y(_3328_),
    .B1(_3319_));
 sg13g2_o21ai_1 _8342_ (.B1(_1632_),
    .Y(_3329_),
    .A1(_1631_),
    .A2(_3328_));
 sg13g2_nand3b_1 _8343_ (.B(_3325_),
    .C(_3329_),
    .Y(_3330_),
    .A_N(_3323_));
 sg13g2_nand2_1 _8344_ (.Y(_3331_),
    .A(_4494_),
    .B(net144));
 sg13g2_xor2_1 _8345_ (.B(_3167_),
    .A(_3331_),
    .X(_3332_));
 sg13g2_nand2_1 _8346_ (.Y(_3333_),
    .A(_3328_),
    .B(_2827_));
 sg13g2_nor2b_1 _8347_ (.A(_3333_),
    .B_N(\i_display.frame_crotchet[1] ),
    .Y(_3334_));
 sg13g2_nand2_1 _8348_ (.Y(_3335_),
    .A(_3167_),
    .B(_4283_));
 sg13g2_xnor2_1 _8349_ (.Y(_3336_),
    .A(_4265_),
    .B(_3198_));
 sg13g2_xor2_1 _8350_ (.B(_3336_),
    .A(_3335_),
    .X(_3337_));
 sg13g2_a221oi_1 _8351_ (.B2(_3337_),
    .C1(_1634_),
    .B1(_3334_),
    .A1(_3176_),
    .Y(_3338_),
    .A2(_3332_));
 sg13g2_a21oi_1 _8352_ (.A1(_3330_),
    .A2(_3338_),
    .Y(_3339_),
    .B1(net127));
 sg13g2_nor2b_1 _8353_ (.A(_3180_),
    .B_N(_3339_),
    .Y(_0106_));
 sg13g2_nand3_1 _8354_ (.B(_3119_),
    .C(_3178_),
    .A(_3116_),
    .Y(_3340_));
 sg13g2_nor2_1 _8355_ (.A(_0026_),
    .B(_3124_),
    .Y(_3341_));
 sg13g2_a21oi_1 _8356_ (.A1(_3198_),
    .A2(_3341_),
    .Y(_3342_),
    .B1(_3169_));
 sg13g2_nand2_1 _8357_ (.Y(_3343_),
    .A(_3337_),
    .B(net144));
 sg13g2_o21ai_1 _8358_ (.B1(_3343_),
    .Y(_3344_),
    .A1(net144),
    .A2(_3198_));
 sg13g2_nand2_1 _8359_ (.Y(_3345_),
    .A(_3336_),
    .B(_3335_));
 sg13g2_o21ai_1 _8360_ (.B1(_3345_),
    .Y(_3346_),
    .A1(_4431_),
    .A2(_3198_));
 sg13g2_xnor2_1 _8361_ (.Y(_3347_),
    .A(_4288_),
    .B(_3280_));
 sg13g2_xor2_1 _8362_ (.B(_3347_),
    .A(_3346_),
    .X(_3348_));
 sg13g2_inv_1 _8363_ (.Y(_3349_),
    .A(_3280_));
 sg13g2_nand3_1 _8364_ (.B(_3349_),
    .C(_3321_),
    .A(_3313_),
    .Y(_3350_));
 sg13g2_nor3_1 _8365_ (.A(_0065_),
    .B(_1632_),
    .C(_3350_),
    .Y(_3351_));
 sg13g2_a221oi_1 _8366_ (.B2(_3348_),
    .C1(_3351_),
    .B1(_3334_),
    .A1(_3176_),
    .Y(_3352_),
    .A2(_3344_));
 sg13g2_a21o_1 _8367_ (.A2(_3169_),
    .A1(_3352_),
    .B1(_2634_),
    .X(_3353_));
 sg13g2_a21oi_1 _8368_ (.A1(_3340_),
    .A2(_3342_),
    .Y(_0107_),
    .B1(_3353_));
 sg13g2_inv_1 _8369_ (.Y(_3354_),
    .A(_3087_));
 sg13g2_o21ai_1 _8370_ (.B1(_3118_),
    .Y(_3355_),
    .A1(_3354_),
    .A2(_3172_));
 sg13g2_a21oi_1 _8371_ (.A1(_3087_),
    .A2(_3089_),
    .Y(_3356_),
    .B1(_3177_));
 sg13g2_inv_1 _8372_ (.Y(_3357_),
    .A(_3125_));
 sg13g2_xnor2_1 _8373_ (.Y(_3358_),
    .A(_3199_),
    .B(_3280_));
 sg13g2_o21ai_1 _8374_ (.B1(_1634_),
    .Y(_3359_),
    .A1(_3357_),
    .A2(_3358_));
 sg13g2_a21oi_1 _8375_ (.A1(_3355_),
    .A2(_3356_),
    .Y(_3360_),
    .B1(_3359_));
 sg13g2_nand3_1 _8376_ (.B(_3087_),
    .C(_3092_),
    .A(_3115_),
    .Y(_3361_));
 sg13g2_nand2_1 _8377_ (.Y(_3362_),
    .A(_3092_),
    .B(_3089_));
 sg13g2_o21ai_1 _8378_ (.B1(_3118_),
    .Y(_3363_),
    .A1(_3354_),
    .A2(_3362_));
 sg13g2_nand3_1 _8379_ (.B(_3363_),
    .C(_3129_),
    .A(_3361_),
    .Y(_3364_));
 sg13g2_nand2_1 _8380_ (.Y(_3365_),
    .A(_3199_),
    .B(net144));
 sg13g2_nand2b_1 _8381_ (.Y(_3366_),
    .B(\i_display.in_line ),
    .A_N(_0024_));
 sg13g2_nand2b_1 _8382_ (.Y(_3367_),
    .B(_3122_),
    .A_N(_0025_));
 sg13g2_nand4_1 _8383_ (.B(_2826_),
    .C(_3366_),
    .A(_3322_),
    .Y(_3368_),
    .D(_3367_));
 sg13g2_buf_1 _8384_ (.A(_3368_),
    .X(_3369_));
 sg13g2_o21ai_1 _8385_ (.B1(_3369_),
    .Y(_3370_),
    .A1(_3322_),
    .A2(_3365_));
 sg13g2_nand2_1 _8386_ (.Y(_3371_),
    .A(_3370_),
    .B(_2826_));
 sg13g2_inv_1 _8387_ (.Y(_3372_),
    .A(_3333_));
 sg13g2_nand2b_1 _8388_ (.Y(_3373_),
    .B(_3372_),
    .A_N(_3343_));
 sg13g2_nor2_1 _8389_ (.A(net144),
    .B(_3280_),
    .Y(_3374_));
 sg13g2_inv_1 _8390_ (.Y(_3375_),
    .A(_3348_));
 sg13g2_nor2_1 _8391_ (.A(_2875_),
    .B(_3375_),
    .Y(_3376_));
 sg13g2_o21ai_1 _8392_ (.B1(_3176_),
    .Y(_3377_),
    .A1(_3374_),
    .A2(_3376_));
 sg13g2_nand3_1 _8393_ (.B(_3373_),
    .C(_3377_),
    .A(_3371_),
    .Y(_3378_));
 sg13g2_o21ai_1 _8394_ (.B1(net134),
    .Y(_3379_),
    .A1(_1634_),
    .A2(_3378_));
 sg13g2_a21oi_1 _8395_ (.A1(_3360_),
    .A2(_3364_),
    .Y(_0108_),
    .B1(_3379_));
 sg13g2_nand3_1 _8396_ (.B(_3363_),
    .C(_3178_),
    .A(_3361_),
    .Y(_3380_));
 sg13g2_nor2_1 _8397_ (.A(_3199_),
    .B(_3349_),
    .Y(_3381_));
 sg13g2_xnor2_1 _8398_ (.Y(_3382_),
    .A(_3381_),
    .B(_3274_));
 sg13g2_a21oi_1 _8399_ (.A1(_3382_),
    .A2(_3125_),
    .Y(_3383_),
    .B1(_3169_));
 sg13g2_o21ai_1 _8400_ (.B1(_3369_),
    .Y(_3384_),
    .A1(_2875_),
    .A2(_3350_));
 sg13g2_nand2_1 _8401_ (.Y(_3385_),
    .A(_3384_),
    .B(_2826_));
 sg13g2_nand2_1 _8402_ (.Y(_3386_),
    .A(_3372_),
    .B(_3376_));
 sg13g2_inv_1 _8403_ (.Y(_3387_),
    .A(_3274_));
 sg13g2_o21ai_1 _8404_ (.B1(_2875_),
    .Y(_3388_),
    .A1(net156),
    .A2(_3387_));
 sg13g2_a21oi_1 _8405_ (.A1(net156),
    .A2(_3387_),
    .Y(_3389_),
    .B1(_3388_));
 sg13g2_nand2_1 _8406_ (.Y(_3390_),
    .A(_3347_),
    .B(_3346_));
 sg13g2_o21ai_1 _8407_ (.B1(_3390_),
    .Y(_3391_),
    .A1(_4463_),
    .A2(_3280_));
 sg13g2_xnor2_1 _8408_ (.Y(_3392_),
    .A(_4350_),
    .B(_3274_));
 sg13g2_nor2_1 _8409_ (.A(_3391_),
    .B(_3392_),
    .Y(_3393_));
 sg13g2_nand2_1 _8410_ (.Y(_3394_),
    .A(_3392_),
    .B(_3391_));
 sg13g2_inv_1 _8411_ (.Y(_3395_),
    .A(_3394_));
 sg13g2_nor3_1 _8412_ (.A(_2875_),
    .B(_3393_),
    .C(_3395_),
    .Y(_3396_));
 sg13g2_o21ai_1 _8413_ (.B1(_3176_),
    .Y(_3397_),
    .A1(_3389_),
    .A2(_3396_));
 sg13g2_nand3_1 _8414_ (.B(_3386_),
    .C(_3397_),
    .A(_3385_),
    .Y(_3398_));
 sg13g2_o21ai_1 _8415_ (.B1(_2690_),
    .Y(_3399_),
    .A1(_1634_),
    .A2(_3398_));
 sg13g2_a21oi_1 _8416_ (.A1(_3380_),
    .A2(_3383_),
    .Y(_0109_),
    .B1(_3399_));
 sg13g2_nand2_1 _8417_ (.Y(_3400_),
    .A(_3092_),
    .B(_3088_));
 sg13g2_nand3_1 _8418_ (.B(_3400_),
    .C(_3086_),
    .A(_3083_),
    .Y(_3401_));
 sg13g2_a21oi_1 _8419_ (.A1(_3118_),
    .A2(_3401_),
    .Y(_3402_),
    .B1(_3177_));
 sg13g2_nand2_1 _8420_ (.Y(_3403_),
    .A(_3087_),
    .B(_3093_));
 sg13g2_nand3_1 _8421_ (.B(_3362_),
    .C(_3086_),
    .A(_3083_),
    .Y(_3404_));
 sg13g2_nand2_1 _8422_ (.Y(_3405_),
    .A(_3403_),
    .B(_3404_));
 sg13g2_nand2_1 _8423_ (.Y(_3406_),
    .A(_3405_),
    .B(_3115_));
 sg13g2_nand2_1 _8424_ (.Y(_3407_),
    .A(_3402_),
    .B(_3406_));
 sg13g2_nor2b_1 _8425_ (.A(_3387_),
    .B_N(_3381_),
    .Y(_3408_));
 sg13g2_nor2_1 _8426_ (.A(_3408_),
    .B(net66),
    .Y(_3409_));
 sg13g2_nor2_1 _8427_ (.A(_3357_),
    .B(_3409_),
    .Y(_3410_));
 sg13g2_nand2_1 _8428_ (.Y(_3411_),
    .A(net66),
    .B(_3408_));
 sg13g2_a21oi_1 _8429_ (.A1(_3410_),
    .A2(_3411_),
    .Y(_3412_),
    .B1(_3169_));
 sg13g2_nand2_1 _8430_ (.Y(_3413_),
    .A(_3407_),
    .B(_3412_));
 sg13g2_nand2_1 _8431_ (.Y(_3414_),
    .A(_3115_),
    .B(_3354_));
 sg13g2_nand2_1 _8432_ (.Y(_3415_),
    .A(_3118_),
    .B(_3404_));
 sg13g2_nand3_1 _8433_ (.B(_3415_),
    .C(_3129_),
    .A(_3414_),
    .Y(_3416_));
 sg13g2_nor2b_1 _8434_ (.A(_3413_),
    .B_N(_3416_),
    .Y(_3417_));
 sg13g2_mux2_1 _8435_ (.A0(_3337_),
    .A1(_3348_),
    .S(_0067_),
    .X(_3418_));
 sg13g2_nand2_1 _8436_ (.Y(_3419_),
    .A(_3199_),
    .B(net156));
 sg13g2_o21ai_1 _8437_ (.B1(_3369_),
    .Y(_3420_),
    .A1(_3322_),
    .A2(_3419_));
 sg13g2_nor2_1 _8438_ (.A(_0067_),
    .B(_3387_),
    .Y(_3421_));
 sg13g2_nand2_1 _8439_ (.Y(_3422_),
    .A(net66),
    .B(_3421_));
 sg13g2_nor2_1 _8440_ (.A(_3421_),
    .B(_3269_),
    .Y(_3423_));
 sg13g2_nor2_1 _8441_ (.A(_1627_),
    .B(_3423_),
    .Y(_3424_));
 sg13g2_xnor2_1 _8442_ (.Y(_3425_),
    .A(net161),
    .B(net66));
 sg13g2_o21ai_1 _8443_ (.B1(_3394_),
    .Y(_3426_),
    .A1(net142),
    .A2(_3274_));
 sg13g2_xnor2_1 _8444_ (.Y(_3427_),
    .A(_3425_),
    .B(_3426_));
 sg13g2_inv_1 _8445_ (.Y(_3428_),
    .A(_3176_));
 sg13g2_a221oi_1 _8446_ (.B2(net144),
    .C1(_3428_),
    .B1(_3427_),
    .A1(_3422_),
    .Y(_3429_),
    .A2(_3424_));
 sg13g2_a221oi_1 _8447_ (.B2(_3329_),
    .C1(_3429_),
    .B1(_3420_),
    .A1(_3372_),
    .Y(_3430_),
    .A2(_3418_));
 sg13g2_a21oi_1 _8448_ (.A1(_3430_),
    .A2(_3169_),
    .Y(_3431_),
    .B1(_2634_));
 sg13g2_nor2b_1 _8449_ (.A(_3417_),
    .B_N(_3431_),
    .Y(_0110_));
 sg13g2_nand3_1 _8450_ (.B(_3415_),
    .C(_3128_),
    .A(_3414_),
    .Y(_3432_));
 sg13g2_xor2_1 _8451_ (.B(_3247_),
    .A(_3409_),
    .X(_3433_));
 sg13g2_a21oi_1 _8452_ (.A1(_3433_),
    .A2(_3125_),
    .Y(_3434_),
    .B1(_3169_));
 sg13g2_inv_1 _8453_ (.Y(_3435_),
    .A(net156));
 sg13g2_o21ai_1 _8454_ (.B1(_3369_),
    .Y(_3436_),
    .A1(_3435_),
    .A2(_3350_));
 sg13g2_xnor2_1 _8455_ (.Y(_3437_),
    .A(_1629_),
    .B(_3422_));
 sg13g2_o21ai_1 _8456_ (.B1(_2875_),
    .Y(_3438_),
    .A1(_3247_),
    .A2(_3437_));
 sg13g2_a21oi_1 _8457_ (.A1(_3247_),
    .A2(_3437_),
    .Y(_3439_),
    .B1(_3438_));
 sg13g2_nand2_1 _8458_ (.Y(_3440_),
    .A(_3426_),
    .B(_3425_));
 sg13g2_o21ai_1 _8459_ (.B1(_3440_),
    .Y(_3441_),
    .A1(net158),
    .A2(net66));
 sg13g2_xnor2_1 _8460_ (.Y(_3442_),
    .A(net159),
    .B(_3247_));
 sg13g2_o21ai_1 _8461_ (.B1(_1627_),
    .Y(_3443_),
    .A1(_3442_),
    .A2(_3441_));
 sg13g2_a21oi_1 _8462_ (.A1(_3441_),
    .A2(_3442_),
    .Y(_3444_),
    .B1(_3443_));
 sg13g2_nor3_1 _8463_ (.A(_3428_),
    .B(_3439_),
    .C(_3444_),
    .Y(_3445_));
 sg13g2_a21oi_1 _8464_ (.A1(_3436_),
    .A2(_2826_),
    .Y(_3446_),
    .B1(_3445_));
 sg13g2_nand4_1 _8465_ (.B(net156),
    .C(_2827_),
    .A(_3328_),
    .Y(_3447_),
    .D(_3348_));
 sg13g2_nand3_1 _8466_ (.B(_3169_),
    .C(_3447_),
    .A(_3446_),
    .Y(_3448_));
 sg13g2_buf_1 _8467_ (.A(_1637_),
    .X(_3449_));
 sg13g2_nand2_1 _8468_ (.Y(_3450_),
    .A(_3448_),
    .B(_3449_));
 sg13g2_a21oi_1 _8469_ (.A1(_3432_),
    .A2(_3434_),
    .Y(_0111_),
    .B1(_3450_));
 sg13g2_nor2_1 _8470_ (.A(net135),
    .B(_1258_),
    .Y(_3451_));
 sg13g2_buf_2 _8471_ (.A(_3451_),
    .X(_3452_));
 sg13g2_inv_1 _8472_ (.Y(_3453_),
    .A(_3452_));
 sg13g2_xor2_1 _8473_ (.B(\i_display.frame_crotchet[0] ),
    .A(_1185_),
    .X(_3454_));
 sg13g2_nor2b_1 _8474_ (.A(_1187_),
    .B_N(_0065_),
    .Y(_3455_));
 sg13g2_nor2_1 _8475_ (.A(_0065_),
    .B(_1188_),
    .Y(_3456_));
 sg13g2_xnor2_1 _8476_ (.Y(_3457_),
    .A(_0067_),
    .B(_1193_));
 sg13g2_nand2_1 _8477_ (.Y(_3458_),
    .A(_1198_),
    .B(_0066_));
 sg13g2_nand2b_1 _8478_ (.Y(_3459_),
    .B(_1197_),
    .A_N(_0066_));
 sg13g2_nand3_1 _8479_ (.B(_3458_),
    .C(_3459_),
    .A(_3457_),
    .Y(_3460_));
 sg13g2_nor4_1 _8480_ (.A(_3454_),
    .B(_3455_),
    .C(_3456_),
    .D(_3460_),
    .Y(_3461_));
 sg13g2_xnor2_1 _8481_ (.Y(_3462_),
    .A(_0054_),
    .B(_1178_));
 sg13g2_xnor2_1 _8482_ (.Y(_3463_),
    .A(_0069_),
    .B(_1176_));
 sg13g2_xnor2_1 _8483_ (.Y(_3464_),
    .A(_0068_),
    .B(_1180_));
 sg13g2_nand4_1 _8484_ (.B(_3462_),
    .C(_3463_),
    .A(_3461_),
    .Y(_3465_),
    .D(_3464_));
 sg13g2_nand2_1 _8485_ (.Y(_3466_),
    .A(_3465_),
    .B(_4414_));
 sg13g2_o21ai_1 _8486_ (.B1(_3466_),
    .Y(_3467_),
    .A1(_4383_),
    .A2(_3465_));
 sg13g2_a21oi_1 _8487_ (.A1(_1208_),
    .A2(_1181_),
    .Y(_3468_),
    .B1(_1263_));
 sg13g2_a22oi_1 _8488_ (.Y(_3469_),
    .B1(_1202_),
    .B2(_3468_),
    .A2(_1276_),
    .A1(_1182_));
 sg13g2_nand3_1 _8489_ (.B(_1202_),
    .C(_1279_),
    .A(_1201_),
    .Y(_3470_));
 sg13g2_o21ai_1 _8490_ (.B1(_3470_),
    .Y(_3471_),
    .A1(_1190_),
    .A2(_3469_));
 sg13g2_o21ai_1 _8491_ (.B1(_1198_),
    .Y(_3472_),
    .A1(_1194_),
    .A2(_1184_));
 sg13g2_a21oi_1 _8492_ (.A1(_1203_),
    .A2(_1194_),
    .Y(_3473_),
    .B1(_1185_));
 sg13g2_a22oi_1 _8493_ (.Y(_3474_),
    .B1(_3472_),
    .B2(_3473_),
    .A2(_1247_),
    .A1(net148));
 sg13g2_nor3_1 _8494_ (.A(_1202_),
    .B(_1188_),
    .C(_3474_),
    .Y(_3475_));
 sg13g2_o21ai_1 _8495_ (.B1(_3465_),
    .Y(_3476_),
    .A1(_3471_),
    .A2(_3475_));
 sg13g2_buf_1 _8496_ (.A(_3476_),
    .X(_3477_));
 sg13g2_nand4_1 _8497_ (.B(net143),
    .C(_1239_),
    .A(_3467_),
    .Y(_3478_),
    .D(_3477_));
 sg13g2_o21ai_1 _8498_ (.B1(_3478_),
    .Y(_0112_),
    .A1(_4414_),
    .A2(_3453_));
 sg13g2_buf_1 _8499_ (.A(net127),
    .X(_3479_));
 sg13g2_a21oi_1 _8500_ (.A1(_1172_),
    .A2(_4413_),
    .Y(_3480_),
    .B1(net160));
 sg13g2_nand2_1 _8501_ (.Y(_3481_),
    .A(_4413_),
    .B(net160));
 sg13g2_a21oi_1 _8502_ (.A1(_3477_),
    .A2(_3481_),
    .Y(_3482_),
    .B1(_1240_));
 sg13g2_nor3_1 _8503_ (.A(_3479_),
    .B(_3480_),
    .C(_3482_),
    .Y(_0113_));
 sg13g2_xnor2_1 _8504_ (.Y(_3483_),
    .A(_4265_),
    .B(_3481_));
 sg13g2_nand3_1 _8505_ (.B(net157),
    .C(_1239_),
    .A(_3477_),
    .Y(_3484_));
 sg13g2_buf_2 _8506_ (.A(_3484_),
    .X(_3485_));
 sg13g2_nand2_1 _8507_ (.Y(_3486_),
    .A(_3452_),
    .B(_4431_));
 sg13g2_o21ai_1 _8508_ (.B1(_3486_),
    .Y(_0114_),
    .A1(_3483_),
    .A2(_3485_));
 sg13g2_nor2_1 _8509_ (.A(_4432_),
    .B(_3481_),
    .Y(_3487_));
 sg13g2_xnor2_1 _8510_ (.Y(_3488_),
    .A(_4393_),
    .B(_3487_));
 sg13g2_nand2_1 _8511_ (.Y(_3489_),
    .A(_3452_),
    .B(net152));
 sg13g2_o21ai_1 _8512_ (.B1(_3489_),
    .Y(_0115_),
    .A1(_3488_),
    .A2(_3485_));
 sg13g2_nor3_1 _8513_ (.A(_4432_),
    .B(_0280_),
    .C(_3481_),
    .Y(_3490_));
 sg13g2_xnor2_1 _8514_ (.Y(_3491_),
    .A(_4351_),
    .B(_3490_));
 sg13g2_nand2_1 _8515_ (.Y(_3492_),
    .A(_3452_),
    .B(net142));
 sg13g2_o21ai_1 _8516_ (.B1(_3492_),
    .Y(_0116_),
    .A1(_3491_),
    .A2(_3485_));
 sg13g2_nand2_1 _8517_ (.Y(_3493_),
    .A(_3490_),
    .B(net142));
 sg13g2_xnor2_1 _8518_ (.Y(_3494_),
    .A(net161),
    .B(_3493_));
 sg13g2_nand2_1 _8519_ (.Y(_3495_),
    .A(_3452_),
    .B(net158));
 sg13g2_o21ai_1 _8520_ (.B1(_3495_),
    .Y(_0117_),
    .A1(_3494_),
    .A2(_3485_));
 sg13g2_nor2_1 _8521_ (.A(_0414_),
    .B(_3493_),
    .Y(_3496_));
 sg13g2_xnor2_1 _8522_ (.Y(_3497_),
    .A(_4343_),
    .B(_3496_));
 sg13g2_nand2_1 _8523_ (.Y(_3498_),
    .A(_3452_),
    .B(net159));
 sg13g2_o21ai_1 _8524_ (.B1(_3498_),
    .Y(_0118_),
    .A1(_3497_),
    .A2(_3485_));
 sg13g2_nand2_1 _8525_ (.Y(_3499_),
    .A(_3496_),
    .B(net159));
 sg13g2_xnor2_1 _8526_ (.Y(_3500_),
    .A(_4575_),
    .B(_3499_));
 sg13g2_nand2_1 _8527_ (.Y(_3501_),
    .A(_3452_),
    .B(_0464_));
 sg13g2_o21ai_1 _8528_ (.B1(_3501_),
    .Y(_0119_),
    .A1(_3500_),
    .A2(_3485_));
 sg13g2_nand3_1 _8529_ (.B(_0464_),
    .C(net159),
    .A(_3496_),
    .Y(_3502_));
 sg13g2_xnor2_1 _8530_ (.Y(_3503_),
    .A(_0306_),
    .B(_3502_));
 sg13g2_nand2_1 _8531_ (.Y(_3504_),
    .A(_3452_),
    .B(_0440_));
 sg13g2_o21ai_1 _8532_ (.B1(_3504_),
    .Y(_0120_),
    .A1(_3503_),
    .A2(_3485_));
 sg13g2_nor2_1 _8533_ (.A(_0441_),
    .B(_3502_),
    .Y(_3505_));
 sg13g2_xnor2_1 _8534_ (.Y(_3506_),
    .A(_0040_),
    .B(_3505_));
 sg13g2_nand3_1 _8535_ (.B(_1477_),
    .C(_3506_),
    .A(_3477_),
    .Y(_3507_));
 sg13g2_o21ai_1 _8536_ (.B1(_3507_),
    .Y(_0121_),
    .A1(_0436_),
    .A2(_3453_));
 sg13g2_nor4_1 _8537_ (.A(_1003_),
    .B(\i_display.i_vga.timing_ver.counter[8] ),
    .C(_0712_),
    .D(\i_display.i_vga.timing_ver.counter[10] ),
    .Y(_3508_));
 sg13g2_nor4_1 _8538_ (.A(_1083_),
    .B(_1023_),
    .C(_1014_),
    .D(_1098_),
    .Y(_3509_));
 sg13g2_nand2_1 _8539_ (.Y(_3510_),
    .A(_1053_),
    .B(_1067_));
 sg13g2_nor2_1 _8540_ (.A(_1042_),
    .B(_3510_),
    .Y(_3511_));
 sg13g2_nand3_1 _8541_ (.B(_3509_),
    .C(_3511_),
    .A(_3508_),
    .Y(_3512_));
 sg13g2_o21ai_1 _8542_ (.B1(_1380_),
    .Y(_3513_),
    .A1(_3512_),
    .A2(_1238_));
 sg13g2_inv_2 _8543_ (.Y(_3514_),
    .A(_3513_));
 sg13g2_nor2_1 _8544_ (.A(_1054_),
    .B(_4243_),
    .Y(_3515_));
 sg13g2_a21oi_1 _8545_ (.A1(_0051_),
    .A2(_4243_),
    .Y(_3516_),
    .B1(_3515_));
 sg13g2_nand2_1 _8546_ (.Y(_0129_),
    .A(_3514_),
    .B(_3516_));
 sg13g2_nor2_1 _8547_ (.A(_3510_),
    .B(_1238_),
    .Y(_3517_));
 sg13g2_inv_1 _8548_ (.Y(_3518_),
    .A(_3517_));
 sg13g2_nor3_1 _8549_ (.A(_1014_),
    .B(_3134_),
    .C(_3518_),
    .Y(_3519_));
 sg13g2_inv_1 _8550_ (.Y(_3520_),
    .A(_3519_));
 sg13g2_nor2_1 _8551_ (.A(_1148_),
    .B(_3520_),
    .Y(_3521_));
 sg13g2_nand2_1 _8552_ (.Y(_3522_),
    .A(_3521_),
    .B(_1003_));
 sg13g2_nor2b_1 _8553_ (.A(_3522_),
    .B_N(_1151_),
    .Y(_3523_));
 sg13g2_nor2_1 _8554_ (.A(_0981_),
    .B(_3522_),
    .Y(_3524_));
 sg13g2_a21oi_1 _8555_ (.A1(_3524_),
    .A2(\i_display.i_vga.timing_ver.counter[9] ),
    .Y(_3525_),
    .B1(\i_display.i_vga.timing_ver.counter[10] ));
 sg13g2_o21ai_1 _8556_ (.B1(_3514_),
    .Y(_0130_),
    .A1(_3523_),
    .A2(_3525_));
 sg13g2_nor2_1 _8557_ (.A(_3148_),
    .B(_1171_),
    .Y(_3526_));
 sg13g2_a21oi_1 _8558_ (.A1(_1067_),
    .A2(_1163_),
    .Y(_3527_),
    .B1(_3526_));
 sg13g2_nand2_1 _8559_ (.Y(_0131_),
    .A(_3514_),
    .B(_3527_));
 sg13g2_xnor2_1 _8560_ (.Y(_3528_),
    .A(_1041_),
    .B(_3517_));
 sg13g2_nand2_1 _8561_ (.Y(_0132_),
    .A(_3528_),
    .B(_3514_));
 sg13g2_nor2_1 _8562_ (.A(_1083_),
    .B(_1237_),
    .Y(_3529_));
 sg13g2_xnor2_1 _8563_ (.Y(_3530_),
    .A(_0052_),
    .B(_3511_));
 sg13g2_a21oi_1 _8564_ (.A1(_3512_),
    .A2(_3530_),
    .Y(_3531_),
    .B1(_1238_));
 sg13g2_nor3_1 _8565_ (.A(_3479_),
    .B(_3529_),
    .C(_3531_),
    .Y(_0133_));
 sg13g2_o21ai_1 _8566_ (.B1(_3520_),
    .Y(_3532_),
    .A1(_1013_),
    .A2(_3517_));
 sg13g2_nor3_1 _8567_ (.A(_3136_),
    .B(_3513_),
    .C(_3532_),
    .Y(_0134_));
 sg13g2_nor2_1 _8568_ (.A(_1023_),
    .B(_3519_),
    .Y(_3533_));
 sg13g2_nor2_1 _8569_ (.A(_1024_),
    .B(_3520_),
    .Y(_3534_));
 sg13g2_o21ai_1 _8570_ (.B1(_3514_),
    .Y(_0135_),
    .A1(_3533_),
    .A2(_3534_));
 sg13g2_nor2_1 _8571_ (.A(\i_display.i_vga.timing_ver.counter[6] ),
    .B(_3534_),
    .Y(_3535_));
 sg13g2_o21ai_1 _8572_ (.B1(_3514_),
    .Y(_0136_),
    .A1(_3521_),
    .A2(_3535_));
 sg13g2_nor2_1 _8573_ (.A(_1003_),
    .B(_3521_),
    .Y(_3536_));
 sg13g2_inv_1 _8574_ (.Y(_3537_),
    .A(_3522_));
 sg13g2_o21ai_1 _8575_ (.B1(_3514_),
    .Y(_0137_),
    .A1(_3536_),
    .A2(_3537_));
 sg13g2_nor2_1 _8576_ (.A(\i_display.i_vga.timing_ver.counter[8] ),
    .B(_3537_),
    .Y(_3538_));
 sg13g2_o21ai_1 _8577_ (.B1(_3514_),
    .Y(_0138_),
    .A1(_3524_),
    .A2(_3538_));
 sg13g2_xnor2_1 _8578_ (.Y(_3539_),
    .A(\i_display.i_vga.timing_ver.counter[9] ),
    .B(_3524_));
 sg13g2_nand2_1 _8579_ (.Y(_0139_),
    .A(_3539_),
    .B(_3449_));
 sg13g2_nand2_1 _8580_ (.Y(_3540_),
    .A(net27),
    .B(_4146_));
 sg13g2_a21oi_1 _8581_ (.A1(_3540_),
    .A2(_1319_),
    .Y(_0143_),
    .B1(net119));
 sg13g2_nand2_1 _8582_ (.Y(_3541_),
    .A(net27),
    .B(_4144_));
 sg13g2_a21oi_1 _8583_ (.A1(_3541_),
    .A2(_1252_),
    .Y(_0144_),
    .B1(net119));
 sg13g2_nand2_1 _8584_ (.Y(_3542_),
    .A(_1167_),
    .B(_0663_));
 sg13g2_nand2b_1 _8585_ (.Y(_3543_),
    .B(net28),
    .A_N(_1220_));
 sg13g2_a21oi_1 _8586_ (.A1(_3542_),
    .A2(_3543_),
    .Y(_0145_),
    .B1(net119));
 sg13g2_nand2_1 _8587_ (.Y(_3544_),
    .A(net27),
    .B(_0667_));
 sg13g2_a21oi_1 _8588_ (.A1(_3544_),
    .A2(_1284_),
    .Y(_0146_),
    .B1(net119));
 sg13g2_nand2_1 _8589_ (.Y(_3545_),
    .A(net27),
    .B(_4158_));
 sg13g2_a21oi_1 _8590_ (.A1(_3545_),
    .A2(_1298_),
    .Y(_0147_),
    .B1(net119));
 sg13g2_nand2_1 _8591_ (.Y(_3546_),
    .A(net27),
    .B(_4157_));
 sg13g2_a21oi_1 _8592_ (.A1(_3546_),
    .A2(_1267_),
    .Y(_0148_),
    .B1(net119));
 sg13g2_nand3_1 _8593_ (.B(_4253_),
    .C(_4178_),
    .A(net28),
    .Y(_3547_));
 sg13g2_xor2_1 _8594_ (.B(_3547_),
    .A(\i_display.x_idx[8] ),
    .X(_3548_));
 sg13g2_nor2_1 _8595_ (.A(_3453_),
    .B(_3548_),
    .Y(_0149_));
 sg13g2_nand2_1 _8596_ (.Y(_0155_),
    .A(_0175_),
    .B(_1618_));
 sg13g2_nand2b_1 _8597_ (.Y(_0156_),
    .B(net133),
    .A_N(_0102_));
 sg13g2_buf_1 _8598_ (.A(net127),
    .X(_3549_));
 sg13g2_nor2_1 _8599_ (.A(_1587_),
    .B(_1586_),
    .Y(_3550_));
 sg13g2_inv_1 _8600_ (.Y(_3551_),
    .A(_1588_));
 sg13g2_nor3_1 _8601_ (.A(_3549_),
    .B(_3550_),
    .C(_3551_),
    .Y(_0157_));
 sg13g2_nor2_1 _8602_ (.A(\i_music.count[11] ),
    .B(_3551_),
    .Y(_3552_));
 sg13g2_nor3_1 _8603_ (.A(net118),
    .B(_1589_),
    .C(_3552_),
    .Y(_0158_));
 sg13g2_nor2_1 _8604_ (.A(\i_music.count[12] ),
    .B(_1589_),
    .Y(_3553_));
 sg13g2_inv_1 _8605_ (.Y(_3554_),
    .A(_1590_));
 sg13g2_nor3_1 _8606_ (.A(_3549_),
    .B(_3553_),
    .C(_3554_),
    .Y(_0159_));
 sg13g2_nor2_1 _8607_ (.A(\i_music.count[13] ),
    .B(_3554_),
    .Y(_3555_));
 sg13g2_nor3_1 _8608_ (.A(net118),
    .B(_1591_),
    .C(_3555_),
    .Y(_0160_));
 sg13g2_nor2_1 _8609_ (.A(\i_music.count[14] ),
    .B(_1591_),
    .Y(_3556_));
 sg13g2_inv_1 _8610_ (.Y(_3557_),
    .A(_1592_));
 sg13g2_nor3_1 _8611_ (.A(net118),
    .B(_3556_),
    .C(_3557_),
    .Y(_0161_));
 sg13g2_nor2_1 _8612_ (.A(\i_music.count[15] ),
    .B(_3557_),
    .Y(_3558_));
 sg13g2_nor3_1 _8613_ (.A(net118),
    .B(_1593_),
    .C(_3558_),
    .Y(_0162_));
 sg13g2_nor2_1 _8614_ (.A(\i_music.count[16] ),
    .B(_1593_),
    .Y(_3559_));
 sg13g2_inv_1 _8615_ (.Y(_3560_),
    .A(_1594_));
 sg13g2_nor3_1 _8616_ (.A(net118),
    .B(_3559_),
    .C(_3560_),
    .Y(_0163_));
 sg13g2_nor2_1 _8617_ (.A(\i_music.count[17] ),
    .B(_3560_),
    .Y(_3561_));
 sg13g2_nor3_1 _8618_ (.A(net118),
    .B(_1595_),
    .C(_3561_),
    .Y(_0164_));
 sg13g2_nor2_1 _8619_ (.A(\i_music.count[18] ),
    .B(_1595_),
    .Y(_3562_));
 sg13g2_inv_1 _8620_ (.Y(_3563_),
    .A(_1596_));
 sg13g2_nor3_1 _8621_ (.A(net118),
    .B(_3562_),
    .C(_3563_),
    .Y(_0165_));
 sg13g2_nor2_1 _8622_ (.A(\i_music.count[19] ),
    .B(_3563_),
    .Y(_3564_));
 sg13g2_nor3_1 _8623_ (.A(net118),
    .B(_1597_),
    .C(_3564_),
    .Y(_0166_));
 sg13g2_nor2_1 _8624_ (.A(net135),
    .B(_3159_),
    .Y(_0167_));
 sg13g2_buf_1 _8625_ (.A(net127),
    .X(_3565_));
 sg13g2_nor2_1 _8626_ (.A(\i_music.count[20] ),
    .B(_1597_),
    .Y(_3566_));
 sg13g2_nor2b_1 _8627_ (.A(_1598_),
    .B_N(\i_music.count[20] ),
    .Y(_3567_));
 sg13g2_nor3_1 _8628_ (.A(net117),
    .B(_3566_),
    .C(_3567_),
    .Y(_0168_));
 sg13g2_nor2_1 _8629_ (.A(_1576_),
    .B(_3567_),
    .Y(_3568_));
 sg13g2_nor3_1 _8630_ (.A(net117),
    .B(_1599_),
    .C(_3568_),
    .Y(_0169_));
 sg13g2_nor2_1 _8631_ (.A(_1600_),
    .B(_1599_),
    .Y(_3569_));
 sg13g2_inv_1 _8632_ (.Y(_3570_),
    .A(_1601_));
 sg13g2_nor3_1 _8633_ (.A(net117),
    .B(_3569_),
    .C(_3570_),
    .Y(_0170_));
 sg13g2_nor2_1 _8634_ (.A(\i_music.count[23] ),
    .B(_3570_),
    .Y(_3571_));
 sg13g2_nor3_1 _8635_ (.A(net117),
    .B(_1602_),
    .C(_3571_),
    .Y(_0171_));
 sg13g2_nor2_1 _8636_ (.A(\i_music.count[24] ),
    .B(_1602_),
    .Y(_3572_));
 sg13g2_nor3_1 _8637_ (.A(net117),
    .B(_3572_),
    .C(_1615_),
    .Y(_0172_));
 sg13g2_inv_1 _8638_ (.Y(_3573_),
    .A(_1191_));
 sg13g2_nand4_1 _8639_ (.B(_1186_),
    .C(_1195_),
    .A(_1611_),
    .Y(_3574_),
    .D(_2031_));
 sg13g2_nor3_1 _8640_ (.A(_3573_),
    .B(_3574_),
    .C(_1598_),
    .Y(_3575_));
 sg13g2_nor2_1 _8641_ (.A(_3574_),
    .B(_1598_),
    .Y(_3576_));
 sg13g2_nor2_1 _8642_ (.A(_1191_),
    .B(_3576_),
    .Y(_3577_));
 sg13g2_nor3_1 _8643_ (.A(net117),
    .B(_3575_),
    .C(_3577_),
    .Y(_0176_));
 sg13g2_a21oi_1 _8644_ (.A1(_1607_),
    .A2(_1191_),
    .Y(_3578_),
    .B1(\crotchet[4] ));
 sg13g2_nand3_1 _8645_ (.B(\crotchet[4] ),
    .C(_1191_),
    .A(_1607_),
    .Y(_3579_));
 sg13g2_inv_1 _8646_ (.Y(_3580_),
    .A(_3579_));
 sg13g2_nor3_1 _8647_ (.A(_3565_),
    .B(_3578_),
    .C(_3580_),
    .Y(_0177_));
 sg13g2_o21ai_1 _8648_ (.B1(net134),
    .Y(_3581_),
    .A1(_0074_),
    .A2(_1530_));
 sg13g2_a21oi_1 _8649_ (.A1(_0074_),
    .A2(_1530_),
    .Y(_0178_),
    .B1(_3581_));
 sg13g2_nor2_1 _8650_ (.A(\crotchet[5] ),
    .B(_3580_),
    .Y(_3582_));
 sg13g2_nand2_1 _8651_ (.Y(_3583_),
    .A(_3580_),
    .B(\crotchet[5] ));
 sg13g2_inv_1 _8652_ (.Y(_3584_),
    .A(_3583_));
 sg13g2_nor3_1 _8653_ (.A(_3565_),
    .B(_3582_),
    .C(_3584_),
    .Y(_0179_));
 sg13g2_inv_1 _8654_ (.Y(_3585_),
    .A(\crotchet[6] ));
 sg13g2_o21ai_1 _8655_ (.B1(_2690_),
    .Y(_3586_),
    .A1(_3585_),
    .A2(_3583_));
 sg13g2_a21oi_1 _8656_ (.A1(_3585_),
    .A2(_3583_),
    .Y(_0180_),
    .B1(_3586_));
 sg13g2_nor2_1 _8657_ (.A(_4239_),
    .B(_4235_),
    .Y(_3587_));
 sg13g2_inv_1 _8658_ (.Y(_3588_),
    .A(_1234_));
 sg13g2_nor3_1 _8659_ (.A(net117),
    .B(_3587_),
    .C(_3588_),
    .Y(_0181_));
 sg13g2_nor2_1 _8660_ (.A(_4238_),
    .B(_3588_),
    .Y(_3589_));
 sg13g2_nor3_1 _8661_ (.A(net117),
    .B(_1235_),
    .C(_3589_),
    .Y(_0182_));
 sg13g2_buf_1 _8662_ (.A(net135),
    .X(_3590_));
 sg13g2_nor2_1 _8663_ (.A(\i_display.i_vga.low_count[5] ),
    .B(_1235_),
    .Y(_3591_));
 sg13g2_nor3_1 _8664_ (.A(net125),
    .B(_3591_),
    .C(_1582_),
    .Y(_0183_));
 sg13g2_nor2_1 _8665_ (.A(_4225_),
    .B(_1582_),
    .Y(_3592_));
 sg13g2_inv_1 _8666_ (.Y(_3593_),
    .A(_1583_));
 sg13g2_nor3_1 _8667_ (.A(net125),
    .B(_3592_),
    .C(_3593_),
    .Y(_0184_));
 sg13g2_nor2_1 _8668_ (.A(\i_display.i_vga.low_count[7] ),
    .B(_3593_),
    .Y(_3594_));
 sg13g2_nor3_1 _8669_ (.A(net125),
    .B(_1584_),
    .C(_3594_),
    .Y(_0185_));
 sg13g2_nor2_1 _8670_ (.A(_4236_),
    .B(_1584_),
    .Y(_3595_));
 sg13g2_inv_1 _8671_ (.Y(_3596_),
    .A(_1585_));
 sg13g2_nor3_1 _8672_ (.A(_3590_),
    .B(_3595_),
    .C(_3596_),
    .Y(_0186_));
 sg13g2_nor2_1 _8673_ (.A(_4237_),
    .B(_3596_),
    .Y(_3597_));
 sg13g2_nor3_1 _8674_ (.A(net125),
    .B(_1586_),
    .C(_3597_),
    .Y(_0187_));
 sg13g2_nand2_1 _8675_ (.Y(_3598_),
    .A(_2332_),
    .B(_1668_));
 sg13g2_nand3_1 _8676_ (.B(_3160_),
    .C(_3598_),
    .A(_2334_),
    .Y(_3599_));
 sg13g2_nand2_1 _8677_ (.Y(_3600_),
    .A(net75),
    .B(_1557_));
 sg13g2_nand2_1 _8678_ (.Y(_3601_),
    .A(net80),
    .B(_1540_));
 sg13g2_buf_2 _8679_ (.A(_3601_),
    .X(_3602_));
 sg13g2_nand2_1 _8680_ (.Y(_3603_),
    .A(net79),
    .B(net78));
 sg13g2_inv_1 _8681_ (.Y(_3604_),
    .A(_3603_));
 sg13g2_buf_1 _8682_ (.A(net78),
    .X(_3605_));
 sg13g2_nor2_1 _8683_ (.A(net79),
    .B(net60),
    .Y(_3606_));
 sg13g2_nor2_1 _8684_ (.A(net73),
    .B(_3606_),
    .Y(_3607_));
 sg13g2_nor2_1 _8685_ (.A(net80),
    .B(net79),
    .Y(_3608_));
 sg13g2_buf_1 _8686_ (.A(_3608_),
    .X(_3609_));
 sg13g2_nand2_1 _8687_ (.Y(_3610_),
    .A(_1531_),
    .B(\i_music.i_sample.t1.genblk1[1].state.Q ));
 sg13g2_inv_1 _8688_ (.Y(_3611_),
    .A(_3610_));
 sg13g2_nor2_1 _8689_ (.A(net65),
    .B(_3611_),
    .Y(_3612_));
 sg13g2_buf_2 _8690_ (.A(_3612_),
    .X(_3613_));
 sg13g2_inv_1 _8691_ (.Y(_3614_),
    .A(_3613_));
 sg13g2_a22oi_1 _8692_ (.Y(_3615_),
    .B1(_3607_),
    .B2(_3614_),
    .A2(_3604_),
    .A1(_3602_));
 sg13g2_o21ai_1 _8693_ (.B1(net67),
    .Y(_3616_),
    .A1(_3600_),
    .A2(_3615_));
 sg13g2_nor2_1 _8694_ (.A(net76),
    .B(_1547_),
    .Y(_3617_));
 sg13g2_nor2_1 _8695_ (.A(_3617_),
    .B(_3604_),
    .Y(_3618_));
 sg13g2_inv_1 _8696_ (.Y(_3619_),
    .A(_3618_));
 sg13g2_nor2_1 _8697_ (.A(net80),
    .B(_1537_),
    .Y(_3620_));
 sg13g2_inv_1 _8698_ (.Y(_3621_),
    .A(_3620_));
 sg13g2_nand2_2 _8699_ (.Y(_3622_),
    .A(net79),
    .B(_1540_));
 sg13g2_nand2_1 _8700_ (.Y(_3623_),
    .A(_3622_),
    .B(net70));
 sg13g2_nor2_1 _8701_ (.A(_1532_),
    .B(_3623_),
    .Y(_3624_));
 sg13g2_a21oi_1 _8702_ (.A1(_3619_),
    .A2(_3621_),
    .Y(_3625_),
    .B1(_3624_));
 sg13g2_buf_1 _8703_ (.A(_1552_),
    .X(_3626_));
 sg13g2_buf_1 _8704_ (.A(net72),
    .X(_3627_));
 sg13g2_buf_1 _8705_ (.A(net74),
    .X(_3628_));
 sg13g2_nand3b_1 _8706_ (.B(net64),
    .C(net63),
    .Y(_3629_),
    .A_N(_3625_));
 sg13g2_nor2_1 _8707_ (.A(_1536_),
    .B(_1540_),
    .Y(_3630_));
 sg13g2_inv_2 _8708_ (.Y(_3631_),
    .A(_3630_));
 sg13g2_nand2_2 _8709_ (.Y(_3632_),
    .A(_3631_),
    .B(net78));
 sg13g2_inv_1 _8710_ (.Y(_3633_),
    .A(_3632_));
 sg13g2_nand2_1 _8711_ (.Y(_3634_),
    .A(net65),
    .B(net76));
 sg13g2_nand2_1 _8712_ (.Y(_3635_),
    .A(_3633_),
    .B(_3634_));
 sg13g2_o21ai_1 _8713_ (.B1(_1548_),
    .Y(_3636_),
    .A1(_1541_),
    .A2(net65));
 sg13g2_nor2_1 _8714_ (.A(_1557_),
    .B(_1553_),
    .Y(_3637_));
 sg13g2_buf_1 _8715_ (.A(_3637_),
    .X(_3638_));
 sg13g2_nand3_1 _8716_ (.B(_3636_),
    .C(net52),
    .A(_3635_),
    .Y(_3639_));
 sg13g2_nand2_1 _8717_ (.Y(_3640_),
    .A(_3619_),
    .B(_3613_));
 sg13g2_inv_1 _8718_ (.Y(_3641_),
    .A(_3623_));
 sg13g2_nand2_1 _8719_ (.Y(_3642_),
    .A(_3641_),
    .B(_1532_));
 sg13g2_nor2_1 _8720_ (.A(_1552_),
    .B(_1557_),
    .Y(_3643_));
 sg13g2_buf_1 _8721_ (.A(_3643_),
    .X(_3644_));
 sg13g2_buf_1 _8722_ (.A(_3644_),
    .X(_3645_));
 sg13g2_nand3_1 _8723_ (.B(_3642_),
    .C(_3645_),
    .A(_3640_),
    .Y(_3646_));
 sg13g2_nand3_1 _8724_ (.B(_3639_),
    .C(_3646_),
    .A(_3629_),
    .Y(_3647_));
 sg13g2_nand2_1 _8725_ (.Y(_3648_),
    .A(_1547_),
    .B(net76));
 sg13g2_nor2_1 _8726_ (.A(net70),
    .B(_3622_),
    .Y(_3649_));
 sg13g2_inv_1 _8727_ (.Y(_3650_),
    .A(_3617_));
 sg13g2_nor2_1 _8728_ (.A(_3650_),
    .B(_3613_),
    .Y(_3651_));
 sg13g2_o21ai_1 _8729_ (.B1(net72),
    .Y(_3652_),
    .A1(_3649_),
    .A2(_3651_));
 sg13g2_o21ai_1 _8730_ (.B1(_3652_),
    .Y(_3653_),
    .A1(_3620_),
    .A2(_3648_));
 sg13g2_inv_2 _8731_ (.Y(_3654_),
    .A(_3602_));
 sg13g2_nor2_1 _8732_ (.A(_1531_),
    .B(_1540_),
    .Y(_3655_));
 sg13g2_buf_1 _8733_ (.A(_3655_),
    .X(_3656_));
 sg13g2_inv_1 _8734_ (.Y(_3657_),
    .A(_3656_));
 sg13g2_nor2_1 _8735_ (.A(_1536_),
    .B(_1546_),
    .Y(_3658_));
 sg13g2_a21oi_1 _8736_ (.A1(net50),
    .A2(_3658_),
    .Y(_3659_),
    .B1(net72));
 sg13g2_o21ai_1 _8737_ (.B1(_3659_),
    .Y(_3660_),
    .A1(_3654_),
    .A2(_3618_));
 sg13g2_nor2_1 _8738_ (.A(net78),
    .B(net50),
    .Y(_3661_));
 sg13g2_inv_1 _8739_ (.Y(_3662_),
    .A(_3661_));
 sg13g2_nand2_2 _8740_ (.Y(_3663_),
    .A(net80),
    .B(net78));
 sg13g2_nand3_1 _8741_ (.B(net72),
    .C(_3663_),
    .A(_3662_),
    .Y(_3664_));
 sg13g2_a21oi_1 _8742_ (.A1(_3660_),
    .A2(_3664_),
    .Y(_3665_),
    .B1(net68));
 sg13g2_a21oi_1 _8743_ (.A1(_3653_),
    .A2(net58),
    .Y(_3666_),
    .B1(_3665_));
 sg13g2_nand2_1 _8744_ (.Y(_3667_),
    .A(_3622_),
    .B(_1546_));
 sg13g2_nor2_1 _8745_ (.A(_3620_),
    .B(_3667_),
    .Y(_3668_));
 sg13g2_a21oi_1 _8746_ (.A1(_3668_),
    .A2(net51),
    .Y(_3669_),
    .B1(_1565_));
 sg13g2_a21oi_1 _8747_ (.A1(_3666_),
    .A2(_3669_),
    .Y(_3670_),
    .B1(net77));
 sg13g2_o21ai_1 _8748_ (.B1(_3670_),
    .Y(_3671_),
    .A1(_3616_),
    .A2(_3647_));
 sg13g2_nor2_1 _8749_ (.A(net60),
    .B(_3621_),
    .Y(_3672_));
 sg13g2_nand2b_1 _8750_ (.Y(_3673_),
    .B(_3633_),
    .A_N(_3672_));
 sg13g2_nand2_2 _8751_ (.Y(_3674_),
    .A(_1542_),
    .B(net80));
 sg13g2_inv_1 _8752_ (.Y(_3675_),
    .A(_3644_));
 sg13g2_a21oi_1 _8753_ (.A1(_3641_),
    .A2(_3674_),
    .Y(_3676_),
    .B1(_3675_));
 sg13g2_a21oi_1 _8754_ (.A1(_3673_),
    .A2(_3676_),
    .Y(_3677_),
    .B1(_1563_));
 sg13g2_nand2_1 _8755_ (.Y(_3678_),
    .A(_1537_),
    .B(net80));
 sg13g2_o21ai_1 _8756_ (.B1(_3642_),
    .Y(_3679_),
    .A1(net59),
    .A2(_3678_));
 sg13g2_nand2_1 _8757_ (.Y(_3680_),
    .A(_3679_),
    .B(_3638_));
 sg13g2_nand2_1 _8758_ (.Y(_3681_),
    .A(_3677_),
    .B(_3680_));
 sg13g2_inv_1 _8759_ (.Y(_3682_),
    .A(_3624_));
 sg13g2_nor2_1 _8760_ (.A(_1537_),
    .B(_3602_),
    .Y(_3683_));
 sg13g2_nor2_1 _8761_ (.A(_1547_),
    .B(_3683_),
    .Y(_3684_));
 sg13g2_nor2_1 _8762_ (.A(_1552_),
    .B(_3684_),
    .Y(_3685_));
 sg13g2_inv_1 _8763_ (.Y(_3686_),
    .A(_3658_));
 sg13g2_nor2_1 _8764_ (.A(net50),
    .B(_3686_),
    .Y(_3687_));
 sg13g2_nor2_1 _8765_ (.A(_3602_),
    .B(_3686_),
    .Y(_3688_));
 sg13g2_a221oi_1 _8766_ (.B2(_3654_),
    .C1(net59),
    .B1(_1537_),
    .A1(_3620_),
    .Y(_3689_),
    .A2(_1543_));
 sg13g2_nor3_1 _8767_ (.A(_3687_),
    .B(_3688_),
    .C(_3689_),
    .Y(_3690_));
 sg13g2_a221oi_1 _8768_ (.B2(net64),
    .C1(net58),
    .B1(_3690_),
    .A1(_3682_),
    .Y(_3691_),
    .A2(_3685_));
 sg13g2_nand2_1 _8769_ (.Y(_3692_),
    .A(_3621_),
    .B(net60));
 sg13g2_nand2_1 _8770_ (.Y(_3693_),
    .A(_3602_),
    .B(_3622_));
 sg13g2_inv_1 _8771_ (.Y(_3694_),
    .A(_3693_));
 sg13g2_nand2_1 _8772_ (.Y(_3695_),
    .A(_3692_),
    .B(_3694_));
 sg13g2_nor2_1 _8773_ (.A(_3600_),
    .B(_3604_),
    .Y(_3696_));
 sg13g2_nor2_2 _8774_ (.A(net60),
    .B(_3611_),
    .Y(_3697_));
 sg13g2_nand2_1 _8775_ (.Y(_3698_),
    .A(_3611_),
    .B(net60));
 sg13g2_nand2_1 _8776_ (.Y(_3699_),
    .A(_3698_),
    .B(net73));
 sg13g2_o21ai_1 _8777_ (.B1(net70),
    .Y(_3700_),
    .A1(_3656_),
    .A2(_3611_));
 sg13g2_o21ai_1 _8778_ (.B1(_3700_),
    .Y(_3701_),
    .A1(_3697_),
    .A2(_3699_));
 sg13g2_a221oi_1 _8779_ (.B2(net52),
    .C1(_1564_),
    .B1(_3701_),
    .A1(_3695_),
    .Y(_3702_),
    .A2(_3696_));
 sg13g2_nor3_1 _8780_ (.A(_3605_),
    .B(_3609_),
    .C(_3654_),
    .Y(_3703_));
 sg13g2_nand2b_1 _8781_ (.Y(_3704_),
    .B(_3699_),
    .A_N(_3703_));
 sg13g2_nor2_1 _8782_ (.A(_1537_),
    .B(net50),
    .Y(_3705_));
 sg13g2_inv_1 _8783_ (.Y(_3706_),
    .A(_3705_));
 sg13g2_nor2_1 _8784_ (.A(_3654_),
    .B(_3667_),
    .Y(_3707_));
 sg13g2_a21oi_1 _8785_ (.A1(_3706_),
    .A2(_3607_),
    .Y(_3708_),
    .B1(_3707_));
 sg13g2_nor3_1 _8786_ (.A(net69),
    .B(net68),
    .C(_3708_),
    .Y(_3709_));
 sg13g2_a21oi_1 _8787_ (.A1(net51),
    .A2(_3704_),
    .Y(_3710_),
    .B1(_3709_));
 sg13g2_a21oi_1 _8788_ (.A1(_3702_),
    .A2(_3710_),
    .Y(_3711_),
    .B1(_1569_));
 sg13g2_o21ai_1 _8789_ (.B1(_3711_),
    .Y(_3712_),
    .A1(_3681_),
    .A2(_3691_));
 sg13g2_nand4_1 _8790_ (.B(net100),
    .C(_3671_),
    .A(net29),
    .Y(_3713_),
    .D(_3712_));
 sg13g2_a21oi_1 _8791_ (.A1(_3599_),
    .A2(_3713_),
    .Y(_0205_),
    .B1(net119));
 sg13g2_inv_2 _8792_ (.Y(_3714_),
    .A(_0167_));
 sg13g2_buf_1 _8793_ (.A(_1563_),
    .X(_3715_));
 sg13g2_nor2_1 _8794_ (.A(_1541_),
    .B(_1537_),
    .Y(_3716_));
 sg13g2_a21oi_1 _8795_ (.A1(net70),
    .A2(_3716_),
    .Y(_3717_),
    .B1(_3688_));
 sg13g2_nor2_1 _8796_ (.A(net79),
    .B(_3674_),
    .Y(_3718_));
 sg13g2_inv_2 _8797_ (.Y(_3719_),
    .A(_3667_));
 sg13g2_nand2b_1 _8798_ (.Y(_3720_),
    .B(_3719_),
    .A_N(_3718_));
 sg13g2_a21oi_1 _8799_ (.A1(_3717_),
    .A2(_3720_),
    .Y(_3721_),
    .B1(_3675_));
 sg13g2_nor2_1 _8800_ (.A(net76),
    .B(_3613_),
    .Y(_3722_));
 sg13g2_buf_1 _8801_ (.A(net73),
    .X(_3723_));
 sg13g2_o21ai_1 _8802_ (.B1(net62),
    .Y(_3724_),
    .A1(_3697_),
    .A2(_3722_));
 sg13g2_inv_1 _8803_ (.Y(_3725_),
    .A(net52));
 sg13g2_a21oi_1 _8804_ (.A1(_3724_),
    .A2(_3682_),
    .Y(_3726_),
    .B1(_3725_));
 sg13g2_nor2_1 _8805_ (.A(_1552_),
    .B(_3633_),
    .Y(_3727_));
 sg13g2_nor2_1 _8806_ (.A(net73),
    .B(_3656_),
    .Y(_3728_));
 sg13g2_a22oi_1 _8807_ (.Y(_3729_),
    .B1(_3614_),
    .B2(_3728_),
    .A2(_3719_),
    .A1(_3692_));
 sg13g2_a221oi_1 _8808_ (.B2(net64),
    .C1(net58),
    .B1(_3729_),
    .A1(net50),
    .Y(_3730_),
    .A2(_3727_));
 sg13g2_nor4_1 _8809_ (.A(net71),
    .B(_3721_),
    .C(_3726_),
    .D(_3730_),
    .Y(_3731_));
 sg13g2_inv_1 _8810_ (.Y(_3732_),
    .A(_3683_));
 sg13g2_nand2_1 _8811_ (.Y(_3733_),
    .A(_3732_),
    .B(_3728_));
 sg13g2_a221oi_1 _8812_ (.B2(net64),
    .C1(net63),
    .B1(_3640_),
    .A1(_3733_),
    .Y(_3734_),
    .A2(_3618_));
 sg13g2_o21ai_1 _8813_ (.B1(net75),
    .Y(_3735_),
    .A1(_3617_),
    .A2(_3613_));
 sg13g2_nor2_2 _8814_ (.A(net76),
    .B(net78),
    .Y(_3736_));
 sg13g2_nor2_1 _8815_ (.A(_3656_),
    .B(_3632_),
    .Y(_3737_));
 sg13g2_inv_1 _8816_ (.Y(_3738_),
    .A(_3737_));
 sg13g2_nand2b_1 _8817_ (.Y(_3739_),
    .B(_3738_),
    .A_N(_3736_));
 sg13g2_inv_1 _8818_ (.Y(_3740_),
    .A(_3739_));
 sg13g2_nor2_1 _8819_ (.A(_3605_),
    .B(_1537_),
    .Y(_3741_));
 sg13g2_buf_1 _8820_ (.A(net72),
    .X(_3742_));
 sg13g2_o21ai_1 _8821_ (.B1(_3742_),
    .Y(_3743_),
    .A1(_3741_),
    .A2(_3668_));
 sg13g2_o21ai_1 _8822_ (.B1(_3743_),
    .Y(_3744_),
    .A1(_3735_),
    .A2(_3740_));
 sg13g2_nor2_1 _8823_ (.A(net58),
    .B(_3744_),
    .Y(_3745_));
 sg13g2_o21ai_1 _8824_ (.B1(net71),
    .Y(_3746_),
    .A1(_3734_),
    .A2(_3745_));
 sg13g2_nand3b_1 _8825_ (.B(net77),
    .C(_3746_),
    .Y(_3747_),
    .A_N(_3731_));
 sg13g2_nand2_1 _8826_ (.Y(_3748_),
    .A(_3619_),
    .B(net50));
 sg13g2_nor2_1 _8827_ (.A(net60),
    .B(_3613_),
    .Y(_3749_));
 sg13g2_inv_1 _8828_ (.Y(_3750_),
    .A(_3749_));
 sg13g2_nand3_1 _8829_ (.B(net59),
    .C(_3674_),
    .A(_3750_),
    .Y(_3751_));
 sg13g2_o21ai_1 _8830_ (.B1(_3751_),
    .Y(_3752_),
    .A1(_3654_),
    .A2(_3748_));
 sg13g2_inv_1 _8831_ (.Y(_3753_),
    .A(_3716_));
 sg13g2_inv_1 _8832_ (.Y(_3754_),
    .A(_3663_));
 sg13g2_a21oi_1 _8833_ (.A1(_3753_),
    .A2(_3754_),
    .Y(_3755_),
    .B1(_3703_));
 sg13g2_a21oi_1 _8834_ (.A1(_3755_),
    .A2(net69),
    .Y(_3756_),
    .B1(net68));
 sg13g2_o21ai_1 _8835_ (.B1(_3756_),
    .Y(_3757_),
    .A1(net69),
    .A2(_3752_));
 sg13g2_o21ai_1 _8836_ (.B1(_3748_),
    .Y(_3758_),
    .A1(_3654_),
    .A2(_3686_));
 sg13g2_nor2_1 _8837_ (.A(net79),
    .B(net50),
    .Y(_3759_));
 sg13g2_inv_1 _8838_ (.Y(_3760_),
    .A(_3759_));
 sg13g2_nand2_1 _8839_ (.Y(_3761_),
    .A(_3684_),
    .B(_3760_));
 sg13g2_o21ai_1 _8840_ (.B1(_3761_),
    .Y(_3762_),
    .A1(_3656_),
    .A2(_3717_));
 sg13g2_a22oi_1 _8841_ (.Y(_3763_),
    .B1(_3638_),
    .B2(_3762_),
    .A2(_3758_),
    .A1(net51));
 sg13g2_nand3_1 _8842_ (.B(net67),
    .C(_3763_),
    .A(_3757_),
    .Y(_3764_));
 sg13g2_nand2_1 _8843_ (.Y(_3765_),
    .A(_3630_),
    .B(net70));
 sg13g2_nand2_1 _8844_ (.Y(_3766_),
    .A(_3765_),
    .B(net72));
 sg13g2_nor3_1 _8845_ (.A(_3654_),
    .B(_3766_),
    .C(_3651_),
    .Y(_3767_));
 sg13g2_a221oi_1 _8846_ (.B2(net62),
    .C1(_3742_),
    .B1(net65),
    .A1(net80),
    .Y(_3768_),
    .A2(net60));
 sg13g2_o21ai_1 _8847_ (.B1(_3628_),
    .Y(_3769_),
    .A1(_3767_),
    .A2(_3768_));
 sg13g2_inv_1 _8848_ (.Y(_3770_),
    .A(_3649_));
 sg13g2_a21oi_1 _8849_ (.A1(_3770_),
    .A2(_3663_),
    .Y(_3771_),
    .B1(_3611_));
 sg13g2_nand2_1 _8850_ (.Y(_3772_),
    .A(_3631_),
    .B(_1548_));
 sg13g2_nor2_1 _8851_ (.A(_3772_),
    .B(_3749_),
    .Y(_3773_));
 sg13g2_o21ai_1 _8852_ (.B1(net52),
    .Y(_3774_),
    .A1(_3771_),
    .A2(_3773_));
 sg13g2_nor2_1 _8853_ (.A(_1549_),
    .B(net50),
    .Y(_3775_));
 sg13g2_o21ai_1 _8854_ (.B1(net51),
    .Y(_3776_),
    .A1(_3688_),
    .A2(_3775_));
 sg13g2_nand4_1 _8855_ (.B(net71),
    .C(_3774_),
    .A(_3769_),
    .Y(_3777_),
    .D(_3776_));
 sg13g2_nand3_1 _8856_ (.B(_1569_),
    .C(_3777_),
    .A(_3764_),
    .Y(_3778_));
 sg13g2_nor2_2 _8857_ (.A(net135),
    .B(_2025_),
    .Y(_3779_));
 sg13g2_nand4_1 _8858_ (.B(_3747_),
    .C(_3778_),
    .A(net29),
    .Y(_3780_),
    .D(_3779_));
 sg13g2_o21ai_1 _8859_ (.B1(_3780_),
    .Y(_0206_),
    .A1(_3714_),
    .A2(_2393_));
 sg13g2_nor2_1 _8860_ (.A(net61),
    .B(net59),
    .Y(_3781_));
 sg13g2_nand2_1 _8861_ (.Y(_3782_),
    .A(_3706_),
    .B(_3732_));
 sg13g2_nor2_1 _8862_ (.A(net60),
    .B(_3614_),
    .Y(_3783_));
 sg13g2_inv_1 _8863_ (.Y(_3784_),
    .A(_3783_));
 sg13g2_a21o_1 _8864_ (.A2(net59),
    .A1(_3784_),
    .B1(_3651_),
    .X(_3785_));
 sg13g2_a22oi_1 _8865_ (.Y(_3786_),
    .B1(net64),
    .B2(_3785_),
    .A2(_3782_),
    .A1(_3781_));
 sg13g2_nand4_1 _8866_ (.B(net61),
    .C(net68),
    .A(_3761_),
    .Y(_3787_),
    .D(_3765_));
 sg13g2_nand2_1 _8867_ (.Y(_3788_),
    .A(_3750_),
    .B(net73));
 sg13g2_nand3_1 _8868_ (.B(_3644_),
    .C(_3662_),
    .A(_3788_),
    .Y(_3789_));
 sg13g2_nand3_1 _8869_ (.B(_3789_),
    .C(_1563_),
    .A(_3787_),
    .Y(_3790_));
 sg13g2_a21oi_1 _8870_ (.A1(_3786_),
    .A2(net63),
    .Y(_3791_),
    .B1(_3790_));
 sg13g2_nand2_1 _8871_ (.Y(_3792_),
    .A(_3631_),
    .B(_3602_));
 sg13g2_a21oi_1 _8872_ (.A1(_3792_),
    .A2(_3663_),
    .Y(_3793_),
    .B1(net61));
 sg13g2_nand2_1 _8873_ (.Y(_3794_),
    .A(_3698_),
    .B(_3634_));
 sg13g2_a221oi_1 _8874_ (.B2(net62),
    .C1(net69),
    .B1(_3794_),
    .A1(_3656_),
    .Y(_3795_),
    .A2(_3658_));
 sg13g2_o21ai_1 _8875_ (.B1(net63),
    .Y(_3796_),
    .A1(_3793_),
    .A2(_3795_));
 sg13g2_nand2_1 _8876_ (.Y(_3797_),
    .A(_3619_),
    .B(_3621_));
 sg13g2_o21ai_1 _8877_ (.B1(_3797_),
    .Y(_3798_),
    .A1(net62),
    .A2(_3722_));
 sg13g2_a221oi_1 _8878_ (.B2(_3741_),
    .C1(_3725_),
    .B1(_3674_),
    .A1(_3754_),
    .Y(_3799_),
    .A2(_3630_));
 sg13g2_a21oi_1 _8879_ (.A1(_3798_),
    .A2(net51),
    .Y(_3800_),
    .B1(_3799_));
 sg13g2_a21oi_1 _8880_ (.A1(_3796_),
    .A2(_3800_),
    .Y(_3801_),
    .B1(net71));
 sg13g2_o21ai_1 _8881_ (.B1(net77),
    .Y(_3802_),
    .A1(_3791_),
    .A2(_3801_));
 sg13g2_nand2_1 _8882_ (.Y(_3803_),
    .A(_3634_),
    .B(_3610_));
 sg13g2_nor2_1 _8883_ (.A(net75),
    .B(_3736_),
    .Y(_3804_));
 sg13g2_inv_1 _8884_ (.Y(_3805_),
    .A(net65));
 sg13g2_nand2_1 _8885_ (.Y(_3806_),
    .A(_3805_),
    .B(_3674_));
 sg13g2_nor2_1 _8886_ (.A(net73),
    .B(_3806_),
    .Y(_3807_));
 sg13g2_nor2_1 _8887_ (.A(net61),
    .B(_3807_),
    .Y(_3808_));
 sg13g2_nand2_1 _8888_ (.Y(_3809_),
    .A(_3668_),
    .B(_3631_));
 sg13g2_a221oi_1 _8889_ (.B2(_3809_),
    .C1(net58),
    .B1(_3808_),
    .A1(_3803_),
    .Y(_3810_),
    .A2(_3804_));
 sg13g2_nor2_1 _8890_ (.A(net62),
    .B(_3631_),
    .Y(_3811_));
 sg13g2_nand2_1 _8891_ (.Y(_3812_),
    .A(_3697_),
    .B(net70));
 sg13g2_a21oi_1 _8892_ (.A1(_3812_),
    .A2(_3699_),
    .Y(_3813_),
    .B1(net65));
 sg13g2_o21ai_1 _8893_ (.B1(net52),
    .Y(_3814_),
    .A1(_3811_),
    .A2(_3813_));
 sg13g2_o21ai_1 _8894_ (.B1(_3733_),
    .Y(_3815_),
    .A1(net59),
    .A2(_3672_));
 sg13g2_a21oi_1 _8895_ (.A1(_3815_),
    .A2(net51),
    .Y(_3816_),
    .B1(net67));
 sg13g2_nand3b_1 _8896_ (.B(_3814_),
    .C(_3816_),
    .Y(_3817_),
    .A_N(_3810_));
 sg13g2_inv_1 _8897_ (.Y(_3818_),
    .A(_3807_));
 sg13g2_a21oi_1 _8898_ (.A1(_3788_),
    .A2(_3818_),
    .Y(_3819_),
    .B1(_3675_));
 sg13g2_nand2_1 _8899_ (.Y(_3820_),
    .A(_3641_),
    .B(_3678_));
 sg13g2_nand3_1 _8900_ (.B(_3770_),
    .C(_3663_),
    .A(_3820_),
    .Y(_3821_));
 sg13g2_inv_1 _8901_ (.Y(_3822_),
    .A(_3727_));
 sg13g2_nand2_1 _8902_ (.Y(_3823_),
    .A(_3822_),
    .B(_1558_));
 sg13g2_nand3_1 _8903_ (.B(_3641_),
    .C(net74),
    .A(_3613_),
    .Y(_3824_));
 sg13g2_a22oi_1 _8904_ (.Y(_3825_),
    .B1(_3823_),
    .B2(_3824_),
    .A2(_3627_),
    .A1(_3821_));
 sg13g2_nand2_1 _8905_ (.Y(_3826_),
    .A(_3784_),
    .B(net73));
 sg13g2_nor2b_1 _8906_ (.A(_3826_),
    .B_N(_3674_),
    .Y(_3827_));
 sg13g2_nor3_1 _8907_ (.A(_3725_),
    .B(_3741_),
    .C(_3827_),
    .Y(_3828_));
 sg13g2_nor3_1 _8908_ (.A(_3819_),
    .B(_3825_),
    .C(_3828_),
    .Y(_3829_));
 sg13g2_nand2_1 _8909_ (.Y(_3830_),
    .A(_3829_),
    .B(net67));
 sg13g2_nand3_1 _8910_ (.B(_3830_),
    .C(_1569_),
    .A(_3817_),
    .Y(_3831_));
 sg13g2_nand4_1 _8911_ (.B(_3779_),
    .C(_3802_),
    .A(net29),
    .Y(_3832_),
    .D(_3831_));
 sg13g2_o21ai_1 _8912_ (.B1(_3832_),
    .Y(_0207_),
    .A1(_3714_),
    .A2(_2462_));
 sg13g2_nand2_1 _8913_ (.Y(_3833_),
    .A(_3736_),
    .B(_3610_));
 sg13g2_o21ai_1 _8914_ (.B1(_3833_),
    .Y(_3834_),
    .A1(_3697_),
    .A2(_3632_));
 sg13g2_a21oi_1 _8915_ (.A1(_3673_),
    .A2(_3686_),
    .Y(_3835_),
    .B1(net75));
 sg13g2_a21oi_1 _8916_ (.A1(_1554_),
    .A2(_3834_),
    .Y(_3836_),
    .B1(_3835_));
 sg13g2_nand3_1 _8917_ (.B(net75),
    .C(_3636_),
    .A(_3826_),
    .Y(_3837_));
 sg13g2_nand2_1 _8918_ (.Y(_3838_),
    .A(_3760_),
    .B(_3719_));
 sg13g2_nand3_1 _8919_ (.B(net72),
    .C(_3820_),
    .A(_3838_),
    .Y(_3839_));
 sg13g2_nand3_1 _8920_ (.B(net74),
    .C(_3839_),
    .A(_3837_),
    .Y(_3840_));
 sg13g2_o21ai_1 _8921_ (.B1(_3840_),
    .Y(_3841_),
    .A1(net63),
    .A2(_3836_));
 sg13g2_nor2b_1 _8922_ (.A(_3715_),
    .B_N(_3841_),
    .Y(_3842_));
 sg13g2_nand3_1 _8923_ (.B(net64),
    .C(_3648_),
    .A(_3724_),
    .Y(_3843_));
 sg13g2_a21oi_1 _8924_ (.A1(_3602_),
    .A2(_3723_),
    .Y(_3844_),
    .B1(net61));
 sg13g2_a21oi_1 _8925_ (.A1(_3844_),
    .A2(_3706_),
    .Y(_3845_),
    .B1(net68));
 sg13g2_a221oi_1 _8926_ (.B2(_3650_),
    .C1(net61),
    .B1(_3806_),
    .A1(net79),
    .Y(_3846_),
    .A2(_3723_));
 sg13g2_nor2_1 _8927_ (.A(net63),
    .B(_3846_),
    .Y(_3847_));
 sg13g2_nor2_1 _8928_ (.A(net65),
    .B(_3648_),
    .Y(_3848_));
 sg13g2_a21oi_1 _8929_ (.A1(_3805_),
    .A2(_3622_),
    .Y(_3849_),
    .B1(net59));
 sg13g2_o21ai_1 _8930_ (.B1(net64),
    .Y(_3850_),
    .A1(_3848_),
    .A2(_3849_));
 sg13g2_a221oi_1 _8931_ (.B2(_3850_),
    .C1(net67),
    .B1(_3847_),
    .A1(_3843_),
    .Y(_3851_),
    .A2(_3845_));
 sg13g2_o21ai_1 _8932_ (.B1(_1569_),
    .Y(_3852_),
    .A1(_3842_),
    .A2(_3851_));
 sg13g2_nand2_1 _8933_ (.Y(_3853_),
    .A(_3794_),
    .B(net70));
 sg13g2_o21ai_1 _8934_ (.B1(net62),
    .Y(_3854_),
    .A1(net76),
    .A2(net65));
 sg13g2_a21oi_1 _8935_ (.A1(_3853_),
    .A2(_3854_),
    .Y(_3855_),
    .B1(_3725_));
 sg13g2_nand2_1 _8936_ (.Y(_3856_),
    .A(_3806_),
    .B(net62));
 sg13g2_a21oi_1 _8937_ (.A1(_3856_),
    .A2(_3833_),
    .Y(_3857_),
    .B1(_3675_));
 sg13g2_nor3_1 _8938_ (.A(net78),
    .B(_3716_),
    .C(_3697_),
    .Y(_3858_));
 sg13g2_a21oi_1 _8939_ (.A1(_3698_),
    .A2(_3719_),
    .Y(_3859_),
    .B1(_3858_));
 sg13g2_a221oi_1 _8940_ (.B2(net64),
    .C1(net68),
    .B1(_3859_),
    .A1(_3751_),
    .Y(_3860_),
    .A2(_3685_));
 sg13g2_nor4_1 _8941_ (.A(net71),
    .B(_3855_),
    .C(_3857_),
    .D(_3860_),
    .Y(_3861_));
 sg13g2_nand2_1 _8942_ (.Y(_3862_),
    .A(_3772_),
    .B(net51));
 sg13g2_nor2_1 _8943_ (.A(_3693_),
    .B(_3632_),
    .Y(_3863_));
 sg13g2_o21ai_1 _8944_ (.B1(net75),
    .Y(_3864_),
    .A1(_3687_),
    .A2(_3863_));
 sg13g2_nand2_1 _8945_ (.Y(_3865_),
    .A(_3737_),
    .B(_3626_));
 sg13g2_a21oi_1 _8946_ (.A1(_3672_),
    .A2(net61),
    .Y(_3866_),
    .B1(_1559_));
 sg13g2_nand3_1 _8947_ (.B(_3865_),
    .C(_3866_),
    .A(_3864_),
    .Y(_3867_));
 sg13g2_o21ai_1 _8948_ (.B1(_3867_),
    .Y(_3868_),
    .A1(_3707_),
    .A2(_3862_));
 sg13g2_nand2_1 _8949_ (.Y(_3869_),
    .A(_3868_),
    .B(net71));
 sg13g2_nand3b_1 _8950_ (.B(net77),
    .C(_3869_),
    .Y(_3870_),
    .A_N(_3861_));
 sg13g2_nand4_1 _8951_ (.B(_3779_),
    .C(_3852_),
    .A(_2546_),
    .Y(_3871_),
    .D(_3870_));
 sg13g2_o21ai_1 _8952_ (.B1(_3871_),
    .Y(_0208_),
    .A1(_3714_),
    .A2(_2507_));
 sg13g2_inv_1 _8953_ (.Y(_3872_),
    .A(_3685_));
 sg13g2_nand2b_1 _8954_ (.Y(_3873_),
    .B(_3732_),
    .A_N(_3772_));
 sg13g2_nand3_1 _8955_ (.B(_3809_),
    .C(net72),
    .A(_3873_),
    .Y(_3874_));
 sg13g2_o21ai_1 _8956_ (.B1(_3874_),
    .Y(_3875_),
    .A1(_3872_),
    .A2(_3858_));
 sg13g2_nand2_1 _8957_ (.Y(_3876_),
    .A(_3875_),
    .B(net74));
 sg13g2_nand4_1 _8958_ (.B(_3610_),
    .C(net52),
    .A(_3632_),
    .Y(_3877_),
    .D(_3663_));
 sg13g2_nand3_1 _8959_ (.B(_3631_),
    .C(_3644_),
    .A(_3657_),
    .Y(_3878_));
 sg13g2_nand3_1 _8960_ (.B(_3877_),
    .C(_3878_),
    .A(_3876_),
    .Y(_3879_));
 sg13g2_nand2_1 _8961_ (.Y(_3880_),
    .A(_3879_),
    .B(net67));
 sg13g2_nor3_1 _8962_ (.A(net69),
    .B(_3641_),
    .C(_3737_),
    .Y(_3881_));
 sg13g2_a21oi_1 _8963_ (.A1(_3765_),
    .A2(net51),
    .Y(_3882_),
    .B1(_1564_));
 sg13g2_o21ai_1 _8964_ (.B1(_3882_),
    .Y(_3883_),
    .A1(_3823_),
    .A2(_3881_));
 sg13g2_nand3_1 _8965_ (.B(net77),
    .C(_3883_),
    .A(_3880_),
    .Y(_3884_));
 sg13g2_nor2_1 _8966_ (.A(_3626_),
    .B(_3719_),
    .Y(_3885_));
 sg13g2_nor3_1 _8967_ (.A(net75),
    .B(_3848_),
    .C(_3619_),
    .Y(_3886_));
 sg13g2_a21oi_1 _8968_ (.A1(_3853_),
    .A2(_3885_),
    .Y(_3887_),
    .B1(_3886_));
 sg13g2_nand2b_1 _8969_ (.Y(_3888_),
    .B(net58),
    .A_N(_3887_));
 sg13g2_nand3_1 _8970_ (.B(net61),
    .C(_3812_),
    .A(_3738_),
    .Y(_3889_));
 sg13g2_nand3b_1 _8971_ (.B(_3889_),
    .C(net74),
    .Y(_3890_),
    .A_N(_3885_));
 sg13g2_nand3_1 _8972_ (.B(net71),
    .C(_3890_),
    .A(_3888_),
    .Y(_3891_));
 sg13g2_a22oi_1 _8973_ (.Y(_3892_),
    .B1(net69),
    .B2(_3661_),
    .A2(net62),
    .A1(_3683_));
 sg13g2_o21ai_1 _8974_ (.B1(net68),
    .Y(_3893_),
    .A1(_3736_),
    .A2(_3606_));
 sg13g2_nand2_1 _8975_ (.Y(_3894_),
    .A(net76),
    .B(net73));
 sg13g2_a21oi_1 _8976_ (.A1(_3894_),
    .A2(net74),
    .Y(_3895_),
    .B1(net69));
 sg13g2_nand2_1 _8977_ (.Y(_3896_),
    .A(_3893_),
    .B(_3895_));
 sg13g2_nand2b_1 _8978_ (.Y(_3897_),
    .B(_3644_),
    .A_N(_3894_));
 sg13g2_nor2_1 _8979_ (.A(_1563_),
    .B(_3811_),
    .Y(_3898_));
 sg13g2_nand4_1 _8980_ (.B(_3896_),
    .C(_3897_),
    .A(_3892_),
    .Y(_3899_),
    .D(_3898_));
 sg13g2_nand3_1 _8981_ (.B(_1569_),
    .C(_3899_),
    .A(_3891_),
    .Y(_3900_));
 sg13g2_nand2_1 _8982_ (.Y(_3901_),
    .A(_3884_),
    .B(_3900_));
 sg13g2_nand3_1 _8983_ (.B(_3779_),
    .C(_3901_),
    .A(net29),
    .Y(_3902_));
 sg13g2_o21ai_1 _8984_ (.B1(_3902_),
    .Y(_0209_),
    .A1(_3714_),
    .A2(_2544_));
 sg13g2_nor2_1 _8985_ (.A(_1564_),
    .B(_3644_),
    .Y(_3903_));
 sg13g2_inv_1 _8986_ (.Y(_3904_),
    .A(_3903_));
 sg13g2_nand2_1 _8987_ (.Y(_3905_),
    .A(_3623_),
    .B(_3627_));
 sg13g2_nor2_1 _8988_ (.A(net58),
    .B(_3905_),
    .Y(_3906_));
 sg13g2_nor2_1 _8989_ (.A(_3904_),
    .B(_3906_),
    .Y(_3907_));
 sg13g2_nor2_1 _8990_ (.A(_3736_),
    .B(_3725_),
    .Y(_3908_));
 sg13g2_a22oi_1 _8991_ (.Y(_3909_),
    .B1(_3645_),
    .B2(_3738_),
    .A2(_3760_),
    .A1(_3908_));
 sg13g2_nand3_1 _8992_ (.B(_1558_),
    .C(_3873_),
    .A(_3865_),
    .Y(_3910_));
 sg13g2_a21oi_1 _8993_ (.A1(_3909_),
    .A2(_3910_),
    .Y(_3911_),
    .B1(_3715_));
 sg13g2_o21ai_1 _8994_ (.B1(net77),
    .Y(_3912_),
    .A1(_3907_),
    .A2(_3911_));
 sg13g2_nor2_1 _8995_ (.A(net69),
    .B(_3740_),
    .Y(_3913_));
 sg13g2_o21ai_1 _8996_ (.B1(net63),
    .Y(_3914_),
    .A1(_3781_),
    .A2(_3913_));
 sg13g2_a22oi_1 _8997_ (.Y(_3915_),
    .B1(net58),
    .B2(_3719_),
    .A2(net52),
    .A1(_3848_));
 sg13g2_nand3_1 _8998_ (.B(net71),
    .C(_3915_),
    .A(_3914_),
    .Y(_3916_));
 sg13g2_o21ai_1 _8999_ (.B1(net52),
    .Y(_3917_),
    .A1(_3649_),
    .A2(_3641_));
 sg13g2_nand2_1 _9000_ (.Y(_3918_),
    .A(_3766_),
    .B(_3628_));
 sg13g2_nand4_1 _9001_ (.B(net67),
    .C(_3897_),
    .A(_3917_),
    .Y(_3919_),
    .D(_3918_));
 sg13g2_nand3_1 _9002_ (.B(_1569_),
    .C(_3919_),
    .A(_3916_),
    .Y(_3920_));
 sg13g2_nand4_1 _9003_ (.B(_3779_),
    .C(_3912_),
    .A(net29),
    .Y(_3921_),
    .D(_3920_));
 sg13g2_o21ai_1 _9004_ (.B1(_3921_),
    .Y(_0210_),
    .A1(_3714_),
    .A2(_2564_));
 sg13g2_a21oi_1 _9005_ (.A1(_1549_),
    .A2(_3694_),
    .Y(_3922_),
    .B1(_3885_));
 sg13g2_a21oi_1 _9006_ (.A1(_3804_),
    .A2(net74),
    .Y(_3923_),
    .B1(_1564_));
 sg13g2_o21ai_1 _9007_ (.B1(_3923_),
    .Y(_3924_),
    .A1(net63),
    .A2(_3922_));
 sg13g2_nand3_1 _9008_ (.B(_1560_),
    .C(_1565_),
    .A(_3905_),
    .Y(_3925_));
 sg13g2_a21o_1 _9009_ (.A2(_3925_),
    .A1(_3924_),
    .B1(_1568_),
    .X(_3926_));
 sg13g2_nor2b_1 _9010_ (.A(_3908_),
    .B_N(_3600_),
    .Y(_3927_));
 sg13g2_a21oi_1 _9011_ (.A1(_3910_),
    .A2(_3927_),
    .Y(_3928_),
    .B1(_1563_));
 sg13g2_o21ai_1 _9012_ (.B1(net77),
    .Y(_3929_),
    .A1(_3903_),
    .A2(_3928_));
 sg13g2_nand3_1 _9013_ (.B(_3926_),
    .C(_3929_),
    .A(_2546_),
    .Y(_3930_));
 sg13g2_nand2_1 _9014_ (.Y(_3931_),
    .A(_3930_),
    .B(_3779_));
 sg13g2_o21ai_1 _9015_ (.B1(_3931_),
    .Y(_0211_),
    .A1(_3714_),
    .A2(_2574_));
 sg13g2_nor2_1 _9016_ (.A(_3714_),
    .B(_2586_),
    .Y(_0212_));
 sg13g2_nor2_1 _9017_ (.A(_3714_),
    .B(_2588_),
    .Y(_0213_));
 sg13g2_a21oi_1 _9018_ (.A1(_1236_),
    .A2(_4228_),
    .Y(\i_display.i_vga.hblank_tmp ),
    .B1(_1233_));
 sg13g2_inv_1 _9019_ (.Y(_3932_),
    .A(_0049_));
 sg13g2_nor2b_1 _9020_ (.A(net122),
    .B_N(_0048_),
    .Y(_3933_));
 sg13g2_nor3_1 _9021_ (.A(_1020_),
    .B(_1010_),
    .C(_3933_),
    .Y(_3934_));
 sg13g2_o21ai_1 _9022_ (.B1(_0048_),
    .Y(_3935_),
    .A1(_4230_),
    .A2(_1080_));
 sg13g2_a21oi_1 _9023_ (.A1(_3934_),
    .A2(_3935_),
    .Y(_3936_),
    .B1(_4227_));
 sg13g2_nor3_1 _9024_ (.A(_3932_),
    .B(_1233_),
    .C(_3936_),
    .Y(\i_display.i_vga.hsync_tmp ));
 sg13g2_nor2b_1 _9025_ (.A(_1232_),
    .B_N(_3147_),
    .Y(_3937_));
 sg13g2_nor2_1 _9026_ (.A(_1083_),
    .B(_1013_),
    .Y(_3938_));
 sg13g2_nor2_1 _9027_ (.A(_3938_),
    .B(_1230_),
    .Y(_3939_));
 sg13g2_o21ai_1 _9028_ (.B1(_1231_),
    .Y(_3940_),
    .A1(_1068_),
    .A2(_0051_));
 sg13g2_and2_1 _9029_ (.A(_3939_),
    .B(_3940_),
    .X(_3941_));
 sg13g2_nand3_1 _9030_ (.B(_1068_),
    .C(_0051_),
    .A(_1231_),
    .Y(_3942_));
 sg13g2_inv_1 _9031_ (.Y(_3943_),
    .A(_1232_));
 sg13g2_a22oi_1 _9032_ (.Y(_3944_),
    .B1(_3184_),
    .B2(_3943_),
    .A2(_3942_),
    .A1(_3939_));
 sg13g2_nor4_1 _9033_ (.A(_0050_),
    .B(_3937_),
    .C(_3941_),
    .D(_3944_),
    .Y(\i_display.i_vga.timing_ver.sync_tmp ));
 sg13g2_nand3_1 _9034_ (.B(_1098_),
    .C(_1004_),
    .A(_3938_),
    .Y(_3945_));
 sg13g2_nor4_1 _9035_ (.A(_1041_),
    .B(_1023_),
    .C(_1228_),
    .D(_3945_),
    .Y(_3946_));
 sg13g2_nand4_1 _9036_ (.B(_0712_),
    .C(_0981_),
    .A(_3946_),
    .Y(_3947_),
    .D(_0051_));
 sg13g2_nand2_1 _9037_ (.Y(\i_display.i_vga.timing_ver.blank ),
    .A(_3947_),
    .B(_1150_));
 sg13g2_nor2b_1 _9038_ (.A(net108),
    .B_N(_0062_),
    .Y(_3948_));
 sg13g2_a21oi_1 _9039_ (.A1(_0063_),
    .A2(net108),
    .Y(_3949_),
    .B1(_3948_));
 sg13g2_nor2_1 _9040_ (.A(_3932_),
    .B(net111),
    .Y(_3950_));
 sg13g2_a21oi_1 _9041_ (.A1(_0070_),
    .A2(net108),
    .Y(_3951_),
    .B1(_3950_));
 sg13g2_inv_1 _9042_ (.Y(_3952_),
    .A(_3951_));
 sg13g2_nor2_1 _9043_ (.A(_3949_),
    .B(_3952_),
    .Y(_3953_));
 sg13g2_nand2_1 _9044_ (.Y(_3954_),
    .A(_3952_),
    .B(_3949_));
 sg13g2_nand2b_1 _9045_ (.Y(_3955_),
    .B(_3954_),
    .A_N(_3953_));
 sg13g2_nor2b_1 _9046_ (.A(_1494_),
    .B_N(_0072_),
    .Y(_3956_));
 sg13g2_a21oi_1 _9047_ (.A1(_0071_),
    .A2(net111),
    .Y(_3957_),
    .B1(_3956_));
 sg13g2_inv_1 _9048_ (.Y(_3958_),
    .A(_0060_));
 sg13g2_buf_1 _9049_ (.A(net115),
    .X(_3959_));
 sg13g2_nor2_1 _9050_ (.A(_3958_),
    .B(net109),
    .Y(_3960_));
 sg13g2_a21oi_1 _9051_ (.A1(_0061_),
    .A2(net111),
    .Y(_3961_),
    .B1(_3960_));
 sg13g2_inv_1 _9052_ (.Y(_3962_),
    .A(_3961_));
 sg13g2_nor2_1 _9053_ (.A(_3957_),
    .B(_3962_),
    .Y(_3963_));
 sg13g2_nand2_1 _9054_ (.Y(_3964_),
    .A(_3962_),
    .B(_3957_));
 sg13g2_inv_1 _9055_ (.Y(_3965_),
    .A(_3964_));
 sg13g2_nor2_1 _9056_ (.A(_3963_),
    .B(_3965_),
    .Y(_3966_));
 sg13g2_nand2_1 _9057_ (.Y(_3967_),
    .A(net111),
    .B(_3932_));
 sg13g2_o21ai_1 _9058_ (.B1(_3967_),
    .Y(_3968_),
    .A1(_0071_),
    .A2(net111));
 sg13g2_nor2b_1 _9059_ (.A(net109),
    .B_N(_0061_),
    .Y(_3969_));
 sg13g2_a21oi_1 _9060_ (.A1(_0062_),
    .A2(net111),
    .Y(_3970_),
    .B1(_3969_));
 sg13g2_inv_1 _9061_ (.Y(_3971_),
    .A(_3970_));
 sg13g2_nor2_1 _9062_ (.A(_3968_),
    .B(_3971_),
    .Y(_3972_));
 sg13g2_nand2_1 _9063_ (.Y(_3973_),
    .A(_3971_),
    .B(_3968_));
 sg13g2_inv_1 _9064_ (.Y(_3974_),
    .A(_3973_));
 sg13g2_nor2_1 _9065_ (.A(_3972_),
    .B(_3974_),
    .Y(_3975_));
 sg13g2_nand2_1 _9066_ (.Y(_3976_),
    .A(_3966_),
    .B(_3975_));
 sg13g2_inv_1 _9067_ (.Y(_3977_),
    .A(_0058_));
 sg13g2_nor2_1 _9068_ (.A(_0056_),
    .B(net115),
    .Y(_3978_));
 sg13g2_a21oi_1 _9069_ (.A1(_3977_),
    .A2(net115),
    .Y(_3979_),
    .B1(_3978_));
 sg13g2_inv_1 _9070_ (.Y(_3980_),
    .A(_0075_));
 sg13g2_nor2_1 _9071_ (.A(_3980_),
    .B(net115),
    .Y(_3981_));
 sg13g2_a21oi_1 _9072_ (.A1(_0074_),
    .A2(net115),
    .Y(_3982_),
    .B1(_3981_));
 sg13g2_inv_1 _9073_ (.Y(_3983_),
    .A(_0076_));
 sg13g2_inv_1 _9074_ (.Y(_3984_),
    .A(_0056_));
 sg13g2_a22oi_1 _9075_ (.Y(_3985_),
    .B1(_3984_),
    .B2(_1493_),
    .A2(_0102_),
    .A1(_3983_));
 sg13g2_o21ai_1 _9076_ (.B1(_3985_),
    .Y(_3986_),
    .A1(_0076_),
    .A2(net109));
 sg13g2_a21oi_1 _9077_ (.A1(_1158_),
    .A2(_3980_),
    .Y(_3987_),
    .B1(_1488_));
 sg13g2_nand4_1 _9078_ (.B(_3984_),
    .C(_3983_),
    .A(net109),
    .Y(_3988_),
    .D(_0102_));
 sg13g2_o21ai_1 _9079_ (.B1(_3988_),
    .Y(_3989_),
    .A1(_3979_),
    .A2(_3982_));
 sg13g2_a21oi_1 _9080_ (.A1(_3986_),
    .A2(_3987_),
    .Y(_3990_),
    .B1(_3989_));
 sg13g2_a21o_1 _9081_ (.A2(_3982_),
    .A1(_3979_),
    .B1(_3990_),
    .X(_3991_));
 sg13g2_nor2b_1 _9082_ (.A(net109),
    .B_N(_0074_),
    .Y(_3992_));
 sg13g2_a21oi_1 _9083_ (.A1(_0048_),
    .A2(_3959_),
    .Y(_3993_),
    .B1(_3992_));
 sg13g2_inv_1 _9084_ (.Y(_3994_),
    .A(_3993_));
 sg13g2_nor2_1 _9085_ (.A(_3977_),
    .B(net109),
    .Y(_3995_));
 sg13g2_a21oi_1 _9086_ (.A1(_0057_),
    .A2(_1494_),
    .Y(_3996_),
    .B1(_3995_));
 sg13g2_nand2_1 _9087_ (.Y(_3997_),
    .A(_3994_),
    .B(_3996_));
 sg13g2_nor2_1 _9088_ (.A(_3996_),
    .B(_3994_),
    .Y(_3998_));
 sg13g2_a21o_1 _9089_ (.A2(_3997_),
    .A1(_3991_),
    .B1(_3998_),
    .X(_3999_));
 sg13g2_nor2b_1 _9090_ (.A(_3959_),
    .B_N(_0073_),
    .Y(_4000_));
 sg13g2_a21oi_1 _9091_ (.A1(_0072_),
    .A2(net111),
    .Y(_4001_),
    .B1(_4000_));
 sg13g2_nand2_1 _9092_ (.Y(_4002_),
    .A(net109),
    .B(_3958_));
 sg13g2_o21ai_1 _9093_ (.B1(_4002_),
    .Y(_4003_),
    .A1(_0059_),
    .A2(net109));
 sg13g2_xor2_1 _9094_ (.B(_4003_),
    .A(_4001_),
    .X(_4004_));
 sg13g2_nor2b_1 _9095_ (.A(net115),
    .B_N(_0057_),
    .Y(_4005_));
 sg13g2_a21oi_1 _9096_ (.A1(_0059_),
    .A2(net115),
    .Y(_4006_),
    .B1(_4005_));
 sg13g2_a21oi_1 _9097_ (.A1(_0073_),
    .A2(_1493_),
    .Y(_4007_),
    .B1(_3933_));
 sg13g2_inv_1 _9098_ (.Y(_4008_),
    .A(_4007_));
 sg13g2_nor2_1 _9099_ (.A(_4006_),
    .B(_4008_),
    .Y(_4009_));
 sg13g2_inv_1 _9100_ (.Y(_4010_),
    .A(_4009_));
 sg13g2_nand2_1 _9101_ (.Y(_4011_),
    .A(_4008_),
    .B(_4006_));
 sg13g2_nand2_1 _9102_ (.Y(_4012_),
    .A(_4010_),
    .B(_4011_));
 sg13g2_nor2_1 _9103_ (.A(_4004_),
    .B(_4012_),
    .Y(_4013_));
 sg13g2_inv_1 _9104_ (.Y(_4014_),
    .A(_4001_));
 sg13g2_nor2_1 _9105_ (.A(_4003_),
    .B(_4014_),
    .Y(_4015_));
 sg13g2_inv_1 _9106_ (.Y(_4016_),
    .A(_4015_));
 sg13g2_o21ai_1 _9107_ (.B1(_4016_),
    .Y(_4017_),
    .A1(_4010_),
    .A2(_4004_));
 sg13g2_a21oi_1 _9108_ (.A1(_3999_),
    .A2(_4013_),
    .Y(_4018_),
    .B1(_4017_));
 sg13g2_a21oi_1 _9109_ (.A1(_3975_),
    .A2(_3965_),
    .Y(_4019_),
    .B1(_3974_));
 sg13g2_o21ai_1 _9110_ (.B1(_4019_),
    .Y(_4020_),
    .A1(_3976_),
    .A2(_4018_));
 sg13g2_xnor2_1 _9111_ (.Y(_4021_),
    .A(_3955_),
    .B(_4020_));
 sg13g2_o21ai_1 _9112_ (.B1(_4011_),
    .Y(_4022_),
    .A1(_4009_),
    .A2(_3999_));
 sg13g2_nor2_1 _9113_ (.A(_4015_),
    .B(_3965_),
    .Y(_4023_));
 sg13g2_o21ai_1 _9114_ (.B1(_4023_),
    .Y(_4024_),
    .A1(_4004_),
    .A2(_4022_));
 sg13g2_nor2b_1 _9115_ (.A(_3963_),
    .B_N(_4024_),
    .Y(_4025_));
 sg13g2_xnor2_1 _9116_ (.Y(_4026_),
    .A(_3975_),
    .B(_4025_));
 sg13g2_nor2_1 _9117_ (.A(_3998_),
    .B(_4012_),
    .Y(_4027_));
 sg13g2_nor2b_1 _9118_ (.A(_4027_),
    .B_N(_3991_),
    .Y(_4028_));
 sg13g2_a21oi_1 _9119_ (.A1(_3997_),
    .A2(_4012_),
    .Y(_4029_),
    .B1(_4027_));
 sg13g2_a21oi_1 _9120_ (.A1(_3991_),
    .A2(_3997_),
    .Y(_4030_),
    .B1(_4029_));
 sg13g2_xnor2_1 _9121_ (.Y(_4031_),
    .A(_3966_),
    .B(_4018_));
 sg13g2_xor2_1 _9122_ (.B(_4022_),
    .A(_4004_),
    .X(_4032_));
 sg13g2_nor4_1 _9123_ (.A(_4028_),
    .B(_4030_),
    .C(_4031_),
    .D(_4032_),
    .Y(_4033_));
 sg13g2_nand2_1 _9124_ (.Y(_4034_),
    .A(_4026_),
    .B(_4033_));
 sg13g2_nor2b_1 _9125_ (.A(net108),
    .B_N(_0070_),
    .Y(_4035_));
 sg13g2_a21oi_1 _9126_ (.A1(_0047_),
    .A2(net108),
    .Y(_4036_),
    .B1(_4035_));
 sg13g2_inv_1 _9127_ (.Y(_4037_),
    .A(_4036_));
 sg13g2_buf_1 _9128_ (.A(\i_music.i_sample.thresh[9] ),
    .X(_4038_));
 sg13g2_mux2_1 _9129_ (.A0(\i_music.i_sample.thresh[8] ),
    .A1(_4038_),
    .S(_1495_),
    .X(_4039_));
 sg13g2_nor2_1 _9130_ (.A(_4037_),
    .B(_4039_),
    .Y(_4040_));
 sg13g2_nand2_1 _9131_ (.Y(_4041_),
    .A(_4039_),
    .B(_4037_));
 sg13g2_nand2b_1 _9132_ (.Y(_4042_),
    .B(_4041_),
    .A_N(_4040_));
 sg13g2_nor2_1 _9133_ (.A(_3953_),
    .B(_4020_),
    .Y(_4043_));
 sg13g2_nor2b_1 _9134_ (.A(_4043_),
    .B_N(_3954_),
    .Y(_4044_));
 sg13g2_xnor2_1 _9135_ (.Y(_4045_),
    .A(_4042_),
    .B(_4044_));
 sg13g2_xor2_1 _9136_ (.B(\i_music.i_sample.thresh[10] ),
    .A(_1587_),
    .X(_4046_));
 sg13g2_xnor2_1 _9137_ (.Y(_4047_),
    .A(_4237_),
    .B(_4038_));
 sg13g2_nor2_1 _9138_ (.A(net108),
    .B(_4047_),
    .Y(_4048_));
 sg13g2_a21oi_1 _9139_ (.A1(_1495_),
    .A2(_4046_),
    .Y(_4049_),
    .B1(_4048_));
 sg13g2_a21oi_1 _9140_ (.A1(_4044_),
    .A2(_4041_),
    .Y(_4050_),
    .B1(_4040_));
 sg13g2_xnor2_1 _9141_ (.Y(_4051_),
    .A(_4049_),
    .B(_4050_));
 sg13g2_nor4_2 _9142_ (.A(_4021_),
    .B(_4034_),
    .C(_4045_),
    .Y(_4052_),
    .D(_4051_));
 sg13g2_nand2_1 _9143_ (.Y(_4053_),
    .A(_4052_),
    .B(net100));
 sg13g2_a21oi_1 _9144_ (.A1(_4053_),
    .A2(net133),
    .Y(\i_music.i_sample.t1.CG.GCLK ),
    .B1(clknet_5_12__leaf_clk));
 sg13g2_nor2_1 _9145_ (.A(\i_music.i_sample.sample_idx[0] ),
    .B(net119),
    .Y(\i_music.i_sample.t1.genblk1[0].state.D ));
 sg13g2_nor2b_1 _9146_ (.A(_2134_),
    .B_N(\i_music.i_sample.thresh[0] ),
    .Y(_4054_));
 sg13g2_xnor2_1 _9147_ (.Y(_4055_),
    .A(_0056_),
    .B(_2123_));
 sg13g2_nand2_1 _9148_ (.Y(_4056_),
    .A(_4054_),
    .B(_4055_));
 sg13g2_nand2_1 _9149_ (.Y(_4057_),
    .A(_2123_),
    .B(\i_music.i_sample.thresh[1] ));
 sg13g2_nand2_1 _9150_ (.Y(_4058_),
    .A(_4056_),
    .B(_4057_));
 sg13g2_nand2_1 _9151_ (.Y(_4059_),
    .A(_2155_),
    .B(_2151_));
 sg13g2_xor2_1 _9152_ (.B(_4059_),
    .A(\i_music.i_sample.thresh[2] ),
    .X(_4060_));
 sg13g2_o21ai_1 _9153_ (.B1(net133),
    .Y(_4061_),
    .A1(_4058_),
    .A2(_4060_));
 sg13g2_nand2_1 _9154_ (.Y(_4062_),
    .A(_4060_),
    .B(_4058_));
 sg13g2_nor2b_1 _9155_ (.A(_4061_),
    .B_N(_4062_),
    .Y(\i_music.i_sample.t1.genblk1[10].state.D ));
 sg13g2_xnor2_1 _9156_ (.Y(_4063_),
    .A(_0057_),
    .B(_2143_));
 sg13g2_nand2_1 _9157_ (.Y(_4064_),
    .A(_4059_),
    .B(_3977_));
 sg13g2_nand2_1 _9158_ (.Y(_4065_),
    .A(_4062_),
    .B(_4064_));
 sg13g2_o21ai_1 _9159_ (.B1(net133),
    .Y(_4066_),
    .A1(_4063_),
    .A2(_4065_));
 sg13g2_nand2_1 _9160_ (.Y(_4067_),
    .A(_4065_),
    .B(_4063_));
 sg13g2_nor2b_1 _9161_ (.A(_4066_),
    .B_N(_4067_),
    .Y(\i_music.i_sample.t1.genblk1[11].state.D ));
 sg13g2_xnor2_1 _9162_ (.Y(_4068_),
    .A(_0059_),
    .B(_2060_));
 sg13g2_nand2_1 _9163_ (.Y(_4069_),
    .A(_2143_),
    .B(\i_music.i_sample.thresh[3] ));
 sg13g2_nand2_1 _9164_ (.Y(_4070_),
    .A(_4067_),
    .B(_4069_));
 sg13g2_o21ai_1 _9165_ (.B1(net133),
    .Y(_4071_),
    .A1(_4068_),
    .A2(_4070_));
 sg13g2_nand2_1 _9166_ (.Y(_4072_),
    .A(_4070_),
    .B(_4068_));
 sg13g2_nor2b_1 _9167_ (.A(_4071_),
    .B_N(_4072_),
    .Y(\i_music.i_sample.t1.genblk1[12].state.D ));
 sg13g2_xnor2_1 _9168_ (.Y(_4073_),
    .A(_0060_),
    .B(_2085_));
 sg13g2_nand2_1 _9169_ (.Y(_4074_),
    .A(_2060_),
    .B(\i_music.i_sample.thresh[4] ));
 sg13g2_nand2_1 _9170_ (.Y(_4075_),
    .A(_4072_),
    .B(_4074_));
 sg13g2_o21ai_1 _9171_ (.B1(net134),
    .Y(_4076_),
    .A1(_4073_),
    .A2(_4075_));
 sg13g2_nand2_1 _9172_ (.Y(_4077_),
    .A(_4075_),
    .B(_4073_));
 sg13g2_nor2b_1 _9173_ (.A(_4076_),
    .B_N(_4077_),
    .Y(\i_music.i_sample.t1.genblk1[13].state.D ));
 sg13g2_xnor2_1 _9174_ (.Y(_4078_),
    .A(_0061_),
    .B(_2095_));
 sg13g2_nand2_1 _9175_ (.Y(_4079_),
    .A(_2085_),
    .B(\i_music.i_sample.thresh[5] ));
 sg13g2_nand2_1 _9176_ (.Y(_4080_),
    .A(_4077_),
    .B(_4079_));
 sg13g2_o21ai_1 _9177_ (.B1(net134),
    .Y(_4081_),
    .A1(_4078_),
    .A2(_4080_));
 sg13g2_nand2_1 _9178_ (.Y(_4082_),
    .A(_4080_),
    .B(_4078_));
 sg13g2_nor2b_1 _9179_ (.A(_4081_),
    .B_N(_4082_),
    .Y(\i_music.i_sample.t1.genblk1[14].state.D ));
 sg13g2_xnor2_1 _9180_ (.Y(_4083_),
    .A(_0062_),
    .B(_2077_));
 sg13g2_nand2_1 _9181_ (.Y(_4084_),
    .A(_2095_),
    .B(\i_music.i_sample.thresh[6] ));
 sg13g2_nand2_1 _9182_ (.Y(_4085_),
    .A(_4082_),
    .B(_4084_));
 sg13g2_o21ai_1 _9183_ (.B1(net134),
    .Y(_4086_),
    .A1(_4083_),
    .A2(_4085_));
 sg13g2_nand2_1 _9184_ (.Y(_4087_),
    .A(_4085_),
    .B(_4083_));
 sg13g2_nor2b_1 _9185_ (.A(_4086_),
    .B_N(_4087_),
    .Y(\i_music.i_sample.t1.genblk1[15].state.D ));
 sg13g2_nand2_1 _9186_ (.Y(_4088_),
    .A(_2077_),
    .B(\i_music.i_sample.thresh[7] ));
 sg13g2_nand2_1 _9187_ (.Y(_4089_),
    .A(_4087_),
    .B(_4088_));
 sg13g2_xnor2_1 _9188_ (.Y(_4090_),
    .A(_0063_),
    .B(_2113_));
 sg13g2_o21ai_1 _9189_ (.B1(net134),
    .Y(_4091_),
    .A1(_4090_),
    .A2(_4089_));
 sg13g2_a21oi_1 _9190_ (.A1(_4089_),
    .A2(_4090_),
    .Y(\i_music.i_sample.t1.genblk1[16].state.D ),
    .B1(_4091_));
 sg13g2_nand2_1 _9191_ (.Y(_4092_),
    .A(_4089_),
    .B(_4090_));
 sg13g2_nand2_1 _9192_ (.Y(_4093_),
    .A(_2113_),
    .B(\i_music.i_sample.thresh[8] ));
 sg13g2_xnor2_1 _9193_ (.Y(_4094_),
    .A(_4038_),
    .B(_2108_));
 sg13g2_a21oi_1 _9194_ (.A1(_4092_),
    .A2(_4093_),
    .Y(_4095_),
    .B1(_4094_));
 sg13g2_and3_1 _9195_ (.X(_4096_),
    .A(_4092_),
    .B(_4093_),
    .C(_4094_));
 sg13g2_nor3_1 _9196_ (.A(_3590_),
    .B(_4095_),
    .C(_4096_),
    .Y(\i_music.i_sample.t1.genblk1[17].state.D ));
 sg13g2_inv_1 _9197_ (.Y(_4097_),
    .A(_4083_));
 sg13g2_o21ai_1 _9198_ (.B1(_4088_),
    .Y(_4098_),
    .A1(_4097_),
    .A2(_4084_));
 sg13g2_nor2b_1 _9199_ (.A(_4094_),
    .B_N(_4090_),
    .Y(_4099_));
 sg13g2_inv_1 _9200_ (.Y(_4100_),
    .A(_4063_));
 sg13g2_o21ai_1 _9201_ (.B1(_4069_),
    .Y(_4101_),
    .A1(_4100_),
    .A2(_4064_));
 sg13g2_and2_1 _9202_ (.A(_4073_),
    .B(_4068_),
    .X(_4102_));
 sg13g2_nand2_1 _9203_ (.Y(_4103_),
    .A(_4101_),
    .B(_4102_));
 sg13g2_nand2b_1 _9204_ (.Y(_4104_),
    .B(_4073_),
    .A_N(_4074_));
 sg13g2_nand3_1 _9205_ (.B(_4104_),
    .C(_4079_),
    .A(_4103_),
    .Y(_4105_));
 sg13g2_and3_1 _9206_ (.X(_4106_),
    .A(_4078_),
    .B(_4083_),
    .C(_4099_));
 sg13g2_nand2_1 _9207_ (.Y(_4107_),
    .A(_2108_),
    .B(_4038_));
 sg13g2_o21ai_1 _9208_ (.B1(_4107_),
    .Y(_4108_),
    .A1(_4094_),
    .A2(_4093_));
 sg13g2_a221oi_1 _9209_ (.B2(_4106_),
    .C1(_4108_),
    .B1(_4105_),
    .A1(_4098_),
    .Y(_4109_),
    .A2(_4099_));
 sg13g2_nor2b_1 _9210_ (.A(_4100_),
    .B_N(_4060_),
    .Y(_4110_));
 sg13g2_nand4_1 _9211_ (.B(_4058_),
    .C(_4102_),
    .A(_4110_),
    .Y(_4111_),
    .D(_4106_));
 sg13g2_xor2_1 _9212_ (.B(_2101_),
    .A(\i_music.i_sample.thresh[10] ),
    .X(_4112_));
 sg13g2_a21oi_1 _9213_ (.A1(_4109_),
    .A2(_4111_),
    .Y(_4113_),
    .B1(_4112_));
 sg13g2_and3_1 _9214_ (.X(_4114_),
    .A(_4109_),
    .B(_4111_),
    .C(_4112_));
 sg13g2_nor3_1 _9215_ (.A(net125),
    .B(_4113_),
    .C(_4114_),
    .Y(\i_music.i_sample.t1.genblk1[18].state.D ));
 sg13g2_nor2_1 _9216_ (.A(\i_music.i_sample.sample_idx[1] ),
    .B(\i_music.i_sample.sample_idx[0] ),
    .Y(_4115_));
 sg13g2_nand2_1 _9217_ (.Y(_4116_),
    .A(\i_music.i_sample.sample_idx[1] ),
    .B(\i_music.i_sample.sample_idx[0] ));
 sg13g2_inv_1 _9218_ (.Y(_4117_),
    .A(_4116_));
 sg13g2_nor3_1 _9219_ (.A(net125),
    .B(_4115_),
    .C(_4117_),
    .Y(\i_music.i_sample.t1.genblk1[1].state.D ));
 sg13g2_nor2_1 _9220_ (.A(\i_music.i_sample.sample_idx[2] ),
    .B(_4117_),
    .Y(_4118_));
 sg13g2_nand2_1 _9221_ (.Y(_4119_),
    .A(_4117_),
    .B(\i_music.i_sample.sample_idx[2] ));
 sg13g2_inv_1 _9222_ (.Y(_4120_),
    .A(_4119_));
 sg13g2_nor3_1 _9223_ (.A(net125),
    .B(_4118_),
    .C(_4120_),
    .Y(\i_music.i_sample.t1.genblk1[2].state.D ));
 sg13g2_nor2_1 _9224_ (.A(\i_music.i_sample.sample_idx[3] ),
    .B(_4120_),
    .Y(_4121_));
 sg13g2_nand2_1 _9225_ (.Y(_4122_),
    .A(_4120_),
    .B(\i_music.i_sample.sample_idx[3] ));
 sg13g2_inv_1 _9226_ (.Y(_4123_),
    .A(_4122_));
 sg13g2_nor3_1 _9227_ (.A(net125),
    .B(_4121_),
    .C(_4123_),
    .Y(\i_music.i_sample.t1.genblk1[3].state.D ));
 sg13g2_nor2_1 _9228_ (.A(\i_music.i_sample.sample_idx[4] ),
    .B(_4123_),
    .Y(_4124_));
 sg13g2_nand2_1 _9229_ (.Y(_4125_),
    .A(_4123_),
    .B(\i_music.i_sample.sample_idx[4] ));
 sg13g2_inv_1 _9230_ (.Y(_4126_),
    .A(_4125_));
 sg13g2_nor3_1 _9231_ (.A(net128),
    .B(_4124_),
    .C(_4126_),
    .Y(\i_music.i_sample.t1.genblk1[4].state.D ));
 sg13g2_nor2_1 _9232_ (.A(\i_music.i_sample.sample_idx[5] ),
    .B(_4126_),
    .Y(_4127_));
 sg13g2_nand2_1 _9233_ (.Y(_4128_),
    .A(_4126_),
    .B(\i_music.i_sample.sample_idx[5] ));
 sg13g2_inv_1 _9234_ (.Y(_4129_),
    .A(_4128_));
 sg13g2_nor3_1 _9235_ (.A(net128),
    .B(_4127_),
    .C(_4129_),
    .Y(\i_music.i_sample.t1.genblk1[5].state.D ));
 sg13g2_nor2_1 _9236_ (.A(\i_music.i_sample.sample_idx[6] ),
    .B(_4129_),
    .Y(_4130_));
 sg13g2_nand2_1 _9237_ (.Y(_4131_),
    .A(_4129_),
    .B(\i_music.i_sample.sample_idx[6] ));
 sg13g2_inv_1 _9238_ (.Y(_4132_),
    .A(_4131_));
 sg13g2_nor3_1 _9239_ (.A(net128),
    .B(_4130_),
    .C(_4132_),
    .Y(\i_music.i_sample.t1.genblk1[6].state.D ));
 sg13g2_nor2b_1 _9240_ (.A(_4131_),
    .B_N(\i_music.i_sample.sample_idx[7] ),
    .Y(_4133_));
 sg13g2_nor2_1 _9241_ (.A(\i_music.i_sample.sample_idx[7] ),
    .B(_4132_),
    .Y(_4134_));
 sg13g2_nor3_1 _9242_ (.A(net128),
    .B(_4133_),
    .C(_4134_),
    .Y(\i_music.i_sample.t1.genblk1[7].state.D ));
 sg13g2_a21oi_1 _9243_ (.A1(_2128_),
    .A2(_2133_),
    .Y(_4135_),
    .B1(\i_music.i_sample.thresh[0] ));
 sg13g2_nor3_1 _9244_ (.A(_1666_),
    .B(_4135_),
    .C(_4054_),
    .Y(\i_music.i_sample.t1.genblk1[8].state.D ));
 sg13g2_o21ai_1 _9245_ (.B1(net134),
    .Y(_4136_),
    .A1(_4055_),
    .A2(_4054_));
 sg13g2_nor2b_1 _9246_ (.A(_4136_),
    .B_N(_4056_),
    .Y(\i_music.i_sample.t1.genblk1[9].state.D ));
 sg13g2_nand2_1 _9247_ (.Y(_4137_),
    .A(_4052_),
    .B(_1485_));
 sg13g2_a21oi_1 _9248_ (.A1(_4137_),
    .A2(net133),
    .Y(\i_music.i_sample.t2.CG.GCLK ),
    .B1(clknet_5_12__leaf_clk));
 sg13g2_nand2_1 _9249_ (.Y(_4138_),
    .A(_4052_),
    .B(_1483_));
 sg13g2_a21oi_1 _9250_ (.A1(_4138_),
    .A2(net133),
    .Y(\i_music.i_sample.t3.CG.GCLK ),
    .B1(clknet_5_6__leaf_clk));
 sg13g2_nand2_1 _9251_ (.Y(_4139_),
    .A(_4052_),
    .B(_1500_));
 sg13g2_a21oi_1 _9252_ (.A1(_4139_),
    .A2(net133),
    .Y(\i_music.i_sample.t4.CG.GCLK ),
    .B1(clknet_5_12__leaf_clk));
 sg13g2_nor2b_1 _9253_ (.A(net131),
    .B_N(\i_display.colour[5] ),
    .Y(net10));
 sg13g2_nor2b_1 _9254_ (.A(net131),
    .B_N(\i_display.colour[3] ),
    .Y(net11));
 sg13g2_nor2b_1 _9255_ (.A(net131),
    .B_N(\i_display.colour[1] ),
    .Y(net12));
 sg13g2_nor2b_1 _9256_ (.A(net131),
    .B_N(\i_display.colour[4] ),
    .Y(net14));
 sg13g2_nor2b_1 _9257_ (.A(_0709_),
    .B_N(\i_display.colour[2] ),
    .Y(net15));
 sg13g2_nor2b_1 _9258_ (.A(_0709_),
    .B_N(\i_display.colour[0] ),
    .Y(net16));
 sg13g2_dfrbp_1 _9259_ (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net180),
    .D(_0000_),
    .Q_N(_4685_),
    .Q(_0024_));
 sg13g2_dfrbp_1 _9260_ (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net181),
    .D(_0001_),
    .Q_N(_4684_),
    .Q(_0025_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _9259__180 (.L_HI(net180));
 sg13g2_buf_1 _9263_ (.A(net166),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9264_ (.A(net167),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9265_ (.A(net168),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9266_ (.A(net169),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9267_ (.A(net170),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9268_ (.A(net171),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9269_ (.A(net172),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9270_ (.A(net182),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9271_ (.A(net173),
    .X(uio_out[0]));
 sg13g2_buf_1 _9272_ (.A(net174),
    .X(uio_out[1]));
 sg13g2_buf_1 _9273_ (.A(net175),
    .X(uio_out[2]));
 sg13g2_buf_1 _9274_ (.A(net176),
    .X(uio_out[3]));
 sg13g2_buf_1 _9275_ (.A(net177),
    .X(uio_out[4]));
 sg13g2_buf_1 _9276_ (.A(net178),
    .X(uio_out[5]));
 sg13g2_buf_1 _9277_ (.A(net179),
    .X(uio_out[6]));
 sg13g2_buf_1 _9278_ (.A(\i_music.i_pwm.pwm ),
    .X(net9));
 sg13g2_buf_1 _9279_ (.A(\i_display.i_vga.timing_ver.sync ),
    .X(net13));
 sg13g2_buf_1 _9280_ (.A(\i_display.hsync ),
    .X(net17));
 sg13g2_dfrbp_1 \i_display.colour[0]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net183),
    .D(_0106_),
    .Q_N(_4683_),
    .Q(\i_display.colour[0] ));
 sg13g2_dfrbp_1 \i_display.colour[1]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3295_clk),
    .RESET_B(net184),
    .D(_0107_),
    .Q_N(_4682_),
    .Q(\i_display.colour[1] ));
 sg13g2_dfrbp_1 \i_display.colour[2]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net185),
    .D(_0108_),
    .Q_N(_4681_),
    .Q(\i_display.colour[2] ));
 sg13g2_dfrbp_1 \i_display.colour[3]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3295_clk),
    .RESET_B(net186),
    .D(_0109_),
    .Q_N(_4680_),
    .Q(\i_display.colour[3] ));
 sg13g2_dfrbp_1 \i_display.colour[4]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3295_clk),
    .RESET_B(net187),
    .D(_0110_),
    .Q_N(_4679_),
    .Q(\i_display.colour[4] ));
 sg13g2_dfrbp_1 \i_display.colour[5]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3295_clk),
    .RESET_B(net188),
    .D(_0111_),
    .Q_N(_4678_),
    .Q(\i_display.colour[5] ));
 sg13g2_dfrbp_1 \i_display.frame[0]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net189),
    .D(_0112_),
    .Q_N(_0096_),
    .Q(\i_display.frame[0] ));
 sg13g2_dfrbp_1 \i_display.frame[1]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_1647_clk),
    .RESET_B(net190),
    .D(_0113_),
    .Q_N(_0090_),
    .Q(\i_display.frame[1] ));
 sg13g2_dfrbp_1 \i_display.frame[2]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net191),
    .D(_0114_),
    .Q_N(_0092_),
    .Q(\i_display.frame[2] ));
 sg13g2_dfrbp_1 \i_display.frame[3]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_1647_clk),
    .RESET_B(net192),
    .D(_0115_),
    .Q_N(_0094_),
    .Q(\i_display.frame[3] ));
 sg13g2_dfrbp_1 \i_display.frame[4]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net193),
    .D(_0116_),
    .Q_N(_0097_),
    .Q(\i_display.frame[4] ));
 sg13g2_dfrbp_1 \i_display.frame[5]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net194),
    .D(_0117_),
    .Q_N(_0099_),
    .Q(\i_display.frame[5] ));
 sg13g2_dfrbp_1 \i_display.frame[6]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net195),
    .D(_0118_),
    .Q_N(_0028_),
    .Q(\i_display.frame[6] ));
 sg13g2_dfrbp_1 \i_display.frame[7]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net196),
    .D(_0119_),
    .Q_N(_0036_),
    .Q(\i_display.frame[7] ));
 sg13g2_dfrbp_1 \i_display.frame[8]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2780_clk),
    .RESET_B(net197),
    .D(_0120_),
    .Q_N(_0038_),
    .Q(\i_display.frame[8] ));
 sg13g2_dfrbp_1 \i_display.frame[9]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_1647_clk),
    .RESET_B(net198),
    .D(_0121_),
    .Q_N(_0040_),
    .Q(\i_display.frame[9] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[0]$_DFFE_PP_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net199),
    .D(_0122_),
    .Q_N(_4677_),
    .Q(\i_display.frame_crotchet[0] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[1]$_DFFE_PP_  (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net200),
    .D(_0123_),
    .Q_N(_0065_),
    .Q(\i_display.frame_crotchet[1] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[2]$_DFFE_PP_  (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net201),
    .D(_0124_),
    .Q_N(_0066_),
    .Q(\i_display.frame_crotchet[2] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[3]$_DFFE_PP_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net202),
    .D(_0125_),
    .Q_N(_0067_),
    .Q(\i_display.frame_crotchet[3] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[4]$_DFFE_PP_  (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net203),
    .D(_0126_),
    .Q_N(_0054_),
    .Q(\i_display.frame_crotchet[4] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[5]$_DFFE_PP_  (.CLK(clknet_level_2_1_3192_clk),
    .RESET_B(net204),
    .D(_0127_),
    .Q_N(_0068_),
    .Q(\i_display.frame_crotchet[5] ));
 sg13g2_dfrbp_1 \i_display.frame_crotchet[6]$_DFFE_PP_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net205),
    .D(_0128_),
    .Q_N(_0069_),
    .Q(\i_display.frame_crotchet[6] ));
 sg13g2_dfrbp_1 \i_display.i_vga.hblank$_DFF_P_  (.CLK(clknet_level_2_1_2883_clk),
    .RESET_B(net206),
    .D(\i_display.i_vga.hblank_tmp ),
    .Q_N(_4686_),
    .Q(\i_display.i_vga.hblank ));
 sg13g2_dfrbp_1 \i_display.i_vga.hsync$_DFF_P_  (.CLK(clknet_level_2_1_1647_clk),
    .RESET_B(net207),
    .D(\i_display.i_vga.hsync_tmp ),
    .Q_N(_4676_),
    .Q(\i_display.hsync ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[0]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2883_clk),
    .RESET_B(net208),
    .D(_0129_),
    .Q_N(_0051_),
    .Q(\i_display.i_vga.timing_ver.counter[0] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[10]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net209),
    .D(_0130_),
    .Q_N(_0050_),
    .Q(\i_display.i_vga.timing_ver.counter[10] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[1]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2883_clk),
    .RESET_B(net210),
    .D(_0131_),
    .Q_N(_4675_),
    .Q(\i_display.i_vga.timing_ver.counter[1] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[2]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net211),
    .D(_0132_),
    .Q_N(_4674_),
    .Q(\i_display.i_vga.timing_ver.counter[2] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net212),
    .D(_0133_),
    .Q_N(_0052_),
    .Q(\i_display.i_vga.timing_ver.counter[3] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net213),
    .D(_0134_),
    .Q_N(_4673_),
    .Q(\i_display.i_vga.timing_ver.counter[4] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[5]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net214),
    .D(_0135_),
    .Q_N(_4672_),
    .Q(\i_display.i_vga.timing_ver.counter[5] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[6]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net215),
    .D(_0136_),
    .Q_N(_4671_),
    .Q(\i_display.i_vga.timing_ver.counter[6] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[7]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net216),
    .D(_0137_),
    .Q_N(_4670_),
    .Q(\i_display.i_vga.timing_ver.counter[7] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[8]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net217),
    .D(_0138_),
    .Q_N(_4669_),
    .Q(\i_display.i_vga.timing_ver.counter[8] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.counter[9]$_SDFFE_PN1P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net218),
    .D(_0139_),
    .Q_N(_4687_),
    .Q(\i_display.i_vga.timing_ver.counter[9] ));
 sg13g2_dfrbp_1 \i_display.i_vga.timing_ver.sync$_DFF_P_  (.CLK(clknet_level_2_1_3295_clk),
    .RESET_B(net219),
    .D(\i_display.i_vga.timing_ver.sync_tmp ),
    .Q_N(_4688_),
    .Q(\i_display.i_vga.timing_ver.sync ));
 sg13g2_dfrbp_1 \i_display.i_vga.vblank$_DFF_P_  (.CLK(clknet_level_2_1_2883_clk),
    .RESET_B(net220),
    .D(\i_display.i_vga.timing_ver.blank ),
    .Q_N(_4668_),
    .Q(\i_display.i_vga.vblank ));
 sg13g2_dfrbp_1 \i_display.in_line$_SDFFE_PP0P_  (.CLK(clknet_level_2_1_1647_clk),
    .RESET_B(net221),
    .D(_0140_),
    .Q_N(_0026_),
    .Q(\i_display.in_line ));
 sg13g2_dfrbp_1 \i_display.x_idx_r[0]$_SDFFE_PP0P_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net222),
    .D(_0141_),
    .Q_N(_0101_),
    .Q(\i_display.x_idx[0] ));
 sg13g2_dfrbp_1 \i_display.x_idx_r[1]$_SDFFE_PP0P_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net223),
    .D(_0142_),
    .Q_N(_4667_),
    .Q(\i_display.x_idx[1] ));
 sg13g2_dfrbp_1 \i_display.y_idx[0]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net224),
    .D(_0143_),
    .Q_N(_0034_),
    .Q(\i_display.x_idx[2] ));
 sg13g2_dfrbp_1 \i_display.y_idx[1]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net225),
    .D(_0144_),
    .Q_N(_0033_),
    .Q(\i_display.x_idx[3] ));
 sg13g2_dfrbp_1 \i_display.y_idx[2]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net226),
    .D(_0145_),
    .Q_N(_0032_),
    .Q(\i_display.x_idx[4] ));
 sg13g2_dfrbp_1 \i_display.y_idx[3]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_1235_clk),
    .RESET_B(net227),
    .D(_0146_),
    .Q_N(_0031_),
    .Q(\i_display.x_idx[5] ));
 sg13g2_dfrbp_1 \i_display.y_idx[4]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_1235_clk),
    .RESET_B(net228),
    .D(_0147_),
    .Q_N(_0087_),
    .Q(\i_display.x_idx[6] ));
 sg13g2_dfrbp_1 \i_display.y_idx[5]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net229),
    .D(_0148_),
    .Q_N(_0030_),
    .Q(\i_display.x_idx[7] ));
 sg13g2_dfrbp_1 \i_display.y_idx[6]$_SDFFE_PN0N_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net230),
    .D(_0149_),
    .Q_N(_0089_),
    .Q(\i_display.x_idx[8] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[0]$_DFF_P_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net231),
    .D(_0011_),
    .Q_N(_0100_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-5] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[1]$_DFF_P_  (.CLK(clknet_level_2_1_720_clk),
    .RESET_B(net232),
    .D(_0012_),
    .Q_N(_0098_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-4] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[2]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net233),
    .D(_0013_),
    .Q_N(_0095_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-3] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[3]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net234),
    .D(_0014_),
    .Q_N(_0093_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-2] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[4]$_DFF_P_  (.CLK(clknet_level_2_1_1235_clk),
    .RESET_B(net235),
    .D(_0015_),
    .Q_N(_0091_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[-1] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[5]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net236),
    .D(_0016_),
    .Q_N(_0088_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[0] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[6]$_DFF_P_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net237),
    .D(_0017_),
    .Q_N(_0027_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[1] ));
 sg13g2_dfrbp_1 \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[7]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net238),
    .D(_0018_),
    .Q_N(_0035_),
    .Q(\i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[2] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[0]$_DFF_P_  (.CLK(clknet_level_2_1_1235_clk),
    .RESET_B(net239),
    .D(_0002_),
    .Q_N(_0029_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[0] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[1]$_DFF_P_  (.CLK(clknet_level_2_1_1235_clk),
    .RESET_B(net240),
    .D(_0003_),
    .Q_N(_0037_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[1] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[2]$_DFF_P_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net241),
    .D(_0004_),
    .Q_N(_0039_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[2] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[3]$_DFF_P_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net242),
    .D(_0005_),
    .Q_N(_0041_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[3] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[4]$_DFF_P_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net243),
    .D(_0006_),
    .Q_N(_0042_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[4] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[5]$_DFF_P_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net244),
    .D(_0007_),
    .Q_N(_0043_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[5] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[6]$_DFF_P_  (.CLK(clknet_level_2_1_1132_clk),
    .RESET_B(net245),
    .D(_0008_),
    .Q_N(_0044_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[6] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[7]$_DFF_P_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net246),
    .D(_0009_),
    .Q_N(_0045_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[7] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[8]$_DFF_P_  (.CLK(clknet_level_2_1_926_clk),
    .RESET_B(net247),
    .D(_0010_),
    .Q_N(_0046_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[8] ));
 sg13g2_dfrbp_1 \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[9]$_SDFF_PP0_  (.CLK(clknet_level_2_1_1544_clk),
    .RESET_B(net248),
    .D(_0150_),
    .Q_N(_4689_),
    .Q(\i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[9] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0]$_DFF_P_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net249),
    .D(_0019_),
    .Q_N(_4666_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10]$_SDFF_PP1_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net250),
    .D(_0151_),
    .Q_N(_4665_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1]$_SDFF_PP1_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net251),
    .D(_0152_),
    .Q_N(_4690_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[2]$_DFF_P_  (.CLK(clknet_level_2_1_2471_clk),
    .RESET_B(net252),
    .D(_0020_),
    .Q_N(_4664_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[2] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3]$_SDFF_PP0_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net253),
    .D(_0153_),
    .Q_N(_4663_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4]$_SDFF_PP1_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net254),
    .D(_0154_),
    .Q_N(_0055_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[5]$_SDFF_PN1_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net255),
    .D(_0155_),
    .Q_N(_4691_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[5] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[6]$_DFF_P_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net256),
    .D(_0021_),
    .Q_N(_4692_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[6] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7]$_DFF_P_  (.CLK(clknet_level_2_1_2574_clk),
    .RESET_B(net257),
    .D(_0022_),
    .Q_N(_4693_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7] ));
 sg13g2_dfrbp_1 \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8]$_DFF_P_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net258),
    .D(_0023_),
    .Q_N(_4662_),
    .Q(\i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8] ));
 sg13g2_dfrbp_1 \i_music.count[0]$_SDFF_PN1_  (.CLK(clknet_level_2_1_823_clk),
    .RESET_B(net259),
    .D(_0156_),
    .Q_N(_0102_),
    .Q(\i_display.i_vga.low_count[0] ));
 sg13g2_dfrbp_1 \i_music.count[10]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net260),
    .D(_0157_),
    .Q_N(_4661_),
    .Q(\i_music.count[10] ));
 sg13g2_dfrbp_1 \i_music.count[11]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net261),
    .D(_0158_),
    .Q_N(_4660_),
    .Q(\i_music.count[11] ));
 sg13g2_dfrbp_1 \i_music.count[12]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2471_clk),
    .RESET_B(net262),
    .D(_0159_),
    .Q_N(_4659_),
    .Q(\i_music.count[12] ));
 sg13g2_dfrbp_1 \i_music.count[13]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net263),
    .D(_0160_),
    .Q_N(_4658_),
    .Q(\i_music.count[13] ));
 sg13g2_dfrbp_1 \i_music.count[14]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net264),
    .D(_0161_),
    .Q_N(_4657_),
    .Q(\i_music.count[14] ));
 sg13g2_dfrbp_1 \i_music.count[15]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net265),
    .D(_0162_),
    .Q_N(_4656_),
    .Q(\i_music.count[15] ));
 sg13g2_dfrbp_1 \i_music.count[16]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net266),
    .D(_0163_),
    .Q_N(_4655_),
    .Q(\i_music.count[16] ));
 sg13g2_dfrbp_1 \i_music.count[17]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net267),
    .D(_0164_),
    .Q_N(_4654_),
    .Q(\i_music.count[17] ));
 sg13g2_dfrbp_1 \i_music.count[18]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net268),
    .D(_0165_),
    .Q_N(_4653_),
    .Q(\i_music.count[18] ));
 sg13g2_dfrbp_1 \i_music.count[19]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2471_clk),
    .RESET_B(net269),
    .D(_0166_),
    .Q_N(_4652_),
    .Q(\i_music.count[19] ));
 sg13g2_dfrbp_1 \i_music.count[1]$_SDFF_PN0_  (.CLK(clknet_level_2_1_823_clk),
    .RESET_B(net270),
    .D(_0167_),
    .Q_N(_0075_),
    .Q(\i_display.i_vga.low_count[1] ));
 sg13g2_dfrbp_1 \i_music.count[20]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2471_clk),
    .RESET_B(net271),
    .D(_0168_),
    .Q_N(_4651_),
    .Q(\i_music.count[20] ));
 sg13g2_dfrbp_1 \i_music.count[21]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net272),
    .D(_0169_),
    .Q_N(_4650_),
    .Q(\i_music.count[21] ));
 sg13g2_dfrbp_1 \i_music.count[22]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net273),
    .D(_0170_),
    .Q_N(_0077_),
    .Q(\i_music.count[22] ));
 sg13g2_dfrbp_1 \i_music.count[23]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2471_clk),
    .RESET_B(net274),
    .D(_0171_),
    .Q_N(_4649_),
    .Q(\i_music.count[23] ));
 sg13g2_dfrbp_1 \i_music.count[24]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2677_clk),
    .RESET_B(net275),
    .D(_0172_),
    .Q_N(_4648_),
    .Q(\i_music.count[24] ));
 sg13g2_dfrbp_1 \i_music.count[25]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net276),
    .D(_0173_),
    .Q_N(_0053_),
    .Q(\crotchet[0] ));
 sg13g2_dfrbp_1 \i_music.count[26]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net277),
    .D(_0174_),
    .Q_N(_4647_),
    .Q(\crotchet[1] ));
 sg13g2_dfrbp_1 \i_music.count[27]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2368_clk),
    .RESET_B(net278),
    .D(_0175_),
    .Q_N(_4646_),
    .Q(\crotchet[2] ));
 sg13g2_dfrbp_1 \i_music.count[28]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net279),
    .D(_0176_),
    .Q_N(_4645_),
    .Q(\crotchet[3] ));
 sg13g2_dfrbp_1 \i_music.count[29]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net280),
    .D(_0177_),
    .Q_N(_4644_),
    .Q(\crotchet[4] ));
 sg13g2_dfrbp_1 \i_music.count[2]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net281),
    .D(_0178_),
    .Q_N(_0074_),
    .Q(\i_display.i_vga.low_count[2] ));
 sg13g2_dfrbp_1 \i_music.count[30]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2986_clk),
    .RESET_B(net282),
    .D(_0179_),
    .Q_N(_4643_),
    .Q(\crotchet[5] ));
 sg13g2_dfrbp_1 \i_music.count[31]$_SDFF_PN0_  (.CLK(clknet_level_2_1_3089_clk),
    .RESET_B(net283),
    .D(_0180_),
    .Q_N(_4642_),
    .Q(\crotchet[6] ));
 sg13g2_dfrbp_1 \i_music.count[3]$_SDFF_PN0_  (.CLK(clknet_level_2_1_2883_clk),
    .RESET_B(net284),
    .D(_0181_),
    .Q_N(_0048_),
    .Q(\i_display.i_vga.low_count[3] ));
 sg13g2_dfrbp_1 \i_music.count[4]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net285),
    .D(_0182_),
    .Q_N(_0073_),
    .Q(\i_display.i_vga.low_count[4] ));
 sg13g2_dfrbp_1 \i_music.count[5]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net286),
    .D(_0183_),
    .Q_N(_0072_),
    .Q(\i_display.i_vga.low_count[5] ));
 sg13g2_dfrbp_1 \i_music.count[6]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net287),
    .D(_0184_),
    .Q_N(_0071_),
    .Q(\i_display.i_vga.low_count[6] ));
 sg13g2_dfrbp_1 \i_music.count[7]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net288),
    .D(_0185_),
    .Q_N(_0049_),
    .Q(\i_display.i_vga.low_count[7] ));
 sg13g2_dfrbp_1 \i_music.count[8]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1338_clk),
    .RESET_B(net289),
    .D(_0186_),
    .Q_N(_0070_),
    .Q(\i_display.i_vga.low_count[8] ));
 sg13g2_dfrbp_1 \i_music.count[9]$_SDFF_PN0_  (.CLK(clknet_level_2_1_1338_clk),
    .RESET_B(net290),
    .D(_0187_),
    .Q_N(_0047_),
    .Q(\i_display.i_vga.low_count[9] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[0]$_SDFF_PP0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net291),
    .D(_0188_),
    .Q_N(_0105_),
    .Q(\i_music.i_pwm.count[0] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[1]$_SDFF_PP0_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net292),
    .D(_0189_),
    .Q_N(_4641_),
    .Q(\i_music.i_pwm.count[1] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[2]$_SDFF_PP0_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net293),
    .D(_0190_),
    .Q_N(_4640_),
    .Q(\i_music.i_pwm.count[2] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[3]$_SDFF_PP0_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net294),
    .D(_0191_),
    .Q_N(_4639_),
    .Q(\i_music.i_pwm.count[3] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[4]$_SDFF_PP0_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net295),
    .D(_0192_),
    .Q_N(_4638_),
    .Q(\i_music.i_pwm.count[4] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[5]$_SDFF_PP0_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net296),
    .D(_0193_),
    .Q_N(_4637_),
    .Q(\i_music.i_pwm.count[5] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[6]$_SDFF_PP0_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net297),
    .D(_0194_),
    .Q_N(_4636_),
    .Q(\i_music.i_pwm.count[6] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.count[7]$_SDFF_PP0_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net298),
    .D(_0195_),
    .Q_N(_4635_),
    .Q(\i_music.i_pwm.count[7] ));
 sg13g2_dfrbp_1 \i_music.i_pwm.pwm$_DFFE_PP_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net299),
    .D(_0196_),
    .Q_N(_4634_),
    .Q(\i_music.i_pwm.pwm ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[0]$_DFFE_PP_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net300),
    .D(_0197_),
    .Q_N(_4633_),
    .Q(\i_music.i_pwm.sample[0] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[1]$_DFFE_PP_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net301),
    .D(_0198_),
    .Q_N(_4632_),
    .Q(\i_music.i_pwm.sample[1] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[2]$_DFFE_PP_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net302),
    .D(_0199_),
    .Q_N(_4631_),
    .Q(\i_music.i_pwm.sample[2] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[3]$_DFFE_PP_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net303),
    .D(_0200_),
    .Q_N(_4630_),
    .Q(\i_music.i_pwm.sample[3] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[4]$_DFFE_PP_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net304),
    .D(_0201_),
    .Q_N(_4629_),
    .Q(\i_music.i_pwm.sample[4] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[5]$_DFFE_PP_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net305),
    .D(_0202_),
    .Q_N(_4628_),
    .Q(\i_music.i_pwm.sample[5] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[6]$_DFFE_PP_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net306),
    .D(_0203_),
    .Q_N(_4627_),
    .Q(\i_music.i_pwm.sample[6] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample[7]$_DFFE_PP_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net307),
    .D(_0204_),
    .Q_N(_4626_),
    .Q(\i_music.i_pwm.sample[7] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[0]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net308),
    .D(_0205_),
    .Q_N(_4625_),
    .Q(\i_music.i_sample.sample_acc[0] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[1]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net309),
    .D(_0206_),
    .Q_N(_4624_),
    .Q(\i_music.i_sample.sample_acc[1] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[2]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net310),
    .D(_0207_),
    .Q_N(_4623_),
    .Q(\i_music.i_sample.sample_acc[2] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[3]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net311),
    .D(_0208_),
    .Q_N(_4622_),
    .Q(\i_music.i_sample.sample_acc[3] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[4]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net312),
    .D(_0209_),
    .Q_N(_4621_),
    .Q(\i_music.i_sample.sample_acc[4] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[5]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net313),
    .D(_0210_),
    .Q_N(_4620_),
    .Q(\i_music.i_sample.sample_acc[5] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[6]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net314),
    .D(_0211_),
    .Q_N(_4619_),
    .Q(\i_music.i_sample.sample_acc[6] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[7]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net315),
    .D(_0212_),
    .Q_N(_0064_),
    .Q(\i_music.i_sample.sample_acc[7] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_acc[8]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net316),
    .D(_0213_),
    .Q_N(_4694_),
    .Q(\i_music.i_sample.sample_acc[8] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[0]$_DFF_P_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net317),
    .D(_0241_),
    .Q_N(_4695_),
    .Q(\i_music.i_sample.sample_idx[0] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[1]$_DFF_P_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net318),
    .D(_0242_),
    .Q_N(_4696_),
    .Q(\i_music.i_sample.sample_idx[1] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[2]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net319),
    .D(_0243_),
    .Q_N(_4697_),
    .Q(\i_music.i_sample.sample_idx[2] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[3]$_DFF_P_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net320),
    .D(_0244_),
    .Q_N(_4698_),
    .Q(\i_music.i_sample.sample_idx[3] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[4]$_DFF_P_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net321),
    .D(_0245_),
    .Q_N(_4699_),
    .Q(\i_music.i_sample.sample_idx[4] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[5]$_DFF_P_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net322),
    .D(_0246_),
    .Q_N(_4700_),
    .Q(\i_music.i_sample.sample_idx[5] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[6]$_DFF_P_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net323),
    .D(_0247_),
    .Q_N(_4701_),
    .Q(\i_music.i_sample.sample_idx[6] ));
 sg13g2_dfrbp_1 \i_music.i_sample.sample_idx[7]$_DFF_P_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net324),
    .D(_0248_),
    .Q_N(_4702_),
    .Q(\i_music.i_sample.sample_idx[7] ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[0].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[0].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[10].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[10].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[11].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[11].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[12].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[12].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[13].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[13].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[14].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[14].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[15].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[15].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[16].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[16].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[17].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[17].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[18].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[18].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[18].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[1].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[1].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[2].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[2].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[3].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[3].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[4].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[4].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[5].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[5].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[6].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[6].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[7].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[7].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[8].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[8].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t1.genblk1[9].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ),
    .Q(\i_music.i_sample.t1.genblk1[9].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[0].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[0].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[10].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[10].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[11].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[11].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[12].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[12].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[13].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[13].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[14].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[14].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[15].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[15].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[16].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[16].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[17].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[17].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[1].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[1].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[2].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[2].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[3].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[3].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[4].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[4].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[5].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[5].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[6].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[6].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[7].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[7].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[8].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[8].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t2.genblk1[9].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ),
    .Q(\i_music.i_sample.t2.genblk1[9].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[0].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[0].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[10].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[10].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[11].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[11].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[12].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[12].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[13].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[13].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[14].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[14].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[15].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[15].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[16].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[16].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[17].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[17].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[1].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[1].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[2].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[2].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[3].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[3].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[4].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[4].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[5].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[5].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[6].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[6].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[7].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[7].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[8].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[8].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t3.genblk1[9].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ),
    .Q(\i_music.i_sample.t3.genblk1[9].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[0].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[0].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[0].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[10].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[10].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[10].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[11].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[11].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[11].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[12].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[12].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[12].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[13].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[13].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[13].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[14].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[14].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[14].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[15].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[15].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[15].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[16].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[16].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[16].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[17].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[17].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[17].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[1].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[1].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[1].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[2].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[2].state.D ),
    .GATE(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[2].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[3].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[3].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[3].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[4].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[4].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[4].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[5].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[5].state.D ),
    .GATE(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[5].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[6].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[6].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[6].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[7].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[7].state.D ),
    .GATE(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[7].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[8].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[8].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[8].state.Q ));
 sg13g2_dlhq_1 \i_music.i_sample.t4.genblk1[9].state.pf.ul.Q$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\i_music.i_sample.t1.genblk1[9].state.D ),
    .GATE(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ),
    .Q(\i_music.i_sample.t4.genblk1[9].state.Q ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[0]$_DFF_P_  (.CLK(clknet_level_2_1_823_clk),
    .RESET_B(net325),
    .D(_0249_),
    .Q_N(_0076_),
    .Q(\i_music.i_sample.thresh[0] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[10]$_DFF_P_  (.CLK(clknet_level_2_1_1441_clk),
    .RESET_B(net326),
    .D(_0250_),
    .Q_N(_4703_),
    .Q(\i_music.i_sample.thresh[10] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[1]$_DFF_P_  (.CLK(clknet_level_2_1_823_clk),
    .RESET_B(net327),
    .D(_0251_),
    .Q_N(_0056_),
    .Q(\i_music.i_sample.thresh[1] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[2]$_DFF_P_  (.CLK(clknet_level_2_1_720_clk),
    .RESET_B(net328),
    .D(_0252_),
    .Q_N(_0058_),
    .Q(\i_music.i_sample.thresh[2] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[3]$_DFF_P_  (.CLK(clknet_level_2_1_720_clk),
    .RESET_B(net329),
    .D(_0253_),
    .Q_N(_0057_),
    .Q(\i_music.i_sample.thresh[3] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[4]$_DFF_P_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net330),
    .D(_0254_),
    .Q_N(_0059_),
    .Q(\i_music.i_sample.thresh[4] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[5]$_DFF_P_  (.CLK(clknet_level_2_1_514_clk),
    .RESET_B(net331),
    .D(_0255_),
    .Q_N(_0060_),
    .Q(\i_music.i_sample.thresh[5] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[6]$_DFF_P_  (.CLK(clknet_level_2_1_720_clk),
    .RESET_B(net332),
    .D(_0256_),
    .Q_N(_0061_),
    .Q(\i_music.i_sample.thresh[6] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[7]$_DFF_P_  (.CLK(clknet_level_2_1_720_clk),
    .RESET_B(net333),
    .D(_0257_),
    .Q_N(_0062_),
    .Q(\i_music.i_sample.thresh[7] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[8]$_DFF_P_  (.CLK(clknet_level_2_1_1338_clk),
    .RESET_B(net334),
    .D(_0258_),
    .Q_N(_0063_),
    .Q(\i_music.i_sample.thresh[8] ));
 sg13g2_dfrbp_1 \i_music.i_sample.thresh[9]$_DFF_P_  (.CLK(clknet_level_2_1_1029_clk),
    .RESET_B(net335),
    .D(_0259_),
    .Q_N(_4618_),
    .Q(\i_music.i_sample.thresh[9] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][0]$_SDFFCE_PP1P_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net336),
    .D(_0214_),
    .Q_N(_0103_),
    .Q(\i_music.violin_note_idx[1][0] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][1]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_823_clk),
    .RESET_B(net337),
    .D(_0215_),
    .Q_N(_0082_),
    .Q(\i_music.violin_note_idx[1][1] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net338),
    .D(_0216_),
    .Q_N(_0083_),
    .Q(\i_music.violin_note_idx[1][2] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net339),
    .D(_0217_),
    .Q_N(_0079_),
    .Q(\i_music.violin_note_idx[1][3] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][4]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net340),
    .D(_0218_),
    .Q_N(_0080_),
    .Q(\i_music.violin_note_idx[1][4] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][5]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net341),
    .D(_0219_),
    .Q_N(_0078_),
    .Q(\i_music.violin_note_idx[1][5] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][6]$_DFFE_PP_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net342),
    .D(_0220_),
    .Q_N(_0081_),
    .Q(\i_music.violin_note_idx[1][6] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][7]$_DFFE_PP_  (.CLK(clknet_level_2_1_2162_clk),
    .RESET_B(net343),
    .D(_0221_),
    .Q_N(_0084_),
    .Q(\i_music.violin_note_idx[1][7] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[1][8]$_DFFE_PP_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net344),
    .D(_0222_),
    .Q_N(_0086_),
    .Q(\i_music.violin_note_idx[1][8] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][0]$_SDFFCE_PP1P_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net345),
    .D(_0223_),
    .Q_N(_0104_),
    .Q(\i_music.violin_note_idx[2][0] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][1]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net346),
    .D(_0224_),
    .Q_N(_4617_),
    .Q(\i_music.violin_note_idx[2][1] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net347),
    .D(_0225_),
    .Q_N(_4616_),
    .Q(\i_music.violin_note_idx[2][2] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][3]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net348),
    .D(_0226_),
    .Q_N(_4615_),
    .Q(\i_music.violin_note_idx[2][3] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][4]$_DFFE_PP_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net349),
    .D(_0227_),
    .Q_N(_4614_),
    .Q(\i_music.violin_note_idx[2][4] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][5]$_DFFE_PP_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net350),
    .D(_0228_),
    .Q_N(_4613_),
    .Q(\i_music.violin_note_idx[2][5] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][6]$_DFFE_PP_  (.CLK(clknet_level_2_1_2265_clk),
    .RESET_B(net351),
    .D(_0229_),
    .Q_N(_4612_),
    .Q(\i_music.violin_note_idx[2][6] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][7]$_DFFE_PP_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net352),
    .D(_0230_),
    .Q_N(_4611_),
    .Q(\i_music.violin_note_idx[2][7] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[2][8]$_DFFE_PP_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net353),
    .D(_0231_),
    .Q_N(_4610_),
    .Q(\i_music.violin_note_idx[2][8] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][0]$_SDFFCE_PP1P_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net354),
    .D(_0232_),
    .Q_N(_4609_),
    .Q(\i_music.violin_note_idx[3][0] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][1]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_1956_clk),
    .RESET_B(net355),
    .D(_0233_),
    .Q_N(_4608_),
    .Q(\i_music.violin_note_idx[3][1] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][2]$_SDFFCE_PN1P_  (.CLK(clknet_level_2_1_617_clk),
    .RESET_B(net356),
    .D(_0234_),
    .Q_N(_4607_),
    .Q(\i_music.violin_note_idx[3][2] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][3]$_SDFFCE_PN0P_  (.CLK(clknet_level_2_1_2059_clk),
    .RESET_B(net357),
    .D(_0235_),
    .Q_N(_4606_),
    .Q(\i_music.violin_note_idx[3][3] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][4]$_DFFE_PP_  (.CLK(clknet_level_2_1_1853_clk),
    .RESET_B(net358),
    .D(_0236_),
    .Q_N(_4605_),
    .Q(\i_music.violin_note_idx[3][4] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][5]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net359),
    .D(_0237_),
    .Q_N(_4604_),
    .Q(\i_music.violin_note_idx[3][5] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][6]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net360),
    .D(_0238_),
    .Q_N(_4603_),
    .Q(\i_music.violin_note_idx[3][6] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][7]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net361),
    .D(_0239_),
    .Q_N(_0085_),
    .Q(\i_music.violin_note_idx[3][7] ));
 sg13g2_dfrbp_1 \i_music.violin_note_idx[3][8]$_DFFE_PP_  (.CLK(clknet_level_2_1_1750_clk),
    .RESET_B(net362),
    .D(_0240_),
    .Q_N(_4602_),
    .Q(\i_music.violin_note_idx[3][8] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[7]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout18 (.A(_1306_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_1226_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1366_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1348_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1333_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1225_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1355_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1314_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1271_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1167_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1242_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2546_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2470_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2468_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2464_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2262_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2475_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2258_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2233_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2201_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_2192_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_2172_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2164_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2755_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2702_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2633_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2272_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2236_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2224_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2220_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2210_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2171_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_3657_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_3645_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_3638_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2247_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2198_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2190_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2183_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2170_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1560_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1549_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1543_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_3742_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_3723_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_3628_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_3627_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_3609_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_3269_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1565_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1559_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1554_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1548_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_3715_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_3626_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_3605_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1558_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1553_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1541_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1568_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1546_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1536_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1531_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_3146_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_4328_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_4534_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_4368_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0705_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0640_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1882_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1814_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1623_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1240_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0704_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_4325_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1798_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1757_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1748_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1745_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1728_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1693_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1681_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1534_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1496_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_4289_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1773_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1741_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1735_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1692_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1680_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1495_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_3959_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1707_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1494_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1483_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2396_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1501_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1493_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_1482_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_3565_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_3549_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_3479_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2644_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1500_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1492_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1486_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_1481_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_3590_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2832_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_2634_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1666_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1499_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1158_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0709_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0649_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_3449_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2690_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1665_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1530_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1193_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1157_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0672_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0667_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0663_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2835_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_1637_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1627_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1489_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1488_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_1308_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1180_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_1178_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0711_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0647_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_4463_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_4294_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_4163_),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_4144_));
 sg13g2_buf_2 fanout156 (.A(_1629_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_1380_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0413_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0410_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_4494_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_4313_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_4158_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_4146_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_4142_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_4140_),
    .X(net165));
 sg13g2_tielo _9263__166 (.L_LO(net166));
 sg13g2_tielo _9264__167 (.L_LO(net167));
 sg13g2_tielo _9265__168 (.L_LO(net168));
 sg13g2_tielo _9266__169 (.L_LO(net169));
 sg13g2_tielo _9267__170 (.L_LO(net170));
 sg13g2_tielo _9268__171 (.L_LO(net171));
 sg13g2_tielo _9269__172 (.L_LO(net172));
 sg13g2_tielo _9271__173 (.L_LO(net173));
 sg13g2_tielo _9272__174 (.L_LO(net174));
 sg13g2_tielo _9273__175 (.L_LO(net175));
 sg13g2_tielo _9274__176 (.L_LO(net176));
 sg13g2_tielo _9275__177 (.L_LO(net177));
 sg13g2_tielo _9276__178 (.L_LO(net178));
 sg13g2_tielo _9277__179 (.L_LO(net179));
 sg13g2_tiehi _9260__181 (.L_HI(net181));
 sg13g2_tiehi _9270__182 (.L_HI(net182));
 sg13g2_tiehi \i_display.colour[0]$_SDFF_PN0__183  (.L_HI(net183));
 sg13g2_tiehi \i_display.colour[1]$_SDFF_PN0__184  (.L_HI(net184));
 sg13g2_tiehi \i_display.colour[2]$_SDFF_PN0__185  (.L_HI(net185));
 sg13g2_tiehi \i_display.colour[3]$_SDFF_PN0__186  (.L_HI(net186));
 sg13g2_tiehi \i_display.colour[4]$_SDFF_PN0__187  (.L_HI(net187));
 sg13g2_tiehi \i_display.colour[5]$_SDFF_PN0__188  (.L_HI(net188));
 sg13g2_tiehi \i_display.frame[0]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \i_display.frame[1]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \i_display.frame[2]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \i_display.frame[3]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \i_display.frame[4]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \i_display.frame[5]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \i_display.frame[6]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \i_display.frame[7]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \i_display.frame[8]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \i_display.frame[9]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \i_display.frame_crotchet[0]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \i_display.frame_crotchet[1]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \i_display.frame_crotchet[2]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \i_display.frame_crotchet[3]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \i_display.frame_crotchet[4]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \i_display.frame_crotchet[5]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \i_display.frame_crotchet[6]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \i_display.i_vga.hblank$_DFF_P__206  (.L_HI(net206));
 sg13g2_tiehi \i_display.i_vga.hsync$_DFF_P__207  (.L_HI(net207));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[0]$_SDFFE_PN1P__208  (.L_HI(net208));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[10]$_SDFFE_PN1P__209  (.L_HI(net209));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[1]$_SDFFE_PN1P__210  (.L_HI(net210));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[2]$_SDFFE_PN1P__211  (.L_HI(net211));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[3]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[4]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[5]$_SDFFE_PN1P__214  (.L_HI(net214));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[6]$_SDFFE_PN1P__215  (.L_HI(net215));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[7]$_SDFFE_PN1P__216  (.L_HI(net216));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[8]$_SDFFE_PN1P__217  (.L_HI(net217));
 sg13g2_tiehi \i_display.i_vga.timing_ver.counter[9]$_SDFFE_PN1P__218  (.L_HI(net218));
 sg13g2_tiehi \i_display.i_vga.timing_ver.sync$_DFF_P__219  (.L_HI(net219));
 sg13g2_tiehi \i_display.i_vga.vblank$_DFF_P__220  (.L_HI(net220));
 sg13g2_tiehi \i_display.in_line$_SDFFE_PP0P__221  (.L_HI(net221));
 sg13g2_tiehi \i_display.x_idx_r[0]$_SDFFE_PP0P__222  (.L_HI(net222));
 sg13g2_tiehi \i_display.x_idx_r[1]$_SDFFE_PP0P__223  (.L_HI(net223));
 sg13g2_tiehi \i_display.y_idx[0]$_SDFFE_PN0N__224  (.L_HI(net224));
 sg13g2_tiehi \i_display.y_idx[1]$_SDFFE_PN0N__225  (.L_HI(net225));
 sg13g2_tiehi \i_display.y_idx[2]$_SDFFE_PN0N__226  (.L_HI(net226));
 sg13g2_tiehi \i_display.y_idx[3]$_SDFFE_PN0N__227  (.L_HI(net227));
 sg13g2_tiehi \i_display.y_idx[4]$_SDFFE_PN0N__228  (.L_HI(net228));
 sg13g2_tiehi \i_display.y_idx[5]$_SDFFE_PN0N__229  (.L_HI(net229));
 sg13g2_tiehi \i_display.y_idx[6]$_SDFFE_PN0N__230  (.L_HI(net230));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[0]$_DFF_P__231  (.L_HI(net231));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[1]$_DFF_P__232  (.L_HI(net232));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[2]$_DFF_P__233  (.L_HI(net233));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[3]$_DFF_P__234  (.L_HI(net234));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[4]$_DFF_P__235  (.L_HI(net235));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[5]$_DFF_P__236  (.L_HI(net236));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[6]$_DFF_P__237  (.L_HI(net237));
 sg13g2_tiehi \i_display.y_offset$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:565$10.$result[7]$_DFF_P__238  (.L_HI(net238));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[0]$_DFF_P__239  (.L_HI(net239));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[1]$_DFF_P__240  (.L_HI(net240));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[2]$_DFF_P__241  (.L_HI(net241));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[3]$_DFF_P__242  (.L_HI(net242));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[4]$_DFF_P__243  (.L_HI(net243));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[5]$_DFF_P__244  (.L_HI(net244));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[6]$_DFF_P__245  (.L_HI(net245));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[7]$_DFF_P__246  (.L_HI(net246));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[8]$_DFF_P__247  (.L_HI(net247));
 sg13g2_tiehi \i_display.y_value$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/display.sv:567$12.$result[9]$_SDFF_PP0__248  (.L_HI(net248));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[0]$_DFF_P__249  (.L_HI(net249));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[10]$_SDFF_PP1__250  (.L_HI(net250));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[1]$_SDFF_PP1__251  (.L_HI(net251));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[2]$_DFF_P__252  (.L_HI(net252));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[3]$_SDFF_PP0__253  (.L_HI(net253));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[4]$_SDFF_PP1__254  (.L_HI(net254));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[5]$_SDFF_PN1__255  (.L_HI(net255));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[6]$_DFF_P__256  (.L_HI(net256));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[7]$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \i_music.cello_rom$func$/home/runner/work/ttihp0p2-demo-canon/ttihp0p2-demo-canon/src/music.v:430$166.$result[8]$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \i_music.count[0]$_SDFF_PN1__259  (.L_HI(net259));
 sg13g2_tiehi \i_music.count[10]$_SDFF_PN0__260  (.L_HI(net260));
 sg13g2_tiehi \i_music.count[11]$_SDFF_PN0__261  (.L_HI(net261));
 sg13g2_tiehi \i_music.count[12]$_SDFF_PN0__262  (.L_HI(net262));
 sg13g2_tiehi \i_music.count[13]$_SDFF_PN0__263  (.L_HI(net263));
 sg13g2_tiehi \i_music.count[14]$_SDFF_PN0__264  (.L_HI(net264));
 sg13g2_tiehi \i_music.count[15]$_SDFF_PN0__265  (.L_HI(net265));
 sg13g2_tiehi \i_music.count[16]$_SDFF_PN0__266  (.L_HI(net266));
 sg13g2_tiehi \i_music.count[17]$_SDFF_PN0__267  (.L_HI(net267));
 sg13g2_tiehi \i_music.count[18]$_SDFF_PN0__268  (.L_HI(net268));
 sg13g2_tiehi \i_music.count[19]$_SDFF_PN0__269  (.L_HI(net269));
 sg13g2_tiehi \i_music.count[1]$_SDFF_PN0__270  (.L_HI(net270));
 sg13g2_tiehi \i_music.count[20]$_SDFF_PN0__271  (.L_HI(net271));
 sg13g2_tiehi \i_music.count[21]$_SDFF_PN0__272  (.L_HI(net272));
 sg13g2_tiehi \i_music.count[22]$_SDFF_PN0__273  (.L_HI(net273));
 sg13g2_tiehi \i_music.count[23]$_SDFF_PN0__274  (.L_HI(net274));
 sg13g2_tiehi \i_music.count[24]$_SDFF_PN0__275  (.L_HI(net275));
 sg13g2_tiehi \i_music.count[25]$_SDFF_PN0__276  (.L_HI(net276));
 sg13g2_tiehi \i_music.count[26]$_SDFF_PN0__277  (.L_HI(net277));
 sg13g2_tiehi \i_music.count[27]$_SDFF_PN0__278  (.L_HI(net278));
 sg13g2_tiehi \i_music.count[28]$_SDFF_PN0__279  (.L_HI(net279));
 sg13g2_tiehi \i_music.count[29]$_SDFF_PN0__280  (.L_HI(net280));
 sg13g2_tiehi \i_music.count[2]$_SDFF_PN0__281  (.L_HI(net281));
 sg13g2_tiehi \i_music.count[30]$_SDFF_PN0__282  (.L_HI(net282));
 sg13g2_tiehi \i_music.count[31]$_SDFF_PN0__283  (.L_HI(net283));
 sg13g2_tiehi \i_music.count[3]$_SDFF_PN0__284  (.L_HI(net284));
 sg13g2_tiehi \i_music.count[4]$_SDFF_PN0__285  (.L_HI(net285));
 sg13g2_tiehi \i_music.count[5]$_SDFF_PN0__286  (.L_HI(net286));
 sg13g2_tiehi \i_music.count[6]$_SDFF_PN0__287  (.L_HI(net287));
 sg13g2_tiehi \i_music.count[7]$_SDFF_PN0__288  (.L_HI(net288));
 sg13g2_tiehi \i_music.count[8]$_SDFF_PN0__289  (.L_HI(net289));
 sg13g2_tiehi \i_music.count[9]$_SDFF_PN0__290  (.L_HI(net290));
 sg13g2_tiehi \i_music.i_pwm.count[0]$_SDFF_PP0__291  (.L_HI(net291));
 sg13g2_tiehi \i_music.i_pwm.count[1]$_SDFF_PP0__292  (.L_HI(net292));
 sg13g2_tiehi \i_music.i_pwm.count[2]$_SDFF_PP0__293  (.L_HI(net293));
 sg13g2_tiehi \i_music.i_pwm.count[3]$_SDFF_PP0__294  (.L_HI(net294));
 sg13g2_tiehi \i_music.i_pwm.count[4]$_SDFF_PP0__295  (.L_HI(net295));
 sg13g2_tiehi \i_music.i_pwm.count[5]$_SDFF_PP0__296  (.L_HI(net296));
 sg13g2_tiehi \i_music.i_pwm.count[6]$_SDFF_PP0__297  (.L_HI(net297));
 sg13g2_tiehi \i_music.i_pwm.count[7]$_SDFF_PP0__298  (.L_HI(net298));
 sg13g2_tiehi \i_music.i_pwm.pwm$_DFFE_PP__299  (.L_HI(net299));
 sg13g2_tiehi \i_music.i_sample.sample[0]$_DFFE_PP__300  (.L_HI(net300));
 sg13g2_tiehi \i_music.i_sample.sample[1]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \i_music.i_sample.sample[2]$_DFFE_PP__302  (.L_HI(net302));
 sg13g2_tiehi \i_music.i_sample.sample[3]$_DFFE_PP__303  (.L_HI(net303));
 sg13g2_tiehi \i_music.i_sample.sample[4]$_DFFE_PP__304  (.L_HI(net304));
 sg13g2_tiehi \i_music.i_sample.sample[5]$_DFFE_PP__305  (.L_HI(net305));
 sg13g2_tiehi \i_music.i_sample.sample[6]$_DFFE_PP__306  (.L_HI(net306));
 sg13g2_tiehi \i_music.i_sample.sample[7]$_DFFE_PP__307  (.L_HI(net307));
 sg13g2_tiehi \i_music.i_sample.sample_acc[0]$_SDFF_PN0__308  (.L_HI(net308));
 sg13g2_tiehi \i_music.i_sample.sample_acc[1]$_SDFF_PN0__309  (.L_HI(net309));
 sg13g2_tiehi \i_music.i_sample.sample_acc[2]$_SDFF_PN0__310  (.L_HI(net310));
 sg13g2_tiehi \i_music.i_sample.sample_acc[3]$_SDFF_PN0__311  (.L_HI(net311));
 sg13g2_tiehi \i_music.i_sample.sample_acc[4]$_SDFF_PN0__312  (.L_HI(net312));
 sg13g2_tiehi \i_music.i_sample.sample_acc[5]$_SDFF_PN0__313  (.L_HI(net313));
 sg13g2_tiehi \i_music.i_sample.sample_acc[6]$_SDFF_PN0__314  (.L_HI(net314));
 sg13g2_tiehi \i_music.i_sample.sample_acc[7]$_SDFF_PN0__315  (.L_HI(net315));
 sg13g2_tiehi \i_music.i_sample.sample_acc[8]$_SDFF_PN0__316  (.L_HI(net316));
 sg13g2_tiehi \i_music.i_sample.sample_idx[0]$_DFF_P__317  (.L_HI(net317));
 sg13g2_tiehi \i_music.i_sample.sample_idx[1]$_DFF_P__318  (.L_HI(net318));
 sg13g2_tiehi \i_music.i_sample.sample_idx[2]$_DFF_P__319  (.L_HI(net319));
 sg13g2_tiehi \i_music.i_sample.sample_idx[3]$_DFF_P__320  (.L_HI(net320));
 sg13g2_tiehi \i_music.i_sample.sample_idx[4]$_DFF_P__321  (.L_HI(net321));
 sg13g2_tiehi \i_music.i_sample.sample_idx[5]$_DFF_P__322  (.L_HI(net322));
 sg13g2_tiehi \i_music.i_sample.sample_idx[6]$_DFF_P__323  (.L_HI(net323));
 sg13g2_tiehi \i_music.i_sample.sample_idx[7]$_DFF_P__324  (.L_HI(net324));
 sg13g2_tiehi \i_music.i_sample.thresh[0]$_DFF_P__325  (.L_HI(net325));
 sg13g2_tiehi \i_music.i_sample.thresh[10]$_DFF_P__326  (.L_HI(net326));
 sg13g2_tiehi \i_music.i_sample.thresh[1]$_DFF_P__327  (.L_HI(net327));
 sg13g2_tiehi \i_music.i_sample.thresh[2]$_DFF_P__328  (.L_HI(net328));
 sg13g2_tiehi \i_music.i_sample.thresh[3]$_DFF_P__329  (.L_HI(net329));
 sg13g2_tiehi \i_music.i_sample.thresh[4]$_DFF_P__330  (.L_HI(net330));
 sg13g2_tiehi \i_music.i_sample.thresh[5]$_DFF_P__331  (.L_HI(net331));
 sg13g2_tiehi \i_music.i_sample.thresh[6]$_DFF_P__332  (.L_HI(net332));
 sg13g2_tiehi \i_music.i_sample.thresh[7]$_DFF_P__333  (.L_HI(net333));
 sg13g2_tiehi \i_music.i_sample.thresh[8]$_DFF_P__334  (.L_HI(net334));
 sg13g2_tiehi \i_music.i_sample.thresh[9]$_DFF_P__335  (.L_HI(net335));
 sg13g2_tiehi \i_music.violin_note_idx[1][0]$_SDFFCE_PP1P__336  (.L_HI(net336));
 sg13g2_tiehi \i_music.violin_note_idx[1][1]$_SDFFCE_PN1P__337  (.L_HI(net337));
 sg13g2_tiehi \i_music.violin_note_idx[1][2]$_SDFFCE_PN1P__338  (.L_HI(net338));
 sg13g2_tiehi \i_music.violin_note_idx[1][3]$_SDFFCE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \i_music.violin_note_idx[1][4]$_DFFE_PP__340  (.L_HI(net340));
 sg13g2_tiehi \i_music.violin_note_idx[1][5]$_DFFE_PP__341  (.L_HI(net341));
 sg13g2_tiehi \i_music.violin_note_idx[1][6]$_DFFE_PP__342  (.L_HI(net342));
 sg13g2_tiehi \i_music.violin_note_idx[1][7]$_DFFE_PP__343  (.L_HI(net343));
 sg13g2_tiehi \i_music.violin_note_idx[1][8]$_DFFE_PP__344  (.L_HI(net344));
 sg13g2_tiehi \i_music.violin_note_idx[2][0]$_SDFFCE_PP1P__345  (.L_HI(net345));
 sg13g2_tiehi \i_music.violin_note_idx[2][1]$_SDFFCE_PN1P__346  (.L_HI(net346));
 sg13g2_tiehi \i_music.violin_note_idx[2][2]$_SDFFCE_PN1P__347  (.L_HI(net347));
 sg13g2_tiehi \i_music.violin_note_idx[2][3]$_SDFFCE_PN1P__348  (.L_HI(net348));
 sg13g2_tiehi \i_music.violin_note_idx[2][4]$_DFFE_PP__349  (.L_HI(net349));
 sg13g2_tiehi \i_music.violin_note_idx[2][5]$_DFFE_PP__350  (.L_HI(net350));
 sg13g2_tiehi \i_music.violin_note_idx[2][6]$_DFFE_PP__351  (.L_HI(net351));
 sg13g2_tiehi \i_music.violin_note_idx[2][7]$_DFFE_PP__352  (.L_HI(net352));
 sg13g2_tiehi \i_music.violin_note_idx[2][8]$_DFFE_PP__353  (.L_HI(net353));
 sg13g2_tiehi \i_music.violin_note_idx[3][0]$_SDFFCE_PP1P__354  (.L_HI(net354));
 sg13g2_tiehi \i_music.violin_note_idx[3][1]$_SDFFCE_PN1P__355  (.L_HI(net355));
 sg13g2_tiehi \i_music.violin_note_idx[3][2]$_SDFFCE_PN1P__356  (.L_HI(net356));
 sg13g2_tiehi \i_music.violin_note_idx[3][3]$_SDFFCE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \i_music.violin_note_idx[3][4]$_DFFE_PP__358  (.L_HI(net358));
 sg13g2_tiehi \i_music.violin_note_idx[3][5]$_DFFE_PP__359  (.L_HI(net359));
 sg13g2_tiehi \i_music.violin_note_idx[3][6]$_DFFE_PP__360  (.L_HI(net360));
 sg13g2_tiehi \i_music.violin_note_idx[3][7]$_DFFE_PP__361  (.L_HI(net361));
 sg13g2_tiehi \i_music.violin_note_idx[3][8]$_DFFE_PP__362  (.L_HI(net362));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_2 clkbuf_level_0_1_10_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_level_0_1_10_clk));
 sg13g2_buf_2 clkbuf_level_1_1_11_clk (.A(clknet_level_0_1_10_clk),
    .X(clknet_level_1_1_11_clk));
 sg13g2_buf_2 clkbuf_level_2_1_12_clk (.A(clknet_level_1_1_11_clk),
    .X(clknet_level_2_1_12_clk));
 sg13g2_buf_2 clkbuf_level_0_1_23_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_level_0_1_23_clk));
 sg13g2_buf_2 clkbuf_level_1_1_24_clk (.A(clknet_level_0_1_23_clk),
    .X(clknet_level_1_1_24_clk));
 sg13g2_buf_2 clkbuf_level_2_1_25_clk (.A(clknet_level_1_1_24_clk),
    .X(clknet_level_2_1_25_clk));
 sg13g2_buf_2 clkbuf_level_0_1_36_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_level_0_1_36_clk));
 sg13g2_buf_2 clkbuf_level_1_1_37_clk (.A(clknet_level_0_1_36_clk),
    .X(clknet_level_1_1_37_clk));
 sg13g2_buf_2 clkbuf_level_2_1_38_clk (.A(clknet_level_1_1_37_clk),
    .X(clknet_level_2_1_38_clk));
 sg13g2_buf_2 clkbuf_level_0_1_49_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_level_0_1_49_clk));
 sg13g2_buf_2 clkbuf_level_1_1_410_clk (.A(clknet_level_0_1_49_clk),
    .X(clknet_level_1_1_410_clk));
 sg13g2_buf_2 clkbuf_level_2_1_411_clk (.A(clknet_level_1_1_410_clk),
    .X(clknet_level_2_1_411_clk));
 sg13g2_buf_2 clkbuf_level_0_1_512_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_level_0_1_512_clk));
 sg13g2_buf_2 clkbuf_level_1_1_513_clk (.A(clknet_level_0_1_512_clk),
    .X(clknet_level_1_1_513_clk));
 sg13g2_buf_2 clkbuf_level_2_1_514_clk (.A(clknet_level_1_1_513_clk),
    .X(clknet_level_2_1_514_clk));
 sg13g2_buf_2 clkbuf_level_0_1_615_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_level_0_1_615_clk));
 sg13g2_buf_2 clkbuf_level_1_1_616_clk (.A(clknet_level_0_1_615_clk),
    .X(clknet_level_1_1_616_clk));
 sg13g2_buf_2 clkbuf_level_2_1_617_clk (.A(clknet_level_1_1_616_clk),
    .X(clknet_level_2_1_617_clk));
 sg13g2_buf_2 clkbuf_level_0_1_718_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_level_0_1_718_clk));
 sg13g2_buf_2 clkbuf_level_1_1_719_clk (.A(clknet_level_0_1_718_clk),
    .X(clknet_level_1_1_719_clk));
 sg13g2_buf_2 clkbuf_level_2_1_720_clk (.A(clknet_level_1_1_719_clk),
    .X(clknet_level_2_1_720_clk));
 sg13g2_buf_2 clkbuf_level_0_1_821_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_level_0_1_821_clk));
 sg13g2_buf_2 clkbuf_level_1_1_822_clk (.A(clknet_level_0_1_821_clk),
    .X(clknet_level_1_1_822_clk));
 sg13g2_buf_2 clkbuf_level_2_1_823_clk (.A(clknet_level_1_1_822_clk),
    .X(clknet_level_2_1_823_clk));
 sg13g2_buf_2 clkbuf_level_0_1_924_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_level_0_1_924_clk));
 sg13g2_buf_2 clkbuf_level_1_1_925_clk (.A(clknet_level_0_1_924_clk),
    .X(clknet_level_1_1_925_clk));
 sg13g2_buf_2 clkbuf_level_2_1_926_clk (.A(clknet_level_1_1_925_clk),
    .X(clknet_level_2_1_926_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1027_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_level_0_1_1027_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1028_clk (.A(clknet_level_0_1_1027_clk),
    .X(clknet_level_1_1_1028_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1029_clk (.A(clknet_level_1_1_1028_clk),
    .X(clknet_level_2_1_1029_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1130_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_level_0_1_1130_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1131_clk (.A(clknet_level_0_1_1130_clk),
    .X(clknet_level_1_1_1131_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1132_clk (.A(clknet_level_1_1_1131_clk),
    .X(clknet_level_2_1_1132_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1233_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_level_0_1_1233_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1234_clk (.A(clknet_level_0_1_1233_clk),
    .X(clknet_level_1_1_1234_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1235_clk (.A(clknet_level_1_1_1234_clk),
    .X(clknet_level_2_1_1235_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1336_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_level_0_1_1336_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1337_clk (.A(clknet_level_0_1_1336_clk),
    .X(clknet_level_1_1_1337_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1338_clk (.A(clknet_level_1_1_1337_clk),
    .X(clknet_level_2_1_1338_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1439_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_level_0_1_1439_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1440_clk (.A(clknet_level_0_1_1439_clk),
    .X(clknet_level_1_1_1440_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1441_clk (.A(clknet_level_1_1_1440_clk),
    .X(clknet_level_2_1_1441_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1542_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_level_0_1_1542_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1543_clk (.A(clknet_level_0_1_1542_clk),
    .X(clknet_level_1_1_1543_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1544_clk (.A(clknet_level_1_1_1543_clk),
    .X(clknet_level_2_1_1544_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1645_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_level_0_1_1645_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1646_clk (.A(clknet_level_0_1_1645_clk),
    .X(clknet_level_1_1_1646_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1647_clk (.A(clknet_level_1_1_1646_clk),
    .X(clknet_level_2_1_1647_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1748_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_level_0_1_1748_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1749_clk (.A(clknet_level_0_1_1748_clk),
    .X(clknet_level_1_1_1749_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1750_clk (.A(clknet_level_1_1_1749_clk),
    .X(clknet_level_2_1_1750_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1851_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_level_0_1_1851_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1852_clk (.A(clknet_level_0_1_1851_clk),
    .X(clknet_level_1_1_1852_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1853_clk (.A(clknet_level_1_1_1852_clk),
    .X(clknet_level_2_1_1853_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1954_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_level_0_1_1954_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1955_clk (.A(clknet_level_0_1_1954_clk),
    .X(clknet_level_1_1_1955_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1956_clk (.A(clknet_level_1_1_1955_clk),
    .X(clknet_level_2_1_1956_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2057_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_level_0_1_2057_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2058_clk (.A(clknet_level_0_1_2057_clk),
    .X(clknet_level_1_1_2058_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2059_clk (.A(clknet_level_1_1_2058_clk),
    .X(clknet_level_2_1_2059_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2160_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_level_0_1_2160_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2161_clk (.A(clknet_level_0_1_2160_clk),
    .X(clknet_level_1_1_2161_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2162_clk (.A(clknet_level_1_1_2161_clk),
    .X(clknet_level_2_1_2162_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2263_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_level_0_1_2263_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2264_clk (.A(clknet_level_0_1_2263_clk),
    .X(clknet_level_1_1_2264_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2265_clk (.A(clknet_level_1_1_2264_clk),
    .X(clknet_level_2_1_2265_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2366_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_level_0_1_2366_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2367_clk (.A(clknet_level_0_1_2366_clk),
    .X(clknet_level_1_1_2367_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2368_clk (.A(clknet_level_1_1_2367_clk),
    .X(clknet_level_2_1_2368_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2469_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_level_0_1_2469_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2470_clk (.A(clknet_level_0_1_2469_clk),
    .X(clknet_level_1_1_2470_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2471_clk (.A(clknet_level_1_1_2470_clk),
    .X(clknet_level_2_1_2471_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2572_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_level_0_1_2572_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2573_clk (.A(clknet_level_0_1_2572_clk),
    .X(clknet_level_1_1_2573_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2574_clk (.A(clknet_level_1_1_2573_clk),
    .X(clknet_level_2_1_2574_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2675_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_level_0_1_2675_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2676_clk (.A(clknet_level_0_1_2675_clk),
    .X(clknet_level_1_1_2676_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2677_clk (.A(clknet_level_1_1_2676_clk),
    .X(clknet_level_2_1_2677_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2778_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_level_0_1_2778_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2779_clk (.A(clknet_level_0_1_2778_clk),
    .X(clknet_level_1_1_2779_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2780_clk (.A(clknet_level_1_1_2779_clk),
    .X(clknet_level_2_1_2780_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2881_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_level_0_1_2881_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2882_clk (.A(clknet_level_0_1_2881_clk),
    .X(clknet_level_1_1_2882_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2883_clk (.A(clknet_level_1_1_2882_clk),
    .X(clknet_level_2_1_2883_clk));
 sg13g2_buf_2 clkbuf_level_0_1_2984_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_level_0_1_2984_clk));
 sg13g2_buf_2 clkbuf_level_1_1_2985_clk (.A(clknet_level_0_1_2984_clk),
    .X(clknet_level_1_1_2985_clk));
 sg13g2_buf_2 clkbuf_level_2_1_2986_clk (.A(clknet_level_1_1_2985_clk),
    .X(clknet_level_2_1_2986_clk));
 sg13g2_buf_2 clkbuf_level_0_1_3087_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_level_0_1_3087_clk));
 sg13g2_buf_2 clkbuf_level_1_1_3088_clk (.A(clknet_level_0_1_3087_clk),
    .X(clknet_level_1_1_3088_clk));
 sg13g2_buf_2 clkbuf_level_2_1_3089_clk (.A(clknet_level_1_1_3088_clk),
    .X(clknet_level_2_1_3089_clk));
 sg13g2_buf_2 clkbuf_level_0_1_3190_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_level_0_1_3190_clk));
 sg13g2_buf_2 clkbuf_level_1_1_3191_clk (.A(clknet_level_0_1_3190_clk),
    .X(clknet_level_1_1_3191_clk));
 sg13g2_buf_2 clkbuf_level_2_1_3192_clk (.A(clknet_level_1_1_3191_clk),
    .X(clknet_level_2_1_3192_clk));
 sg13g2_buf_2 clkbuf_level_0_1_3293_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_level_0_1_3293_clk));
 sg13g2_buf_2 clkbuf_level_1_1_3294_clk (.A(clknet_level_0_1_3293_clk),
    .X(clknet_level_1_1_3294_clk));
 sg13g2_buf_2 clkbuf_level_2_1_3295_clk (.A(clknet_level_1_1_3294_clk),
    .X(clknet_level_2_1_3295_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_1 \clkbuf_0_i_music.i_sample.t1.CG.GCLK  (.A(\i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_0__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_1__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_2__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_3__f_i_music.i_sample.t1.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t1.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_2 clkload2 (.A(\clknet_2_3__leaf_i_music.i_sample.t1.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_0_i_music.i_sample.t2.CG.GCLK  (.A(\i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_0__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_1__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_2__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_3__f_i_music.i_sample.t2.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t2.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 clkload3 (.A(\clknet_2_1__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_2 clkload4 (.A(\clknet_2_3__leaf_i_music.i_sample.t2.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_0_i_music.i_sample.t3.CG.GCLK  (.A(\i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_0__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_1__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_2__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_3__f_i_music.i_sample.t3.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t3.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 clkload5 (.A(\clknet_2_1__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_2 clkload6 (.A(\clknet_2_3__leaf_i_music.i_sample.t3.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_0_i_music.i_sample.t4.CG.GCLK  (.A(\i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_0_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_0__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_0__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_1__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_2__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_2__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_1 \clkbuf_2_3__f_i_music.i_sample.t4.CG.GCLK  (.A(\clknet_0_i_music.i_sample.t4.CG.GCLK ),
    .X(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 clkload7 (.A(\clknet_2_1__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_buf_2 clkload8 (.A(\clknet_2_3__leaf_i_music.i_sample.t4.CG.GCLK ));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_34 ();
 sg13g2_fill_1 FILLER_0_71 ();
 sg13g2_decap_8 FILLER_0_92 ();
 sg13g2_decap_8 FILLER_0_99 ();
 sg13g2_fill_2 FILLER_0_106 ();
 sg13g2_fill_1 FILLER_0_108 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_decap_4 FILLER_0_253 ();
 sg13g2_fill_1 FILLER_0_257 ();
 sg13g2_fill_1 FILLER_0_268 ();
 sg13g2_fill_2 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_274 ();
 sg13g2_fill_1 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_4 FILLER_0_301 ();
 sg13g2_fill_1 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_fill_2 FILLER_0_327 ();
 sg13g2_fill_1 FILLER_0_329 ();
 sg13g2_decap_4 FILLER_0_335 ();
 sg13g2_fill_2 FILLER_0_342 ();
 sg13g2_fill_1 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_fill_2 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_fill_2 FILLER_0_385 ();
 sg13g2_fill_1 FILLER_0_387 ();
 sg13g2_fill_1 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_16 ();
 sg13g2_fill_2 FILLER_1_96 ();
 sg13g2_fill_1 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_4 FILLER_1_198 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_decap_4 FILLER_1_229 ();
 sg13g2_fill_1 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_257 ();
 sg13g2_fill_1 FILLER_1_264 ();
 sg13g2_fill_2 FILLER_1_270 ();
 sg13g2_fill_1 FILLER_1_335 ();
 sg13g2_fill_2 FILLER_1_351 ();
 sg13g2_fill_1 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_16 ();
 sg13g2_fill_1 FILLER_2_47 ();
 sg13g2_decap_4 FILLER_2_100 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_134 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_fill_2 FILLER_2_148 ();
 sg13g2_fill_1 FILLER_2_150 ();
 sg13g2_fill_2 FILLER_2_164 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_186 ();
 sg13g2_fill_2 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_223 ();
 sg13g2_fill_1 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_4 FILLER_2_249 ();
 sg13g2_decap_4 FILLER_2_270 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_332 ();
 sg13g2_decap_4 FILLER_2_338 ();
 sg13g2_fill_2 FILLER_2_342 ();
 sg13g2_decap_4 FILLER_2_352 ();
 sg13g2_fill_2 FILLER_2_356 ();
 sg13g2_decap_4 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_4 FILLER_2_389 ();
 sg13g2_fill_2 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_36 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_82 ();
 sg13g2_fill_2 FILLER_3_101 ();
 sg13g2_fill_1 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_4 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_222 ();
 sg13g2_fill_1 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_261 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_270 ();
 sg13g2_fill_2 FILLER_3_298 ();
 sg13g2_fill_1 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_348 ();
 sg13g2_decap_4 FILLER_3_386 ();
 sg13g2_fill_2 FILLER_3_397 ();
 sg13g2_fill_1 FILLER_3_399 ();
 sg13g2_fill_1 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_11 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_fill_1 FILLER_4_22 ();
 sg13g2_fill_1 FILLER_4_32 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_fill_1 FILLER_4_100 ();
 sg13g2_fill_2 FILLER_4_145 ();
 sg13g2_fill_1 FILLER_4_161 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_180 ();
 sg13g2_fill_1 FILLER_4_186 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_fill_2 FILLER_4_321 ();
 sg13g2_fill_1 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_332 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_364 ();
 sg13g2_fill_1 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_405 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_15 ();
 sg13g2_fill_1 FILLER_5_38 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_1 FILLER_5_147 ();
 sg13g2_fill_1 FILLER_5_162 ();
 sg13g2_fill_2 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_fill_2 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_4 FILLER_5_242 ();
 sg13g2_decap_4 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_310 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_decap_4 FILLER_5_339 ();
 sg13g2_fill_2 FILLER_5_343 ();
 sg13g2_fill_1 FILLER_5_357 ();
 sg13g2_fill_1 FILLER_5_386 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_fill_2 FILLER_6_15 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_1 FILLER_6_51 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_fill_1 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_136 ();
 sg13g2_decap_4 FILLER_6_186 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_fill_1 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_fill_2 FILLER_6_258 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_fill_2 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_327 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_fill_2 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_fill_1 FILLER_6_352 ();
 sg13g2_decap_4 FILLER_6_356 ();
 sg13g2_decap_4 FILLER_6_374 ();
 sg13g2_fill_1 FILLER_6_378 ();
 sg13g2_fill_1 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_388 ();
 sg13g2_fill_1 FILLER_6_395 ();
 sg13g2_fill_2 FILLER_6_400 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_7_8 ();
 sg13g2_fill_2 FILLER_7_12 ();
 sg13g2_decap_4 FILLER_7_24 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_decap_4 FILLER_7_96 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_decap_4 FILLER_7_197 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_207 ();
 sg13g2_fill_1 FILLER_7_220 ();
 sg13g2_decap_4 FILLER_7_259 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_298 ();
 sg13g2_fill_2 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_333 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_4 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_fill_2 FILLER_7_381 ();
 sg13g2_fill_1 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_409 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_1 FILLER_8_19 ();
 sg13g2_fill_2 FILLER_8_24 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_fill_1 FILLER_8_37 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_62 ();
 sg13g2_decap_4 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_fill_1 FILLER_8_106 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_2 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_224 ();
 sg13g2_decap_4 FILLER_8_237 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_decap_8 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_304 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_fill_2 FILLER_8_324 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_decap_4 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_8_383 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_16 ();
 sg13g2_fill_2 FILLER_9_33 ();
 sg13g2_fill_1 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_decap_4 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_fill_2 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_decap_4 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_312 ();
 sg13g2_fill_2 FILLER_9_326 ();
 sg13g2_decap_4 FILLER_9_332 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_fill_1 FILLER_9_354 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_2 FILLER_9_395 ();
 sg13g2_fill_1 FILLER_9_397 ();
 sg13g2_fill_1 FILLER_9_402 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_1 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_fill_1 FILLER_10_43 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_decap_4 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_2 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_decap_4 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_decap_4 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_fill_2 FILLER_10_382 ();
 sg13g2_fill_1 FILLER_10_384 ();
 sg13g2_fill_2 FILLER_10_389 ();
 sg13g2_fill_1 FILLER_10_391 ();
 sg13g2_fill_2 FILLER_10_399 ();
 sg13g2_fill_1 FILLER_10_401 ();
 sg13g2_fill_2 FILLER_10_414 ();
 sg13g2_fill_1 FILLER_10_416 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_4 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_8 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_4 FILLER_11_134 ();
 sg13g2_fill_1 FILLER_11_138 ();
 sg13g2_fill_1 FILLER_11_144 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_185 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_202 ();
 sg13g2_fill_1 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_4 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_decap_4 FILLER_11_359 ();
 sg13g2_fill_2 FILLER_11_377 ();
 sg13g2_fill_1 FILLER_11_379 ();
 sg13g2_decap_4 FILLER_11_384 ();
 sg13g2_fill_2 FILLER_11_388 ();
 sg13g2_fill_1 FILLER_11_394 ();
 sg13g2_fill_2 FILLER_11_410 ();
 sg13g2_fill_1 FILLER_11_412 ();
 sg13g2_decap_4 FILLER_11_425 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_27 ();
 sg13g2_fill_1 FILLER_12_37 ();
 sg13g2_fill_2 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_151 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_2 FILLER_12_371 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_12_410 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_13 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_decap_4 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_240 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_316 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_1 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_371 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_decap_4 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_12 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_fill_2 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_50 ();
 sg13g2_fill_1 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_decap_4 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_379 ();
 sg13g2_fill_1 FILLER_14_394 ();
 sg13g2_fill_2 FILLER_14_399 ();
 sg13g2_fill_1 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_414 ();
 sg13g2_fill_1 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_fill_1 FILLER_15_15 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_287 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_352 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_376 ();
 sg13g2_fill_1 FILLER_15_386 ();
 sg13g2_fill_1 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_18 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_59 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_103 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_fill_2 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_decap_4 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_356 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_1 FILLER_17_22 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_decap_4 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_decap_4 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_4 FILLER_17_397 ();
 sg13g2_fill_2 FILLER_17_413 ();
 sg13g2_fill_2 FILLER_17_423 ();
 sg13g2_fill_1 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_17 ();
 sg13g2_fill_2 FILLER_18_47 ();
 sg13g2_fill_1 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_fill_1 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_decap_4 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_367 ();
 sg13g2_decap_4 FILLER_18_378 ();
 sg13g2_fill_2 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_18_388 ();
 sg13g2_fill_1 FILLER_18_390 ();
 sg13g2_fill_2 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_406 ();
 sg13g2_decap_4 FILLER_18_411 ();
 sg13g2_fill_1 FILLER_18_415 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_13 ();
 sg13g2_fill_2 FILLER_19_19 ();
 sg13g2_fill_2 FILLER_19_44 ();
 sg13g2_fill_1 FILLER_19_51 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_decap_4 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_103 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_114 ();
 sg13g2_decap_4 FILLER_19_124 ();
 sg13g2_decap_4 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_decap_4 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_decap_4 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_fill_1 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_415 ();
 sg13g2_fill_1 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_fill_2 FILLER_20_33 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_106 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_fill_2 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_decap_4 FILLER_20_391 ();
 sg13g2_fill_2 FILLER_20_395 ();
 sg13g2_decap_4 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_417 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_8 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_fill_1 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_285 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_363 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_decap_4 FILLER_22_360 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_1 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_22_412 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_15 ();
 sg13g2_fill_1 FILLER_23_25 ();
 sg13g2_fill_2 FILLER_23_50 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_4 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_418 ();
 sg13g2_fill_1 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_fill_2 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_decap_4 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_373 ();
 sg13g2_decap_4 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_414 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_fill_2 FILLER_25_409 ();
 sg13g2_decap_4 FILLER_25_415 ();
 sg13g2_fill_1 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_25_424 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_decap_4 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_decap_4 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_424 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_decap_4 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_fill_2 FILLER_27_398 ();
 sg13g2_fill_1 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_6 ();
 sg13g2_fill_1 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_decap_4 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_28_413 ();
 sg13g2_fill_1 FILLER_28_415 ();
 sg13g2_fill_1 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_decap_4 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_29_415 ();
 sg13g2_fill_1 FILLER_29_423 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_402 ();
 sg13g2_fill_1 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_414 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_2 FILLER_31_403 ();
 sg13g2_decap_4 FILLER_31_411 ();
 sg13g2_fill_2 FILLER_31_415 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_5 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_decap_4 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_370 ();
 sg13g2_fill_1 FILLER_32_372 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_10 ();
 sg13g2_fill_1 FILLER_33_12 ();
 sg13g2_fill_2 FILLER_33_33 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_fill_2 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_decap_4 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_decap_4 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_1 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_decap_4 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_decap_4 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_decap_4 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_decap_4 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_decap_4 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_4 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_decap_4 FILLER_35_393 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_417 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_2 FILLER_36_48 ();
 sg13g2_decap_8 FILLER_36_62 ();
 sg13g2_decap_4 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_decap_4 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_417 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_2 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_decap_4 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_2 FILLER_37_394 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_fill_1 FILLER_37_420 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_38_31 ();
 sg13g2_decap_8 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_86 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_decap_4 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_fill_1 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_422 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_15 ();
 sg13g2_fill_2 FILLER_39_19 ();
 sg13g2_fill_1 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_41 ();
 sg13g2_fill_1 FILLER_39_87 ();
 sg13g2_fill_2 FILLER_39_116 ();
 sg13g2_fill_1 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_215 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_248 ();
 sg13g2_fill_2 FILLER_39_262 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_279 ();
 sg13g2_decap_4 FILLER_39_286 ();
 sg13g2_fill_1 FILLER_39_290 ();
 sg13g2_fill_2 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_333 ();
 sg13g2_fill_1 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_342 ();
 sg13g2_decap_4 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_353 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_39_422 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_fill_1 FILLER_40_50 ();
 sg13g2_fill_2 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_76 ();
 sg13g2_fill_2 FILLER_40_99 ();
 sg13g2_fill_2 FILLER_40_148 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_fill_2 FILLER_40_166 ();
 sg13g2_fill_1 FILLER_40_176 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_281 ();
 sg13g2_fill_1 FILLER_40_293 ();
 sg13g2_fill_1 FILLER_40_298 ();
 sg13g2_fill_2 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_334 ();
 sg13g2_fill_1 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_fill_2 FILLER_40_428 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_15 ();
 sg13g2_fill_2 FILLER_41_22 ();
 sg13g2_fill_2 FILLER_41_92 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_fill_2 FILLER_41_112 ();
 sg13g2_fill_1 FILLER_41_114 ();
 sg13g2_fill_2 FILLER_41_120 ();
 sg13g2_fill_2 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_143 ();
 sg13g2_fill_2 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_206 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_decap_4 FILLER_41_244 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_323 ();
 sg13g2_fill_1 FILLER_41_328 ();
 sg13g2_fill_1 FILLER_41_333 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_decap_4 FILLER_41_386 ();
 sg13g2_fill_1 FILLER_41_390 ();
 sg13g2_fill_1 FILLER_41_400 ();
 sg13g2_fill_1 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_42_26 ();
 sg13g2_decap_4 FILLER_42_33 ();
 sg13g2_decap_4 FILLER_42_72 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_1 FILLER_42_99 ();
 sg13g2_fill_2 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_180 ();
 sg13g2_fill_1 FILLER_42_193 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_2 FILLER_42_238 ();
 sg13g2_fill_2 FILLER_42_244 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_fill_2 FILLER_42_252 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_fill_2 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_decap_4 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_322 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_decap_4 FILLER_42_353 ();
 sg13g2_fill_1 FILLER_42_357 ();
 sg13g2_fill_2 FILLER_42_362 ();
 sg13g2_decap_4 FILLER_42_394 ();
 sg13g2_fill_1 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_422 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_15 ();
 sg13g2_decap_4 FILLER_43_27 ();
 sg13g2_fill_2 FILLER_43_31 ();
 sg13g2_fill_2 FILLER_43_45 ();
 sg13g2_fill_1 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_52 ();
 sg13g2_fill_1 FILLER_43_54 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_70 ();
 sg13g2_decap_4 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_fill_2 FILLER_43_103 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_157 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_205 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_245 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_275 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_fill_2 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_338 ();
 sg13g2_decap_4 FILLER_43_351 ();
 sg13g2_decap_8 FILLER_43_384 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_5 ();
 sg13g2_fill_2 FILLER_44_16 ();
 sg13g2_fill_2 FILLER_44_22 ();
 sg13g2_fill_2 FILLER_44_29 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_175 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_215 ();
 sg13g2_fill_2 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_234 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_fill_1 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_288 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_decap_8 FILLER_44_337 ();
 sg13g2_decap_4 FILLER_44_344 ();
 sg13g2_decap_4 FILLER_44_353 ();
 sg13g2_fill_2 FILLER_44_362 ();
 sg13g2_decap_4 FILLER_44_372 ();
 sg13g2_fill_2 FILLER_44_384 ();
 sg13g2_fill_2 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_2 FILLER_44_397 ();
 sg13g2_fill_1 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_fill_2 FILLER_45_113 ();
 sg13g2_fill_2 FILLER_45_146 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_fill_1 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_254 ();
 sg13g2_decap_4 FILLER_45_364 ();
 sg13g2_fill_2 FILLER_45_368 ();
 sg13g2_fill_2 FILLER_45_374 ();
 sg13g2_fill_1 FILLER_45_376 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_fill_1 FILLER_46_9 ();
 sg13g2_fill_2 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_fill_2 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_134 ();
 sg13g2_fill_1 FILLER_46_139 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_fill_1 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_238 ();
 sg13g2_decap_4 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_259 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_2 FILLER_46_297 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_fill_2 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_343 ();
 sg13g2_fill_2 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_387 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_414 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_1 FILLER_47_29 ();
 sg13g2_fill_1 FILLER_47_47 ();
 sg13g2_decap_8 FILLER_47_66 ();
 sg13g2_decap_4 FILLER_47_73 ();
 sg13g2_fill_1 FILLER_47_77 ();
 sg13g2_decap_4 FILLER_47_149 ();
 sg13g2_fill_2 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_170 ();
 sg13g2_fill_1 FILLER_47_225 ();
 sg13g2_fill_1 FILLER_47_230 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_decap_4 FILLER_47_248 ();
 sg13g2_decap_4 FILLER_47_256 ();
 sg13g2_fill_2 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_332 ();
 sg13g2_decap_4 FILLER_47_337 ();
 sg13g2_fill_1 FILLER_47_341 ();
 sg13g2_decap_4 FILLER_47_354 ();
 sg13g2_fill_2 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_369 ();
 sg13g2_fill_2 FILLER_47_404 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_fill_1 FILLER_47_421 ();
 sg13g2_fill_2 FILLER_48_16 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_4 FILLER_48_66 ();
 sg13g2_fill_2 FILLER_48_70 ();
 sg13g2_decap_4 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_99 ();
 sg13g2_fill_1 FILLER_48_118 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_159 ();
 sg13g2_fill_2 FILLER_48_165 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_fill_2 FILLER_48_279 ();
 sg13g2_fill_2 FILLER_48_310 ();
 sg13g2_fill_1 FILLER_48_312 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_decap_4 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_fill_1 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_412 ();
 sg13g2_fill_1 FILLER_48_414 ();
 sg13g2_decap_4 FILLER_48_419 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_fill_2 FILLER_49_31 ();
 sg13g2_fill_2 FILLER_49_60 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_fill_1 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_fill_1 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_fill_2 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_167 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_1 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_186 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_fill_2 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_208 ();
 sg13g2_fill_2 FILLER_49_218 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_fill_2 FILLER_49_232 ();
 sg13g2_decap_4 FILLER_49_239 ();
 sg13g2_decap_4 FILLER_49_247 ();
 sg13g2_fill_2 FILLER_49_251 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_fill_1 FILLER_49_334 ();
 sg13g2_fill_2 FILLER_49_427 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_12 ();
 sg13g2_fill_2 FILLER_50_38 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_1 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_59 ();
 sg13g2_fill_1 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_142 ();
 sg13g2_fill_1 FILLER_50_144 ();
 sg13g2_fill_2 FILLER_50_162 ();
 sg13g2_fill_1 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_183 ();
 sg13g2_fill_1 FILLER_50_189 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_fill_2 FILLER_50_235 ();
 sg13g2_fill_2 FILLER_50_263 ();
 sg13g2_decap_4 FILLER_50_274 ();
 sg13g2_fill_1 FILLER_50_311 ();
 sg13g2_fill_2 FILLER_50_321 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_2 FILLER_50_331 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_1 FILLER_50_387 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_424 ();
 sg13g2_fill_1 FILLER_51_5 ();
 sg13g2_fill_1 FILLER_51_19 ();
 sg13g2_fill_1 FILLER_51_25 ();
 sg13g2_fill_1 FILLER_51_39 ();
 sg13g2_fill_1 FILLER_51_48 ();
 sg13g2_fill_1 FILLER_51_54 ();
 sg13g2_decap_4 FILLER_51_75 ();
 sg13g2_fill_2 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_fill_2 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_fill_1 FILLER_51_125 ();
 sg13g2_fill_1 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_174 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_fill_1 FILLER_51_187 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_fill_1 FILLER_51_199 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_decap_4 FILLER_51_214 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_226 ();
 sg13g2_fill_1 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_233 ();
 sg13g2_fill_2 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_245 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_290 ();
 sg13g2_decap_4 FILLER_51_295 ();
 sg13g2_fill_2 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_357 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_fill_2 FILLER_51_373 ();
 sg13g2_decap_8 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_387 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_fill_2 FILLER_52_12 ();
 sg13g2_fill_1 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_55 ();
 sg13g2_decap_8 FILLER_52_67 ();
 sg13g2_fill_1 FILLER_52_74 ();
 sg13g2_decap_4 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_fill_2 FILLER_52_88 ();
 sg13g2_fill_2 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_163 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_fill_1 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_2 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_decap_4 FILLER_52_386 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_425 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_81 ();
 sg13g2_fill_1 FILLER_53_83 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_fill_1 FILLER_53_245 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_fill_1 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_fill_1 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_317 ();
 sg13g2_fill_2 FILLER_53_339 ();
 sg13g2_fill_1 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_fill_1 FILLER_53_412 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_1 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_45 ();
 sg13g2_fill_1 FILLER_54_60 ();
 sg13g2_fill_2 FILLER_54_66 ();
 sg13g2_decap_4 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_80 ();
 sg13g2_decap_4 FILLER_54_87 ();
 sg13g2_decap_4 FILLER_54_95 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_104 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_1 FILLER_54_134 ();
 sg13g2_fill_1 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_164 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_241 ();
 sg13g2_fill_1 FILLER_54_265 ();
 sg13g2_fill_1 FILLER_54_270 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_283 ();
 sg13g2_fill_1 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_fill_1 FILLER_54_349 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_fill_1 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_389 ();
 sg13g2_fill_1 FILLER_54_391 ();
 sg13g2_fill_1 FILLER_54_407 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_fill_2 FILLER_54_427 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_58 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_117 ();
 sg13g2_fill_1 FILLER_55_119 ();
 sg13g2_fill_1 FILLER_55_125 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_153 ();
 sg13g2_fill_1 FILLER_55_167 ();
 sg13g2_fill_1 FILLER_55_172 ();
 sg13g2_fill_1 FILLER_55_199 ();
 sg13g2_fill_1 FILLER_55_226 ();
 sg13g2_fill_2 FILLER_55_253 ();
 sg13g2_fill_1 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_276 ();
 sg13g2_decap_4 FILLER_55_300 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_decap_4 FILLER_55_327 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_341 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_decap_8 FILLER_55_384 ();
 sg13g2_fill_1 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_419 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_2 FILLER_56_61 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_72 ();
 sg13g2_decap_4 FILLER_56_87 ();
 sg13g2_decap_4 FILLER_56_109 ();
 sg13g2_fill_1 FILLER_56_142 ();
 sg13g2_fill_1 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_156 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_fill_2 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_2 FILLER_56_215 ();
 sg13g2_fill_2 FILLER_56_230 ();
 sg13g2_fill_2 FILLER_56_236 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_fill_2 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_275 ();
 sg13g2_decap_4 FILLER_56_284 ();
 sg13g2_fill_2 FILLER_56_303 ();
 sg13g2_fill_2 FILLER_56_325 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_395 ();
 sg13g2_decap_4 FILLER_56_400 ();
 sg13g2_fill_1 FILLER_56_404 ();
 sg13g2_fill_2 FILLER_56_421 ();
 sg13g2_fill_2 FILLER_56_427 ();
 sg13g2_fill_1 FILLER_56_429 ();
 sg13g2_fill_1 FILLER_57_10 ();
 sg13g2_fill_1 FILLER_57_31 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_63 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_decap_8 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_fill_2 FILLER_57_117 ();
 sg13g2_fill_1 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_149 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_decap_4 FILLER_57_187 ();
 sg13g2_fill_2 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_324 ();
 sg13g2_fill_1 FILLER_57_329 ();
 sg13g2_decap_4 FILLER_57_338 ();
 sg13g2_fill_2 FILLER_57_342 ();
 sg13g2_decap_4 FILLER_57_356 ();
 sg13g2_fill_1 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_fill_2 FILLER_57_386 ();
 sg13g2_fill_2 FILLER_57_393 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_58_41 ();
 sg13g2_fill_1 FILLER_58_60 ();
 sg13g2_fill_2 FILLER_58_65 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_fill_1 FILLER_58_79 ();
 sg13g2_fill_1 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_90 ();
 sg13g2_fill_2 FILLER_58_96 ();
 sg13g2_fill_2 FILLER_58_103 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_fill_2 FILLER_58_113 ();
 sg13g2_decap_4 FILLER_58_144 ();
 sg13g2_fill_2 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_158 ();
 sg13g2_fill_1 FILLER_58_172 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_fill_2 FILLER_58_210 ();
 sg13g2_decap_4 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_1 FILLER_58_268 ();
 sg13g2_fill_1 FILLER_58_275 ();
 sg13g2_fill_2 FILLER_58_286 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_349 ();
 sg13g2_fill_2 FILLER_58_355 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_decap_8 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_386 ();
 sg13g2_fill_1 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_409 ();
 sg13g2_fill_1 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_5 ();
 sg13g2_fill_2 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_29 ();
 sg13g2_fill_2 FILLER_59_41 ();
 sg13g2_fill_1 FILLER_59_48 ();
 sg13g2_fill_1 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_136 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_145 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_157 ();
 sg13g2_fill_2 FILLER_59_196 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_fill_2 FILLER_59_312 ();
 sg13g2_fill_1 FILLER_59_314 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_332 ();
 sg13g2_fill_1 FILLER_59_352 ();
 sg13g2_fill_2 FILLER_59_356 ();
 sg13g2_fill_2 FILLER_59_393 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_fill_2 FILLER_59_428 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_10 ();
 sg13g2_fill_1 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_30 ();
 sg13g2_fill_1 FILLER_60_40 ();
 sg13g2_fill_1 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_61 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_decap_4 FILLER_60_89 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_decap_4 FILLER_60_109 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_fill_1 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_125 ();
 sg13g2_fill_1 FILLER_60_144 ();
 sg13g2_fill_2 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_278 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_2 FILLER_60_300 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_decap_4 FILLER_60_363 ();
 sg13g2_fill_1 FILLER_60_378 ();
 sg13g2_decap_4 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_390 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_4 FILLER_61_15 ();
 sg13g2_fill_2 FILLER_61_40 ();
 sg13g2_fill_1 FILLER_61_46 ();
 sg13g2_fill_2 FILLER_61_80 ();
 sg13g2_fill_2 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_194 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_fill_2 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_319 ();
 sg13g2_fill_2 FILLER_61_338 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_370 ();
 sg13g2_fill_2 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_390 ();
 sg13g2_fill_1 FILLER_61_395 ();
 sg13g2_fill_1 FILLER_61_400 ();
 sg13g2_fill_1 FILLER_61_404 ();
 sg13g2_fill_2 FILLER_61_410 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_fill_1 FILLER_62_10 ();
 sg13g2_fill_1 FILLER_62_15 ();
 sg13g2_fill_2 FILLER_62_29 ();
 sg13g2_fill_2 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_61 ();
 sg13g2_fill_2 FILLER_62_66 ();
 sg13g2_fill_1 FILLER_62_86 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_fill_2 FILLER_62_144 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_fill_2 FILLER_62_165 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_fill_1 FILLER_62_212 ();
 sg13g2_fill_2 FILLER_62_262 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_296 ();
 sg13g2_fill_2 FILLER_62_300 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_313 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_359 ();
 sg13g2_decap_4 FILLER_62_365 ();
 sg13g2_fill_2 FILLER_62_378 ();
 sg13g2_fill_2 FILLER_62_387 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_418 ();
 sg13g2_fill_2 FILLER_62_428 ();
 sg13g2_fill_1 FILLER_63_9 ();
 sg13g2_fill_1 FILLER_63_74 ();
 sg13g2_fill_1 FILLER_63_80 ();
 sg13g2_fill_1 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_142 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_fill_2 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_178 ();
 sg13g2_fill_2 FILLER_63_220 ();
 sg13g2_fill_2 FILLER_63_226 ();
 sg13g2_decap_4 FILLER_63_231 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_2 FILLER_63_241 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_1 FILLER_63_280 ();
 sg13g2_fill_1 FILLER_63_284 ();
 sg13g2_fill_1 FILLER_63_316 ();
 sg13g2_fill_2 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_329 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_fill_2 FILLER_63_359 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_374 ();
 sg13g2_fill_2 FILLER_63_381 ();
 sg13g2_fill_1 FILLER_63_383 ();
 sg13g2_fill_1 FILLER_63_392 ();
 sg13g2_fill_1 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_fill_2 FILLER_63_418 ();
 sg13g2_fill_1 FILLER_63_420 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_fill_1 FILLER_64_29 ();
 sg13g2_fill_1 FILLER_64_40 ();
 sg13g2_decap_4 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_89 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_114 ();
 sg13g2_fill_1 FILLER_64_119 ();
 sg13g2_fill_1 FILLER_64_129 ();
 sg13g2_fill_2 FILLER_64_187 ();
 sg13g2_fill_2 FILLER_64_192 ();
 sg13g2_fill_2 FILLER_64_198 ();
 sg13g2_fill_2 FILLER_64_204 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_fill_1 FILLER_64_290 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_305 ();
 sg13g2_fill_1 FILLER_64_312 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_337 ();
 sg13g2_fill_2 FILLER_64_351 ();
 sg13g2_fill_2 FILLER_64_369 ();
 sg13g2_fill_1 FILLER_64_371 ();
 sg13g2_fill_1 FILLER_64_375 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_fill_1 FILLER_64_388 ();
 sg13g2_fill_2 FILLER_64_394 ();
 sg13g2_fill_2 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_5 ();
 sg13g2_fill_2 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_52 ();
 sg13g2_fill_2 FILLER_65_57 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_2 FILLER_65_90 ();
 sg13g2_fill_2 FILLER_65_96 ();
 sg13g2_fill_2 FILLER_65_127 ();
 sg13g2_fill_2 FILLER_65_166 ();
 sg13g2_fill_1 FILLER_65_168 ();
 sg13g2_fill_2 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_fill_2 FILLER_65_245 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_318 ();
 sg13g2_fill_2 FILLER_65_323 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_fill_1 FILLER_65_341 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_fill_1 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_366 ();
 sg13g2_fill_1 FILLER_65_372 ();
 sg13g2_fill_2 FILLER_65_385 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_65_421 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_33 ();
 sg13g2_fill_1 FILLER_66_79 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_2 FILLER_66_106 ();
 sg13g2_fill_2 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_134 ();
 sg13g2_fill_1 FILLER_66_144 ();
 sg13g2_fill_2 FILLER_66_149 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_fill_2 FILLER_66_162 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_180 ();
 sg13g2_fill_2 FILLER_66_185 ();
 sg13g2_fill_1 FILLER_66_191 ();
 sg13g2_fill_1 FILLER_66_210 ();
 sg13g2_decap_4 FILLER_66_222 ();
 sg13g2_fill_2 FILLER_66_226 ();
 sg13g2_fill_2 FILLER_66_232 ();
 sg13g2_fill_1 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_260 ();
 sg13g2_fill_1 FILLER_66_287 ();
 sg13g2_fill_1 FILLER_66_296 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_310 ();
 sg13g2_fill_2 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_1 FILLER_66_397 ();
 sg13g2_fill_1 FILLER_66_403 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_13 ();
 sg13g2_fill_1 FILLER_67_23 ();
 sg13g2_fill_1 FILLER_67_34 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_61 ();
 sg13g2_fill_2 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_95 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_133 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_176 ();
 sg13g2_fill_1 FILLER_67_187 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_349 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_399 ();
 sg13g2_fill_1 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_6 ();
 sg13g2_fill_1 FILLER_68_12 ();
 sg13g2_fill_1 FILLER_68_27 ();
 sg13g2_fill_2 FILLER_68_43 ();
 sg13g2_fill_2 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_91 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_fill_2 FILLER_68_123 ();
 sg13g2_fill_1 FILLER_68_129 ();
 sg13g2_fill_2 FILLER_68_134 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_fill_2 FILLER_68_182 ();
 sg13g2_fill_2 FILLER_68_204 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_1 FILLER_68_233 ();
 sg13g2_fill_1 FILLER_68_237 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_fill_1 FILLER_68_256 ();
 sg13g2_fill_2 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_268 ();
 sg13g2_fill_2 FILLER_68_274 ();
 sg13g2_fill_1 FILLER_68_276 ();
 sg13g2_fill_1 FILLER_68_308 ();
 sg13g2_fill_1 FILLER_68_313 ();
 sg13g2_fill_1 FILLER_68_322 ();
 sg13g2_fill_1 FILLER_68_350 ();
 sg13g2_fill_2 FILLER_68_356 ();
 sg13g2_fill_1 FILLER_68_376 ();
 sg13g2_fill_2 FILLER_68_390 ();
 sg13g2_fill_1 FILLER_68_400 ();
 sg13g2_fill_1 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_fill_1 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_fill_1 FILLER_69_13 ();
 sg13g2_fill_1 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_33 ();
 sg13g2_fill_1 FILLER_69_38 ();
 sg13g2_fill_1 FILLER_69_43 ();
 sg13g2_fill_2 FILLER_69_59 ();
 sg13g2_fill_1 FILLER_69_94 ();
 sg13g2_fill_1 FILLER_69_118 ();
 sg13g2_fill_1 FILLER_69_245 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_4 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_333 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_fill_2 FILLER_69_353 ();
 sg13g2_fill_2 FILLER_69_359 ();
 sg13g2_fill_2 FILLER_69_365 ();
 sg13g2_fill_1 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_373 ();
 sg13g2_fill_2 FILLER_69_379 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_fill_2 FILLER_69_392 ();
 sg13g2_fill_2 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_410 ();
 sg13g2_fill_1 FILLER_69_420 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_fill_1 FILLER_70_29 ();
 sg13g2_fill_2 FILLER_70_33 ();
 sg13g2_fill_1 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_decap_8 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_158 ();
 sg13g2_fill_1 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_2 FILLER_70_337 ();
 sg13g2_fill_2 FILLER_70_374 ();
 sg13g2_fill_1 FILLER_70_379 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_fill_1 FILLER_70_405 ();
 sg13g2_fill_2 FILLER_70_410 ();
 sg13g2_fill_1 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_417 ();
 sg13g2_decap_4 FILLER_70_426 ();
 sg13g2_fill_1 FILLER_71_31 ();
 sg13g2_fill_1 FILLER_71_36 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_66 ();
 sg13g2_fill_1 FILLER_71_75 ();
 sg13g2_decap_4 FILLER_71_163 ();
 sg13g2_fill_1 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_201 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_238 ();
 sg13g2_fill_2 FILLER_71_290 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_decap_8 FILLER_71_297 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_fill_1 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_314 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_334 ();
 sg13g2_decap_4 FILLER_71_360 ();
 sg13g2_decap_8 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_1 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_22 ();
 sg13g2_fill_1 FILLER_72_28 ();
 sg13g2_fill_1 FILLER_72_34 ();
 sg13g2_fill_1 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_110 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_fill_1 FILLER_72_214 ();
 sg13g2_decap_4 FILLER_72_266 ();
 sg13g2_fill_1 FILLER_72_301 ();
 sg13g2_fill_1 FILLER_72_308 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_2 FILLER_72_340 ();
 sg13g2_fill_2 FILLER_72_370 ();
 sg13g2_fill_2 FILLER_72_416 ();
 sg13g2_fill_2 FILLER_73_12 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_79 ();
 sg13g2_fill_1 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_89 ();
 sg13g2_fill_1 FILLER_73_103 ();
 sg13g2_fill_2 FILLER_73_142 ();
 sg13g2_fill_1 FILLER_73_191 ();
 sg13g2_fill_2 FILLER_73_212 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_2 FILLER_73_261 ();
 sg13g2_fill_1 FILLER_73_263 ();
 sg13g2_fill_1 FILLER_73_329 ();
 sg13g2_decap_4 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_356 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_decap_4 FILLER_73_375 ();
 sg13g2_fill_1 FILLER_73_383 ();
 sg13g2_fill_2 FILLER_73_388 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_fill_2 FILLER_73_416 ();
 sg13g2_fill_1 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_89 ();
 sg13g2_fill_1 FILLER_74_158 ();
 sg13g2_fill_1 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_329 ();
 sg13g2_fill_2 FILLER_74_348 ();
 sg13g2_fill_1 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_decap_4 FILLER_74_418 ();
 sg13g2_fill_1 FILLER_74_422 ();
 sg13g2_fill_2 FILLER_74_427 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_fill_2 FILLER_75_31 ();
 sg13g2_fill_2 FILLER_75_59 ();
 sg13g2_fill_2 FILLER_75_69 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_211 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_1 FILLER_75_224 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_fill_1 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_249 ();
 sg13g2_fill_2 FILLER_75_259 ();
 sg13g2_fill_2 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_fill_2 FILLER_75_304 ();
 sg13g2_fill_1 FILLER_75_336 ();
 sg13g2_fill_1 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_decap_4 FILLER_75_363 ();
 sg13g2_fill_1 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_422 ();
 sg13g2_fill_2 FILLER_75_428 ();
 sg13g2_fill_1 FILLER_76_26 ();
 sg13g2_fill_2 FILLER_76_62 ();
 sg13g2_fill_1 FILLER_76_133 ();
 sg13g2_fill_2 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_251 ();
 sg13g2_fill_1 FILLER_76_352 ();
 sg13g2_fill_1 FILLER_76_357 ();
 sg13g2_fill_1 FILLER_76_362 ();
 sg13g2_fill_2 FILLER_76_376 ();
 sg13g2_fill_1 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_decap_4 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_410 ();
 sg13g2_fill_2 FILLER_76_428 ();
 sg13g2_fill_2 FILLER_77_41 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_fill_2 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_2 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_233 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_316 ();
 sg13g2_fill_1 FILLER_77_331 ();
 sg13g2_decap_4 FILLER_77_335 ();
 sg13g2_fill_1 FILLER_77_339 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_358 ();
 sg13g2_fill_1 FILLER_77_362 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_fill_1 FILLER_77_383 ();
 sg13g2_fill_1 FILLER_77_389 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_fill_1 FILLER_77_398 ();
 sg13g2_fill_1 FILLER_77_407 ();
 sg13g2_fill_2 FILLER_77_413 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_78_47 ();
 sg13g2_fill_2 FILLER_78_73 ();
 sg13g2_fill_1 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_157 ();
 sg13g2_fill_1 FILLER_78_162 ();
 sg13g2_fill_1 FILLER_78_172 ();
 sg13g2_fill_2 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_209 ();
 sg13g2_fill_2 FILLER_78_316 ();
 sg13g2_fill_1 FILLER_78_325 ();
 sg13g2_decap_4 FILLER_78_331 ();
 sg13g2_fill_1 FILLER_78_392 ();
 sg13g2_fill_1 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_411 ();
 sg13g2_fill_2 FILLER_78_416 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_fill_2 FILLER_79_31 ();
 sg13g2_fill_1 FILLER_79_93 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_168 ();
 sg13g2_fill_2 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_384 ();
 sg13g2_fill_1 FILLER_79_416 ();
 sg13g2_decap_4 FILLER_79_426 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_66 ();
 sg13g2_fill_2 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_91 ();
 sg13g2_fill_2 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_394 ();
 sg13g2_fill_1 FILLER_80_419 ();
 sg13g2_fill_2 FILLER_80_427 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
