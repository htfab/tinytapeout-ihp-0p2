module tt_um_dlmiles_tt05_i2c_bert (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire clknet_0_clk;
 wire net110;
 wire \i2c_bert.div12[0] ;
 wire \i2c_bert.div12[10] ;
 wire \i2c_bert.div12[11] ;
 wire \i2c_bert.div12[1] ;
 wire \i2c_bert.div12[2] ;
 wire \i2c_bert.div12[3] ;
 wire \i2c_bert.div12[4] ;
 wire \i2c_bert.div12[5] ;
 wire \i2c_bert.div12[6] ;
 wire \i2c_bert.div12[7] ;
 wire \i2c_bert.div12[8] ;
 wire \i2c_bert.div12[9] ;
 wire \i2c_bert.i2c.clockGate.sel ;
 wire \i2c_bert.i2c.fsm_bitCount[0] ;
 wire \i2c_bert.i2c.fsm_bitCount[1] ;
 wire \i2c_bert.i2c.fsm_bitCount[2] ;
 wire \i2c_bert.i2c.fsm_stateReg[0] ;
 wire \i2c_bert.i2c.fsm_stateReg[1] ;
 wire \i2c_bert.i2c.fsm_stateReg[2] ;
 wire \i2c_bert.i2c.fsm_stateReg[3] ;
 wire \i2c_bert.i2c.fsm_wantStart ;
 wire \i2c_bert.i2c.io_bus_sclOe ;
 wire \i2c_bert.i2c.io_bus_sclOut ;
 wire \i2c_bert.i2c.io_bus_sdaOe ;
 wire \i2c_bert.i2c.io_bus_sdaOut ;
 wire \i2c_bert.i2c.io_canStretch ;
 wire \i2c_bert.i2c.io_data8rx[0] ;
 wire \i2c_bert.i2c.io_data8rx[1] ;
 wire \i2c_bert.i2c.io_data8rx[2] ;
 wire \i2c_bert.i2c.io_data8rx[3] ;
 wire \i2c_bert.i2c.io_data8rx[4] ;
 wire \i2c_bert.i2c.io_data8rx[5] ;
 wire \i2c_bert.i2c.io_data8rx[6] ;
 wire \i2c_bert.i2c.io_data8rx[7] ;
 wire \i2c_bert.i2c.io_pushPullMode ;
 wire \i2c_bert.i2c.io_sclMode[1] ;
 wire \i2c_bert.i2c.io_sclMode[2] ;
 wire \i2c_bert.i2c.io_sdaSignal ;
 wire \i2c_bert.i2c.io_timerAutobaud ;
 wire \i2c_bert.i2c.io_wantReset ;
 wire \i2c_bert.i2c.rst_n ;
 wire \i2c_bert.i2c.scl ;
 wire \i2c_bert.i2c.sclAndNor3.io_b ;
 wire \i2c_bert.i2c.sclAndNor3.io_c ;
 wire \i2c_bert.i2c.sclAndNor3.io_o ;
 wire \i2c_bert.i2c.sclAndNor5.io_d ;
 wire \i2c_bert.i2c.sclAndNor5.io_e ;
 wire \i2c_bert.i2c.sclAndNor5.io_o ;
 wire \i2c_bert.i2c.scl_regNext ;
 wire \i2c_bert.i2c.sdaAndNor3.io_b ;
 wire \i2c_bert.i2c.sdaAndNor3.io_c ;
 wire \i2c_bert.i2c.sdaAndNor3.io_o ;
 wire \i2c_bert.i2c.sdaAndNor5.io_d ;
 wire \i2c_bert.i2c.sdaAndNor5.io_e ;
 wire \i2c_bert.i2c.sdaAndNor5.io_o ;
 wire \i2c_bert.i2c.sda_regNext ;
 wire \i2c_bert.latched[16] ;
 wire \i2c_bert.latched[17] ;
 wire \i2c_bert.latched[18] ;
 wire \i2c_bert.latched[19] ;
 wire \i2c_bert.latched[20] ;
 wire \i2c_bert.latched[21] ;
 wire \i2c_bert.latched[22] ;
 wire \i2c_bert.latched[23] ;
 wire \i2c_bert.latched[24] ;
 wire \i2c_bert.latched[25] ;
 wire \i2c_bert.latched[26] ;
 wire \i2c_bert.latched[27] ;
 wire \i2c_bert.latched[28] ;
 wire \i2c_bert.latched[29] ;
 wire \i2c_bert.latched[30] ;
 wire \i2c_bert.latched[31] ;
 wire \i2c_bert.myState_1._zz__zz_io_data8tx[0] ;
 wire \i2c_bert.myState_1._zz__zz_io_data8tx[1] ;
 wire \i2c_bert.myState_1._zz__zz_io_data8tx[2] ;
 wire \i2c_bert.myState_1._zz__zz_io_data8tx[3] ;
 wire \i2c_bert.myState_1.alu_1.acc[0] ;
 wire \i2c_bert.myState_1.alu_1.acc[1] ;
 wire \i2c_bert.myState_1.alu_1.acc[2] ;
 wire \i2c_bert.myState_1.alu_1.acc[3] ;
 wire \i2c_bert.myState_1.alu_1.acc[4] ;
 wire \i2c_bert.myState_1.alu_1.acc[5] ;
 wire \i2c_bert.myState_1.alu_1.acc[6] ;
 wire \i2c_bert.myState_1.alu_1.acc[7] ;
 wire \i2c_bert.myState_1.alu_1.io_op[0] ;
 wire \i2c_bert.myState_1.alu_1.io_op[1] ;
 wire \i2c_bert.myState_1.cmd7[0] ;
 wire \i2c_bert.myState_1.cmd7[3] ;
 wire \i2c_bert.myState_1.cmd7[4] ;
 wire \i2c_bert.myState_1.cmd7[5] ;
 wire \i2c_bert.myState_1.cmd7[6] ;
 wire \i2c_bert.myState_1.counter[0] ;
 wire \i2c_bert.myState_1.counter[10] ;
 wire \i2c_bert.myState_1.counter[11] ;
 wire \i2c_bert.myState_1.counter[1] ;
 wire \i2c_bert.myState_1.counter[2] ;
 wire \i2c_bert.myState_1.counter[3] ;
 wire \i2c_bert.myState_1.counter[4] ;
 wire \i2c_bert.myState_1.counter[5] ;
 wire \i2c_bert.myState_1.counter[6] ;
 wire \i2c_bert.myState_1.counter[7] ;
 wire \i2c_bert.myState_1.counter[8] ;
 wire \i2c_bert.myState_1.counter[9] ;
 wire \i2c_bert.myState_1.fsmPhase_stateReg[1] ;
 wire \i2c_bert.myState_1.fsmPhase_stateReg[2] ;
 wire \i2c_bert.myState_1.fsmPhase_stateReg[3] ;
 wire \i2c_bert.myState_1.fsmPhase_stateReg[5] ;
 wire \i2c_bert.myState_1.io_timerEndstop[0] ;
 wire \i2c_bert.myState_1.io_timerEndstop[1] ;
 wire \i2c_bert.myState_1.io_timerEndstop[2] ;
 wire \i2c_bert.myState_1.io_timerEndstop[3] ;
 wire \i2c_bert.myState_1.io_timerEndstop[4] ;
 wire \i2c_bert.myState_1.io_timerEndstop[5] ;
 wire \i2c_bert.myState_1.io_timerEndstop[6] ;
 wire \i2c_bert.myState_1.io_timerEndstop[7] ;
 wire \i2c_bert.myState_1.led8[0] ;
 wire \i2c_bert.myState_1.led8[1] ;
 wire \i2c_bert.myState_1.led8[2] ;
 wire \i2c_bert.myState_1.led8[3] ;
 wire \i2c_bert.myState_1.led8[4] ;
 wire \i2c_bert.myState_1.led8[5] ;
 wire \i2c_bert.myState_1.led8[6] ;
 wire \i2c_bert.myState_1.led8[7] ;
 wire \i2c_bert.myState_1.len12[10] ;
 wire \i2c_bert.myState_1.len12[11] ;
 wire \i2c_bert.myState_1.len12[4] ;
 wire \i2c_bert.myState_1.len12[5] ;
 wire \i2c_bert.myState_1.len12[6] ;
 wire \i2c_bert.myState_1.len12[7] ;
 wire \i2c_bert.myState_1.len12[8] ;
 wire \i2c_bert.myState_1.len12[9] ;
 wire \i2c_bert.myState_1.readWriteBit ;
 wire \i2c_bert.powerOnSense.D ;
 wire \i2c_bert.powerOnSense.GATE ;
 wire \i2c_bert.powerOnSense.Q ;
 wire \i2c_bert.powerOnSenseCaptured.GATE ;
 wire \i2c_bert.powerOnSenseCaptured.Q ;
 wire \i2c_bert.timer_1.ticker_count[0] ;
 wire \i2c_bert.timer_1.ticker_count[10] ;
 wire \i2c_bert.timer_1.ticker_count[11] ;
 wire \i2c_bert.timer_1.ticker_count[1] ;
 wire \i2c_bert.timer_1.ticker_count[2] ;
 wire \i2c_bert.timer_1.ticker_count[3] ;
 wire \i2c_bert.timer_1.ticker_count[4] ;
 wire \i2c_bert.timer_1.ticker_count[5] ;
 wire \i2c_bert.timer_1.ticker_count[6] ;
 wire \i2c_bert.timer_1.ticker_count[7] ;
 wire \i2c_bert.timer_1.ticker_count[8] ;
 wire \i2c_bert.timer_1.ticker_count[9] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[0] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[1] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[2] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[3] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[4] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[5] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[6] ;
 wire \i2c_bert.timer_1.ticker_endstopTmpL[7] ;
 wire \i2c_bert.timer_1.ticker_timerSampleTickState ;
 wire \i2c_bert.timer_1.ticker_timerSampleTickState_regNext ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_1 _1259_ (.Y(_0764_),
    .A(\i2c_bert.myState_1.readWriteBit ));
 sg13g2_a22oi_1 _1260_ (.Y(_0765_),
    .B1(_0763_),
    .B2(_0764_),
    .A2(_0761_),
    .A1(_0754_));
 sg13g2_buf_1 _1261_ (.A(net87),
    .X(_0766_));
 sg13g2_inv_1 _1262_ (.Y(_0767_),
    .A(_0620_));
 sg13g2_buf_1 _1263_ (.A(_0608_),
    .X(_0768_));
 sg13g2_and2_1 _1264_ (.A(net73),
    .B(_0628_),
    .X(_0769_));
 sg13g2_nor4_1 _1265_ (.A(\i2c_bert.i2c.io_wantReset ),
    .B(net50),
    .C(_0767_),
    .D(_0769_),
    .Y(_0770_));
 sg13g2_a21oi_1 _1266_ (.A1(_0025_),
    .A2(net50),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_nor3_1 _1267_ (.A(net85),
    .B(_0638_),
    .C(_0620_),
    .Y(_0772_));
 sg13g2_o21ai_1 _1268_ (.B1(_0689_),
    .Y(_0773_),
    .A1(_0709_),
    .A2(_0772_));
 sg13g2_o21ai_1 _1269_ (.B1(_0773_),
    .Y(_0774_),
    .A1(_0594_),
    .A2(_0771_));
 sg13g2_nand2_1 _1270_ (.Y(_0775_),
    .A(net74),
    .B(_0774_));
 sg13g2_o21ai_1 _1271_ (.B1(_0775_),
    .Y(_0005_),
    .A1(_0595_),
    .A2(_0765_));
 sg13g2_nand3_1 _1272_ (.B(_0025_),
    .C(_0605_),
    .A(net79),
    .Y(_0776_));
 sg13g2_a21oi_1 _1273_ (.A1(_0593_),
    .A2(_0776_),
    .Y(_0002_),
    .B1(_0582_));
 sg13g2_nor2_1 _1274_ (.A(_0648_),
    .B(_0656_),
    .Y(_0777_));
 sg13g2_o21ai_1 _1275_ (.B1(_0755_),
    .Y(_0778_),
    .A1(_0664_),
    .A2(_0777_));
 sg13g2_and4_1 _1276_ (.A(net79),
    .B(\i2c_bert.i2c.io_sdaSignal ),
    .C(net49),
    .D(_0778_),
    .X(_0779_));
 sg13g2_a21oi_1 _1277_ (.A1(\i2c_bert.myState_1.readWriteBit ),
    .A2(_0763_),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_nand2b_1 _1278_ (.Y(_0781_),
    .B(_0721_),
    .A_N(_0717_));
 sg13g2_nor2_1 _1279_ (.A(\i2c_bert.i2c.io_wantReset ),
    .B(_0743_),
    .Y(_0782_));
 sg13g2_nand4_1 _1280_ (.B(_0724_),
    .C(_0781_),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[1] ),
    .Y(_0783_),
    .D(_0782_));
 sg13g2_o21ai_1 _1281_ (.B1(_0783_),
    .Y(_0001_),
    .A1(_0595_),
    .A2(_0780_));
 sg13g2_o21ai_1 _1282_ (.B1(_0020_),
    .Y(_0784_),
    .A1(net76),
    .A2(_0730_));
 sg13g2_inv_1 _1283_ (.Y(_0785_),
    .A(_0584_));
 sg13g2_nand2_2 _1284_ (.Y(_0786_),
    .A(_0785_),
    .B(\i2c_bert.i2c.fsm_stateReg[0] ));
 sg13g2_buf_1 _1285_ (.A(_0586_),
    .X(_0787_));
 sg13g2_inv_1 _1286_ (.Y(_0788_),
    .A(_0587_));
 sg13g2_nor2_2 _1287_ (.A(net72),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_a21oi_1 _1288_ (.A1(_0745_),
    .A2(_0789_),
    .Y(_0790_),
    .B1(_0737_));
 sg13g2_nor2_1 _1289_ (.A(_0786_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nor4_1 _1290_ (.A(_0555_),
    .B(_0581_),
    .C(_0784_),
    .D(_0791_),
    .Y(_0792_));
 sg13g2_nand2_1 _1291_ (.Y(_0793_),
    .A(\i2c_bert.timer_1.ticker_count[11] ),
    .B(\i2c_bert.i2c.io_timerAutobaud ));
 sg13g2_nor3_1 _1292_ (.A(\i2c_bert.myState_1._zz__zz_io_data8tx[3] ),
    .B(\i2c_bert.timer_1.ticker_count[11] ),
    .C(\i2c_bert.i2c.io_timerAutobaud ),
    .Y(_0794_));
 sg13g2_and2_1 _1293_ (.A(\i2c_bert.myState_1._zz__zz_io_data8tx[3] ),
    .B(\i2c_bert.timer_1.ticker_count[11] ),
    .X(_0795_));
 sg13g2_buf_1 _1294_ (.A(\i2c_bert.timer_1.ticker_count[9] ),
    .X(_0796_));
 sg13g2_xnor2_1 _1295_ (.Y(_0797_),
    .A(\i2c_bert.myState_1._zz__zz_io_data8tx[1] ),
    .B(_0796_));
 sg13g2_buf_2 _1296_ (.A(\i2c_bert.timer_1.ticker_count[8] ),
    .X(_0798_));
 sg13g2_xnor2_1 _1297_ (.Y(_0799_),
    .A(\i2c_bert.myState_1._zz__zz_io_data8tx[0] ),
    .B(_0798_));
 sg13g2_xnor2_1 _1298_ (.Y(_0800_),
    .A(\i2c_bert.myState_1.io_timerEndstop[2] ),
    .B(\i2c_bert.timer_1.ticker_count[2] ));
 sg13g2_nand3_1 _1299_ (.B(_0799_),
    .C(_0800_),
    .A(_0797_),
    .Y(_0801_));
 sg13g2_xnor2_1 _1300_ (.Y(_0802_),
    .A(\i2c_bert.myState_1._zz__zz_io_data8tx[2] ),
    .B(\i2c_bert.timer_1.ticker_count[10] ));
 sg13g2_xnor2_1 _1301_ (.Y(_0803_),
    .A(\i2c_bert.myState_1.io_timerEndstop[6] ),
    .B(\i2c_bert.timer_1.ticker_count[6] ));
 sg13g2_xnor2_1 _1302_ (.Y(_0804_),
    .A(\i2c_bert.myState_1.io_timerEndstop[7] ),
    .B(\i2c_bert.timer_1.ticker_count[7] ));
 sg13g2_buf_2 _1303_ (.A(\i2c_bert.timer_1.ticker_count[4] ),
    .X(_0805_));
 sg13g2_xnor2_1 _1304_ (.Y(_0806_),
    .A(\i2c_bert.myState_1.io_timerEndstop[4] ),
    .B(_0805_));
 sg13g2_nand4_1 _1305_ (.B(_0803_),
    .C(_0804_),
    .A(_0802_),
    .Y(_0807_),
    .D(_0806_));
 sg13g2_buf_2 _1306_ (.A(\i2c_bert.timer_1.ticker_count[0] ),
    .X(_0808_));
 sg13g2_xnor2_1 _1307_ (.Y(_0809_),
    .A(\i2c_bert.myState_1.io_timerEndstop[0] ),
    .B(_0808_));
 sg13g2_xnor2_1 _1308_ (.Y(_0810_),
    .A(\i2c_bert.myState_1.io_timerEndstop[3] ),
    .B(\i2c_bert.timer_1.ticker_count[3] ));
 sg13g2_buf_2 _1309_ (.A(\i2c_bert.timer_1.ticker_count[5] ),
    .X(_0811_));
 sg13g2_xnor2_1 _1310_ (.Y(_0812_),
    .A(\i2c_bert.myState_1.io_timerEndstop[5] ),
    .B(_0811_));
 sg13g2_buf_2 _1311_ (.A(\i2c_bert.timer_1.ticker_count[1] ),
    .X(_0813_));
 sg13g2_xnor2_1 _1312_ (.Y(_0814_),
    .A(\i2c_bert.myState_1.io_timerEndstop[1] ),
    .B(_0813_));
 sg13g2_nand4_1 _1313_ (.B(_0810_),
    .C(_0812_),
    .A(_0809_),
    .Y(_0815_),
    .D(_0814_));
 sg13g2_nor3_1 _1314_ (.A(_0801_),
    .B(_0807_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_o21ai_1 _1315_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0794_),
    .A2(_0795_));
 sg13g2_nand2_1 _1316_ (.Y(_0818_),
    .A(_0793_),
    .B(_0817_));
 sg13g2_or2_1 _1317_ (.X(_0819_),
    .B(_0818_),
    .A(_0792_));
 sg13g2_nor2_1 _1318_ (.A(_0785_),
    .B(_0787_),
    .Y(_0820_));
 sg13g2_buf_1 _1319_ (.A(_0587_),
    .X(_0821_));
 sg13g2_xor2_1 _1320_ (.B(net71),
    .A(net76),
    .X(_0822_));
 sg13g2_nor2_2 _1321_ (.A(_0730_),
    .B(_0786_),
    .Y(_0823_));
 sg13g2_a21o_1 _1322_ (.A2(_0822_),
    .A1(_0820_),
    .B1(_0823_),
    .X(_0824_));
 sg13g2_buf_1 _1323_ (.A(_0824_),
    .X(_0825_));
 sg13g2_o21ai_1 _1324_ (.B1(_0825_),
    .Y(_0826_),
    .A1(net53),
    .A2(_0602_));
 sg13g2_nand2_1 _1325_ (.Y(_0827_),
    .A(net53),
    .B(_0739_));
 sg13g2_a21oi_1 _1326_ (.A1(_0826_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(_0028_));
 sg13g2_buf_1 _1327_ (.A(_0597_),
    .X(_0829_));
 sg13g2_buf_2 _1328_ (.A(_0019_),
    .X(_0830_));
 sg13g2_and2_1 _1329_ (.A(_0539_),
    .B(_0028_),
    .X(_0831_));
 sg13g2_a21oi_1 _1330_ (.A1(_0540_),
    .A2(_0830_),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_o21ai_1 _1331_ (.B1(_0733_),
    .Y(_0833_),
    .A1(net55),
    .A2(_0832_));
 sg13g2_nand2_1 _1332_ (.Y(_0834_),
    .A(_0598_),
    .B(_0788_));
 sg13g2_nor2_1 _1333_ (.A(_0787_),
    .B(_0028_),
    .Y(_0835_));
 sg13g2_a21oi_1 _1334_ (.A1(net72),
    .A2(_0540_),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_nand2_1 _1335_ (.Y(_0837_),
    .A(net76),
    .B(_0587_));
 sg13g2_o21ai_1 _1336_ (.B1(_0837_),
    .Y(_0838_),
    .A1(_0834_),
    .A2(_0836_));
 sg13g2_buf_1 _1337_ (.A(_0736_),
    .X(_0839_));
 sg13g2_nor3_1 _1338_ (.A(net64),
    .B(net70),
    .C(net72),
    .Y(_0840_));
 sg13g2_o21ai_1 _1339_ (.B1(net70),
    .Y(_0841_),
    .A1(net72),
    .A2(net77));
 sg13g2_nand2b_1 _1340_ (.Y(_0842_),
    .B(_0841_),
    .A_N(_0840_));
 sg13g2_a22oi_1 _1341_ (.Y(_0843_),
    .B1(_0842_),
    .B2(net71),
    .A2(_0838_),
    .A1(net64));
 sg13g2_nand3_1 _1342_ (.B(_0833_),
    .C(_0843_),
    .A(_0593_),
    .Y(_0844_));
 sg13g2_nor4_2 _1343_ (.A(\i2c_bert.i2c.fsm_wantStart ),
    .B(_0819_),
    .C(_0828_),
    .Y(_0845_),
    .D(_0844_));
 sg13g2_nor2_1 _1344_ (.A(_0584_),
    .B(_0736_),
    .Y(_0846_));
 sg13g2_nand2_2 _1345_ (.Y(_0847_),
    .A(_0737_),
    .B(_0846_));
 sg13g2_nor3_1 _1346_ (.A(net77),
    .B(_0670_),
    .C(_0847_),
    .Y(_0848_));
 sg13g2_nor2_1 _1347_ (.A(_0024_),
    .B(_0738_),
    .Y(_0849_));
 sg13g2_mux2_1 _1348_ (.A0(_0848_),
    .A1(_0849_),
    .S(_0741_),
    .X(_0850_));
 sg13g2_nor2_1 _1349_ (.A(_0598_),
    .B(net71),
    .Y(_0851_));
 sg13g2_inv_1 _1350_ (.Y(_0852_),
    .A(_0586_));
 sg13g2_nand3_1 _1351_ (.B(_0852_),
    .C(_0725_),
    .A(net76),
    .Y(_0853_));
 sg13g2_a21oi_1 _1352_ (.A1(_0730_),
    .A2(_0853_),
    .Y(_0854_),
    .B1(net64));
 sg13g2_a21oi_1 _1353_ (.A1(\i2c_bert.i2c.io_canStretch ),
    .A2(\i2c_bert.myState_1.readWriteBit ),
    .Y(_0855_),
    .B1(\i2c_bert.myState_1.fsmPhase_stateReg[1] ));
 sg13g2_a21oi_1 _1354_ (.A1(net71),
    .A2(_0855_),
    .Y(_0856_),
    .B1(net64));
 sg13g2_nor3_1 _1355_ (.A(net70),
    .B(net72),
    .C(_0856_),
    .Y(_0857_));
 sg13g2_nor3_1 _1356_ (.A(_0851_),
    .B(_0854_),
    .C(_0857_),
    .Y(_0858_));
 sg13g2_nor2_1 _1357_ (.A(_0850_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_nor2_1 _1358_ (.A(net53),
    .B(_0602_),
    .Y(_0860_));
 sg13g2_nand2_1 _1359_ (.Y(_0861_),
    .A(_0860_),
    .B(_0825_));
 sg13g2_a21oi_1 _1360_ (.A1(net64),
    .A2(net70),
    .Y(_0862_),
    .B1(net72));
 sg13g2_nand2b_1 _1361_ (.Y(_0863_),
    .B(_0846_),
    .A_N(_0589_));
 sg13g2_o21ai_1 _1362_ (.B1(_0863_),
    .Y(_0864_),
    .A1(_0788_),
    .A2(_0862_));
 sg13g2_a21oi_1 _1363_ (.A1(_0859_),
    .A2(_0861_),
    .Y(_0865_),
    .B1(_0864_));
 sg13g2_nor2_1 _1364_ (.A(_0540_),
    .B(_0597_),
    .Y(_0866_));
 sg13g2_nand3b_1 _1365_ (.B(\i2c_bert.i2c.scl ),
    .C(_0581_),
    .Y(_0867_),
    .A_N(_0020_));
 sg13g2_a22oi_1 _1366_ (.Y(_0868_),
    .B1(_0867_),
    .B2(_0590_),
    .A2(_0866_),
    .A1(_0733_));
 sg13g2_nor2_1 _1367_ (.A(net77),
    .B(_0847_),
    .Y(_0869_));
 sg13g2_inv_1 _1368_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_a21oi_1 _1369_ (.A1(_0670_),
    .A2(net55),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_nor4_1 _1370_ (.A(_0825_),
    .B(_0850_),
    .C(_0858_),
    .D(_0871_),
    .Y(_0872_));
 sg13g2_a21oi_1 _1371_ (.A1(_0868_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(_0024_));
 sg13g2_inv_1 _1372_ (.Y(_0874_),
    .A(_0021_));
 sg13g2_nor3_1 _1373_ (.A(_0874_),
    .B(_0792_),
    .C(_0818_),
    .Y(_0875_));
 sg13g2_o21ai_1 _1374_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0865_),
    .A2(_0873_));
 sg13g2_buf_1 _1375_ (.A(_0876_),
    .X(_0877_));
 sg13g2_o21ai_1 _1376_ (.B1(_0733_),
    .Y(_0878_),
    .A1(_0539_),
    .A2(_0745_));
 sg13g2_nand2_1 _1377_ (.Y(_0879_),
    .A(_0738_),
    .B(_0878_));
 sg13g2_a22oi_1 _1378_ (.Y(_0880_),
    .B1(_0879_),
    .B2(net53),
    .A2(_0837_),
    .A1(_0820_));
 sg13g2_nor2_1 _1379_ (.A(net70),
    .B(net71),
    .Y(_0881_));
 sg13g2_nor3_1 _1380_ (.A(_0741_),
    .B(_0602_),
    .C(_0881_),
    .Y(_0882_));
 sg13g2_nand3_1 _1381_ (.B(net76),
    .C(_0737_),
    .A(_0785_),
    .Y(_0883_));
 sg13g2_nor2b_1 _1382_ (.A(_0830_),
    .B_N(\i2c_bert.i2c.io_canStretch ),
    .Y(_0884_));
 sg13g2_o21ai_1 _1383_ (.B1(_0855_),
    .Y(_0885_),
    .A1(_0726_),
    .A2(_0884_));
 sg13g2_or4_1 _1384_ (.A(\i2c_bert.i2c.io_canStretch ),
    .B(_0730_),
    .C(_0732_),
    .D(_0885_),
    .X(_0886_));
 sg13g2_o21ai_1 _1385_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0602_),
    .A2(_0883_));
 sg13g2_o21ai_1 _1386_ (.B1(_0852_),
    .Y(_0888_),
    .A1(_0732_),
    .A2(_0885_));
 sg13g2_nand2_1 _1387_ (.Y(_0889_),
    .A(net76),
    .B(_0586_));
 sg13g2_o21ai_1 _1388_ (.B1(_0589_),
    .Y(_0890_),
    .A1(_0022_),
    .A2(_0889_));
 sg13g2_o21ai_1 _1389_ (.B1(_0837_),
    .Y(_0891_),
    .A1(net76),
    .A2(_0852_));
 sg13g2_mux2_1 _1390_ (.A0(_0890_),
    .A1(_0891_),
    .S(net64),
    .X(_0892_));
 sg13g2_a21o_1 _1391_ (.A2(_0888_),
    .A1(_0821_),
    .B1(_0892_),
    .X(_0893_));
 sg13g2_a221oi_1 _1392_ (.B2(_0887_),
    .C1(_0893_),
    .B1(net55),
    .A1(\i2c_bert.i2c.scl ),
    .Y(_0894_),
    .A2(_0592_));
 sg13g2_o21ai_1 _1393_ (.B1(_0894_),
    .Y(_0895_),
    .A1(_0880_),
    .A2(_0882_));
 sg13g2_a21oi_1 _1394_ (.A1(_0821_),
    .A2(_0888_),
    .Y(_0896_),
    .B1(_0892_));
 sg13g2_nand2_1 _1395_ (.Y(_0897_),
    .A(net55),
    .B(_0887_));
 sg13g2_nand4_1 _1396_ (.B(_0593_),
    .C(_0896_),
    .A(_0022_),
    .Y(_0898_),
    .D(_0897_));
 sg13g2_nand2_1 _1397_ (.Y(_0899_),
    .A(_0022_),
    .B(_0864_));
 sg13g2_nand4_1 _1398_ (.B(_0895_),
    .C(_0898_),
    .A(_0875_),
    .Y(_0900_),
    .D(_0899_));
 sg13g2_buf_2 _1399_ (.A(_0900_),
    .X(_0901_));
 sg13g2_nand3_1 _1400_ (.B(_0877_),
    .C(_0901_),
    .A(_0845_),
    .Y(_0902_));
 sg13g2_nand2_1 _1401_ (.Y(_0903_),
    .A(_0583_),
    .B(_0902_));
 sg13g2_o21ai_1 _1402_ (.B1(_0877_),
    .Y(_0904_),
    .A1(_0845_),
    .A2(_0901_));
 sg13g2_and2_1 _1403_ (.A(_0583_),
    .B(_0904_),
    .X(_0905_));
 sg13g2_o21ai_1 _1404_ (.B1(_0738_),
    .Y(_0906_),
    .A1(_0830_),
    .A2(_0847_));
 sg13g2_a22oi_1 _1405_ (.Y(_0907_),
    .B1(_0589_),
    .B2(net64),
    .A2(_0725_),
    .A1(net71));
 sg13g2_nand2b_1 _1406_ (.Y(_0908_),
    .B(net70),
    .A_N(_0907_));
 sg13g2_nand2_1 _1407_ (.Y(_0909_),
    .A(net72),
    .B(net71));
 sg13g2_nand3_1 _1408_ (.B(_0909_),
    .C(_0863_),
    .A(_0908_),
    .Y(_0910_));
 sg13g2_or4_1 _1409_ (.A(net53),
    .B(_0602_),
    .C(_0906_),
    .D(_0910_),
    .X(_0911_));
 sg13g2_nor3_1 _1410_ (.A(_0539_),
    .B(_0830_),
    .C(_0847_),
    .Y(_0912_));
 sg13g2_o21ai_1 _1411_ (.B1(_0906_),
    .Y(_0913_),
    .A1(net55),
    .A2(_0912_));
 sg13g2_a21oi_1 _1412_ (.A1(_0820_),
    .A2(_0822_),
    .Y(_0914_),
    .B1(_0823_));
 sg13g2_nand3b_1 _1413_ (.B(_0913_),
    .C(_0914_),
    .Y(_0915_),
    .A_N(_0910_));
 sg13g2_nand2_1 _1414_ (.Y(_0916_),
    .A(_0911_),
    .B(_0915_));
 sg13g2_nand2_1 _1415_ (.Y(_0917_),
    .A(_0852_),
    .B(net71));
 sg13g2_nor2_1 _1416_ (.A(_0786_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_inv_1 _1417_ (.Y(_0919_),
    .A(_0017_));
 sg13g2_a21oi_1 _1418_ (.A1(net77),
    .A2(_0918_),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_a22oi_1 _1419_ (.Y(_0921_),
    .B1(_0920_),
    .B2(_0913_),
    .A2(_0916_),
    .A1(_0868_));
 sg13g2_nand2_1 _1420_ (.Y(_0922_),
    .A(net78),
    .B(_0921_));
 sg13g2_nor3_1 _1421_ (.A(\i2c_bert.i2c.fsm_wantStart ),
    .B(_0819_),
    .C(_0922_),
    .Y(_0038_));
 sg13g2_mux2_1 _1422_ (.A0(_0903_),
    .A1(_0905_),
    .S(_0038_),
    .X(_0000_));
 sg13g2_buf_1 _1423_ (.A(net3),
    .X(_0923_));
 sg13g2_mux2_1 _1424_ (.A0(_0813_),
    .A1(\i2c_bert.timer_1.ticker_count[2] ),
    .S(_0923_),
    .X(_0924_));
 sg13g2_inv_1 _1425_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_nor2b_1 _1426_ (.A(net4),
    .B_N(_0923_),
    .Y(_0926_));
 sg13g2_a22oi_1 _1427_ (.Y(\i2c_bert.timer_1.ticker_timerSampleTickState ),
    .B1(_0926_),
    .B2(_0007_),
    .A2(_0925_),
    .A1(net4));
 sg13g2_nand2_1 _1428_ (.Y(_0927_),
    .A(net4),
    .B(\i2c_bert.timer_1.ticker_timerSampleTickState_regNext ));
 sg13g2_nand2_1 _1429_ (.Y(_0928_),
    .A(\i2c_bert.timer_1.ticker_timerSampleTickState ),
    .B(_0927_));
 sg13g2_buf_1 _1430_ (.A(_0928_),
    .X(_0929_));
 sg13g2_nand2_1 _1431_ (.Y(_0930_),
    .A(\i2c_bert.i2c.sclAndNor3.io_b ),
    .B(net57));
 sg13g2_o21ai_1 _1432_ (.B1(_0930_),
    .Y(_0042_),
    .A1(_0540_),
    .A2(net57));
 sg13g2_mux2_1 _1433_ (.A0(\i2c_bert.i2c.sclAndNor3.io_b ),
    .A1(\i2c_bert.i2c.sclAndNor3.io_c ),
    .S(net57),
    .X(_0043_));
 sg13g2_mux2_1 _1434_ (.A0(\i2c_bert.i2c.sclAndNor3.io_c ),
    .A1(\i2c_bert.i2c.sclAndNor5.io_d ),
    .S(net57),
    .X(_0044_));
 sg13g2_mux2_1 _1435_ (.A0(\i2c_bert.i2c.sclAndNor5.io_d ),
    .A1(\i2c_bert.i2c.sclAndNor5.io_e ),
    .S(net57),
    .X(_0045_));
 sg13g2_nand2_1 _1436_ (.Y(_0931_),
    .A(\i2c_bert.i2c.sdaAndNor3.io_b ),
    .B(net57));
 sg13g2_o21ai_1 _1437_ (.B1(_0931_),
    .Y(_0048_),
    .A1(_0573_),
    .A2(net57));
 sg13g2_nand2_1 _1438_ (.Y(_0932_),
    .A(net88),
    .B(net57));
 sg13g2_o21ai_1 _1439_ (.B1(_0932_),
    .Y(_0049_),
    .A1(_0567_),
    .A2(_0929_));
 sg13g2_mux2_1 _1440_ (.A0(net88),
    .A1(_0558_),
    .S(_0929_),
    .X(_0050_));
 sg13g2_mux2_1 _1441_ (.A0(_0558_),
    .A1(_0560_),
    .S(_0928_),
    .X(_0051_));
 sg13g2_nand2b_1 _1442_ (.Y(_0933_),
    .B(_0851_),
    .A_N(_0599_));
 sg13g2_a21oi_2 _1443_ (.B1(_0732_),
    .Y(_0934_),
    .A2(_0917_),
    .A1(_0730_));
 sg13g2_nand2b_1 _1444_ (.Y(_0935_),
    .B(_0934_),
    .A_N(_0855_));
 sg13g2_nand2_1 _1445_ (.Y(_0936_),
    .A(_0933_),
    .B(_0847_));
 sg13g2_nor2_1 _1446_ (.A(_0830_),
    .B(_0847_),
    .Y(_0937_));
 sg13g2_a221oi_1 _1447_ (.B2(net53),
    .C1(_0937_),
    .B1(_0936_),
    .A1(_0933_),
    .Y(_0938_),
    .A2(_0935_));
 sg13g2_buf_1 _1448_ (.A(_0938_),
    .X(_0939_));
 sg13g2_buf_1 _1449_ (.A(_0939_),
    .X(_0940_));
 sg13g2_buf_1 _1450_ (.A(\i2c_bert.myState_1.alu_1.acc[0] ),
    .X(_0941_));
 sg13g2_nor3_2 _1451_ (.A(_0026_),
    .B(_0617_),
    .C(_0674_),
    .Y(_0942_));
 sg13g2_nand2_1 _1452_ (.Y(_0943_),
    .A(_0614_),
    .B(_0942_));
 sg13g2_nand2_2 _1453_ (.Y(_0944_),
    .A(_0031_),
    .B(_0943_));
 sg13g2_nand2_1 _1454_ (.Y(_0945_),
    .A(_0631_),
    .B(_0674_));
 sg13g2_inv_1 _1455_ (.Y(_0946_),
    .A(_0031_));
 sg13g2_a21oi_2 _1456_ (.B1(_0946_),
    .Y(_0947_),
    .A2(_0945_),
    .A1(_0618_));
 sg13g2_mux2_1 _1457_ (.A0(\i2c_bert.myState_1.io_timerEndstop[0] ),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[0] ),
    .S(net67),
    .X(_0948_));
 sg13g2_a22oi_1 _1458_ (.Y(_0949_),
    .B1(_0947_),
    .B2(_0948_),
    .A2(_0944_),
    .A1(net95));
 sg13g2_nor3_2 _1459_ (.A(_0610_),
    .B(_0611_),
    .C(_0619_),
    .Y(_0950_));
 sg13g2_inv_1 _1460_ (.Y(_0951_),
    .A(net86));
 sg13g2_nor3_1 _1461_ (.A(_0951_),
    .B(_0611_),
    .C(_0619_),
    .Y(_0952_));
 sg13g2_buf_1 _1462_ (.A(_0952_),
    .X(_0953_));
 sg13g2_a22oi_1 _1463_ (.Y(_0954_),
    .B1(net56),
    .B2(\i2c_bert.myState_1.len12[4] ),
    .A2(_0950_),
    .A1(net90));
 sg13g2_and3_1 _1464_ (.X(_0955_),
    .A(net66),
    .B(_0710_),
    .C(_0942_));
 sg13g2_buf_1 _1465_ (.A(_0955_),
    .X(_0956_));
 sg13g2_nor2_2 _1466_ (.A(_0619_),
    .B(_0674_),
    .Y(_0957_));
 sg13g2_buf_2 _1467_ (.A(_0621_),
    .X(_0958_));
 sg13g2_mux4_1 _1468_ (.S0(net73),
    .A0(net90),
    .A1(\i2c_bert.div12[4] ),
    .A2(\i2c_bert.latched[16] ),
    .A3(\i2c_bert.latched[24] ),
    .S1(net69),
    .X(_0959_));
 sg13g2_a22oi_1 _1469_ (.Y(_0960_),
    .B1(_0957_),
    .B2(_0959_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[0] ));
 sg13g2_nand3_1 _1470_ (.B(_0954_),
    .C(_0960_),
    .A(_0949_),
    .Y(_0961_));
 sg13g2_nor2_2 _1471_ (.A(_0823_),
    .B(_0934_),
    .Y(_0962_));
 sg13g2_and2_1 _1472_ (.A(\i2c_bert.i2c.io_sdaSignal ),
    .B(_0962_),
    .X(_0963_));
 sg13g2_a221oi_1 _1473_ (.B2(_0961_),
    .C1(_0963_),
    .B1(_0934_),
    .A1(\i2c_bert.i2c.io_data8rx[7] ),
    .Y(_0964_),
    .A2(_0823_));
 sg13g2_nor2_1 _1474_ (.A(net75),
    .B(net48),
    .Y(_0965_));
 sg13g2_a21oi_1 _1475_ (.A1(net48),
    .A2(_0964_),
    .Y(_0052_),
    .B1(_0965_));
 sg13g2_buf_1 _1476_ (.A(\i2c_bert.myState_1.alu_1.acc[1] ),
    .X(_0966_));
 sg13g2_mux2_1 _1477_ (.A0(\i2c_bert.myState_1.io_timerEndstop[1] ),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[1] ),
    .S(net67),
    .X(_0967_));
 sg13g2_a22oi_1 _1478_ (.Y(_0968_),
    .B1(_0947_),
    .B2(_0967_),
    .A2(_0944_),
    .A1(net94));
 sg13g2_a22oi_1 _1479_ (.Y(_0969_),
    .B1(net56),
    .B2(\i2c_bert.myState_1.len12[5] ),
    .A2(_0950_),
    .A1(_0527_));
 sg13g2_mux4_1 _1480_ (.S0(net73),
    .A0(net91),
    .A1(\i2c_bert.div12[5] ),
    .A2(\i2c_bert.latched[17] ),
    .A3(\i2c_bert.latched[25] ),
    .S1(net69),
    .X(_0970_));
 sg13g2_a22oi_1 _1481_ (.Y(_0971_),
    .B1(_0957_),
    .B2(_0970_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[1] ));
 sg13g2_nand3_1 _1482_ (.B(_0969_),
    .C(_0971_),
    .A(_0968_),
    .Y(_0972_));
 sg13g2_nor2_1 _1483_ (.A(_0661_),
    .B(_0883_),
    .Y(_0973_));
 sg13g2_a221oi_1 _1484_ (.B2(_0934_),
    .C1(_0973_),
    .B1(_0972_),
    .A1(net75),
    .Y(_0974_),
    .A2(_0962_));
 sg13g2_nor2_1 _1485_ (.A(net82),
    .B(net48),
    .Y(_0975_));
 sg13g2_a21oi_1 _1486_ (.A1(net48),
    .A2(_0974_),
    .Y(_0053_),
    .B1(_0975_));
 sg13g2_buf_1 _1487_ (.A(\i2c_bert.myState_1.alu_1.acc[2] ),
    .X(_0976_));
 sg13g2_mux2_1 _1488_ (.A0(\i2c_bert.myState_1.io_timerEndstop[2] ),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[2] ),
    .S(net67),
    .X(_0977_));
 sg13g2_a22oi_1 _1489_ (.Y(_0978_),
    .B1(_0947_),
    .B2(_0977_),
    .A2(_0944_),
    .A1(net93));
 sg13g2_a22oi_1 _1490_ (.Y(_0979_),
    .B1(net56),
    .B2(\i2c_bert.myState_1.len12[6] ),
    .A2(_0950_),
    .A1(net89));
 sg13g2_mux4_1 _1491_ (.S0(net73),
    .A0(net89),
    .A1(\i2c_bert.div12[6] ),
    .A2(\i2c_bert.latched[18] ),
    .A3(\i2c_bert.latched[26] ),
    .S1(net69),
    .X(_0980_));
 sg13g2_a22oi_1 _1492_ (.Y(_0981_),
    .B1(_0957_),
    .B2(_0980_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[2] ));
 sg13g2_nand3_1 _1493_ (.B(_0979_),
    .C(_0981_),
    .A(_0978_),
    .Y(_0982_));
 sg13g2_nor2_1 _1494_ (.A(_0010_),
    .B(_0883_),
    .Y(_0983_));
 sg13g2_a221oi_1 _1495_ (.B2(_0934_),
    .C1(_0983_),
    .B1(_0982_),
    .A1(_0643_),
    .Y(_0984_),
    .A2(_0962_));
 sg13g2_nor2_1 _1496_ (.A(net63),
    .B(net48),
    .Y(_0985_));
 sg13g2_a21oi_1 _1497_ (.A1(net48),
    .A2(_0984_),
    .Y(_0054_),
    .B1(_0985_));
 sg13g2_mux2_1 _1498_ (.A0(\i2c_bert.myState_1.io_timerEndstop[3] ),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[3] ),
    .S(_0609_),
    .X(_0986_));
 sg13g2_a22oi_1 _1499_ (.Y(_0987_),
    .B1(_0947_),
    .B2(_0986_),
    .A2(_0944_),
    .A1(\i2c_bert.myState_1.alu_1.acc[3] ));
 sg13g2_buf_2 _1500_ (.A(\i2c_bert.i2c.io_pushPullMode ),
    .X(_0988_));
 sg13g2_a22oi_1 _1501_ (.Y(_0989_),
    .B1(net56),
    .B2(\i2c_bert.myState_1.len12[7] ),
    .A2(_0950_),
    .A1(_0988_));
 sg13g2_mux4_1 _1502_ (.S0(net73),
    .A0(_0988_),
    .A1(\i2c_bert.div12[7] ),
    .A2(\i2c_bert.latched[19] ),
    .A3(\i2c_bert.latched[27] ),
    .S1(net69),
    .X(_0990_));
 sg13g2_a22oi_1 _1503_ (.Y(_0991_),
    .B1(_0957_),
    .B2(_0990_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[3] ));
 sg13g2_nand3_1 _1504_ (.B(_0989_),
    .C(_0991_),
    .A(_0987_),
    .Y(_0992_));
 sg13g2_buf_2 _1505_ (.A(_0011_),
    .X(_0993_));
 sg13g2_nor2_1 _1506_ (.A(_0993_),
    .B(_0883_),
    .Y(_0994_));
 sg13g2_a221oi_1 _1507_ (.B2(_0934_),
    .C1(_0994_),
    .B1(_0992_),
    .A1(net63),
    .Y(_0995_),
    .A2(_0962_));
 sg13g2_nor2_1 _1508_ (.A(net81),
    .B(_0940_),
    .Y(_0996_));
 sg13g2_a21oi_1 _1509_ (.A1(_0940_),
    .A2(_0995_),
    .Y(_0055_),
    .B1(_0996_));
 sg13g2_o21ai_1 _1510_ (.B1(_0846_),
    .Y(_0997_),
    .A1(_0737_),
    .A2(_0789_));
 sg13g2_buf_1 _1511_ (.A(_0997_),
    .X(_0998_));
 sg13g2_nor2b_1 _1512_ (.A(_0609_),
    .B_N(_0947_),
    .Y(_0999_));
 sg13g2_buf_1 _1513_ (.A(\i2c_bert.myState_1.alu_1.acc[4] ),
    .X(_1000_));
 sg13g2_inv_1 _1514_ (.Y(_1001_),
    .A(net92));
 sg13g2_a21oi_2 _1515_ (.B1(_0946_),
    .Y(_1002_),
    .A2(_0942_),
    .A1(net65));
 sg13g2_mux4_1 _1516_ (.S0(net69),
    .A0(\i2c_bert.div12[0] ),
    .A1(\i2c_bert.latched[20] ),
    .A2(\i2c_bert.div12[8] ),
    .A3(\i2c_bert.latched[28] ),
    .S1(net73),
    .X(_1003_));
 sg13g2_a22oi_1 _1517_ (.Y(_1004_),
    .B1(_0957_),
    .B2(_1003_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[4] ));
 sg13g2_o21ai_1 _1518_ (.B1(_1004_),
    .Y(_1005_),
    .A1(_1001_),
    .A2(_1002_));
 sg13g2_a221oi_1 _1519_ (.B2(\i2c_bert.myState_1.io_timerEndstop[4] ),
    .C1(_1005_),
    .B1(_0999_),
    .A1(\i2c_bert.myState_1.len12[8] ),
    .Y(_1006_),
    .A2(net56));
 sg13g2_inv_1 _1520_ (.Y(_1007_),
    .A(_0012_));
 sg13g2_a22oi_1 _1521_ (.Y(_1008_),
    .B1(_0962_),
    .B2(net81),
    .A2(_0823_),
    .A1(_1007_));
 sg13g2_o21ai_1 _1522_ (.B1(_1008_),
    .Y(_1009_),
    .A1(_0998_),
    .A2(_1006_));
 sg13g2_mux2_1 _1523_ (.A0(_0649_),
    .A1(_1009_),
    .S(net48),
    .X(_0056_));
 sg13g2_buf_2 _1524_ (.A(\i2c_bert.myState_1.alu_1.acc[5] ),
    .X(_1010_));
 sg13g2_inv_2 _1525_ (.Y(_1011_),
    .A(_1010_));
 sg13g2_mux4_1 _1526_ (.S0(net69),
    .A0(\i2c_bert.div12[1] ),
    .A1(\i2c_bert.latched[21] ),
    .A2(\i2c_bert.div12[9] ),
    .A3(\i2c_bert.latched[29] ),
    .S1(net73),
    .X(_1012_));
 sg13g2_a22oi_1 _1527_ (.Y(_1013_),
    .B1(_0957_),
    .B2(_1012_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[5] ));
 sg13g2_o21ai_1 _1528_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1011_),
    .A2(_1002_));
 sg13g2_a221oi_1 _1529_ (.B2(\i2c_bert.myState_1.io_timerEndstop[5] ),
    .C1(_1014_),
    .B1(_0999_),
    .A1(\i2c_bert.myState_1.len12[9] ),
    .Y(_1015_),
    .A2(net56));
 sg13g2_buf_2 _1530_ (.A(_0013_),
    .X(_1016_));
 sg13g2_inv_1 _1531_ (.Y(_1017_),
    .A(_1016_));
 sg13g2_a22oi_1 _1532_ (.Y(_1018_),
    .B1(_0962_),
    .B2(net80),
    .A2(_0823_),
    .A1(_1017_));
 sg13g2_o21ai_1 _1533_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_0998_),
    .A2(_1015_));
 sg13g2_mux2_1 _1534_ (.A0(net84),
    .A1(_1019_),
    .S(net48),
    .X(_0057_));
 sg13g2_mux4_1 _1535_ (.S0(_0958_),
    .A0(\i2c_bert.div12[2] ),
    .A1(\i2c_bert.latched[22] ),
    .A2(\i2c_bert.div12[10] ),
    .A3(\i2c_bert.latched[30] ),
    .S1(_0768_),
    .X(_1020_));
 sg13g2_a22oi_1 _1536_ (.Y(_1021_),
    .B1(_0957_),
    .B2(_1020_),
    .A2(_0956_),
    .A1(\i2c_bert.myState_1.led8[6] ));
 sg13g2_o21ai_1 _1537_ (.B1(_1021_),
    .Y(_1022_),
    .A1(_0014_),
    .A2(_1002_));
 sg13g2_a221oi_1 _1538_ (.B2(\i2c_bert.myState_1.io_timerEndstop[6] ),
    .C1(_1022_),
    .B1(_0999_),
    .A1(\i2c_bert.myState_1.len12[10] ),
    .Y(_1023_),
    .A2(net56));
 sg13g2_buf_2 _1539_ (.A(_0015_),
    .X(_1024_));
 sg13g2_inv_1 _1540_ (.Y(_1025_),
    .A(_1024_));
 sg13g2_a22oi_1 _1541_ (.Y(_1026_),
    .B1(_0962_),
    .B2(net84),
    .A2(_0823_),
    .A1(_1025_));
 sg13g2_o21ai_1 _1542_ (.B1(_1026_),
    .Y(_1027_),
    .A1(_0998_),
    .A2(_1023_));
 sg13g2_mux2_1 _1543_ (.A0(net83),
    .A1(_1027_),
    .S(_0939_),
    .X(_0058_));
 sg13g2_mux4_1 _1544_ (.S0(_0958_),
    .A0(\i2c_bert.div12[3] ),
    .A1(\i2c_bert.latched[23] ),
    .A2(\i2c_bert.div12[11] ),
    .A3(\i2c_bert.latched[31] ),
    .S1(_0768_),
    .X(_1028_));
 sg13g2_a22oi_1 _1545_ (.Y(_1029_),
    .B1(_0957_),
    .B2(_1028_),
    .A2(net58),
    .A1(\i2c_bert.myState_1.led8[7] ));
 sg13g2_o21ai_1 _1546_ (.B1(_1029_),
    .Y(_1030_),
    .A1(_0016_),
    .A2(_1002_));
 sg13g2_a221oi_1 _1547_ (.B2(\i2c_bert.myState_1.io_timerEndstop[7] ),
    .C1(_1030_),
    .B1(_0999_),
    .A1(\i2c_bert.myState_1.len12[11] ),
    .Y(_1031_),
    .A2(_0953_));
 sg13g2_inv_1 _1548_ (.Y(_1032_),
    .A(_0009_));
 sg13g2_a22oi_1 _1549_ (.Y(_1033_),
    .B1(_0962_),
    .B2(_0641_),
    .A2(_0823_),
    .A1(_1032_));
 sg13g2_o21ai_1 _1550_ (.B1(_1033_),
    .Y(_1034_),
    .A1(_0998_),
    .A2(_1031_));
 sg13g2_mux2_1 _1551_ (.A0(\i2c_bert.i2c.io_data8rx[7] ),
    .A1(_1034_),
    .S(_0939_),
    .X(_0059_));
 sg13g2_nor2_1 _1552_ (.A(net62),
    .B(_0755_),
    .Y(_1035_));
 sg13g2_nor2b_1 _1553_ (.A(net62),
    .B_N(net79),
    .Y(_1036_));
 sg13g2_nand2_1 _1554_ (.Y(_1037_),
    .A(_0669_),
    .B(net50));
 sg13g2_o21ai_1 _1555_ (.B1(_1037_),
    .Y(_1038_),
    .A1(_0763_),
    .A2(_1036_));
 sg13g2_buf_1 _1556_ (.A(_1038_),
    .X(_1039_));
 sg13g2_mux2_1 _1557_ (.A0(_1035_),
    .A1(net85),
    .S(net47),
    .X(_0069_));
 sg13g2_nor2_1 _1558_ (.A(_0762_),
    .B(_0644_),
    .Y(_1040_));
 sg13g2_buf_1 _1559_ (.A(net66),
    .X(_1041_));
 sg13g2_mux2_1 _1560_ (.A0(_1040_),
    .A1(_1041_),
    .S(net47),
    .X(_0070_));
 sg13g2_nor3_1 _1561_ (.A(net62),
    .B(net63),
    .C(_1038_),
    .Y(_1042_));
 sg13g2_a21oi_1 _1562_ (.A1(_0710_),
    .A2(_1039_),
    .Y(_0071_),
    .B1(_1042_));
 sg13g2_nor2_1 _1563_ (.A(net62),
    .B(net81),
    .Y(_1043_));
 sg13g2_nand2_1 _1564_ (.Y(_1044_),
    .A(net86),
    .B(net47));
 sg13g2_o21ai_1 _1565_ (.B1(_1044_),
    .Y(_0072_),
    .A1(net47),
    .A2(_1043_));
 sg13g2_nor3_1 _1566_ (.A(net62),
    .B(net80),
    .C(_1038_),
    .Y(_1045_));
 sg13g2_a21oi_1 _1567_ (.A1(_0612_),
    .A2(_1039_),
    .Y(_0073_),
    .B1(_1045_));
 sg13g2_nor2_1 _1568_ (.A(net62),
    .B(net84),
    .Y(_1046_));
 sg13g2_nand2_1 _1569_ (.Y(_1047_),
    .A(\i2c_bert.myState_1.cmd7[5] ),
    .B(net47));
 sg13g2_o21ai_1 _1570_ (.B1(_1047_),
    .Y(_0074_),
    .A1(net47),
    .A2(_1046_));
 sg13g2_nor2_1 _1571_ (.A(net62),
    .B(net83),
    .Y(_1048_));
 sg13g2_nand2_1 _1572_ (.Y(_1049_),
    .A(\i2c_bert.myState_1.cmd7[6] ),
    .B(net47));
 sg13g2_o21ai_1 _1573_ (.B1(_1049_),
    .Y(_0075_),
    .A1(net47),
    .A2(_1048_));
 sg13g2_nor2_1 _1574_ (.A(net74),
    .B(net95),
    .Y(_1050_));
 sg13g2_a21oi_1 _1575_ (.A1(net74),
    .A2(\i2c_bert.powerOnSense.D ),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_nand3_1 _1576_ (.B(net55),
    .C(_0603_),
    .A(net87),
    .Y(_1052_));
 sg13g2_buf_2 _1577_ (.A(_1052_),
    .X(_1053_));
 sg13g2_nor3_1 _1578_ (.A(net75),
    .B(_0644_),
    .C(net63),
    .Y(_1054_));
 sg13g2_nand4_1 _1579_ (.B(_0655_),
    .C(_0754_),
    .A(_0663_),
    .Y(_1055_),
    .D(_1054_));
 sg13g2_nor2b_1 _1580_ (.A(net79),
    .B_N(_0606_),
    .Y(_1056_));
 sg13g2_o21ai_1 _1581_ (.B1(_1056_),
    .Y(_1057_),
    .A1(_0030_),
    .A2(net49));
 sg13g2_nand2_1 _1582_ (.Y(_1058_),
    .A(_1055_),
    .B(_1057_));
 sg13g2_o21ai_1 _1583_ (.B1(_1058_),
    .Y(_1059_),
    .A1(net58),
    .A2(_1053_));
 sg13g2_buf_1 _1584_ (.A(_1059_),
    .X(_1060_));
 sg13g2_mux2_1 _1585_ (.A0(_1051_),
    .A1(\i2c_bert.myState_1.led8[0] ),
    .S(net37),
    .X(_0088_));
 sg13g2_nand2_1 _1586_ (.Y(_1061_),
    .A(_0766_),
    .B(net75));
 sg13g2_nand2b_1 _1587_ (.Y(_1062_),
    .B(net94),
    .A_N(net68));
 sg13g2_and2_1 _1588_ (.A(_1061_),
    .B(_1062_),
    .X(_1063_));
 sg13g2_nand2_1 _1589_ (.Y(_1064_),
    .A(\i2c_bert.myState_1.led8[1] ),
    .B(net37));
 sg13g2_o21ai_1 _1590_ (.B1(_1064_),
    .Y(_0089_),
    .A1(net37),
    .A2(_1063_));
 sg13g2_nand2_1 _1591_ (.Y(_1065_),
    .A(net68),
    .B(_0643_));
 sg13g2_nand2b_1 _1592_ (.Y(_1066_),
    .B(net93),
    .A_N(net68));
 sg13g2_and2_1 _1593_ (.A(_1065_),
    .B(_1066_),
    .X(_1067_));
 sg13g2_nand2_1 _1594_ (.Y(_1068_),
    .A(\i2c_bert.myState_1.led8[2] ),
    .B(net37));
 sg13g2_o21ai_1 _1595_ (.B1(_1068_),
    .Y(_0090_),
    .A1(net37),
    .A2(_1067_));
 sg13g2_inv_1 _1596_ (.Y(_1069_),
    .A(\i2c_bert.myState_1.alu_1.acc[3] ));
 sg13g2_nand2_1 _1597_ (.Y(_1070_),
    .A(_0607_),
    .B(net63));
 sg13g2_o21ai_1 _1598_ (.B1(_1070_),
    .Y(_1071_),
    .A1(net74),
    .A2(_1069_));
 sg13g2_mux2_1 _1599_ (.A0(_1071_),
    .A1(\i2c_bert.myState_1.led8[3] ),
    .S(net37),
    .X(_0091_));
 sg13g2_nand2_1 _1600_ (.Y(_1072_),
    .A(net68),
    .B(_0646_));
 sg13g2_nand2b_1 _1601_ (.Y(_1073_),
    .B(net92),
    .A_N(_0607_));
 sg13g2_and2_1 _1602_ (.A(_1072_),
    .B(_1073_),
    .X(_1074_));
 sg13g2_nand2_1 _1603_ (.Y(_1075_),
    .A(\i2c_bert.myState_1.led8[4] ),
    .B(_1060_));
 sg13g2_o21ai_1 _1604_ (.B1(_1075_),
    .Y(_0092_),
    .A1(_1060_),
    .A2(_1074_));
 sg13g2_nand2_1 _1605_ (.Y(_1076_),
    .A(net68),
    .B(net80));
 sg13g2_o21ai_1 _1606_ (.B1(_1076_),
    .Y(_1077_),
    .A1(net74),
    .A2(_1011_));
 sg13g2_mux2_1 _1607_ (.A0(_1077_),
    .A1(\i2c_bert.myState_1.led8[5] ),
    .S(net37),
    .X(_0093_));
 sg13g2_buf_2 _1608_ (.A(\i2c_bert.myState_1.alu_1.acc[6] ),
    .X(_1078_));
 sg13g2_inv_1 _1609_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_nand2_1 _1610_ (.Y(_1080_),
    .A(net68),
    .B(net84));
 sg13g2_o21ai_1 _1611_ (.B1(_1080_),
    .Y(_1081_),
    .A1(net74),
    .A2(_1079_));
 sg13g2_mux2_1 _1612_ (.A0(_1081_),
    .A1(\i2c_bert.myState_1.led8[6] ),
    .S(net37),
    .X(_0094_));
 sg13g2_inv_2 _1613_ (.Y(_1082_),
    .A(\i2c_bert.myState_1.alu_1.acc[7] ));
 sg13g2_nand2_1 _1614_ (.Y(_1083_),
    .A(net68),
    .B(_0641_));
 sg13g2_o21ai_1 _1615_ (.B1(_1083_),
    .Y(_1084_),
    .A1(_0766_),
    .A2(_1082_));
 sg13g2_mux2_1 _1616_ (.A0(_1084_),
    .A1(\i2c_bert.myState_1.led8[7] ),
    .S(_1059_),
    .X(_0095_));
 sg13g2_nor4_1 _1617_ (.A(_0747_),
    .B(_0640_),
    .C(net83),
    .D(_0651_),
    .Y(_1085_));
 sg13g2_a21oi_1 _1618_ (.A1(_0663_),
    .A2(_0665_),
    .Y(_1086_),
    .B1(_1085_));
 sg13g2_a21oi_1 _1619_ (.A1(_0663_),
    .A2(_0648_),
    .Y(_1087_),
    .B1(net75));
 sg13g2_o21ai_1 _1620_ (.B1(_1087_),
    .Y(_1088_),
    .A1(net82),
    .A2(_1086_));
 sg13g2_nor2_1 _1621_ (.A(net75),
    .B(_0653_),
    .Y(_1089_));
 sg13g2_nor3_1 _1622_ (.A(_0640_),
    .B(_0009_),
    .C(_0651_),
    .Y(_1090_));
 sg13g2_nand4_1 _1623_ (.B(_0655_),
    .C(_0656_),
    .A(_0661_),
    .Y(_1091_),
    .D(_0657_));
 sg13g2_nor2_1 _1624_ (.A(net52),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_a221oi_1 _1625_ (.B2(_1090_),
    .C1(_1092_),
    .B1(_1089_),
    .A1(net52),
    .Y(_1093_),
    .A2(_1088_));
 sg13g2_inv_1 _1626_ (.Y(_1094_),
    .A(_1093_));
 sg13g2_xnor2_1 _1627_ (.Y(_1095_),
    .A(\i2c_bert.myState_1.len12[4] ),
    .B(net52));
 sg13g2_xnor2_1 _1628_ (.Y(_1096_),
    .A(\i2c_bert.myState_1.len12[10] ),
    .B(net84));
 sg13g2_xnor2_1 _1629_ (.Y(_1097_),
    .A(\i2c_bert.myState_1.len12[8] ),
    .B(net81));
 sg13g2_xnor2_1 _1630_ (.Y(_1098_),
    .A(\i2c_bert.myState_1.len12[9] ),
    .B(net80));
 sg13g2_xor2_1 _1631_ (.B(net75),
    .A(\i2c_bert.myState_1.len12[5] ),
    .X(_1099_));
 sg13g2_xor2_1 _1632_ (.B(net82),
    .A(\i2c_bert.myState_1.len12[6] ),
    .X(_1100_));
 sg13g2_xor2_1 _1633_ (.B(net83),
    .A(\i2c_bert.myState_1.len12[11] ),
    .X(_1101_));
 sg13g2_xor2_1 _1634_ (.B(net63),
    .A(\i2c_bert.myState_1.len12[7] ),
    .X(_1102_));
 sg13g2_nand4_1 _1635_ (.B(_1100_),
    .C(_1101_),
    .A(_1099_),
    .Y(_1103_),
    .D(_1102_));
 sg13g2_nor4_1 _1636_ (.A(_1096_),
    .B(_1097_),
    .C(_1098_),
    .D(_1103_),
    .Y(_1104_));
 sg13g2_nand3b_1 _1637_ (.B(_1095_),
    .C(_1104_),
    .Y(_1105_),
    .A_N(_0950_));
 sg13g2_nand3_1 _1638_ (.B(_0632_),
    .C(_1105_),
    .A(net74),
    .Y(_1106_));
 sg13g2_o21ai_1 _1639_ (.B1(_1106_),
    .Y(_1107_),
    .A1(net74),
    .A2(_1094_));
 sg13g2_nor3_1 _1640_ (.A(_0767_),
    .B(_0628_),
    .C(_1053_),
    .Y(_1108_));
 sg13g2_nor2b_1 _1641_ (.A(net73),
    .B_N(_0629_),
    .Y(_1109_));
 sg13g2_nor2_1 _1642_ (.A(_0031_),
    .B(_0705_),
    .Y(_1110_));
 sg13g2_nor3_1 _1643_ (.A(_0772_),
    .B(_1109_),
    .C(_1110_),
    .Y(_1111_));
 sg13g2_a21oi_1 _1644_ (.A1(net49),
    .A2(_1111_),
    .Y(_1112_),
    .B1(_0030_));
 sg13g2_nor2_1 _1645_ (.A(_1108_),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_nand4_1 _1646_ (.B(_1037_),
    .C(_1055_),
    .A(_0726_),
    .Y(_1114_),
    .D(_1113_));
 sg13g2_mux2_1 _1647_ (.A0(_1107_),
    .A1(\i2c_bert.myState_1.readWriteBit ),
    .S(_1114_),
    .X(_0104_));
 sg13g2_nand4_1 _1648_ (.B(_0608_),
    .C(net49),
    .A(net87),
    .Y(_1115_),
    .D(_0629_));
 sg13g2_buf_2 _1649_ (.A(_1115_),
    .X(_1116_));
 sg13g2_nor2_1 _1650_ (.A(_0785_),
    .B(net70),
    .Y(_1117_));
 sg13g2_nand3_1 _1651_ (.B(_0789_),
    .C(_0860_),
    .A(_1117_),
    .Y(_1118_));
 sg13g2_buf_2 _1652_ (.A(_1118_),
    .X(_1119_));
 sg13g2_and3_1 _1653_ (.X(_1120_),
    .A(_0583_),
    .B(_1116_),
    .C(_1119_));
 sg13g2_buf_1 _1654_ (.A(_1120_),
    .X(_1121_));
 sg13g2_buf_1 _1655_ (.A(_1121_),
    .X(_1122_));
 sg13g2_buf_1 _1656_ (.A(_1119_),
    .X(_1123_));
 sg13g2_buf_1 _1657_ (.A(_1119_),
    .X(_1124_));
 sg13g2_buf_1 _1658_ (.A(_1116_),
    .X(_1125_));
 sg13g2_buf_1 _1659_ (.A(_1116_),
    .X(_1126_));
 sg13g2_nand2_1 _1660_ (.Y(_1127_),
    .A(\i2c_bert.div12[0] ),
    .B(_1126_));
 sg13g2_o21ai_1 _1661_ (.B1(_1127_),
    .Y(_1128_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[0] ),
    .A2(net44));
 sg13g2_nand2_1 _1662_ (.Y(_1129_),
    .A(net45),
    .B(_1128_));
 sg13g2_o21ai_1 _1663_ (.B1(_1129_),
    .Y(_1130_),
    .A1(_0808_),
    .A2(net46));
 sg13g2_nand2_1 _1664_ (.Y(_1131_),
    .A(\i2c_bert.myState_1.io_timerEndstop[0] ),
    .B(net36));
 sg13g2_o21ai_1 _1665_ (.B1(_1131_),
    .Y(_0105_),
    .A1(net36),
    .A2(_1130_));
 sg13g2_nand2_1 _1666_ (.Y(_1132_),
    .A(\i2c_bert.div12[10] ),
    .B(net43));
 sg13g2_o21ai_1 _1667_ (.B1(_1132_),
    .Y(_1133_),
    .A1(net82),
    .A2(net44));
 sg13g2_nor2_1 _1668_ (.A(\i2c_bert.timer_1.ticker_count[10] ),
    .B(_1119_),
    .Y(_1134_));
 sg13g2_a21oi_1 _1669_ (.A1(_1123_),
    .A2(_1133_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_buf_1 _1670_ (.A(_1121_),
    .X(_1136_));
 sg13g2_mux2_1 _1671_ (.A0(_1135_),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[2] ),
    .S(net35),
    .X(_0106_));
 sg13g2_nand2_1 _1672_ (.Y(_1137_),
    .A(\i2c_bert.div12[11] ),
    .B(net43));
 sg13g2_o21ai_1 _1673_ (.B1(_1137_),
    .Y(_1138_),
    .A1(net63),
    .A2(net44));
 sg13g2_nor2_1 _1674_ (.A(\i2c_bert.timer_1.ticker_count[11] ),
    .B(_1119_),
    .Y(_1139_));
 sg13g2_a21oi_1 _1675_ (.A1(net45),
    .A2(_1138_),
    .Y(_1140_),
    .B1(_1139_));
 sg13g2_mux2_1 _1676_ (.A0(_1140_),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[3] ),
    .S(net35),
    .X(_0107_));
 sg13g2_nand2_1 _1677_ (.Y(_1141_),
    .A(\i2c_bert.div12[1] ),
    .B(net43));
 sg13g2_o21ai_1 _1678_ (.B1(_1141_),
    .Y(_1142_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[1] ),
    .A2(net44));
 sg13g2_nand2_1 _1679_ (.Y(_1143_),
    .A(net45),
    .B(_1142_));
 sg13g2_o21ai_1 _1680_ (.B1(_1143_),
    .Y(_1144_),
    .A1(_0813_),
    .A2(net46));
 sg13g2_nand2_1 _1681_ (.Y(_1145_),
    .A(\i2c_bert.myState_1.io_timerEndstop[1] ),
    .B(_1136_));
 sg13g2_o21ai_1 _1682_ (.B1(_1145_),
    .Y(_0108_),
    .A1(_1122_),
    .A2(_1144_));
 sg13g2_nand2_1 _1683_ (.Y(_1146_),
    .A(\i2c_bert.div12[2] ),
    .B(_1126_));
 sg13g2_o21ai_1 _1684_ (.B1(_1146_),
    .Y(_1147_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[2] ),
    .A2(net44));
 sg13g2_nand2_1 _1685_ (.Y(_1148_),
    .A(net45),
    .B(_1147_));
 sg13g2_o21ai_1 _1686_ (.B1(_1148_),
    .Y(_1149_),
    .A1(\i2c_bert.timer_1.ticker_count[2] ),
    .A2(net46));
 sg13g2_nand2_1 _1687_ (.Y(_1150_),
    .A(\i2c_bert.myState_1.io_timerEndstop[2] ),
    .B(net35));
 sg13g2_o21ai_1 _1688_ (.B1(_1150_),
    .Y(_0109_),
    .A1(net36),
    .A2(_1149_));
 sg13g2_nand2_1 _1689_ (.Y(_1151_),
    .A(\i2c_bert.div12[3] ),
    .B(net43));
 sg13g2_o21ai_1 _1690_ (.B1(_1151_),
    .Y(_1152_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[3] ),
    .A2(net44));
 sg13g2_nand2_1 _1691_ (.Y(_1153_),
    .A(net45),
    .B(_1152_));
 sg13g2_o21ai_1 _1692_ (.B1(_1153_),
    .Y(_1154_),
    .A1(\i2c_bert.timer_1.ticker_count[3] ),
    .A2(net46));
 sg13g2_nand2_1 _1693_ (.Y(_1155_),
    .A(\i2c_bert.myState_1.io_timerEndstop[3] ),
    .B(net35));
 sg13g2_o21ai_1 _1694_ (.B1(_1155_),
    .Y(_0110_),
    .A1(net36),
    .A2(_1154_));
 sg13g2_nand2_1 _1695_ (.Y(_1156_),
    .A(\i2c_bert.div12[4] ),
    .B(_1116_));
 sg13g2_o21ai_1 _1696_ (.B1(_1156_),
    .Y(_1157_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[4] ),
    .A2(_1125_));
 sg13g2_nand2_1 _1697_ (.Y(_1158_),
    .A(net45),
    .B(_1157_));
 sg13g2_o21ai_1 _1698_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_0805_),
    .A2(net46));
 sg13g2_nand2_1 _1699_ (.Y(_1160_),
    .A(\i2c_bert.myState_1.io_timerEndstop[4] ),
    .B(net35));
 sg13g2_o21ai_1 _1700_ (.B1(_1160_),
    .Y(_0111_),
    .A1(net36),
    .A2(_1159_));
 sg13g2_nand2_1 _1701_ (.Y(_1161_),
    .A(\i2c_bert.div12[5] ),
    .B(_1116_));
 sg13g2_o21ai_1 _1702_ (.B1(_1161_),
    .Y(_1162_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[5] ),
    .A2(_1125_));
 sg13g2_nand2_1 _1703_ (.Y(_1163_),
    .A(_1124_),
    .B(_1162_));
 sg13g2_o21ai_1 _1704_ (.B1(_1163_),
    .Y(_1164_),
    .A1(_0811_),
    .A2(net46));
 sg13g2_nand2_1 _1705_ (.Y(_1165_),
    .A(\i2c_bert.myState_1.io_timerEndstop[5] ),
    .B(net35));
 sg13g2_o21ai_1 _1706_ (.B1(_1165_),
    .Y(_0112_),
    .A1(net36),
    .A2(_1164_));
 sg13g2_nand2_1 _1707_ (.Y(_1166_),
    .A(\i2c_bert.div12[6] ),
    .B(_1116_));
 sg13g2_o21ai_1 _1708_ (.B1(_1166_),
    .Y(_1167_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[6] ),
    .A2(net43));
 sg13g2_nand2_1 _1709_ (.Y(_0137_),
    .A(net45),
    .B(_1167_));
 sg13g2_o21ai_1 _1710_ (.B1(_0137_),
    .Y(_0138_),
    .A1(\i2c_bert.timer_1.ticker_count[6] ),
    .A2(net46));
 sg13g2_nand2_1 _1711_ (.Y(_0139_),
    .A(\i2c_bert.myState_1.io_timerEndstop[6] ),
    .B(_1136_));
 sg13g2_o21ai_1 _1712_ (.B1(_0139_),
    .Y(_0113_),
    .A1(_1122_),
    .A2(_0138_));
 sg13g2_nand2_1 _1713_ (.Y(_0140_),
    .A(\i2c_bert.div12[7] ),
    .B(_1116_));
 sg13g2_o21ai_1 _1714_ (.B1(_0140_),
    .Y(_0141_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[7] ),
    .A2(net43));
 sg13g2_nand2_1 _1715_ (.Y(_0142_),
    .A(_1124_),
    .B(_0141_));
 sg13g2_o21ai_1 _1716_ (.B1(_0142_),
    .Y(_0143_),
    .A1(\i2c_bert.timer_1.ticker_count[7] ),
    .A2(_1123_));
 sg13g2_nand2_1 _1717_ (.Y(_0144_),
    .A(\i2c_bert.myState_1.io_timerEndstop[7] ),
    .B(net35));
 sg13g2_o21ai_1 _1718_ (.B1(_0144_),
    .Y(_0114_),
    .A1(net36),
    .A2(_0143_));
 sg13g2_nand3b_1 _1719_ (.B(net43),
    .C(_0582_),
    .Y(_0145_),
    .A_N(\i2c_bert.div12[8] ));
 sg13g2_o21ai_1 _1720_ (.B1(_0145_),
    .Y(_0146_),
    .A1(net52),
    .A2(net44));
 sg13g2_mux2_1 _1721_ (.A0(_0798_),
    .A1(_0146_),
    .S(_1119_),
    .X(_0147_));
 sg13g2_a21o_1 _1722_ (.A2(net36),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[0] ),
    .B1(_0147_),
    .X(_0115_));
 sg13g2_nand2_1 _1723_ (.Y(_0148_),
    .A(\i2c_bert.div12[9] ),
    .B(net43));
 sg13g2_o21ai_1 _1724_ (.B1(_0148_),
    .Y(_0149_),
    .A1(_0750_),
    .A2(net44));
 sg13g2_nor2_1 _1725_ (.A(_0796_),
    .B(_1119_),
    .Y(_0150_));
 sg13g2_a21oi_1 _1726_ (.A1(net45),
    .A2(_0149_),
    .Y(_0151_),
    .B1(_0150_));
 sg13g2_mux2_1 _1727_ (.A0(_0151_),
    .A1(\i2c_bert.myState_1._zz__zz_io_data8tx[1] ),
    .S(net35),
    .X(_0116_));
 sg13g2_nand2b_1 _1728_ (.Y(_0152_),
    .B(_1109_),
    .A_N(_1053_));
 sg13g2_buf_1 _1729_ (.A(_0152_),
    .X(_0153_));
 sg13g2_nand2_1 _1730_ (.Y(_0154_),
    .A(\i2c_bert.timer_1.ticker_endstopTmpL[0] ),
    .B(net42));
 sg13g2_o21ai_1 _1731_ (.B1(_0154_),
    .Y(_0129_),
    .A1(\i2c_bert.powerOnSense.D ),
    .A2(net42));
 sg13g2_nand2_1 _1732_ (.Y(_0155_),
    .A(\i2c_bert.timer_1.ticker_endstopTmpL[1] ),
    .B(net42));
 sg13g2_o21ai_1 _1733_ (.B1(_0155_),
    .Y(_0130_),
    .A1(_0755_),
    .A2(net42));
 sg13g2_nand2_1 _1734_ (.Y(_0156_),
    .A(\i2c_bert.timer_1.ticker_endstopTmpL[2] ),
    .B(net42));
 sg13g2_o21ai_1 _1735_ (.B1(_0156_),
    .Y(_0131_),
    .A1(_0644_),
    .A2(net42));
 sg13g2_mux2_1 _1736_ (.A0(_0747_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[3] ),
    .S(net42),
    .X(_0132_));
 sg13g2_mux2_1 _1737_ (.A0(net81),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[4] ),
    .S(net42),
    .X(_0133_));
 sg13g2_mux2_1 _1738_ (.A0(_0649_),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[5] ),
    .S(_0153_),
    .X(_0134_));
 sg13g2_mux2_1 _1739_ (.A0(net84),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[6] ),
    .S(_0153_),
    .X(_0135_));
 sg13g2_mux2_1 _1740_ (.A0(net83),
    .A1(\i2c_bert.timer_1.ticker_endstopTmpL[7] ),
    .S(_0152_),
    .X(_0136_));
 sg13g2_nand2_1 _1741_ (.Y(_0157_),
    .A(_0829_),
    .B(_0937_));
 sg13g2_nand2b_1 _1742_ (.Y(_0158_),
    .B(_0998_),
    .A_N(_0590_));
 sg13g2_o21ai_1 _1743_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_0539_),
    .A2(_0847_));
 sg13g2_nand2_1 _1744_ (.Y(_0160_),
    .A(_0742_),
    .B(_0159_));
 sg13g2_a21o_1 _1745_ (.A2(_0825_),
    .A1(_0602_),
    .B1(_0158_),
    .X(_0161_));
 sg13g2_nand4_1 _1746_ (.B(_0157_),
    .C(_0160_),
    .A(_0868_),
    .Y(_0162_),
    .D(_0161_));
 sg13g2_buf_1 _1747_ (.A(_0162_),
    .X(_0163_));
 sg13g2_nand2b_1 _1748_ (.Y(_0164_),
    .B(_0825_),
    .A_N(_0163_));
 sg13g2_nand2_1 _1749_ (.Y(_0165_),
    .A(_0600_),
    .B(_0163_));
 sg13g2_o21ai_1 _1750_ (.B1(_0165_),
    .Y(_0166_),
    .A1(_0600_),
    .A2(_0164_));
 sg13g2_nand2_1 _1751_ (.Y(_0167_),
    .A(_1117_),
    .B(_0789_));
 sg13g2_a221oi_1 _1752_ (.B2(_0913_),
    .C1(_0901_),
    .B1(_0920_),
    .A1(_0868_),
    .Y(_0168_),
    .A2(_0916_));
 sg13g2_nand4_1 _1753_ (.B(_0877_),
    .C(_0167_),
    .A(_0845_),
    .Y(_0169_),
    .D(_0168_));
 sg13g2_and2_1 _1754_ (.A(_0166_),
    .B(_0169_),
    .X(_0032_));
 sg13g2_nand2b_1 _1755_ (.Y(_0170_),
    .B(_0600_),
    .A_N(\i2c_bert.i2c.fsm_bitCount[1] ));
 sg13g2_nor2_1 _1756_ (.A(_0600_),
    .B(_0914_),
    .Y(_0171_));
 sg13g2_o21ai_1 _1757_ (.B1(\i2c_bert.i2c.fsm_bitCount[1] ),
    .Y(_0172_),
    .A1(_0163_),
    .A2(_0171_));
 sg13g2_o21ai_1 _1758_ (.B1(_0172_),
    .Y(_0173_),
    .A1(_0164_),
    .A2(_0170_));
 sg13g2_and2_1 _1759_ (.A(_0169_),
    .B(_0173_),
    .X(_0033_));
 sg13g2_nand2_1 _1760_ (.Y(_0174_),
    .A(\i2c_bert.i2c.fsm_bitCount[1] ),
    .B(_0600_));
 sg13g2_nand2_1 _1761_ (.Y(_0175_),
    .A(_0018_),
    .B(_0174_));
 sg13g2_nand3_1 _1762_ (.B(_0825_),
    .C(_0175_),
    .A(_0602_),
    .Y(_0176_));
 sg13g2_nand2_1 _1763_ (.Y(_0177_),
    .A(\i2c_bert.i2c.fsm_bitCount[2] ),
    .B(_0163_));
 sg13g2_o21ai_1 _1764_ (.B1(_0177_),
    .Y(_0178_),
    .A1(_0163_),
    .A2(_0176_));
 sg13g2_and2_1 _1765_ (.A(_0169_),
    .B(_0178_),
    .X(_0034_));
 sg13g2_nand2_1 _1766_ (.Y(_0179_),
    .A(_0877_),
    .B(_0901_));
 sg13g2_nor4_1 _1767_ (.A(_0582_),
    .B(_0038_),
    .C(_0845_),
    .D(_0179_),
    .Y(_0039_));
 sg13g2_inv_1 _1768_ (.Y(_0180_),
    .A(\i2c_bert.i2c.sclAndNor3.io_o ));
 sg13g2_o21ai_1 _1769_ (.B1(_0539_),
    .Y(_0181_),
    .A1(\i2c_bert.i2c.sclAndNor3.io_o ),
    .A2(_0534_));
 sg13g2_o21ai_1 _1770_ (.B1(_0181_),
    .Y(_0040_),
    .A1(_0180_),
    .A2(_0542_));
 sg13g2_nand2_1 _1771_ (.Y(_0182_),
    .A(\i2c_bert.i2c.io_timerAutobaud ),
    .B(net46));
 sg13g2_nand2b_1 _1772_ (.Y(_0183_),
    .B(_0583_),
    .A_N(_0818_));
 sg13g2_a21oi_1 _1773_ (.A1(_0169_),
    .A2(_0182_),
    .Y(_0060_),
    .B1(_0183_));
 sg13g2_nor3_1 _1774_ (.A(net66),
    .B(_0943_),
    .C(_1053_),
    .Y(_0184_));
 sg13g2_buf_1 _1775_ (.A(_0184_),
    .X(_0185_));
 sg13g2_a21oi_1 _1776_ (.A1(_0552_),
    .A2(_0553_),
    .Y(_0186_),
    .B1(\i2c_bert.i2c.scl_regNext ));
 sg13g2_nand3_1 _1777_ (.B(_0613_),
    .C(_0614_),
    .A(net87),
    .Y(_0187_));
 sg13g2_inv_1 _1778_ (.Y(_0188_),
    .A(_0187_));
 sg13g2_nand4_1 _1779_ (.B(_0603_),
    .C(_0942_),
    .A(_0186_),
    .Y(_0189_),
    .D(_0188_));
 sg13g2_a21o_1 _1780_ (.A2(_0551_),
    .A1(_0538_),
    .B1(_0189_),
    .X(_0190_));
 sg13g2_buf_2 _1781_ (.A(_0190_),
    .X(_0191_));
 sg13g2_buf_8 _1782_ (.A(_0191_),
    .X(_0192_));
 sg13g2_nand2_2 _1783_ (.Y(_0193_),
    .A(net52),
    .B(net51));
 sg13g2_nor2_2 _1784_ (.A(_1002_),
    .B(_1053_),
    .Y(_0194_));
 sg13g2_nand2b_1 _1785_ (.Y(_0195_),
    .B(_0194_),
    .A_N(_0193_));
 sg13g2_o21ai_1 _1786_ (.B1(_0195_),
    .Y(_0196_),
    .A1(net95),
    .A2(_0185_));
 sg13g2_or3_1 _1787_ (.A(net66),
    .B(_0943_),
    .C(_1053_),
    .X(_0197_));
 sg13g2_buf_1 _1788_ (.A(_0197_),
    .X(_0198_));
 sg13g2_nand3_1 _1789_ (.B(net95),
    .C(_0193_),
    .A(net65),
    .Y(_0199_));
 sg13g2_nand2b_1 _1790_ (.Y(_0200_),
    .B(net40),
    .A_N(_0199_));
 sg13g2_o21ai_1 _1791_ (.B1(_0200_),
    .Y(_0201_),
    .A1(_0193_),
    .A2(net40));
 sg13g2_a21oi_1 _1792_ (.A1(_0193_),
    .A2(_0194_),
    .Y(_0202_),
    .B1(net95));
 sg13g2_nand4_1 _1793_ (.B(_0581_),
    .C(net55),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[2] ),
    .Y(_0203_),
    .D(_0603_));
 sg13g2_nand3_1 _1794_ (.B(_0648_),
    .C(_1089_),
    .A(_0663_),
    .Y(_0204_));
 sg13g2_nor2_1 _1795_ (.A(_0203_),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_nor2_2 _1796_ (.A(_0582_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_nand2b_1 _1797_ (.Y(_0207_),
    .B(_0206_),
    .A_N(_0202_));
 sg13g2_a221oi_1 _1798_ (.B2(_0194_),
    .C1(_0207_),
    .B1(_0201_),
    .A1(_0615_),
    .Y(_0061_),
    .A2(_0196_));
 sg13g2_buf_1 _1799_ (.A(net65),
    .X(_0208_));
 sg13g2_nand3_1 _1800_ (.B(net95),
    .C(_0193_),
    .A(net66),
    .Y(_0209_));
 sg13g2_a21oi_1 _1801_ (.A1(_0538_),
    .A2(_0551_),
    .Y(_0210_),
    .B1(_0189_));
 sg13g2_buf_1 _1802_ (.A(_0210_),
    .X(_0211_));
 sg13g2_nor2_2 _1803_ (.A(_0661_),
    .B(net54),
    .Y(_0212_));
 sg13g2_xnor2_1 _1804_ (.Y(_0213_),
    .A(net94),
    .B(_0212_));
 sg13g2_nand4_1 _1805_ (.B(net40),
    .C(_0212_),
    .A(net94),
    .Y(_0214_),
    .D(_0209_));
 sg13g2_o21ai_1 _1806_ (.B1(_0214_),
    .Y(_0215_),
    .A1(_0209_),
    .A2(_0213_));
 sg13g2_a21o_1 _1807_ (.A2(_0212_),
    .A1(net94),
    .B1(net65),
    .X(_0216_));
 sg13g2_o21ai_1 _1808_ (.B1(_0216_),
    .Y(_0217_),
    .A1(net94),
    .A2(_0212_));
 sg13g2_nand2b_1 _1809_ (.Y(_0218_),
    .B(_0199_),
    .A_N(net94));
 sg13g2_a21oi_1 _1810_ (.A1(net40),
    .A2(_0218_),
    .Y(_0219_),
    .B1(_0212_));
 sg13g2_a221oi_1 _1811_ (.B2(_0634_),
    .C1(_0219_),
    .B1(_0217_),
    .A1(net60),
    .Y(_0220_),
    .A2(_0215_));
 sg13g2_nand2_1 _1812_ (.Y(_0221_),
    .A(_0194_),
    .B(_0220_));
 sg13g2_nand2b_1 _1813_ (.Y(_0222_),
    .B(_0944_),
    .A_N(_1053_));
 sg13g2_buf_1 _1814_ (.A(_0222_),
    .X(_0223_));
 sg13g2_nand2_1 _1815_ (.Y(_0224_),
    .A(_0966_),
    .B(net39));
 sg13g2_o21ai_1 _1816_ (.B1(_0583_),
    .Y(_0225_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_a21oi_1 _1817_ (.A1(_0221_),
    .A2(_0224_),
    .Y(_0062_),
    .B1(_0225_));
 sg13g2_nand2_1 _1818_ (.Y(_0226_),
    .A(_0538_),
    .B(_0551_));
 sg13g2_inv_1 _1819_ (.Y(_0227_),
    .A(_0189_));
 sg13g2_o21ai_1 _1820_ (.B1(_0941_),
    .Y(_0228_),
    .A1(_0566_),
    .A2(_0579_));
 sg13g2_nand2_1 _1821_ (.Y(_0229_),
    .A(net14),
    .B(\i2c_bert.myState_1.alu_1.acc[0] ));
 sg13g2_a21oi_1 _1822_ (.A1(_0568_),
    .A2(_0572_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_nor2_1 _1823_ (.A(\i2c_bert.myState_1.alu_1.acc[1] ),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_a221oi_1 _1824_ (.B2(_0231_),
    .C1(_0661_),
    .B1(_0228_),
    .A1(_0226_),
    .Y(_0232_),
    .A2(_0227_));
 sg13g2_buf_2 _1825_ (.A(_0232_),
    .X(_0233_));
 sg13g2_nand2_1 _1826_ (.Y(_0234_),
    .A(net95),
    .B(\i2c_bert.myState_1.alu_1.acc[1] ));
 sg13g2_a21oi_2 _1827_ (.B1(_0234_),
    .Y(_0235_),
    .A2(_0191_),
    .A1(_0581_));
 sg13g2_or2_1 _1828_ (.X(_0236_),
    .B(_0235_),
    .A(_0233_));
 sg13g2_nand2_1 _1829_ (.Y(_0237_),
    .A(net61),
    .B(_0236_));
 sg13g2_inv_1 _1830_ (.Y(_0238_),
    .A(_0010_));
 sg13g2_nand2_1 _1831_ (.Y(_0239_),
    .A(_0238_),
    .B(_0192_));
 sg13g2_nor2_1 _1832_ (.A(net41),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_nand4_1 _1833_ (.B(net93),
    .C(_0237_),
    .A(_0208_),
    .Y(_0241_),
    .D(_0240_));
 sg13g2_mux2_1 _1834_ (.A0(_0240_),
    .A1(_0239_),
    .S(net93),
    .X(_0242_));
 sg13g2_nand4_1 _1835_ (.B(_0208_),
    .C(_0236_),
    .A(net61),
    .Y(_0243_),
    .D(_0242_));
 sg13g2_and2_1 _1836_ (.A(net65),
    .B(_0236_),
    .X(_0244_));
 sg13g2_o21ai_1 _1837_ (.B1(_0198_),
    .Y(_0245_),
    .A1(net93),
    .A2(_0244_));
 sg13g2_and3_1 _1838_ (.X(_0246_),
    .A(\i2c_bert.myState_1.alu_1.acc[2] ),
    .B(_0238_),
    .C(_0191_));
 sg13g2_nand2b_1 _1839_ (.Y(_0247_),
    .B(_0239_),
    .A_N(net93));
 sg13g2_o21ai_1 _1840_ (.B1(_0247_),
    .Y(_0248_),
    .A1(net65),
    .A2(_0246_));
 sg13g2_a22oi_1 _1841_ (.Y(_0249_),
    .B1(_0248_),
    .B2(_0634_),
    .A2(_0245_),
    .A1(_0239_));
 sg13g2_nand4_1 _1842_ (.B(_0241_),
    .C(_0243_),
    .A(_0194_),
    .Y(_0250_),
    .D(_0249_));
 sg13g2_nand2_1 _1843_ (.Y(_0251_),
    .A(_0976_),
    .B(net39));
 sg13g2_a21oi_1 _1844_ (.A1(_0250_),
    .A2(_0251_),
    .Y(_0063_),
    .B1(_0225_));
 sg13g2_or3_1 _1845_ (.A(_0233_),
    .B(_0235_),
    .C(_0246_),
    .X(_0252_));
 sg13g2_and2_1 _1846_ (.A(_0247_),
    .B(_0252_),
    .X(_0253_));
 sg13g2_nor3_2 _1847_ (.A(_1069_),
    .B(_0993_),
    .C(net54),
    .Y(_0254_));
 sg13g2_a21o_1 _1848_ (.A2(_0253_),
    .A1(net61),
    .B1(_0254_),
    .X(_0255_));
 sg13g2_nor2_2 _1849_ (.A(_0993_),
    .B(_0210_),
    .Y(_0256_));
 sg13g2_xnor2_1 _1850_ (.Y(_0257_),
    .A(\i2c_bert.myState_1.alu_1.acc[3] ),
    .B(_0256_));
 sg13g2_nand3_1 _1851_ (.B(_0253_),
    .C(_0257_),
    .A(_1041_),
    .Y(_0258_));
 sg13g2_nand3_1 _1852_ (.B(_0255_),
    .C(_0258_),
    .A(net60),
    .Y(_0259_));
 sg13g2_o21ai_1 _1853_ (.B1(_1069_),
    .Y(_0260_),
    .A1(_0993_),
    .A2(net54));
 sg13g2_o21ai_1 _1854_ (.B1(_0260_),
    .Y(_0261_),
    .A1(net60),
    .A2(_0254_));
 sg13g2_nand2_1 _1855_ (.Y(_0262_),
    .A(_0194_),
    .B(net40));
 sg13g2_a21oi_1 _1856_ (.A1(_0634_),
    .A2(_0261_),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_a21o_1 _1857_ (.A2(_0253_),
    .A1(net60),
    .B1(_0260_),
    .X(_0264_));
 sg13g2_nand3_1 _1858_ (.B(_0263_),
    .C(_0264_),
    .A(_0259_),
    .Y(_0265_));
 sg13g2_a22oi_1 _1859_ (.Y(_0266_),
    .B1(net41),
    .B2(_0256_),
    .A2(net39),
    .A1(\i2c_bert.myState_1.alu_1.acc[3] ));
 sg13g2_a21oi_1 _1860_ (.A1(_0265_),
    .A2(_0266_),
    .Y(_0064_),
    .B1(_0225_));
 sg13g2_a21oi_1 _1861_ (.A1(_1007_),
    .A2(_0191_),
    .Y(_0267_),
    .B1(net92));
 sg13g2_and3_1 _1862_ (.X(_0268_),
    .A(_0247_),
    .B(_0252_),
    .C(_0260_));
 sg13g2_o21ai_1 _1863_ (.B1(net60),
    .Y(_0269_),
    .A1(_0254_),
    .A2(_0268_));
 sg13g2_nand2_1 _1864_ (.Y(_0270_),
    .A(_0267_),
    .B(_0269_));
 sg13g2_nor2_1 _1865_ (.A(_1001_),
    .B(_0012_),
    .Y(_0271_));
 sg13g2_a21oi_1 _1866_ (.A1(net51),
    .A2(_0271_),
    .Y(_0272_),
    .B1(net60));
 sg13g2_o21ai_1 _1867_ (.B1(_0634_),
    .Y(_0273_),
    .A1(_0267_),
    .A2(_0272_));
 sg13g2_nand2_1 _1868_ (.Y(_0274_),
    .A(_1007_),
    .B(_0192_));
 sg13g2_a21oi_1 _1869_ (.A1(net41),
    .A2(_0274_),
    .Y(_0275_),
    .B1(net39));
 sg13g2_nand4_1 _1870_ (.B(_0270_),
    .C(_0273_),
    .A(_0206_),
    .Y(_0276_),
    .D(_0275_));
 sg13g2_nor3_1 _1871_ (.A(net92),
    .B(net41),
    .C(_0274_),
    .Y(_0277_));
 sg13g2_a21oi_1 _1872_ (.A1(net92),
    .A2(_0274_),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_nor2_1 _1873_ (.A(_0012_),
    .B(net54),
    .Y(_0279_));
 sg13g2_nand3_1 _1874_ (.B(net40),
    .C(_0279_),
    .A(net92),
    .Y(_0280_));
 sg13g2_o21ai_1 _1875_ (.B1(net61),
    .Y(_0281_),
    .A1(_0254_),
    .A2(_0268_));
 sg13g2_mux2_1 _1876_ (.A0(_0278_),
    .A1(_0280_),
    .S(_0281_),
    .X(_0282_));
 sg13g2_nor2_1 _1877_ (.A(_0710_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_nand3_1 _1878_ (.B(net39),
    .C(_0206_),
    .A(net92),
    .Y(_0284_));
 sg13g2_o21ai_1 _1879_ (.B1(_0284_),
    .Y(_0065_),
    .A1(_0276_),
    .A2(_0283_));
 sg13g2_nor4_2 _1880_ (.A(_0233_),
    .B(_0235_),
    .C(_0246_),
    .Y(_0285_),
    .D(_0256_));
 sg13g2_nand2_1 _1881_ (.Y(_0286_),
    .A(_0010_),
    .B(_0993_));
 sg13g2_a21oi_1 _1882_ (.A1(net51),
    .A2(_0286_),
    .Y(_0287_),
    .B1(\i2c_bert.myState_1.alu_1.acc[2] ));
 sg13g2_or3_1 _1883_ (.A(_1069_),
    .B(_0267_),
    .C(_0287_),
    .X(_0288_));
 sg13g2_buf_1 _1884_ (.A(_0288_),
    .X(_0289_));
 sg13g2_inv_1 _1885_ (.Y(_0290_),
    .A(_0271_));
 sg13g2_o21ai_1 _1886_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0285_),
    .A2(_0289_));
 sg13g2_a21o_1 _1887_ (.A2(_0012_),
    .A1(_1001_),
    .B1(_0993_),
    .X(_0292_));
 sg13g2_nand3b_1 _1888_ (.B(_0252_),
    .C(_0247_),
    .Y(_0293_),
    .A_N(_0292_));
 sg13g2_nor2b_1 _1889_ (.A(_0291_),
    .B_N(_0293_),
    .Y(_0294_));
 sg13g2_and4_1 _1890_ (.A(_0829_),
    .B(_0603_),
    .C(_0942_),
    .D(_0188_),
    .X(_0295_));
 sg13g2_a21oi_1 _1891_ (.A1(_0290_),
    .A2(_0293_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_mux2_1 _1892_ (.A0(_0294_),
    .A1(_0296_),
    .S(_1011_),
    .X(_0297_));
 sg13g2_nor2_1 _1893_ (.A(_1017_),
    .B(net41),
    .Y(_0298_));
 sg13g2_nor2_1 _1894_ (.A(_0285_),
    .B(_0289_),
    .Y(_0299_));
 sg13g2_nand2_1 _1895_ (.Y(_0300_),
    .A(_1010_),
    .B(net54));
 sg13g2_nor2_1 _1896_ (.A(_1016_),
    .B(net54),
    .Y(_0301_));
 sg13g2_nor2_1 _1897_ (.A(_1010_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nand2_1 _1898_ (.Y(_0303_),
    .A(_0299_),
    .B(_0302_));
 sg13g2_o21ai_1 _1899_ (.B1(_0303_),
    .Y(_0304_),
    .A1(_0299_),
    .A2(_0300_));
 sg13g2_a22oi_1 _1900_ (.Y(_0305_),
    .B1(_0304_),
    .B2(net40),
    .A2(_0298_),
    .A1(_0297_));
 sg13g2_xnor2_1 _1901_ (.Y(_0306_),
    .A(_1011_),
    .B(_0294_));
 sg13g2_inv_1 _1902_ (.Y(_0307_),
    .A(_0301_));
 sg13g2_o21ai_1 _1903_ (.B1(_0307_),
    .Y(_0308_),
    .A1(_0615_),
    .A2(net41));
 sg13g2_nor2_1 _1904_ (.A(_0615_),
    .B(_0307_),
    .Y(_0309_));
 sg13g2_a22oi_1 _1905_ (.Y(_0310_),
    .B1(_0309_),
    .B2(_0194_),
    .A2(_0308_),
    .A1(_1010_));
 sg13g2_nor2_1 _1906_ (.A(_1011_),
    .B(_1016_),
    .Y(_0311_));
 sg13g2_o21ai_1 _1907_ (.B1(_0677_),
    .Y(_0312_),
    .A1(net61),
    .A2(_0311_));
 sg13g2_inv_1 _1908_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_a22oi_1 _1909_ (.Y(_0314_),
    .B1(net41),
    .B2(_0301_),
    .A2(net39),
    .A1(_1010_));
 sg13g2_o21ai_1 _1910_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0310_),
    .A2(_0313_));
 sg13g2_a21oi_1 _1911_ (.A1(_0301_),
    .A2(_0306_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_nor2_1 _1912_ (.A(_0718_),
    .B(net39),
    .Y(_0317_));
 sg13g2_o21ai_1 _1913_ (.B1(_0206_),
    .Y(_0318_),
    .A1(_0315_),
    .A2(_0317_));
 sg13g2_a21oi_1 _1914_ (.A1(_0305_),
    .A2(_0316_),
    .Y(_0066_),
    .B1(_0318_));
 sg13g2_nor3_1 _1915_ (.A(net66),
    .B(_1078_),
    .C(_1024_),
    .Y(_0319_));
 sg13g2_nand2_1 _1916_ (.Y(_0320_),
    .A(_1011_),
    .B(_1016_));
 sg13g2_a21oi_1 _1917_ (.A1(_0271_),
    .A2(_0320_),
    .Y(_0321_),
    .B1(_0311_));
 sg13g2_xnor2_1 _1918_ (.Y(_0322_),
    .A(_1078_),
    .B(_1024_));
 sg13g2_nor3_1 _1919_ (.A(_0634_),
    .B(_0321_),
    .C(_0322_),
    .Y(_0323_));
 sg13g2_or2_1 _1920_ (.X(_0324_),
    .B(_0323_),
    .A(_0319_));
 sg13g2_nor3_1 _1921_ (.A(net66),
    .B(_1079_),
    .C(_1025_),
    .Y(_0325_));
 sg13g2_a21oi_1 _1922_ (.A1(net51),
    .A2(_0324_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_nor2_1 _1923_ (.A(_0710_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nor2_1 _1924_ (.A(_1024_),
    .B(net54),
    .Y(_0328_));
 sg13g2_nand2b_1 _1925_ (.Y(_0329_),
    .B(_0328_),
    .A_N(_0014_));
 sg13g2_o21ai_1 _1926_ (.B1(net61),
    .Y(_0330_),
    .A1(_1078_),
    .A2(_0328_));
 sg13g2_a21oi_1 _1927_ (.A1(_0329_),
    .A2(_0330_),
    .Y(_0331_),
    .B1(_0677_));
 sg13g2_nor3_1 _1928_ (.A(_0262_),
    .B(_0327_),
    .C(_0331_),
    .Y(_0332_));
 sg13g2_nand2_1 _1929_ (.Y(_0333_),
    .A(_0328_),
    .B(_0321_));
 sg13g2_a21oi_1 _1930_ (.A1(_1024_),
    .A2(_0321_),
    .Y(_0334_),
    .B1(_0211_));
 sg13g2_nor3_1 _1931_ (.A(_1011_),
    .B(_1016_),
    .C(_0211_),
    .Y(_0335_));
 sg13g2_xnor2_1 _1932_ (.Y(_0336_),
    .A(net92),
    .B(_0279_));
 sg13g2_nor3_1 _1933_ (.A(_0302_),
    .B(_0335_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_o21ai_1 _1934_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0254_),
    .A2(_0268_));
 sg13g2_xnor2_1 _1935_ (.Y(_0339_),
    .A(_1078_),
    .B(_0338_));
 sg13g2_mux2_1 _1936_ (.A0(_0333_),
    .A1(_0334_),
    .S(_0339_),
    .X(_0340_));
 sg13g2_o21ai_1 _1937_ (.B1(_0206_),
    .Y(_0341_),
    .A1(net40),
    .A2(_0328_));
 sg13g2_a21o_1 _1938_ (.A2(_0223_),
    .A1(_1079_),
    .B1(_0341_),
    .X(_0342_));
 sg13g2_a21o_1 _1939_ (.A2(_0332_),
    .A1(_0718_),
    .B1(_0342_),
    .X(_0343_));
 sg13g2_a21oi_1 _1940_ (.A1(_0332_),
    .A2(_0340_),
    .Y(_0067_),
    .B1(_0343_));
 sg13g2_nor2_1 _1941_ (.A(_1010_),
    .B(_1016_),
    .Y(_0344_));
 sg13g2_nor4_1 _1942_ (.A(_1011_),
    .B(_1078_),
    .C(_1017_),
    .D(_1024_),
    .Y(_0345_));
 sg13g2_a21oi_1 _1943_ (.A1(_0322_),
    .A2(_0344_),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_nor2_1 _1944_ (.A(net54),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_nand2_1 _1945_ (.Y(_0348_),
    .A(_1016_),
    .B(_1024_));
 sg13g2_nand2_1 _1946_ (.Y(_0349_),
    .A(_1010_),
    .B(_1078_));
 sg13g2_a21oi_1 _1947_ (.A1(net51),
    .A2(_0348_),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_or2_1 _1948_ (.X(_0351_),
    .B(_0350_),
    .A(_0347_));
 sg13g2_nand2_1 _1949_ (.Y(_0352_),
    .A(_1032_),
    .B(net51));
 sg13g2_nand2_1 _1950_ (.Y(_0353_),
    .A(_0311_),
    .B(_0322_));
 sg13g2_o21ai_1 _1951_ (.B1(_0353_),
    .Y(_0354_),
    .A1(_0014_),
    .A2(_1024_));
 sg13g2_or2_1 _1952_ (.X(_0355_),
    .B(_0354_),
    .A(_0352_));
 sg13g2_nor2_1 _1953_ (.A(_0351_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_and3_1 _1954_ (.X(_0357_),
    .A(net95),
    .B(_0966_),
    .C(_0976_));
 sg13g2_a221oi_1 _1955_ (.B2(_0193_),
    .C1(_0246_),
    .B1(_0357_),
    .A1(net93),
    .Y(_0358_),
    .A2(_0233_));
 sg13g2_o21ai_1 _1956_ (.B1(_0238_),
    .Y(_0359_),
    .A1(_0233_),
    .A2(_0235_));
 sg13g2_a221oi_1 _1957_ (.B2(_0359_),
    .C1(_0292_),
    .B1(_0358_),
    .A1(_0226_),
    .Y(_0360_),
    .A2(_0227_));
 sg13g2_nand2_1 _1958_ (.Y(_0361_),
    .A(net51),
    .B(_0271_));
 sg13g2_o21ai_1 _1959_ (.B1(_0361_),
    .Y(_0362_),
    .A1(_0285_),
    .A2(_0289_));
 sg13g2_nor3_1 _1960_ (.A(_0355_),
    .B(_0360_),
    .C(_0362_),
    .Y(_0363_));
 sg13g2_o21ai_1 _1961_ (.B1(_1082_),
    .Y(_0364_),
    .A1(_0356_),
    .A2(_0363_));
 sg13g2_nor3_1 _1962_ (.A(_0285_),
    .B(_0289_),
    .C(_0349_),
    .Y(_0365_));
 sg13g2_xnor2_1 _1963_ (.Y(_0366_),
    .A(_1082_),
    .B(_0365_));
 sg13g2_nand3_1 _1964_ (.B(_1032_),
    .C(_0351_),
    .A(\i2c_bert.myState_1.alu_1.acc[7] ),
    .Y(_0367_));
 sg13g2_a21oi_1 _1965_ (.A1(_0295_),
    .A2(_0365_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_nand2b_1 _1966_ (.Y(_0369_),
    .B(_0293_),
    .A_N(_0291_));
 sg13g2_a22oi_1 _1967_ (.Y(_0370_),
    .B1(_0368_),
    .B2(_0369_),
    .A2(_0366_),
    .A1(_0295_));
 sg13g2_a22oi_1 _1968_ (.Y(_0371_),
    .B1(net41),
    .B2(_0352_),
    .A2(net39),
    .A1(_1082_));
 sg13g2_nand2_1 _1969_ (.Y(_0372_),
    .A(_0206_),
    .B(_0371_));
 sg13g2_or2_1 _1970_ (.X(_0373_),
    .B(_0372_),
    .A(_0718_));
 sg13g2_a21oi_1 _1971_ (.A1(_0364_),
    .A2(_0370_),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_inv_1 _1972_ (.Y(_0375_),
    .A(_0372_));
 sg13g2_nand2_1 _1973_ (.Y(_0376_),
    .A(_1082_),
    .B(_0352_));
 sg13g2_nor2_1 _1974_ (.A(_0016_),
    .B(_0352_),
    .Y(_0377_));
 sg13g2_a21oi_1 _1975_ (.A1(net61),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_xor2_1 _1976_ (.B(_0009_),
    .A(\i2c_bert.myState_1.alu_1.acc[7] ),
    .X(_0379_));
 sg13g2_nand4_1 _1977_ (.B(net51),
    .C(_0379_),
    .A(_0676_),
    .Y(_0380_),
    .D(_0354_));
 sg13g2_o21ai_1 _1978_ (.B1(_0380_),
    .Y(_0381_),
    .A1(net61),
    .A2(_0379_));
 sg13g2_a21oi_1 _1979_ (.A1(net60),
    .A2(_0381_),
    .Y(_0382_),
    .B1(_0262_));
 sg13g2_o21ai_1 _1980_ (.B1(_0382_),
    .Y(_0383_),
    .A1(net60),
    .A2(_0378_));
 sg13g2_nor3_1 _1981_ (.A(_1032_),
    .B(_0718_),
    .C(_0372_),
    .Y(_0384_));
 sg13g2_nor2_1 _1982_ (.A(_1082_),
    .B(_0354_),
    .Y(_0385_));
 sg13g2_o21ai_1 _1983_ (.B1(_0351_),
    .Y(_0386_),
    .A1(_0360_),
    .A2(_0362_));
 sg13g2_mux2_1 _1984_ (.A0(_1082_),
    .A1(_0385_),
    .S(_0386_),
    .X(_0387_));
 sg13g2_a22oi_1 _1985_ (.Y(_0388_),
    .B1(_0384_),
    .B2(_0387_),
    .A2(_0383_),
    .A1(_0375_));
 sg13g2_nand2b_1 _1986_ (.Y(_0068_),
    .B(_0388_),
    .A_N(_0374_));
 sg13g2_buf_1 _1987_ (.A(_0687_),
    .X(_0389_));
 sg13g2_nor2_1 _1988_ (.A(net59),
    .B(_0845_),
    .Y(_0035_));
 sg13g2_nor2_1 _1989_ (.A(net59),
    .B(_0901_),
    .Y(_0036_));
 sg13g2_nor2_1 _1990_ (.A(net59),
    .B(_0877_),
    .Y(_0037_));
 sg13g2_inv_1 _1991_ (.Y(_0390_),
    .A(\i2c_bert.i2c.sclAndNor5.io_o ));
 sg13g2_nand3_1 _1992_ (.B(\i2c_bert.i2c.sclAndNor5.io_d ),
    .C(_0534_),
    .A(\i2c_bert.i2c.sclAndNor5.io_e ),
    .Y(_0391_));
 sg13g2_nand2_1 _1993_ (.Y(_0392_),
    .A(_0542_),
    .B(_0544_));
 sg13g2_a21oi_1 _1994_ (.A1(\i2c_bert.i2c.sclAndNor5.io_o ),
    .A2(_0392_),
    .Y(_0393_),
    .B1(_0539_));
 sg13g2_a21oi_1 _1995_ (.A1(_0390_),
    .A2(_0391_),
    .Y(_0041_),
    .B1(_0393_));
 sg13g2_nand2_1 _1996_ (.Y(_0394_),
    .A(\i2c_bert.i2c.sdaAndNor3.io_o ),
    .B(_0570_));
 sg13g2_o21ai_1 _1997_ (.B1(net14),
    .Y(_0395_),
    .A1(\i2c_bert.i2c.sdaAndNor3.io_o ),
    .A2(_0577_));
 sg13g2_nand2_1 _1998_ (.Y(_0046_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_inv_1 _1999_ (.Y(_0396_),
    .A(\i2c_bert.i2c.sdaAndNor5.io_o ));
 sg13g2_nor3_1 _2000_ (.A(_0558_),
    .B(_0560_),
    .C(_0570_),
    .Y(_0397_));
 sg13g2_and3_1 _2001_ (.X(_0398_),
    .A(_0558_),
    .B(_0560_),
    .C(_0577_));
 sg13g2_o21ai_1 _2002_ (.B1(net14),
    .Y(_0399_),
    .A1(\i2c_bert.i2c.sdaAndNor5.io_o ),
    .A2(_0398_));
 sg13g2_o21ai_1 _2003_ (.B1(_0399_),
    .Y(_0047_),
    .A1(_0396_),
    .A2(_0397_));
 sg13g2_nor2_1 _2004_ (.A(_0029_),
    .B(net50),
    .Y(_0400_));
 sg13g2_nor2_1 _2005_ (.A(net77),
    .B(_0707_),
    .Y(_0401_));
 sg13g2_nor2_1 _2006_ (.A(\i2c_bert.myState_1.fsmPhase_stateReg[2] ),
    .B(_0707_),
    .Y(_0402_));
 sg13g2_nor2_1 _2007_ (.A(net49),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_a221oi_1 _2008_ (.B2(_0029_),
    .C1(_0403_),
    .B1(_0401_),
    .A1(_0668_),
    .Y(_0404_),
    .A2(_0400_));
 sg13g2_buf_1 _2009_ (.A(_0404_),
    .X(_0405_));
 sg13g2_nor2_1 _2010_ (.A(_0830_),
    .B(_0705_),
    .Y(_0406_));
 sg13g2_nor2_1 _2011_ (.A(_0707_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_nor3_1 _2012_ (.A(net67),
    .B(_0401_),
    .C(_0407_),
    .Y(_0408_));
 sg13g2_nand2_1 _2013_ (.Y(_0409_),
    .A(net38),
    .B(_0408_));
 sg13g2_nand2b_1 _2014_ (.Y(_0410_),
    .B(net67),
    .A_N(net38));
 sg13g2_nand3_1 _2015_ (.B(_0409_),
    .C(_0410_),
    .A(net78),
    .Y(_0076_));
 sg13g2_a21o_1 _2016_ (.A2(_0407_),
    .A1(net38),
    .B1(_0687_),
    .X(_0411_));
 sg13g2_buf_1 _2017_ (.A(_0411_),
    .X(_0412_));
 sg13g2_and2_1 _2018_ (.A(_0608_),
    .B(_0621_),
    .X(_0413_));
 sg13g2_buf_1 _2019_ (.A(_0413_),
    .X(_0414_));
 sg13g2_nand3_1 _2020_ (.B(\i2c_bert.myState_1.counter[4] ),
    .C(\i2c_bert.myState_1.counter[5] ),
    .A(_0625_),
    .Y(_0415_));
 sg13g2_nand2_1 _2021_ (.Y(_0416_),
    .A(_0624_),
    .B(\i2c_bert.myState_1.counter[6] ));
 sg13g2_nor2_1 _2022_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_and2_1 _2023_ (.A(\i2c_bert.myState_1.counter[7] ),
    .B(_0417_),
    .X(_0418_));
 sg13g2_and4_1 _2024_ (.A(\i2c_bert.myState_1.counter[8] ),
    .B(net38),
    .C(_0414_),
    .D(_0418_),
    .X(_0419_));
 sg13g2_nand2_1 _2025_ (.Y(_0420_),
    .A(\i2c_bert.myState_1.counter[9] ),
    .B(_0419_));
 sg13g2_xor2_1 _2026_ (.B(_0420_),
    .A(\i2c_bert.myState_1.counter[10] ),
    .X(_0421_));
 sg13g2_nor2_1 _2027_ (.A(_0412_),
    .B(_0421_),
    .Y(_0077_));
 sg13g2_nand3_1 _2028_ (.B(\i2c_bert.myState_1.counter[10] ),
    .C(_0419_),
    .A(\i2c_bert.myState_1.counter[9] ),
    .Y(_0422_));
 sg13g2_xor2_1 _2029_ (.B(_0422_),
    .A(\i2c_bert.myState_1.counter[11] ),
    .X(_0423_));
 sg13g2_nor2_1 _2030_ (.A(_0412_),
    .B(_0423_),
    .Y(_0078_));
 sg13g2_o21ai_1 _2031_ (.B1(_0405_),
    .Y(_0424_),
    .A1(net67),
    .A2(_0407_));
 sg13g2_nor2_1 _2032_ (.A(net69),
    .B(_0407_),
    .Y(_0425_));
 sg13g2_and2_1 _2033_ (.A(net67),
    .B(_0405_),
    .X(_0426_));
 sg13g2_a22oi_1 _2034_ (.Y(_0427_),
    .B1(_0425_),
    .B2(_0426_),
    .A2(_0424_),
    .A1(net69));
 sg13g2_nor2_1 _2035_ (.A(net59),
    .B(_0427_),
    .Y(_0079_));
 sg13g2_nand2_1 _2036_ (.Y(_0428_),
    .A(net38),
    .B(_0414_));
 sg13g2_xor2_1 _2037_ (.B(_0428_),
    .A(_0624_),
    .X(_0429_));
 sg13g2_nor2_1 _2038_ (.A(net34),
    .B(_0429_),
    .Y(_0080_));
 sg13g2_and3_1 _2039_ (.X(_0430_),
    .A(_0624_),
    .B(net38),
    .C(_0414_));
 sg13g2_buf_1 _2040_ (.A(_0430_),
    .X(_0431_));
 sg13g2_xnor2_1 _2041_ (.Y(_0432_),
    .A(_0625_),
    .B(_0431_));
 sg13g2_nor2_1 _2042_ (.A(net34),
    .B(_0432_),
    .Y(_0081_));
 sg13g2_nand2_1 _2043_ (.Y(_0433_),
    .A(_0625_),
    .B(_0431_));
 sg13g2_xor2_1 _2044_ (.B(_0433_),
    .A(\i2c_bert.myState_1.counter[4] ),
    .X(_0434_));
 sg13g2_nor2_1 _2045_ (.A(net34),
    .B(_0434_),
    .Y(_0082_));
 sg13g2_nand3_1 _2046_ (.B(\i2c_bert.myState_1.counter[4] ),
    .C(_0431_),
    .A(_0625_),
    .Y(_0435_));
 sg13g2_xor2_1 _2047_ (.B(_0435_),
    .A(\i2c_bert.myState_1.counter[5] ),
    .X(_0436_));
 sg13g2_nor2_1 _2048_ (.A(net34),
    .B(_0436_),
    .Y(_0083_));
 sg13g2_nand2b_1 _2049_ (.Y(_0437_),
    .B(_0431_),
    .A_N(_0415_));
 sg13g2_xor2_1 _2050_ (.B(_0437_),
    .A(\i2c_bert.myState_1.counter[6] ),
    .X(_0438_));
 sg13g2_nor2_1 _2051_ (.A(net34),
    .B(_0438_),
    .Y(_0084_));
 sg13g2_nand3_1 _2052_ (.B(_0414_),
    .C(_0417_),
    .A(net38),
    .Y(_0439_));
 sg13g2_xor2_1 _2053_ (.B(_0439_),
    .A(\i2c_bert.myState_1.counter[7] ),
    .X(_0440_));
 sg13g2_nor2_1 _2054_ (.A(net34),
    .B(_0440_),
    .Y(_0085_));
 sg13g2_nand3_1 _2055_ (.B(_0414_),
    .C(_0418_),
    .A(net38),
    .Y(_0441_));
 sg13g2_xor2_1 _2056_ (.B(_0441_),
    .A(\i2c_bert.myState_1.counter[8] ),
    .X(_0442_));
 sg13g2_nor2_1 _2057_ (.A(net34),
    .B(_0442_),
    .Y(_0086_));
 sg13g2_xnor2_1 _2058_ (.Y(_0443_),
    .A(\i2c_bert.myState_1.counter[9] ),
    .B(_0419_));
 sg13g2_nor2_1 _2059_ (.A(net34),
    .B(_0443_),
    .Y(_0087_));
 sg13g2_and2_1 _2060_ (.A(_0606_),
    .B(_0203_),
    .X(_0444_));
 sg13g2_nand2_1 _2061_ (.Y(_0445_),
    .A(net79),
    .B(\i2c_bert.i2c.io_sdaSignal ));
 sg13g2_nand3_1 _2062_ (.B(net56),
    .C(_0445_),
    .A(net49),
    .Y(_0446_));
 sg13g2_nand3b_1 _2063_ (.B(_0030_),
    .C(_0605_),
    .Y(_0447_),
    .A_N(net79));
 sg13g2_nand3_1 _2064_ (.B(_0446_),
    .C(_0447_),
    .A(net87),
    .Y(_0448_));
 sg13g2_o21ai_1 _2065_ (.B1(_0448_),
    .Y(_0449_),
    .A1(_0205_),
    .A2(_0444_));
 sg13g2_buf_1 _2066_ (.A(_0449_),
    .X(_0450_));
 sg13g2_buf_1 _2067_ (.A(_0450_),
    .X(_0451_));
 sg13g2_nor3_1 _2068_ (.A(_0030_),
    .B(net52),
    .C(_0450_),
    .Y(_0452_));
 sg13g2_a21oi_1 _2069_ (.A1(\i2c_bert.myState_1.len12[4] ),
    .A2(net33),
    .Y(_0453_),
    .B1(_0452_));
 sg13g2_nor2_1 _2070_ (.A(net59),
    .B(_0453_),
    .Y(_0096_));
 sg13g2_nand2_1 _2071_ (.Y(_0454_),
    .A(\i2c_bert.myState_1.len12[5] ),
    .B(_0450_));
 sg13g2_o21ai_1 _2072_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_1061_),
    .A2(net33));
 sg13g2_and2_1 _2073_ (.A(net78),
    .B(_0455_),
    .X(_0097_));
 sg13g2_nand2_1 _2074_ (.Y(_0456_),
    .A(\i2c_bert.myState_1.len12[6] ),
    .B(_0450_));
 sg13g2_o21ai_1 _2075_ (.B1(_0456_),
    .Y(_0457_),
    .A1(_1065_),
    .A2(_0451_));
 sg13g2_and2_1 _2076_ (.A(net78),
    .B(_0457_),
    .X(_0098_));
 sg13g2_nor2_1 _2077_ (.A(_1070_),
    .B(net33),
    .Y(_0458_));
 sg13g2_a21oi_1 _2078_ (.A1(\i2c_bert.myState_1.len12[7] ),
    .A2(net33),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_nor2_1 _2079_ (.A(net59),
    .B(_0459_),
    .Y(_0099_));
 sg13g2_nand2_1 _2080_ (.Y(_0460_),
    .A(\i2c_bert.myState_1.len12[8] ),
    .B(_0450_));
 sg13g2_o21ai_1 _2081_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_1072_),
    .A2(_0451_));
 sg13g2_and2_1 _2082_ (.A(net78),
    .B(_0461_),
    .X(_0100_));
 sg13g2_nor2_1 _2083_ (.A(_1076_),
    .B(net33),
    .Y(_0462_));
 sg13g2_a21oi_1 _2084_ (.A1(\i2c_bert.myState_1.len12[9] ),
    .A2(net33),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_nor2_1 _2085_ (.A(net59),
    .B(_0463_),
    .Y(_0101_));
 sg13g2_nor2_1 _2086_ (.A(_1080_),
    .B(_0450_),
    .Y(_0464_));
 sg13g2_a21oi_1 _2087_ (.A1(\i2c_bert.myState_1.len12[10] ),
    .A2(net33),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nor2_1 _2088_ (.A(net59),
    .B(_0465_),
    .Y(_0102_));
 sg13g2_nor2_1 _2089_ (.A(_1083_),
    .B(_0450_),
    .Y(_0466_));
 sg13g2_a21oi_1 _2090_ (.A1(\i2c_bert.myState_1.len12[11] ),
    .A2(net33),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_nor2_1 _2091_ (.A(_0389_),
    .B(_0467_),
    .Y(_0103_));
 sg13g2_and2_1 _2092_ (.A(_0686_),
    .B(_0007_),
    .X(_0468_));
 sg13g2_nor2_1 _2093_ (.A(_0808_),
    .B(_0687_),
    .Y(_0469_));
 sg13g2_o21ai_1 _2094_ (.B1(net64),
    .Y(_0470_),
    .A1(net70),
    .A2(net72));
 sg13g2_nand2_1 _2095_ (.Y(_0471_),
    .A(_0889_),
    .B(_0470_));
 sg13g2_o21ai_1 _2096_ (.B1(_0585_),
    .Y(_0472_),
    .A1(_0830_),
    .A2(_0786_));
 sg13g2_a22oi_1 _2097_ (.Y(_0473_),
    .B1(_0472_),
    .B2(_0789_),
    .A2(_0471_),
    .A1(_0788_));
 sg13g2_nand2b_1 _2098_ (.Y(_0474_),
    .B(net53),
    .A_N(_0878_));
 sg13g2_nand3_1 _2099_ (.B(_0473_),
    .C(_0474_),
    .A(\i2c_bert.powerOnSenseCaptured.Q ),
    .Y(_0475_));
 sg13g2_and2_1 _2100_ (.A(\i2c_bert.powerOnSenseCaptured.Q ),
    .B(_0167_),
    .X(_0476_));
 sg13g2_nand4_1 _2101_ (.B(_0877_),
    .C(_0168_),
    .A(_0845_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_nand2_1 _2102_ (.Y(_0478_),
    .A(_0475_),
    .B(_0477_));
 sg13g2_mux2_1 _2103_ (.A0(_0468_),
    .A1(_0469_),
    .S(_0478_),
    .X(_0117_));
 sg13g2_nand3_1 _2104_ (.B(_0475_),
    .C(_0477_),
    .A(net78),
    .Y(_0479_));
 sg13g2_buf_1 _2105_ (.A(_0479_),
    .X(_0480_));
 sg13g2_inv_1 _2106_ (.Y(_0481_),
    .A(\i2c_bert.timer_1.ticker_count[7] ));
 sg13g2_inv_1 _2107_ (.Y(_0482_),
    .A(\i2c_bert.timer_1.ticker_count[3] ));
 sg13g2_nand3_1 _2108_ (.B(_0813_),
    .C(\i2c_bert.timer_1.ticker_count[2] ),
    .A(_0808_),
    .Y(_0483_));
 sg13g2_nor2_2 _2109_ (.A(_0482_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nand4_1 _2110_ (.B(_0811_),
    .C(\i2c_bert.timer_1.ticker_count[6] ),
    .A(_0805_),
    .Y(_0485_),
    .D(_0484_));
 sg13g2_nor2_2 _2111_ (.A(_0481_),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_nand3_1 _2112_ (.B(_0796_),
    .C(_0486_),
    .A(_0798_),
    .Y(_0487_));
 sg13g2_xor2_1 _2113_ (.B(_0487_),
    .A(\i2c_bert.timer_1.ticker_count[10] ),
    .X(_0488_));
 sg13g2_nor2_1 _2114_ (.A(net32),
    .B(_0488_),
    .Y(_0118_));
 sg13g2_nand4_1 _2115_ (.B(_0796_),
    .C(\i2c_bert.timer_1.ticker_count[10] ),
    .A(_0798_),
    .Y(_0489_),
    .D(_0486_));
 sg13g2_xor2_1 _2116_ (.B(_0489_),
    .A(\i2c_bert.timer_1.ticker_count[11] ),
    .X(_0490_));
 sg13g2_nor2_1 _2117_ (.A(net32),
    .B(_0490_),
    .Y(_0119_));
 sg13g2_xnor2_1 _2118_ (.Y(_0491_),
    .A(_0808_),
    .B(_0813_));
 sg13g2_nor2_1 _2119_ (.A(_0389_),
    .B(_0491_),
    .Y(_0120_));
 sg13g2_nand2_1 _2120_ (.Y(_0492_),
    .A(_0808_),
    .B(_0813_));
 sg13g2_xnor2_1 _2121_ (.Y(_0493_),
    .A(_0008_),
    .B(_0492_));
 sg13g2_nor2_1 _2122_ (.A(_0687_),
    .B(_0493_),
    .Y(_0121_));
 sg13g2_xnor2_1 _2123_ (.Y(_0494_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_nor2_1 _2124_ (.A(net32),
    .B(_0494_),
    .Y(_0122_));
 sg13g2_xnor2_1 _2125_ (.Y(_0495_),
    .A(_0805_),
    .B(_0484_));
 sg13g2_nor2_1 _2126_ (.A(net32),
    .B(_0495_),
    .Y(_0123_));
 sg13g2_nand2_1 _2127_ (.Y(_0496_),
    .A(_0805_),
    .B(_0484_));
 sg13g2_xor2_1 _2128_ (.B(_0496_),
    .A(_0811_),
    .X(_0497_));
 sg13g2_nor2_1 _2129_ (.A(net32),
    .B(_0497_),
    .Y(_0124_));
 sg13g2_nand3_1 _2130_ (.B(_0811_),
    .C(_0484_),
    .A(_0805_),
    .Y(_0498_));
 sg13g2_xor2_1 _2131_ (.B(_0498_),
    .A(\i2c_bert.timer_1.ticker_count[6] ),
    .X(_0499_));
 sg13g2_nor2_1 _2132_ (.A(_0480_),
    .B(_0499_),
    .Y(_0125_));
 sg13g2_xnor2_1 _2133_ (.Y(_0500_),
    .A(_0481_),
    .B(_0485_));
 sg13g2_nor2_1 _2134_ (.A(net32),
    .B(_0500_),
    .Y(_0126_));
 sg13g2_xnor2_1 _2135_ (.Y(_0501_),
    .A(_0798_),
    .B(_0486_));
 sg13g2_nor2_1 _2136_ (.A(net32),
    .B(_0501_),
    .Y(_0127_));
 sg13g2_nand2_1 _2137_ (.Y(_0502_),
    .A(_0798_),
    .B(_0486_));
 sg13g2_xor2_1 _2138_ (.B(_0502_),
    .A(_0796_),
    .X(_0503_));
 sg13g2_nor2_1 _2139_ (.A(net32),
    .B(_0503_),
    .Y(_0128_));
 sg13g2_o21ai_1 _2140_ (.B1(_0937_),
    .Y(_0504_),
    .A1(_0762_),
    .A2(_0988_));
 sg13g2_inv_1 _2141_ (.Y(_0505_),
    .A(_0918_));
 sg13g2_o21ai_1 _2142_ (.B1(_0505_),
    .Y(\i2c_bert.i2c.io_bus_sclOe ),
    .A1(_0866_),
    .A2(_0504_));
 sg13g2_nand2_1 _2143_ (.Y(_0506_),
    .A(_0539_),
    .B(_0742_));
 sg13g2_nor2_1 _2144_ (.A(_0745_),
    .B(_0847_),
    .Y(_0507_));
 sg13g2_a21oi_1 _2145_ (.A1(_0506_),
    .A2(_0507_),
    .Y(\i2c_bert.i2c.io_bus_sclOut ),
    .B1(_0918_));
 sg13g2_a21oi_1 _2146_ (.A1(_0670_),
    .A2(net55),
    .Y(_0508_),
    .B1(_0866_));
 sg13g2_a21oi_1 _2147_ (.A1(_0869_),
    .A2(_0508_),
    .Y(_0509_),
    .B1(_0791_));
 sg13g2_nand2b_1 _2148_ (.Y(_0510_),
    .B(net77),
    .A_N(_0988_));
 sg13g2_nand4_1 _2149_ (.B(_0728_),
    .C(_0789_),
    .A(_0839_),
    .Y(_0511_),
    .D(_0510_));
 sg13g2_a21o_1 _2150_ (.A2(\i2c_bert.i2c.io_data8rx[7] ),
    .A1(_0839_),
    .B1(_0730_),
    .X(_0512_));
 sg13g2_a21o_1 _2151_ (.A2(_0510_),
    .A1(_0728_),
    .B1(_0866_),
    .X(_0513_));
 sg13g2_o21ai_1 _2152_ (.B1(_0513_),
    .Y(_0514_),
    .A1(_0988_),
    .A2(_0506_));
 sg13g2_a221oi_1 _2153_ (.B2(_0733_),
    .C1(_0735_),
    .B1(_0514_),
    .A1(_0511_),
    .Y(_0515_),
    .A2(_0512_));
 sg13g2_nor2_1 _2154_ (.A(_0988_),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_nor2_1 _2155_ (.A(_0509_),
    .B(_0516_),
    .Y(\i2c_bert.i2c.io_bus_sdaOe ));
 sg13g2_a21oi_1 _2156_ (.A1(_0785_),
    .A2(_0737_),
    .Y(_0517_),
    .B1(_0918_));
 sg13g2_a21oi_1 _2157_ (.A1(_0988_),
    .A2(_0517_),
    .Y(\i2c_bert.i2c.io_bus_sdaOut ),
    .B1(_0515_));
 sg13g2_nor2b_1 _2158_ (.A(_0006_),
    .B_N(_0008_),
    .Y(_0518_));
 sg13g2_nor2_1 _2159_ (.A(_0923_),
    .B(_0008_),
    .Y(_0519_));
 sg13g2_a22oi_1 _2160_ (.Y(_0520_),
    .B1(_0519_),
    .B2(_0007_),
    .A2(_0518_),
    .A1(_0923_));
 sg13g2_or2_1 _2161_ (.X(_0521_),
    .B(_0520_),
    .A(_0813_));
 sg13g2_inv_1 _2162_ (.Y(_0522_),
    .A(_0805_));
 sg13g2_nor4_1 _2163_ (.A(\i2c_bert.timer_1.ticker_count[2] ),
    .B(\i2c_bert.timer_1.ticker_count[3] ),
    .C(_0522_),
    .D(_0923_),
    .Y(_0523_));
 sg13g2_and4_1 _2164_ (.A(_0522_),
    .B(_0811_),
    .C(_0923_),
    .D(_0006_),
    .X(_0524_));
 sg13g2_o21ai_1 _2165_ (.B1(net4),
    .Y(_0525_),
    .A1(_0523_),
    .A2(_0524_));
 sg13g2_o21ai_1 _2166_ (.B1(_0525_),
    .Y(\i2c_bert.powerOnSenseCaptured.GATE ),
    .A1(net4),
    .A2(_0521_));
 sg13g2_nor2b_1 _2167_ (.A(\i2c_bert.powerOnSenseCaptured.Q ),
    .B_N(\i2c_bert.powerOnSenseCaptured.GATE ),
    .Y(\i2c_bert.powerOnSense.GATE ));
 sg13g2_buf_4 _2168_ (.X(_0526_),
    .A(net10));
 sg13g2_mux2_1 _2169_ (.A0(\i2c_bert.myState_1.led8[0] ),
    .A1(_0941_),
    .S(_0526_),
    .X(net24));
 sg13g2_mux2_1 _2170_ (.A0(\i2c_bert.myState_1.led8[1] ),
    .A1(net94),
    .S(_0526_),
    .X(net25));
 sg13g2_mux2_1 _2171_ (.A0(\i2c_bert.myState_1.led8[2] ),
    .A1(net93),
    .S(_0526_),
    .X(net26));
 sg13g2_mux2_1 _2172_ (.A0(\i2c_bert.myState_1.led8[3] ),
    .A1(\i2c_bert.myState_1.alu_1.acc[3] ),
    .S(_0526_),
    .X(net27));
 sg13g2_mux2_1 _2173_ (.A0(\i2c_bert.myState_1.led8[4] ),
    .A1(_1000_),
    .S(_0526_),
    .X(net28));
 sg13g2_mux2_1 _2174_ (.A0(\i2c_bert.myState_1.led8[5] ),
    .A1(_1010_),
    .S(_0526_),
    .X(net29));
 sg13g2_mux2_1 _2175_ (.A0(\i2c_bert.myState_1.led8[6] ),
    .A1(_1078_),
    .S(_0526_),
    .X(net30));
 sg13g2_mux2_1 _2176_ (.A0(\i2c_bert.myState_1.led8[7] ),
    .A1(\i2c_bert.myState_1.alu_1.acc[7] ),
    .S(_0526_),
    .X(net31));
 sg13g2_buf_1 _2177_ (.A(\i2c_bert.i2c.io_sclMode[1] ),
    .X(_0527_));
 sg13g2_buf_1 _2178_ (.A(\i2c_bert.i2c.clockGate.sel ),
    .X(_0528_));
 sg13g2_or2_1 _2179_ (.X(_0529_),
    .B(\i2c_bert.i2c.sclAndNor3.io_o ),
    .A(\i2c_bert.i2c.io_sclMode[2] ));
 sg13g2_buf_1 _2180_ (.A(\i2c_bert.i2c.io_sclMode[2] ),
    .X(_0530_));
 sg13g2_nor2_1 _2181_ (.A(net90),
    .B(net89),
    .Y(_0531_));
 sg13g2_a22oi_1 _2182_ (.Y(_0532_),
    .B1(_0531_),
    .B2(\i2c_bert.i2c.sclAndNor3.io_c ),
    .A2(_0529_),
    .A1(net90));
 sg13g2_nor2b_1 _2183_ (.A(_0528_),
    .B_N(\i2c_bert.i2c.io_sclMode[2] ),
    .Y(_0533_));
 sg13g2_and2_1 _2184_ (.A(\i2c_bert.i2c.sclAndNor3.io_b ),
    .B(\i2c_bert.i2c.sclAndNor3.io_c ),
    .X(_0534_));
 sg13g2_nor2b_1 _2185_ (.A(_0530_),
    .B_N(\i2c_bert.i2c.clockGate.sel ),
    .Y(_0535_));
 sg13g2_a221oi_1 _2186_ (.B2(_0535_),
    .C1(net91),
    .B1(_0534_),
    .A1(\i2c_bert.i2c.sclAndNor5.io_e ),
    .Y(_0536_),
    .A2(_0533_));
 sg13g2_a21o_1 _2187_ (.A2(_0532_),
    .A1(net91),
    .B1(_0536_),
    .X(_0537_));
 sg13g2_buf_1 _2188_ (.A(_0537_),
    .X(_0538_));
 sg13g2_buf_2 _2189_ (.A(net13),
    .X(_0539_));
 sg13g2_inv_2 _2190_ (.Y(_0540_),
    .A(_0539_));
 sg13g2_nand2_1 _2191_ (.Y(_0541_),
    .A(\i2c_bert.i2c.sclAndNor5.io_e ),
    .B(\i2c_bert.i2c.sclAndNor5.io_d ));
 sg13g2_nor2_1 _2192_ (.A(\i2c_bert.i2c.sclAndNor3.io_b ),
    .B(\i2c_bert.i2c.sclAndNor3.io_c ),
    .Y(_0542_));
 sg13g2_nand3_1 _2193_ (.B(_0541_),
    .C(_0542_),
    .A(_0540_),
    .Y(_0543_));
 sg13g2_nor2_1 _2194_ (.A(\i2c_bert.i2c.sclAndNor5.io_e ),
    .B(\i2c_bert.i2c.sclAndNor5.io_d ),
    .Y(_0544_));
 sg13g2_nand2_1 _2195_ (.Y(_0545_),
    .A(net90),
    .B(net89));
 sg13g2_nor3_1 _2196_ (.A(\i2c_bert.i2c.io_sclMode[1] ),
    .B(_0544_),
    .C(_0545_),
    .Y(_0546_));
 sg13g2_xnor2_1 _2197_ (.Y(_0547_),
    .A(\i2c_bert.i2c.io_sclMode[1] ),
    .B(net89));
 sg13g2_nor2_1 _2198_ (.A(_0528_),
    .B(_0540_),
    .Y(_0548_));
 sg13g2_nor4_1 _2199_ (.A(net91),
    .B(net89),
    .C(_0540_),
    .D(_0542_),
    .Y(_0549_));
 sg13g2_a221oi_1 _2200_ (.B2(_0548_),
    .C1(_0549_),
    .B1(_0547_),
    .A1(_0543_),
    .Y(_0550_),
    .A2(_0546_));
 sg13g2_buf_2 _2201_ (.A(_0550_),
    .X(_0551_));
 sg13g2_and2_1 _2202_ (.A(net90),
    .B(net89),
    .X(_0552_));
 sg13g2_nor2b_1 _2203_ (.A(\i2c_bert.i2c.sclAndNor5.io_o ),
    .B_N(\i2c_bert.i2c.io_sclMode[1] ),
    .Y(_0553_));
 sg13g2_and2_1 _2204_ (.A(_0552_),
    .B(_0553_),
    .X(_0554_));
 sg13g2_a21o_1 _2205_ (.A2(_0551_),
    .A1(_0538_),
    .B1(_0554_),
    .X(_0555_));
 sg13g2_inv_2 _2206_ (.Y(\i2c_bert.i2c.scl ),
    .A(_0555_));
 sg13g2_nor2_1 _2207_ (.A(net14),
    .B(\i2c_bert.i2c.sdaAndNor3.io_b ),
    .Y(_0556_));
 sg13g2_buf_1 _2208_ (.A(\i2c_bert.i2c.sdaAndNor3.io_c ),
    .X(_0557_));
 sg13g2_buf_2 _2209_ (.A(\i2c_bert.i2c.sdaAndNor5.io_d ),
    .X(_0558_));
 sg13g2_nor2_1 _2210_ (.A(net88),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_buf_2 _2211_ (.A(\i2c_bert.i2c.sdaAndNor5.io_e ),
    .X(_0560_));
 sg13g2_a21oi_1 _2212_ (.A1(net88),
    .A2(_0558_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_or3_1 _2213_ (.A(_0556_),
    .B(_0559_),
    .C(_0561_),
    .X(_0562_));
 sg13g2_nand3_1 _2214_ (.B(_0558_),
    .C(_0560_),
    .A(net88),
    .Y(_0563_));
 sg13g2_nor3_1 _2215_ (.A(net88),
    .B(_0558_),
    .C(_0560_),
    .Y(_0564_));
 sg13g2_or3_1 _2216_ (.A(net91),
    .B(_0545_),
    .C(_0564_),
    .X(_0565_));
 sg13g2_a21oi_2 _2217_ (.B1(_0565_),
    .Y(_0566_),
    .A2(_0563_),
    .A1(_0562_));
 sg13g2_inv_1 _2218_ (.Y(_0567_),
    .A(\i2c_bert.i2c.sdaAndNor3.io_b ));
 sg13g2_or4_1 _2219_ (.A(net91),
    .B(_0567_),
    .C(_0545_),
    .D(_0564_),
    .X(_0568_));
 sg13g2_inv_1 _2220_ (.Y(_0569_),
    .A(net90));
 sg13g2_or2_1 _2221_ (.X(_0570_),
    .B(net88),
    .A(\i2c_bert.i2c.sdaAndNor3.io_b ));
 sg13g2_nor2_1 _2222_ (.A(net91),
    .B(net89),
    .Y(_0571_));
 sg13g2_a22oi_1 _2223_ (.Y(_0572_),
    .B1(_0570_),
    .B2(_0571_),
    .A2(_0547_),
    .A1(_0569_));
 sg13g2_inv_1 _2224_ (.Y(_0573_),
    .A(net14));
 sg13g2_a21oi_1 _2225_ (.A1(_0568_),
    .A2(_0572_),
    .Y(_0574_),
    .B1(_0573_));
 sg13g2_mux2_1 _2226_ (.A0(\i2c_bert.i2c.sdaAndNor3.io_o ),
    .A1(\i2c_bert.i2c.sdaAndNor5.io_o ),
    .S(_0530_),
    .X(_0575_));
 sg13g2_a22oi_1 _2227_ (.Y(_0576_),
    .B1(_0575_),
    .B2(net90),
    .A2(_0531_),
    .A1(net88));
 sg13g2_and2_1 _2228_ (.A(\i2c_bert.i2c.sdaAndNor3.io_b ),
    .B(_0557_),
    .X(_0577_));
 sg13g2_a221oi_1 _2229_ (.B2(_0577_),
    .C1(_0527_),
    .B1(_0535_),
    .A1(_0560_),
    .Y(_0578_),
    .A2(_0533_));
 sg13g2_a21oi_2 _2230_ (.B1(_0578_),
    .Y(_0579_),
    .A2(_0576_),
    .A1(net91));
 sg13g2_nor3_1 _2231_ (.A(_0566_),
    .B(_0574_),
    .C(_0579_),
    .Y(_0580_));
 sg13g2_buf_2 _2232_ (.A(_0580_),
    .X(_0581_));
 sg13g2_inv_2 _2233_ (.Y(\i2c_bert.i2c.io_sdaSignal ),
    .A(_0581_));
 sg13g2_buf_2 _2234_ (.A(_0023_),
    .X(_0582_));
 sg13g2_inv_1 _2235_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_buf_2 _2236_ (.A(\i2c_bert.i2c.fsm_stateReg[1] ),
    .X(_0584_));
 sg13g2_nand2b_1 _2237_ (.Y(_0585_),
    .B(_0584_),
    .A_N(\i2c_bert.i2c.fsm_stateReg[0] ));
 sg13g2_buf_2 _2238_ (.A(\i2c_bert.i2c.fsm_stateReg[2] ),
    .X(_0586_));
 sg13g2_buf_2 _2239_ (.A(\i2c_bert.i2c.fsm_stateReg[3] ),
    .X(_0587_));
 sg13g2_or2_1 _2240_ (.X(_0588_),
    .B(_0587_),
    .A(_0586_));
 sg13g2_buf_1 _2241_ (.A(_0588_),
    .X(_0589_));
 sg13g2_nor2_1 _2242_ (.A(_0585_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_nand2b_1 _2243_ (.Y(_0591_),
    .B(_0590_),
    .A_N(_0020_));
 sg13g2_nor4_2 _2244_ (.A(_0566_),
    .B(_0574_),
    .C(_0579_),
    .Y(_0592_),
    .D(_0591_));
 sg13g2_nand2_2 _2245_ (.Y(_0593_),
    .A(\i2c_bert.i2c.scl ),
    .B(_0592_));
 sg13g2_nand2_1 _2246_ (.Y(_0594_),
    .A(_0583_),
    .B(_0593_));
 sg13g2_or2_1 _2247_ (.X(_0595_),
    .B(_0594_),
    .A(\i2c_bert.i2c.io_wantReset ));
 sg13g2_or2_1 _2248_ (.X(_0596_),
    .B(_0554_),
    .A(\i2c_bert.i2c.scl_regNext ));
 sg13g2_a21oi_2 _2249_ (.B1(_0596_),
    .Y(_0597_),
    .A2(_0551_),
    .A1(_0538_));
 sg13g2_inv_1 _2250_ (.Y(_0598_),
    .A(\i2c_bert.i2c.fsm_stateReg[0] ));
 sg13g2_xnor2_1 _2251_ (.Y(_0599_),
    .A(_0584_),
    .B(_0586_));
 sg13g2_buf_8 _2252_ (.A(\i2c_bert.i2c.fsm_bitCount[0] ),
    .X(_0600_));
 sg13g2_nand3b_1 _2253_ (.B(_0600_),
    .C(\i2c_bert.i2c.fsm_bitCount[1] ),
    .Y(_0601_),
    .A_N(_0018_));
 sg13g2_buf_2 _2254_ (.A(_0601_),
    .X(_0602_));
 sg13g2_nor4_2 _2255_ (.A(_0598_),
    .B(_0587_),
    .C(_0599_),
    .Y(_0603_),
    .D(_0602_));
 sg13g2_nand2_1 _2256_ (.Y(_0604_),
    .A(_0597_),
    .B(_0603_));
 sg13g2_buf_1 _2257_ (.A(_0604_),
    .X(_0605_));
 sg13g2_buf_1 _2258_ (.A(\i2c_bert.myState_1.fsmPhase_stateReg[5] ),
    .X(_0606_));
 sg13g2_buf_1 _2259_ (.A(net87),
    .X(_0607_));
 sg13g2_buf_1 _2260_ (.A(\i2c_bert.myState_1.counter[0] ),
    .X(_0608_));
 sg13g2_buf_1 _2261_ (.A(_0608_),
    .X(_0609_));
 sg13g2_buf_1 _2262_ (.A(\i2c_bert.myState_1.cmd7[3] ),
    .X(_0610_));
 sg13g2_buf_2 _2263_ (.A(\i2c_bert.myState_1.cmd7[4] ),
    .X(_0611_));
 sg13g2_inv_1 _2264_ (.Y(_0612_),
    .A(_0611_));
 sg13g2_buf_2 _2265_ (.A(\i2c_bert.myState_1.alu_1.io_op[0] ),
    .X(_0613_));
 sg13g2_buf_2 _2266_ (.A(\i2c_bert.myState_1.alu_1.io_op[1] ),
    .X(_0614_));
 sg13g2_nor2_2 _2267_ (.A(_0613_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_buf_1 _2268_ (.A(\i2c_bert.myState_1.cmd7[0] ),
    .X(_0616_));
 sg13g2_nand2b_1 _2269_ (.Y(_0617_),
    .B(\i2c_bert.myState_1.cmd7[5] ),
    .A_N(net85));
 sg13g2_nor2_2 _2270_ (.A(_0026_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_nand2_2 _2271_ (.Y(_0619_),
    .A(_0615_),
    .B(_0618_));
 sg13g2_nor3_1 _2272_ (.A(net86),
    .B(_0612_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_buf_1 _2273_ (.A(\i2c_bert.myState_1.counter[1] ),
    .X(_0621_));
 sg13g2_nor2_1 _2274_ (.A(\i2c_bert.myState_1.counter[10] ),
    .B(\i2c_bert.myState_1.counter[11] ),
    .Y(_0622_));
 sg13g2_nor4_1 _2275_ (.A(\i2c_bert.myState_1.counter[6] ),
    .B(\i2c_bert.myState_1.counter[7] ),
    .C(\i2c_bert.myState_1.counter[8] ),
    .D(\i2c_bert.myState_1.counter[9] ),
    .Y(_0623_));
 sg13g2_buf_1 _2276_ (.A(\i2c_bert.myState_1.counter[2] ),
    .X(_0624_));
 sg13g2_buf_2 _2277_ (.A(\i2c_bert.myState_1.counter[3] ),
    .X(_0625_));
 sg13g2_nor4_1 _2278_ (.A(_0624_),
    .B(_0625_),
    .C(\i2c_bert.myState_1.counter[4] ),
    .D(\i2c_bert.myState_1.counter[5] ),
    .Y(_0626_));
 sg13g2_nand3_1 _2279_ (.B(_0623_),
    .C(_0626_),
    .A(_0622_),
    .Y(_0627_));
 sg13g2_nor2_1 _2280_ (.A(_0621_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_and2_1 _2281_ (.A(_0620_),
    .B(_0628_),
    .X(_0629_));
 sg13g2_mux2_1 _2282_ (.A0(\i2c_bert.myState_1.cmd7[6] ),
    .A1(_0026_),
    .S(\i2c_bert.myState_1.cmd7[5] ),
    .X(_0630_));
 sg13g2_nand2_1 _2283_ (.Y(_0631_),
    .A(_0612_),
    .B(_0615_));
 sg13g2_nor4_1 _2284_ (.A(net85),
    .B(net86),
    .C(_0630_),
    .D(_0631_),
    .Y(_0632_));
 sg13g2_xor2_1 _2285_ (.B(_0613_),
    .A(_0611_),
    .X(_0633_));
 sg13g2_inv_2 _2286_ (.Y(_0634_),
    .A(_0613_));
 sg13g2_nand3_1 _2287_ (.B(_0634_),
    .C(_0614_),
    .A(_0611_),
    .Y(_0635_));
 sg13g2_o21ai_1 _2288_ (.B1(_0635_),
    .Y(_0636_),
    .A1(_0614_),
    .A2(_0633_));
 sg13g2_nand3_1 _2289_ (.B(_0636_),
    .C(_0618_),
    .A(net86),
    .Y(_0637_));
 sg13g2_nand2b_1 _2290_ (.Y(_0638_),
    .B(_0637_),
    .A_N(_0632_));
 sg13g2_a21o_1 _2291_ (.A2(_0629_),
    .A1(net67),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_buf_1 _2292_ (.A(\i2c_bert.i2c.io_data8rx[5] ),
    .X(_0640_));
 sg13g2_buf_1 _2293_ (.A(\i2c_bert.i2c.io_data8rx[6] ),
    .X(_0641_));
 sg13g2_nand2_1 _2294_ (.Y(_0642_),
    .A(net84),
    .B(net83));
 sg13g2_buf_1 _2295_ (.A(\i2c_bert.i2c.io_data8rx[1] ),
    .X(_0643_));
 sg13g2_inv_1 _2296_ (.Y(_0644_),
    .A(net82));
 sg13g2_buf_1 _2297_ (.A(\i2c_bert.i2c.io_data8rx[2] ),
    .X(_0645_));
 sg13g2_buf_1 _2298_ (.A(\i2c_bert.i2c.io_data8rx[3] ),
    .X(_0646_));
 sg13g2_and2_1 _2299_ (.A(_0646_),
    .B(\i2c_bert.i2c.io_data8rx[4] ),
    .X(_0647_));
 sg13g2_buf_2 _2300_ (.A(_0647_),
    .X(_0648_));
 sg13g2_buf_1 _2301_ (.A(\i2c_bert.i2c.io_data8rx[4] ),
    .X(_0649_));
 sg13g2_or2_1 _2302_ (.X(_0650_),
    .B(net80),
    .A(net81));
 sg13g2_buf_1 _2303_ (.A(_0650_),
    .X(_0651_));
 sg13g2_o21ai_1 _2304_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_0645_),
    .A2(_0648_));
 sg13g2_or2_1 _2305_ (.X(_0653_),
    .B(_0645_),
    .A(net82));
 sg13g2_a22oi_1 _2306_ (.Y(_0654_),
    .B1(_0653_),
    .B2(_0648_),
    .A2(_0652_),
    .A1(_0644_));
 sg13g2_nor2_1 _2307_ (.A(net81),
    .B(net80),
    .Y(_0655_));
 sg13g2_nor2_1 _2308_ (.A(net82),
    .B(_0645_),
    .Y(_0656_));
 sg13g2_nor2_1 _2309_ (.A(net84),
    .B(net83),
    .Y(_0657_));
 sg13g2_nand3_1 _2310_ (.B(_0656_),
    .C(_0657_),
    .A(_0655_),
    .Y(_0658_));
 sg13g2_o21ai_1 _2311_ (.B1(_0658_),
    .Y(_0659_),
    .A1(_0642_),
    .A2(_0654_));
 sg13g2_and2_1 _2312_ (.A(_0581_),
    .B(_0659_),
    .X(_0660_));
 sg13g2_buf_2 _2313_ (.A(_0027_),
    .X(_0661_));
 sg13g2_and2_1 _2314_ (.A(\i2c_bert.i2c.io_data8rx[5] ),
    .B(net83),
    .X(_0662_));
 sg13g2_buf_1 _2315_ (.A(_0662_),
    .X(_0663_));
 sg13g2_nand2_1 _2316_ (.Y(_0664_),
    .A(_0661_),
    .B(_0663_));
 sg13g2_nand2_1 _2317_ (.Y(_0665_),
    .A(_0645_),
    .B(_0651_));
 sg13g2_a21oi_1 _2318_ (.A1(_0644_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0648_));
 sg13g2_nor3_1 _2319_ (.A(_0581_),
    .B(_0664_),
    .C(_0666_),
    .Y(_0667_));
 sg13g2_nor3_1 _2320_ (.A(\i2c_bert.i2c.io_data8rx[0] ),
    .B(_0660_),
    .C(_0667_),
    .Y(_0668_));
 sg13g2_buf_1 _2321_ (.A(\i2c_bert.myState_1.fsmPhase_stateReg[2] ),
    .X(_0669_));
 sg13g2_inv_1 _2322_ (.Y(_0670_),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[1] ));
 sg13g2_xnor2_1 _2323_ (.Y(_0671_),
    .A(net86),
    .B(_0621_));
 sg13g2_nand2_1 _2324_ (.Y(_0672_),
    .A(_0608_),
    .B(_0671_));
 sg13g2_o21ai_1 _2325_ (.B1(_0611_),
    .Y(_0673_),
    .A1(_0627_),
    .A2(_0672_));
 sg13g2_nand2_2 _2326_ (.Y(_0674_),
    .A(net86),
    .B(_0611_));
 sg13g2_inv_1 _2327_ (.Y(_0675_),
    .A(_0674_));
 sg13g2_buf_1 _2328_ (.A(_0613_),
    .X(_0676_));
 sg13g2_buf_1 _2329_ (.A(_0614_),
    .X(_0677_));
 sg13g2_xor2_1 _2330_ (.B(net65),
    .A(net66),
    .X(_0678_));
 sg13g2_a22oi_1 _2331_ (.Y(_0679_),
    .B1(_0675_),
    .B2(_0678_),
    .A2(_0673_),
    .A1(_0615_));
 sg13g2_nand3_1 _2332_ (.B(\i2c_bert.myState_1.cmd7[5] ),
    .C(\i2c_bert.myState_1.cmd7[6] ),
    .A(\i2c_bert.myState_1.readWriteBit ),
    .Y(_0680_));
 sg13g2_nor4_1 _2333_ (.A(_0670_),
    .B(net85),
    .C(_0679_),
    .D(_0680_),
    .Y(_0681_));
 sg13g2_a221oi_1 _2334_ (.B2(net79),
    .C1(_0681_),
    .B1(_0668_),
    .A1(net68),
    .Y(_0682_),
    .A2(_0639_));
 sg13g2_inv_1 _2335_ (.Y(_0683_),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[3] ));
 sg13g2_o21ai_1 _2336_ (.B1(_0683_),
    .Y(_0684_),
    .A1(net50),
    .A2(_0682_));
 sg13g2_nand2b_1 _2337_ (.Y(_0685_),
    .B(_0684_),
    .A_N(_0595_));
 sg13g2_buf_1 _2338_ (.A(\i2c_bert.i2c.rst_n ),
    .X(_0686_));
 sg13g2_inv_1 _2339_ (.Y(_0687_),
    .A(_0686_));
 sg13g2_and2_1 _2340_ (.A(\i2c_bert.i2c.scl ),
    .B(_0592_),
    .X(_0688_));
 sg13g2_nor4_1 _2341_ (.A(_0687_),
    .B(\i2c_bert.i2c.io_wantReset ),
    .C(_0688_),
    .D(net50),
    .Y(_0689_));
 sg13g2_xnor2_1 _2342_ (.Y(_0690_),
    .A(_0621_),
    .B(_0611_));
 sg13g2_xnor2_1 _2343_ (.Y(_0691_),
    .A(\i2c_bert.myState_1.len12[11] ),
    .B(\i2c_bert.myState_1.counter[11] ));
 sg13g2_xnor2_1 _2344_ (.Y(_0692_),
    .A(\i2c_bert.myState_1.len12[5] ),
    .B(\i2c_bert.myState_1.counter[5] ));
 sg13g2_xnor2_1 _2345_ (.Y(_0693_),
    .A(_0624_),
    .B(\i2c_bert.myState_1.cmd7[5] ));
 sg13g2_nand4_1 _2346_ (.B(_0691_),
    .C(_0692_),
    .A(_0690_),
    .Y(_0694_),
    .D(_0693_));
 sg13g2_xnor2_1 _2347_ (.Y(_0695_),
    .A(\i2c_bert.myState_1.len12[4] ),
    .B(\i2c_bert.myState_1.counter[4] ));
 sg13g2_xnor2_1 _2348_ (.Y(_0696_),
    .A(\i2c_bert.myState_1.len12[7] ),
    .B(\i2c_bert.myState_1.counter[7] ));
 sg13g2_xnor2_1 _2349_ (.Y(_0697_),
    .A(_0625_),
    .B(\i2c_bert.myState_1.cmd7[6] ));
 sg13g2_xnor2_1 _2350_ (.Y(_0698_),
    .A(\i2c_bert.myState_1.len12[9] ),
    .B(\i2c_bert.myState_1.counter[9] ));
 sg13g2_nand4_1 _2351_ (.B(_0696_),
    .C(_0697_),
    .A(_0695_),
    .Y(_0699_),
    .D(_0698_));
 sg13g2_xnor2_1 _2352_ (.Y(_0700_),
    .A(_0608_),
    .B(net86));
 sg13g2_xnor2_1 _2353_ (.Y(_0701_),
    .A(\i2c_bert.myState_1.len12[10] ),
    .B(\i2c_bert.myState_1.counter[10] ));
 sg13g2_xnor2_1 _2354_ (.Y(_0702_),
    .A(\i2c_bert.myState_1.len12[8] ),
    .B(\i2c_bert.myState_1.counter[8] ));
 sg13g2_xnor2_1 _2355_ (.Y(_0703_),
    .A(\i2c_bert.myState_1.len12[6] ),
    .B(\i2c_bert.myState_1.counter[6] ));
 sg13g2_nand4_1 _2356_ (.B(_0701_),
    .C(_0702_),
    .A(_0700_),
    .Y(_0704_),
    .D(_0703_));
 sg13g2_nor3_2 _2357_ (.A(_0694_),
    .B(_0699_),
    .C(_0704_),
    .Y(_0705_));
 sg13g2_or2_1 _2358_ (.X(_0706_),
    .B(net87),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[1] ));
 sg13g2_buf_1 _2359_ (.A(_0706_),
    .X(_0707_));
 sg13g2_nand4_1 _2360_ (.B(_0689_),
    .C(_0705_),
    .A(net85),
    .Y(_0708_),
    .D(_0707_));
 sg13g2_nor2b_1 _2361_ (.A(_0705_),
    .B_N(net85),
    .Y(_0709_));
 sg13g2_inv_1 _2362_ (.Y(_0710_),
    .A(_0614_));
 sg13g2_nand2_1 _2363_ (.Y(_0711_),
    .A(_0634_),
    .B(_0710_));
 sg13g2_nor4_1 _2364_ (.A(_0582_),
    .B(net85),
    .C(_0711_),
    .D(_0680_),
    .Y(_0712_));
 sg13g2_nor2b_1 _2365_ (.A(_0673_),
    .B_N(_0712_),
    .Y(_0713_));
 sg13g2_a21oi_1 _2366_ (.A1(net78),
    .A2(_0709_),
    .Y(_0714_),
    .B1(_0713_));
 sg13g2_and2_1 _2367_ (.A(_0597_),
    .B(_0603_),
    .X(_0715_));
 sg13g2_buf_1 _2368_ (.A(_0715_),
    .X(_0716_));
 sg13g2_o21ai_1 _2369_ (.B1(net49),
    .Y(_0717_),
    .A1(_0688_),
    .A2(_0714_));
 sg13g2_nand2_2 _2370_ (.Y(_0718_),
    .A(_0676_),
    .B(net65));
 sg13g2_a21oi_1 _2371_ (.A1(_0711_),
    .A2(_0674_),
    .Y(_0719_),
    .B1(_0680_));
 sg13g2_a21oi_1 _2372_ (.A1(_0718_),
    .A2(_0719_),
    .Y(_0720_),
    .B1(_0616_));
 sg13g2_nand3_1 _2373_ (.B(_0593_),
    .C(_0720_),
    .A(net78),
    .Y(_0721_));
 sg13g2_nor3_1 _2374_ (.A(\i2c_bert.i2c.io_wantReset ),
    .B(net50),
    .C(_0721_),
    .Y(_0722_));
 sg13g2_a21o_1 _2375_ (.A2(_0717_),
    .A1(_0025_),
    .B1(_0722_),
    .X(_0723_));
 sg13g2_nand2_1 _2376_ (.Y(_0724_),
    .A(_0594_),
    .B(net50));
 sg13g2_buf_1 _2377_ (.A(\i2c_bert.i2c.io_canStretch ),
    .X(_0725_));
 sg13g2_or2_1 _2378_ (.X(_0726_),
    .B(\i2c_bert.myState_1.fsmPhase_stateReg[2] ),
    .A(net87));
 sg13g2_nor3_1 _2379_ (.A(net77),
    .B(\i2c_bert.myState_1.fsmPhase_stateReg[1] ),
    .C(_0726_),
    .Y(_0727_));
 sg13g2_o21ai_1 _2380_ (.B1(_0727_),
    .Y(_0728_),
    .A1(\i2c_bert.myState_1.readWriteBit ),
    .A2(_0683_));
 sg13g2_nand2b_1 _2381_ (.Y(_0729_),
    .B(_0586_),
    .A_N(_0587_));
 sg13g2_buf_2 _2382_ (.A(_0729_),
    .X(_0730_));
 sg13g2_or2_1 _2383_ (.X(_0731_),
    .B(\i2c_bert.i2c.fsm_stateReg[0] ),
    .A(_0584_));
 sg13g2_buf_1 _2384_ (.A(_0731_),
    .X(_0732_));
 sg13g2_nor2_2 _2385_ (.A(_0730_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nand2b_1 _2386_ (.Y(_0734_),
    .B(_0733_),
    .A_N(_0728_));
 sg13g2_buf_1 _2387_ (.A(_0584_),
    .X(_0735_));
 sg13g2_buf_1 _2388_ (.A(\i2c_bert.i2c.fsm_stateReg[0] ),
    .X(_0736_));
 sg13g2_nor2b_2 _2389_ (.A(_0587_),
    .B_N(_0586_),
    .Y(_0737_));
 sg13g2_nand3_1 _2390_ (.B(net76),
    .C(_0737_),
    .A(_0735_),
    .Y(_0738_));
 sg13g2_inv_1 _2391_ (.Y(_0739_),
    .A(_0738_));
 sg13g2_nand2_1 _2392_ (.Y(_0740_),
    .A(\i2c_bert.i2c.io_sdaSignal ),
    .B(_0739_));
 sg13g2_a21o_1 _2393_ (.A2(_0551_),
    .A1(_0538_),
    .B1(_0596_),
    .X(_0741_));
 sg13g2_buf_8 _2394_ (.A(_0741_),
    .X(_0742_));
 sg13g2_a21oi_1 _2395_ (.A1(_0734_),
    .A2(_0740_),
    .Y(_0743_),
    .B1(net53));
 sg13g2_nand4_1 _2396_ (.B(_0723_),
    .C(_0724_),
    .A(\i2c_bert.myState_1.fsmPhase_stateReg[1] ),
    .Y(_0744_),
    .D(_0743_));
 sg13g2_nand3_1 _2397_ (.B(_0708_),
    .C(_0744_),
    .A(_0685_),
    .Y(_0003_));
 sg13g2_inv_1 _2398_ (.Y(_0745_),
    .A(\i2c_bert.i2c.io_canStretch ));
 sg13g2_or3_1 _2399_ (.A(_0745_),
    .B(\i2c_bert.i2c.io_wantReset ),
    .C(_0705_),
    .X(_0746_));
 sg13g2_buf_1 _2400_ (.A(_0645_),
    .X(_0747_));
 sg13g2_nand2_1 _2401_ (.Y(_0748_),
    .A(_0025_),
    .B(net63));
 sg13g2_nor4_1 _2402_ (.A(net82),
    .B(_0642_),
    .C(_0651_),
    .D(_0748_),
    .Y(_0749_));
 sg13g2_buf_1 _2403_ (.A(\i2c_bert.i2c.io_data8rx[0] ),
    .X(_0750_));
 sg13g2_nand2_1 _2404_ (.Y(_0751_),
    .A(_0661_),
    .B(\i2c_bert.i2c.io_sdaSignal ));
 sg13g2_o21ai_1 _2405_ (.B1(_0751_),
    .Y(_0752_),
    .A1(net75),
    .A2(\i2c_bert.i2c.io_sdaSignal ));
 sg13g2_nand4_1 _2406_ (.B(net49),
    .C(_0749_),
    .A(net79),
    .Y(_0753_),
    .D(_0752_));
 sg13g2_a21oi_1 _2407_ (.A1(_0746_),
    .A2(_0753_),
    .Y(_0004_),
    .B1(_0594_));
 sg13g2_buf_1 _2408_ (.A(_0581_),
    .X(\i2c_bert.powerOnSense.D ));
 sg13g2_and3_1 _2409_ (.X(_0754_),
    .A(_0669_),
    .B(net52),
    .C(_0716_));
 sg13g2_inv_1 _2410_ (.Y(_0755_),
    .A(_0750_));
 sg13g2_nand2b_1 _2411_ (.Y(_0756_),
    .B(_0657_),
    .A_N(net80));
 sg13g2_a21oi_1 _2412_ (.A1(_0642_),
    .A2(_0756_),
    .Y(_0757_),
    .B1(net81));
 sg13g2_nor2_1 _2413_ (.A(net80),
    .B(_0642_),
    .Y(_0758_));
 sg13g2_o21ai_1 _2414_ (.B1(_0656_),
    .Y(_0759_),
    .A1(_0757_),
    .A2(_0758_));
 sg13g2_nand3_1 _2415_ (.B(_0648_),
    .C(_0653_),
    .A(_0663_),
    .Y(_0760_));
 sg13g2_nand3_1 _2416_ (.B(_0759_),
    .C(_0760_),
    .A(_0755_),
    .Y(_0761_));
 sg13g2_buf_1 _2417_ (.A(net77),
    .X(_0762_));
 sg13g2_and2_1 _2418_ (.A(net62),
    .B(_0705_),
    .X(_0763_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2428__110 (.L_HI(net110));
 sg13g2_buf_1 _2421_ (.A(net100),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2422_ (.A(net101),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2423_ (.A(\i2c_bert.i2c.io_bus_sclOe ),
    .X(net19));
 sg13g2_buf_1 _2424_ (.A(\i2c_bert.i2c.io_bus_sdaOe ),
    .X(net20));
 sg13g2_buf_1 _2425_ (.A(net102),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2426_ (.A(net103),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2427_ (.A(net104),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2428_ (.A(net110),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2429_ (.A(net105),
    .X(uio_out[0]));
 sg13g2_buf_1 _2430_ (.A(net106),
    .X(uio_out[1]));
 sg13g2_buf_1 _2431_ (.A(\i2c_bert.i2c.io_bus_sclOut ),
    .X(net21));
 sg13g2_buf_1 _2432_ (.A(\i2c_bert.i2c.io_bus_sdaOut ),
    .X(net22));
 sg13g2_buf_1 _2433_ (.A(net107),
    .X(uio_out[4]));
 sg13g2_buf_1 _2434_ (.A(net108),
    .X(uio_out[5]));
 sg13g2_buf_1 _2435_ (.A(net109),
    .X(uio_out[6]));
 sg13g2_buf_1 _2436_ (.A(\i2c_bert.powerOnSense.Q ),
    .X(net23));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_bitCount[0]$_SDFFE_PP0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net111),
    .D(_0032_),
    .Q_N(_1249_),
    .Q(\i2c_bert.i2c.fsm_bitCount[0] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_bitCount[1]$_SDFFE_PP0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net112),
    .D(_0033_),
    .Q_N(_1248_),
    .Q(\i2c_bert.i2c.fsm_bitCount[1] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_bitCount[2]$_SDFFE_PP0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net113),
    .D(_0034_),
    .Q_N(_0018_),
    .Q(\i2c_bert.i2c.fsm_bitCount[2] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_stateReg[0]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net114),
    .D(_0035_),
    .Q_N(_0028_),
    .Q(\i2c_bert.i2c.fsm_stateReg[0] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_stateReg[1]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net115),
    .D(_0036_),
    .Q_N(_0022_),
    .Q(\i2c_bert.i2c.fsm_stateReg[1] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_stateReg[2]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net116),
    .D(_0037_),
    .Q_N(_0024_),
    .Q(\i2c_bert.i2c.fsm_stateReg[2] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_stateReg[3]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net117),
    .D(_0038_),
    .Q_N(_0017_),
    .Q(\i2c_bert.i2c.fsm_stateReg[3] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.fsm_wantStart$_DFF_P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net118),
    .D(_0000_),
    .Q_N(_0021_),
    .Q(\i2c_bert.i2c.fsm_wantStart ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.io_wantReset$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net119),
    .D(_0039_),
    .Q_N(_0025_),
    .Q(\i2c_bert.i2c.io_wantReset ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclAndNor3.state$_SDFFE_PP0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net120),
    .D(_0040_),
    .Q_N(_1247_),
    .Q(\i2c_bert.i2c.sclAndNor3.io_o ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclAndNor5.state$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net121),
    .D(_0041_),
    .Q_N(_1246_),
    .Q(\i2c_bert.i2c.sclAndNor5.io_o ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclHistory5_1$_DFFE_PP_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net122),
    .D(_0042_),
    .Q_N(_1245_),
    .Q(\i2c_bert.i2c.sclAndNor3.io_b ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclHistory5_2$_DFFE_PP_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net123),
    .D(_0043_),
    .Q_N(_1244_),
    .Q(\i2c_bert.i2c.sclAndNor3.io_c ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclHistory5_3$_DFFE_PP_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net124),
    .D(_0044_),
    .Q_N(_1243_),
    .Q(\i2c_bert.i2c.sclAndNor5.io_d ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sclHistory5_4$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net125),
    .D(_0045_),
    .Q_N(_1250_),
    .Q(\i2c_bert.i2c.sclAndNor5.io_e ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.scl_regNext$_DFF_P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net126),
    .D(\i2c_bert.i2c.scl ),
    .Q_N(_1242_),
    .Q(\i2c_bert.i2c.scl_regNext ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaAndNor3.state$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net127),
    .D(_0046_),
    .Q_N(_1241_),
    .Q(\i2c_bert.i2c.sdaAndNor3.io_o ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaAndNor5.state$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net128),
    .D(_0047_),
    .Q_N(_1240_),
    .Q(\i2c_bert.i2c.sdaAndNor5.io_o ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaHistory5_1$_DFFE_PP_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net129),
    .D(_0048_),
    .Q_N(_1239_),
    .Q(\i2c_bert.i2c.sdaAndNor3.io_b ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaHistory5_2$_DFFE_PP_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net130),
    .D(_0049_),
    .Q_N(_1238_),
    .Q(\i2c_bert.i2c.sdaAndNor3.io_c ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaHistory5_3$_DFFE_PP_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net131),
    .D(_0050_),
    .Q_N(_1237_),
    .Q(\i2c_bert.i2c.sdaAndNor5.io_d ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sdaHistory5_4$_DFFE_PP_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net132),
    .D(_0051_),
    .Q_N(_1251_),
    .Q(\i2c_bert.i2c.sdaAndNor5.io_e ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.sda_regNext$_DFF_P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net133),
    .D(\i2c_bert.i2c.io_sdaSignal ),
    .Q_N(_0020_),
    .Q(\i2c_bert.i2c.sda_regNext ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[0]$_DFFE_PP_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net134),
    .D(_0052_),
    .Q_N(_0027_),
    .Q(\i2c_bert.i2c.io_data8rx[0] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[1]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net135),
    .D(_0053_),
    .Q_N(_0010_),
    .Q(\i2c_bert.i2c.io_data8rx[1] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[2]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net136),
    .D(_0054_),
    .Q_N(_0011_),
    .Q(\i2c_bert.i2c.io_data8rx[2] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[3]$_DFFE_PP_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net137),
    .D(_0055_),
    .Q_N(_0012_),
    .Q(\i2c_bert.i2c.io_data8rx[3] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[4]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0056_),
    .Q_N(_0013_),
    .Q(\i2c_bert.i2c.io_data8rx[4] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[5]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net139),
    .D(_0057_),
    .Q_N(_0015_),
    .Q(\i2c_bert.i2c.io_data8rx[5] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[6]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net140),
    .D(_0058_),
    .Q_N(_0009_),
    .Q(\i2c_bert.i2c.io_data8rx[6] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.shifter[7]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net141),
    .D(_0059_),
    .Q_N(_1236_),
    .Q(\i2c_bert.i2c.io_data8rx[7] ));
 sg13g2_dfrbp_1 \i2c_bert.i2c.timerAutobaud$_SDFFE_PP0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net142),
    .D(_0060_),
    .Q_N(_1235_),
    .Q(\i2c_bert.i2c.io_timerAutobaud ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[0]$_SDFFE_PP0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net143),
    .D(_0061_),
    .Q_N(_1234_),
    .Q(\i2c_bert.myState_1.alu_1.acc[0] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[1]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net144),
    .D(_0062_),
    .Q_N(_1233_),
    .Q(\i2c_bert.myState_1.alu_1.acc[1] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[2]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(_0063_),
    .Q_N(_1232_),
    .Q(\i2c_bert.myState_1.alu_1.acc[2] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[3]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net146),
    .D(_0064_),
    .Q_N(_1231_),
    .Q(\i2c_bert.myState_1.alu_1.acc[3] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[4]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net147),
    .D(_0065_),
    .Q_N(_1230_),
    .Q(\i2c_bert.myState_1.alu_1.acc[4] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[5]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net148),
    .D(_0066_),
    .Q_N(_1229_),
    .Q(\i2c_bert.myState_1.alu_1.acc[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[6]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net149),
    .D(_0067_),
    .Q_N(_0014_),
    .Q(\i2c_bert.myState_1.alu_1.acc[6] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.alu_1.acc[7]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net150),
    .D(_0068_),
    .Q_N(_0016_),
    .Q(\i2c_bert.myState_1.alu_1.acc[7] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net151),
    .D(_0069_),
    .Q_N(_0031_),
    .Q(\i2c_bert.myState_1.cmd7[0] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net152),
    .D(_0070_),
    .Q_N(_1228_),
    .Q(\i2c_bert.myState_1.alu_1.io_op[0] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[2]$_SDFFCE_PP1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net153),
    .D(_0071_),
    .Q_N(_1227_),
    .Q(\i2c_bert.myState_1.alu_1.io_op[1] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[3]$_SDFFCE_PP1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net154),
    .D(_0072_),
    .Q_N(_1226_),
    .Q(\i2c_bert.myState_1.cmd7[3] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[4]$_SDFFCE_PP1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net155),
    .D(_0073_),
    .Q_N(_1225_),
    .Q(\i2c_bert.myState_1.cmd7[4] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[5]$_SDFFCE_PP1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net156),
    .D(_0074_),
    .Q_N(_1224_),
    .Q(\i2c_bert.myState_1.cmd7[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.cmd7[6]$_SDFFCE_PP1P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net157),
    .D(_0075_),
    .Q_N(_0026_),
    .Q(\i2c_bert.myState_1.cmd7[6] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[0]$_SDFFE_PN1P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net158),
    .D(_0076_),
    .Q_N(_1223_),
    .Q(\i2c_bert.myState_1.counter[0] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[10]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net159),
    .D(_0077_),
    .Q_N(_1222_),
    .Q(\i2c_bert.myState_1.counter[10] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[11]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net160),
    .D(_0078_),
    .Q_N(_1221_),
    .Q(\i2c_bert.myState_1.counter[11] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net161),
    .D(_0079_),
    .Q_N(_1220_),
    .Q(\i2c_bert.myState_1.counter[1] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net162),
    .D(_0080_),
    .Q_N(_1219_),
    .Q(\i2c_bert.myState_1.counter[2] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net163),
    .D(_0081_),
    .Q_N(_1218_),
    .Q(\i2c_bert.myState_1.counter[3] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net164),
    .D(_0082_),
    .Q_N(_1217_),
    .Q(\i2c_bert.myState_1.counter[4] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net165),
    .D(_0083_),
    .Q_N(_1216_),
    .Q(\i2c_bert.myState_1.counter[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net166),
    .D(_0084_),
    .Q_N(_1215_),
    .Q(\i2c_bert.myState_1.counter[6] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net167),
    .D(_0085_),
    .Q_N(_1214_),
    .Q(\i2c_bert.myState_1.counter[7] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net168),
    .D(_0086_),
    .Q_N(_1213_),
    .Q(\i2c_bert.myState_1.counter[8] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.counter[9]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net169),
    .D(_0087_),
    .Q_N(_1252_),
    .Q(\i2c_bert.myState_1.counter[9] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.fsmPhase_stateReg[1]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net170),
    .D(_0001_),
    .Q_N(_1253_),
    .Q(\i2c_bert.myState_1.fsmPhase_stateReg[1] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.fsmPhase_stateReg[2]$_DFF_P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net171),
    .D(_0002_),
    .Q_N(_0029_),
    .Q(\i2c_bert.myState_1.fsmPhase_stateReg[2] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.fsmPhase_stateReg[3]$_DFF_P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net172),
    .D(_0003_),
    .Q_N(_1254_),
    .Q(\i2c_bert.myState_1.fsmPhase_stateReg[3] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.fsmPhase_stateReg[4]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net173),
    .D(_0004_),
    .Q_N(_0019_),
    .Q(\i2c_bert.i2c.io_canStretch ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.fsmPhase_stateReg[5]$_DFF_P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net174),
    .D(_0005_),
    .Q_N(_0030_),
    .Q(\i2c_bert.myState_1.fsmPhase_stateReg[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[0]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net175),
    .D(_0088_),
    .Q_N(_1212_),
    .Q(\i2c_bert.myState_1.led8[0] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[1]$_DFFE_PP_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net176),
    .D(_0089_),
    .Q_N(_1211_),
    .Q(\i2c_bert.myState_1.led8[1] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[2]$_DFFE_PP_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net177),
    .D(_0090_),
    .Q_N(_1210_),
    .Q(\i2c_bert.myState_1.led8[2] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[3]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net178),
    .D(_0091_),
    .Q_N(_1209_),
    .Q(\i2c_bert.myState_1.led8[3] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[4]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net179),
    .D(_0092_),
    .Q_N(_1208_),
    .Q(\i2c_bert.myState_1.led8[4] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[5]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net180),
    .D(_0093_),
    .Q_N(_1207_),
    .Q(\i2c_bert.myState_1.led8[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[6]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net181),
    .D(_0094_),
    .Q_N(_1206_),
    .Q(\i2c_bert.myState_1.led8[6] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.led8[7]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net182),
    .D(_0095_),
    .Q_N(_1205_),
    .Q(\i2c_bert.myState_1.led8[7] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[0]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net183),
    .D(_0096_),
    .Q_N(_1204_),
    .Q(\i2c_bert.myState_1.len12[4] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[1]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net184),
    .D(_0097_),
    .Q_N(_1203_),
    .Q(\i2c_bert.myState_1.len12[5] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[2]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net185),
    .D(_0098_),
    .Q_N(_1202_),
    .Q(\i2c_bert.myState_1.len12[6] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[3]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net186),
    .D(_0099_),
    .Q_N(_1201_),
    .Q(\i2c_bert.myState_1.len12[7] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[4]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net187),
    .D(_0100_),
    .Q_N(_1200_),
    .Q(\i2c_bert.myState_1.len12[8] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[5]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net188),
    .D(_0101_),
    .Q_N(_1199_),
    .Q(\i2c_bert.myState_1.len12[9] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[6]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net189),
    .D(_0102_),
    .Q_N(_1198_),
    .Q(\i2c_bert.myState_1.len12[10] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.len8[7]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net190),
    .D(_0103_),
    .Q_N(_1197_),
    .Q(\i2c_bert.myState_1.len12[11] ));
 sg13g2_dfrbp_1 \i2c_bert.myState_1.readWriteBit$_DFFE_PP_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net191),
    .D(_0104_),
    .Q_N(_1196_),
    .Q(\i2c_bert.myState_1.readWriteBit ));
 sg13g2_dlhrq_1 \i2c_bert.powerOnSense.genblk1.dlhrq_1  (.D(net52),
    .GATE(\i2c_bert.powerOnSense.GATE ),
    .RESET_B(\i2c_bert.i2c.rst_n ),
    .Q(\i2c_bert.powerOnSense.Q ));
 sg13g2_dlhrq_1 \i2c_bert.powerOnSenseCaptured.genblk1.dlhrq_1  (.D(net192),
    .GATE(\i2c_bert.powerOnSenseCaptured.GATE ),
    .RESET_B(\i2c_bert.i2c.rst_n ),
    .Q(\i2c_bert.powerOnSenseCaptured.Q ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[0]$_DFFE_PP_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net193),
    .D(_0105_),
    .Q_N(_1195_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[0] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[10]$_DFFE_PP_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net194),
    .D(_0106_),
    .Q_N(_1194_),
    .Q(\i2c_bert.myState_1._zz__zz_io_data8tx[2] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[11]$_DFFE_PP_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net195),
    .D(_0107_),
    .Q_N(_1193_),
    .Q(\i2c_bert.myState_1._zz__zz_io_data8tx[3] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[1]$_DFFE_PP_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net196),
    .D(_0108_),
    .Q_N(_1192_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[1] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[2]$_DFFE_PP_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net197),
    .D(_0109_),
    .Q_N(_1191_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[2] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[3]$_DFFE_PP_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net198),
    .D(_0110_),
    .Q_N(_1190_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[3] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[4]$_DFFE_PP_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net199),
    .D(_0111_),
    .Q_N(_1189_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[4] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[5]$_DFFE_PP_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net200),
    .D(_0112_),
    .Q_N(_1188_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[5] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[6]$_DFFE_PP_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net201),
    .D(_0113_),
    .Q_N(_1187_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[6] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[7]$_DFFE_PP_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net202),
    .D(_0114_),
    .Q_N(_1186_),
    .Q(\i2c_bert.myState_1.io_timerEndstop[7] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[8]$_DFFE_PP_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net203),
    .D(_0115_),
    .Q_N(_1185_),
    .Q(\i2c_bert.myState_1._zz__zz_io_data8tx[0] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.endstop[9]$_DFFE_PP_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net204),
    .D(_0116_),
    .Q_N(_1184_),
    .Q(\i2c_bert.myState_1._zz__zz_io_data8tx[1] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[0]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(_0117_),
    .Q_N(_0007_),
    .Q(\i2c_bert.timer_1.ticker_count[0] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[10]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net206),
    .D(_0118_),
    .Q_N(_1183_),
    .Q(\i2c_bert.timer_1.ticker_count[10] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[11]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net207),
    .D(_0119_),
    .Q_N(_1182_),
    .Q(\i2c_bert.timer_1.ticker_count[11] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[1]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net208),
    .D(_0120_),
    .Q_N(_1181_),
    .Q(\i2c_bert.timer_1.ticker_count[1] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[2]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net209),
    .D(_0121_),
    .Q_N(_0008_),
    .Q(\i2c_bert.timer_1.ticker_count[2] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[3]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net210),
    .D(_0122_),
    .Q_N(_0006_),
    .Q(\i2c_bert.timer_1.ticker_count[3] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[4]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net211),
    .D(_0123_),
    .Q_N(_1180_),
    .Q(\i2c_bert.timer_1.ticker_count[4] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[5]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net212),
    .D(_0124_),
    .Q_N(_1179_),
    .Q(\i2c_bert.timer_1.ticker_count[5] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[6]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net213),
    .D(_0125_),
    .Q_N(_1178_),
    .Q(\i2c_bert.timer_1.ticker_count[6] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[7]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net214),
    .D(_0126_),
    .Q_N(_1177_),
    .Q(\i2c_bert.timer_1.ticker_count[7] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[8]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net215),
    .D(_0127_),
    .Q_N(_1176_),
    .Q(\i2c_bert.timer_1.ticker_count[8] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_count[9]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net216),
    .D(_0128_),
    .Q_N(_1175_),
    .Q(\i2c_bert.timer_1.ticker_count[9] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[0]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net217),
    .D(_0129_),
    .Q_N(_1174_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[0] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[1]$_DFFE_PP_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net218),
    .D(_0130_),
    .Q_N(_1173_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[1] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[2]$_DFFE_PP_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net219),
    .D(_0131_),
    .Q_N(_1172_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[2] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[3]$_DFFE_PP_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net220),
    .D(_0132_),
    .Q_N(_1171_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[3] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[4]$_DFFE_PP_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net221),
    .D(_0133_),
    .Q_N(_1170_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[4] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[5]$_DFFE_PP_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net222),
    .D(_0134_),
    .Q_N(_1169_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[5] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[6]$_DFFE_PP_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net223),
    .D(_0135_),
    .Q_N(_1168_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[6] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_endstopTmpL[7]$_DFFE_PP_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net224),
    .D(_0136_),
    .Q_N(_1255_),
    .Q(\i2c_bert.timer_1.ticker_endstopTmpL[7] ));
 sg13g2_dfrbp_1 \i2c_bert.timer_1.ticker_timerSampleTickState_regNext$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net225),
    .D(\i2c_bert.timer_1.ticker_timerSampleTickState ),
    .Q_N(_1256_),
    .Q(\i2c_bert.timer_1.ticker_timerSampleTickState_regNext ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net3),
    .GATE_N(net98),
    .RESET_B(net226),
    .Q(\i2c_bert.latched[16] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net4),
    .GATE_N(net98),
    .RESET_B(net227),
    .Q(\i2c_bert.latched[17] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net5),
    .GATE_N(net98),
    .RESET_B(net228),
    .Q(\i2c_bert.latched[18] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net6),
    .GATE_N(net99),
    .RESET_B(net229),
    .Q(\i2c_bert.latched[19] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net7),
    .GATE_N(net99),
    .RESET_B(net230),
    .Q(\i2c_bert.latched[20] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net8),
    .GATE_N(net99),
    .RESET_B(net231),
    .Q(\i2c_bert.latched[21] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net9),
    .GATE_N(net98),
    .RESET_B(net232),
    .Q(\i2c_bert.latched[22] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_ui_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net10),
    .GATE_N(net99),
    .RESET_B(net233),
    .Q(\i2c_bert.latched[23] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net11),
    .GATE_N(net98),
    .RESET_B(net234),
    .Q(\i2c_bert.latched[24] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net12),
    .GATE_N(net98),
    .RESET_B(net235),
    .Q(\i2c_bert.latched[25] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net13),
    .GATE_N(net98),
    .RESET_B(net236),
    .Q(\i2c_bert.latched[26] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net14),
    .GATE_N(net99),
    .RESET_B(net237),
    .Q(\i2c_bert.latched[27] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net15),
    .GATE_N(net99),
    .RESET_B(net238),
    .Q(\i2c_bert.latched[28] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net16),
    .GATE_N(net99),
    .RESET_B(net239),
    .Q(\i2c_bert.latched[29] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net17),
    .GATE_N(net98),
    .RESET_B(net240),
    .Q(\i2c_bert.latched[30] ));
 sg13g2_dllrq_1 \latched_config.latched_ena_uio_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net18),
    .GATE_N(net99),
    .RESET_B(net241),
    .Q(\i2c_bert.latched[31] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net3),
    .GATE_N(net96),
    .RESET_B(net242),
    .Q(\i2c_bert.i2c.clockGate.sel ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net4),
    .GATE_N(net97),
    .RESET_B(net243),
    .Q(\i2c_bert.i2c.io_sclMode[1] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net5),
    .GATE_N(net97),
    .RESET_B(net244),
    .Q(\i2c_bert.i2c.io_sclMode[2] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net6),
    .GATE_N(net96),
    .RESET_B(net245),
    .Q(\i2c_bert.i2c.io_pushPullMode ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net7),
    .GATE_N(net96),
    .RESET_B(net246),
    .Q(\i2c_bert.div12[0] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net8),
    .GATE_N(net96),
    .RESET_B(net247),
    .Q(\i2c_bert.div12[1] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net9),
    .GATE_N(net97),
    .RESET_B(net248),
    .Q(\i2c_bert.div12[2] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_ui_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net10),
    .GATE_N(net96),
    .RESET_B(net249),
    .Q(\i2c_bert.div12[3] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net11),
    .GATE_N(net97),
    .RESET_B(net250),
    .Q(\i2c_bert.div12[4] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net12),
    .GATE_N(net97),
    .RESET_B(net251),
    .Q(\i2c_bert.div12[5] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net13),
    .GATE_N(net97),
    .RESET_B(net252),
    .Q(\i2c_bert.div12[6] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net14),
    .GATE_N(net2),
    .RESET_B(net253),
    .Q(\i2c_bert.div12[7] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net15),
    .GATE_N(net96),
    .RESET_B(net254),
    .Q(\i2c_bert.div12[8] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net16),
    .GATE_N(net96),
    .RESET_B(net255),
    .Q(\i2c_bert.div12[9] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net17),
    .GATE_N(net97),
    .RESET_B(net256),
    .Q(\i2c_bert.div12[10] ));
 sg13g2_dllrq_1 \latched_config.latched_rst_n_uio_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(net18),
    .GATE_N(net96),
    .RESET_B(net257),
    .Q(\i2c_bert.div12[11] ));
 sg13g2_dfrbp_1 \rst_n_sync$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net258),
    .D(net97),
    .Q_N(_0023_),
    .Q(\i2c_bert.i2c.rst_n ));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[6]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(uio_in[7]),
    .X(net18));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[7]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[0]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[1]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[2]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[3]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[4]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[5]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[6]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout32 (.A(_0480_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0451_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0412_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1136_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1122_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1060_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0405_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0223_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0198_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0185_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0153_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1126_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1125_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1124_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1123_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1039_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0940_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0716_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0605_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0192_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(\i2c_bert.powerOnSense.D ),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0742_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0211_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0829_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0953_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0929_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0956_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0389_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0208_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1041_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0762_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0747_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0735_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0677_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0676_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0609_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0607_),
    .X(net68));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(_0958_));
 sg13g2_buf_2 fanout70 (.A(_0839_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0821_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0787_),
    .X(net72));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_0768_));
 sg13g2_buf_2 fanout74 (.A(_0766_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0750_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0736_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0725_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0686_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0669_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0649_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0646_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0643_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0641_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0640_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0616_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0610_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0606_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0557_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0530_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0528_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0527_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1000_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0976_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0966_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0941_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net2),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(net2),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net1),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net1),
    .X(net99));
 sg13g2_tielo _2421__100 (.L_LO(net100));
 sg13g2_tielo _2422__101 (.L_LO(net101));
 sg13g2_tielo _2425__102 (.L_LO(net102));
 sg13g2_tielo _2426__103 (.L_LO(net103));
 sg13g2_tielo _2427__104 (.L_LO(net104));
 sg13g2_tielo _2429__105 (.L_LO(net105));
 sg13g2_tielo _2430__106 (.L_LO(net106));
 sg13g2_tielo _2433__107 (.L_LO(net107));
 sg13g2_tielo _2434__108 (.L_LO(net108));
 sg13g2_tielo _2435__109 (.L_LO(net109));
 sg13g2_tiehi \i2c_bert.i2c.fsm_bitCount[0]$_SDFFE_PP0P__111  (.L_HI(net111));
 sg13g2_tiehi \i2c_bert.i2c.fsm_bitCount[1]$_SDFFE_PP0P__112  (.L_HI(net112));
 sg13g2_tiehi \i2c_bert.i2c.fsm_bitCount[2]$_SDFFE_PP0P__113  (.L_HI(net113));
 sg13g2_tiehi \i2c_bert.i2c.fsm_stateReg[0]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \i2c_bert.i2c.fsm_stateReg[1]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \i2c_bert.i2c.fsm_stateReg[2]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \i2c_bert.i2c.fsm_stateReg[3]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \i2c_bert.i2c.fsm_wantStart$_DFF_P__118  (.L_HI(net118));
 sg13g2_tiehi \i2c_bert.i2c.io_wantReset$_SDFF_PP0__119  (.L_HI(net119));
 sg13g2_tiehi \i2c_bert.i2c.sclAndNor3.state$_SDFFE_PP0P__120  (.L_HI(net120));
 sg13g2_tiehi \i2c_bert.i2c.sclAndNor5.state$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \i2c_bert.i2c.sclHistory5_1$_DFFE_PP__122  (.L_HI(net122));
 sg13g2_tiehi \i2c_bert.i2c.sclHistory5_2$_DFFE_PP__123  (.L_HI(net123));
 sg13g2_tiehi \i2c_bert.i2c.sclHistory5_3$_DFFE_PP__124  (.L_HI(net124));
 sg13g2_tiehi \i2c_bert.i2c.sclHistory5_4$_DFFE_PP__125  (.L_HI(net125));
 sg13g2_tiehi \i2c_bert.i2c.scl_regNext$_DFF_P__126  (.L_HI(net126));
 sg13g2_tiehi \i2c_bert.i2c.sdaAndNor3.state$_SDFFE_PN0N__127  (.L_HI(net127));
 sg13g2_tiehi \i2c_bert.i2c.sdaAndNor5.state$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \i2c_bert.i2c.sdaHistory5_1$_DFFE_PP__129  (.L_HI(net129));
 sg13g2_tiehi \i2c_bert.i2c.sdaHistory5_2$_DFFE_PP__130  (.L_HI(net130));
 sg13g2_tiehi \i2c_bert.i2c.sdaHistory5_3$_DFFE_PP__131  (.L_HI(net131));
 sg13g2_tiehi \i2c_bert.i2c.sdaHistory5_4$_DFFE_PP__132  (.L_HI(net132));
 sg13g2_tiehi \i2c_bert.i2c.sda_regNext$_DFF_P__133  (.L_HI(net133));
 sg13g2_tiehi \i2c_bert.i2c.shifter[0]$_DFFE_PP__134  (.L_HI(net134));
 sg13g2_tiehi \i2c_bert.i2c.shifter[1]$_DFFE_PP__135  (.L_HI(net135));
 sg13g2_tiehi \i2c_bert.i2c.shifter[2]$_DFFE_PP__136  (.L_HI(net136));
 sg13g2_tiehi \i2c_bert.i2c.shifter[3]$_DFFE_PP__137  (.L_HI(net137));
 sg13g2_tiehi \i2c_bert.i2c.shifter[4]$_DFFE_PP__138  (.L_HI(net138));
 sg13g2_tiehi \i2c_bert.i2c.shifter[5]$_DFFE_PP__139  (.L_HI(net139));
 sg13g2_tiehi \i2c_bert.i2c.shifter[6]$_DFFE_PP__140  (.L_HI(net140));
 sg13g2_tiehi \i2c_bert.i2c.shifter[7]$_DFFE_PP__141  (.L_HI(net141));
 sg13g2_tiehi \i2c_bert.i2c.timerAutobaud$_SDFFE_PP0P__142  (.L_HI(net142));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[0]$_SDFFE_PP0P__143  (.L_HI(net143));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[1]$_SDFFE_PP0P__144  (.L_HI(net144));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[2]$_SDFFE_PP0P__145  (.L_HI(net145));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[3]$_SDFFE_PP0P__146  (.L_HI(net146));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[4]$_SDFFE_PP0P__147  (.L_HI(net147));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[5]$_SDFFE_PP0P__148  (.L_HI(net148));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[6]$_SDFFE_PP0P__149  (.L_HI(net149));
 sg13g2_tiehi \i2c_bert.myState_1.alu_1.acc[7]$_SDFFE_PP0P__150  (.L_HI(net150));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[0]$_SDFFCE_PP0P__151  (.L_HI(net151));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[1]$_SDFFCE_PP0P__152  (.L_HI(net152));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[2]$_SDFFCE_PP1P__153  (.L_HI(net153));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[3]$_SDFFCE_PP1P__154  (.L_HI(net154));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[4]$_SDFFCE_PP1P__155  (.L_HI(net155));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[5]$_SDFFCE_PP1P__156  (.L_HI(net156));
 sg13g2_tiehi \i2c_bert.myState_1.cmd7[6]$_SDFFCE_PP1P__157  (.L_HI(net157));
 sg13g2_tiehi \i2c_bert.myState_1.counter[0]$_SDFFE_PN1P__158  (.L_HI(net158));
 sg13g2_tiehi \i2c_bert.myState_1.counter[10]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \i2c_bert.myState_1.counter[11]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \i2c_bert.myState_1.counter[1]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \i2c_bert.myState_1.counter[2]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \i2c_bert.myState_1.counter[3]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \i2c_bert.myState_1.counter[4]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \i2c_bert.myState_1.counter[5]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \i2c_bert.myState_1.counter[6]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \i2c_bert.myState_1.counter[7]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \i2c_bert.myState_1.counter[8]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \i2c_bert.myState_1.counter[9]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \i2c_bert.myState_1.fsmPhase_stateReg[1]$_DFF_P__170  (.L_HI(net170));
 sg13g2_tiehi \i2c_bert.myState_1.fsmPhase_stateReg[2]$_DFF_P__171  (.L_HI(net171));
 sg13g2_tiehi \i2c_bert.myState_1.fsmPhase_stateReg[3]$_DFF_P__172  (.L_HI(net172));
 sg13g2_tiehi \i2c_bert.myState_1.fsmPhase_stateReg[4]$_DFF_P__173  (.L_HI(net173));
 sg13g2_tiehi \i2c_bert.myState_1.fsmPhase_stateReg[5]$_DFF_P__174  (.L_HI(net174));
 sg13g2_tiehi \i2c_bert.myState_1.led8[0]$_DFFE_PP__175  (.L_HI(net175));
 sg13g2_tiehi \i2c_bert.myState_1.led8[1]$_DFFE_PP__176  (.L_HI(net176));
 sg13g2_tiehi \i2c_bert.myState_1.led8[2]$_DFFE_PP__177  (.L_HI(net177));
 sg13g2_tiehi \i2c_bert.myState_1.led8[3]$_DFFE_PP__178  (.L_HI(net178));
 sg13g2_tiehi \i2c_bert.myState_1.led8[4]$_DFFE_PP__179  (.L_HI(net179));
 sg13g2_tiehi \i2c_bert.myState_1.led8[5]$_DFFE_PP__180  (.L_HI(net180));
 sg13g2_tiehi \i2c_bert.myState_1.led8[6]$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \i2c_bert.myState_1.led8[7]$_DFFE_PP__182  (.L_HI(net182));
 sg13g2_tiehi \i2c_bert.myState_1.len8[0]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \i2c_bert.myState_1.len8[1]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \i2c_bert.myState_1.len8[2]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \i2c_bert.myState_1.len8[3]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \i2c_bert.myState_1.len8[4]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \i2c_bert.myState_1.len8[5]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \i2c_bert.myState_1.len8[6]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \i2c_bert.myState_1.len8[7]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \i2c_bert.myState_1.readWriteBit$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \i2c_bert.powerOnSenseCaptured.genblk1.dlhrq_1_192  (.L_HI(net192));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[0]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[10]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[11]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[1]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[2]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[3]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[4]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[5]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[6]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[7]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[8]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \i2c_bert.timer_1.endstop[9]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[0]$_SDFF_PN0__205  (.L_HI(net205));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[10]$_SDFF_PN0__206  (.L_HI(net206));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[11]$_SDFF_PN0__207  (.L_HI(net207));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[1]$_SDFF_PN0__208  (.L_HI(net208));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[2]$_SDFF_PN0__209  (.L_HI(net209));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[3]$_SDFF_PN0__210  (.L_HI(net210));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[4]$_SDFF_PN0__211  (.L_HI(net211));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[5]$_SDFF_PN0__212  (.L_HI(net212));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[6]$_SDFF_PN0__213  (.L_HI(net213));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[7]$_SDFF_PN0__214  (.L_HI(net214));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[8]$_SDFF_PN0__215  (.L_HI(net215));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_count[9]$_SDFF_PN0__216  (.L_HI(net216));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[0]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[1]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[2]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[3]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[4]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[5]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[6]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_endstopTmpL[7]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \i2c_bert.timer_1.ticker_timerSampleTickState_regNext$_DFF_P__225  (.L_HI(net225));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N_226  (.L_HI(net226));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N_227  (.L_HI(net227));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N_228  (.L_HI(net228));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N_229  (.L_HI(net229));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N_230  (.L_HI(net230));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N_231  (.L_HI(net231));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N_232  (.L_HI(net232));
 sg13g2_tiehi \latched_config.latched_ena_ui_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N_233  (.L_HI(net233));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N_234  (.L_HI(net234));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N_235  (.L_HI(net235));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N_236  (.L_HI(net236));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N_237  (.L_HI(net237));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N_238  (.L_HI(net238));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N_239  (.L_HI(net239));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N_240  (.L_HI(net240));
 sg13g2_tiehi \latched_config.latched_ena_uio_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N_241  (.L_HI(net241));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N_242  (.L_HI(net242));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N_243  (.L_HI(net243));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N_244  (.L_HI(net244));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N_245  (.L_HI(net245));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N_246  (.L_HI(net246));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N_247  (.L_HI(net247));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N_248  (.L_HI(net248));
 sg13g2_tiehi \latched_config.latched_rst_n_ui_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N_249  (.L_HI(net249));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[0]$_DLATCH_N_._TECHMAP_DLATCH_N_250  (.L_HI(net250));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[1]$_DLATCH_N_._TECHMAP_DLATCH_N_251  (.L_HI(net251));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[2]$_DLATCH_N_._TECHMAP_DLATCH_N_252  (.L_HI(net252));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[3]$_DLATCH_N_._TECHMAP_DLATCH_N_253  (.L_HI(net253));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[4]$_DLATCH_N_._TECHMAP_DLATCH_N_254  (.L_HI(net254));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[5]$_DLATCH_N_._TECHMAP_DLATCH_N_255  (.L_HI(net255));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[6]$_DLATCH_N_._TECHMAP_DLATCH_N_256  (.L_HI(net256));
 sg13g2_tiehi \latched_config.latched_rst_n_uio_in[7]$_DLATCH_N_._TECHMAP_DLATCH_N_257  (.L_HI(net257));
 sg13g2_tiehi \rst_n_sync$_DFF_P__258  (.L_HI(net258));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_4 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_4 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_404 ();
 sg13g2_decap_8 FILLER_19_411 ();
 sg13g2_decap_8 FILLER_19_418 ();
 sg13g2_decap_4 FILLER_19_425 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_decap_4 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_8 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_20_412 ();
 sg13g2_decap_8 FILLER_20_419 ();
 sg13g2_decap_4 FILLER_20_426 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_decap_4 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_4 FILLER_21_424 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_4 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_4 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_4 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_4 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_260 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_4 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_243 ();
 sg13g2_decap_4 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_decap_4 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_decap_4 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_decap_4 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_decap_8 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_8 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_211 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_4 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_305 ();
 sg13g2_decap_4 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_4 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_4 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_8 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_4 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_8 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_32_412 ();
 sg13g2_decap_8 FILLER_32_419 ();
 sg13g2_decap_4 FILLER_32_426 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_decap_8 FILLER_33_283 ();
 sg13g2_decap_4 FILLER_33_290 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_4 FILLER_33_371 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_decap_4 FILLER_33_392 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_decap_4 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_decap_4 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_decap_4 FILLER_35_165 ();
 sg13g2_decap_4 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_decap_4 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_decap_4 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_8 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_decap_4 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_decap_4 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_decap_4 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_4 FILLER_37_211 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_4 FILLER_37_311 ();
 sg13g2_decap_4 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_4 FILLER_38_112 ();
 sg13g2_fill_1 FILLER_38_120 ();
 sg13g2_decap_8 FILLER_38_125 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_4 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_376 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_4 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_149 ();
 sg13g2_decap_8 FILLER_39_156 ();
 sg13g2_decap_8 FILLER_39_163 ();
 sg13g2_decap_8 FILLER_39_170 ();
 sg13g2_decap_4 FILLER_39_177 ();
 sg13g2_fill_1 FILLER_39_181 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_232 ();
 sg13g2_decap_4 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_fill_2 FILLER_39_259 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_fill_2 FILLER_39_266 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_290 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_decap_4 FILLER_39_307 ();
 sg13g2_fill_1 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_338 ();
 sg13g2_fill_2 FILLER_39_345 ();
 sg13g2_fill_1 FILLER_39_352 ();
 sg13g2_decap_4 FILLER_39_372 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_39_409 ();
 sg13g2_decap_8 FILLER_39_414 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_112 ();
 sg13g2_decap_4 FILLER_40_120 ();
 sg13g2_decap_8 FILLER_40_128 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_173 ();
 sg13g2_decap_4 FILLER_40_180 ();
 sg13g2_fill_1 FILLER_40_184 ();
 sg13g2_decap_8 FILLER_40_193 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_208 ();
 sg13g2_decap_8 FILLER_40_215 ();
 sg13g2_fill_2 FILLER_40_222 ();
 sg13g2_fill_1 FILLER_40_227 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_240 ();
 sg13g2_fill_1 FILLER_40_250 ();
 sg13g2_decap_4 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_decap_4 FILLER_40_270 ();
 sg13g2_fill_2 FILLER_40_274 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_4 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_298 ();
 sg13g2_fill_2 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_decap_8 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_344 ();
 sg13g2_decap_4 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_355 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_422 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_4 FILLER_41_105 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_137 ();
 sg13g2_decap_8 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_2 FILLER_41_172 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_4 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_decap_4 FILLER_41_299 ();
 sg13g2_fill_1 FILLER_41_316 ();
 sg13g2_decap_4 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_381 ();
 sg13g2_decap_4 FILLER_41_388 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_402 ();
 sg13g2_decap_8 FILLER_41_409 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_4 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_decap_8 FILLER_42_125 ();
 sg13g2_decap_8 FILLER_42_132 ();
 sg13g2_decap_4 FILLER_42_139 ();
 sg13g2_fill_2 FILLER_42_170 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_decap_4 FILLER_42_178 ();
 sg13g2_fill_2 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_210 ();
 sg13g2_fill_2 FILLER_42_218 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_fill_1 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_284 ();
 sg13g2_decap_4 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_decap_8 FILLER_42_302 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_decap_8 FILLER_42_316 ();
 sg13g2_decap_4 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_350 ();
 sg13g2_decap_4 FILLER_42_361 ();
 sg13g2_decap_8 FILLER_42_421 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_4 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_137 ();
 sg13g2_decap_4 FILLER_43_153 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_209 ();
 sg13g2_fill_1 FILLER_43_211 ();
 sg13g2_fill_1 FILLER_43_237 ();
 sg13g2_fill_1 FILLER_43_249 ();
 sg13g2_fill_2 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_274 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_decap_4 FILLER_43_368 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_fill_1 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_43_410 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_decap_4 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_fill_2 FILLER_44_126 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_decap_4 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_decap_8 FILLER_44_163 ();
 sg13g2_decap_8 FILLER_44_183 ();
 sg13g2_decap_8 FILLER_44_190 ();
 sg13g2_decap_8 FILLER_44_197 ();
 sg13g2_fill_1 FILLER_44_204 ();
 sg13g2_fill_2 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_211 ();
 sg13g2_fill_1 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_233 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_decap_4 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_decap_4 FILLER_44_313 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_decap_4 FILLER_44_323 ();
 sg13g2_decap_4 FILLER_44_332 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_363 ();
 sg13g2_decap_4 FILLER_44_370 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_fill_2 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_decap_8 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_44_414 ();
 sg13g2_decap_8 FILLER_44_421 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_4 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_130 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_fill_2 FILLER_45_160 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_fill_2 FILLER_45_182 ();
 sg13g2_fill_1 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_fill_2 FILLER_45_223 ();
 sg13g2_decap_4 FILLER_45_255 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_decap_4 FILLER_45_274 ();
 sg13g2_decap_4 FILLER_45_283 ();
 sg13g2_fill_2 FILLER_45_287 ();
 sg13g2_decap_4 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_1 FILLER_45_374 ();
 sg13g2_fill_1 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_416 ();
 sg13g2_decap_8 FILLER_45_423 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_1 FILLER_46_152 ();
 sg13g2_decap_8 FILLER_46_186 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_decap_4 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_204 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_4 FILLER_46_229 ();
 sg13g2_fill_2 FILLER_46_233 ();
 sg13g2_decap_4 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_253 ();
 sg13g2_fill_1 FILLER_46_260 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_276 ();
 sg13g2_decap_4 FILLER_46_287 ();
 sg13g2_fill_1 FILLER_46_291 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_fill_2 FILLER_46_323 ();
 sg13g2_fill_1 FILLER_46_340 ();
 sg13g2_fill_2 FILLER_46_345 ();
 sg13g2_decap_4 FILLER_46_360 ();
 sg13g2_fill_2 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_418 ();
 sg13g2_decap_4 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_4 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_fill_2 FILLER_47_175 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_decap_4 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_fill_2 FILLER_47_203 ();
 sg13g2_fill_1 FILLER_47_205 ();
 sg13g2_decap_4 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_fill_1 FILLER_47_262 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_287 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_fill_1 FILLER_47_299 ();
 sg13g2_decap_8 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_317 ();
 sg13g2_decap_4 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_47_409 ();
 sg13g2_decap_8 FILLER_47_416 ();
 sg13g2_decap_8 FILLER_47_423 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_4 FILLER_48_105 ();
 sg13g2_fill_2 FILLER_48_109 ();
 sg13g2_fill_1 FILLER_48_136 ();
 sg13g2_fill_1 FILLER_48_141 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_186 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_2 FILLER_48_229 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_fill_1 FILLER_48_247 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_fill_2 FILLER_48_339 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_4 FILLER_48_357 ();
 sg13g2_fill_1 FILLER_48_395 ();
 sg13g2_decap_4 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_48_411 ();
 sg13g2_decap_8 FILLER_48_418 ();
 sg13g2_decap_4 FILLER_48_425 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_fill_2 FILLER_49_123 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_181 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_decap_4 FILLER_49_222 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_4 FILLER_49_245 ();
 sg13g2_fill_2 FILLER_49_249 ();
 sg13g2_decap_4 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_265 ();
 sg13g2_decap_4 FILLER_49_309 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_decap_8 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_decap_8 FILLER_49_348 ();
 sg13g2_fill_2 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_4 FILLER_49_386 ();
 sg13g2_fill_1 FILLER_49_390 ();
 sg13g2_fill_1 FILLER_49_401 ();
 sg13g2_decap_8 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_4 FILLER_50_112 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_fill_1 FILLER_50_159 ();
 sg13g2_fill_1 FILLER_50_165 ();
 sg13g2_decap_8 FILLER_50_174 ();
 sg13g2_decap_8 FILLER_50_181 ();
 sg13g2_decap_4 FILLER_50_188 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_207 ();
 sg13g2_decap_8 FILLER_50_214 ();
 sg13g2_decap_8 FILLER_50_221 ();
 sg13g2_decap_8 FILLER_50_228 ();
 sg13g2_decap_8 FILLER_50_235 ();
 sg13g2_decap_4 FILLER_50_242 ();
 sg13g2_decap_4 FILLER_50_260 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_decap_4 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_fill_2 FILLER_50_334 ();
 sg13g2_decap_4 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_fill_1 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_fill_2 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_412 ();
 sg13g2_decap_8 FILLER_50_419 ();
 sg13g2_decap_4 FILLER_50_426 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_160 ();
 sg13g2_decap_8 FILLER_51_174 ();
 sg13g2_decap_4 FILLER_51_186 ();
 sg13g2_fill_2 FILLER_51_204 ();
 sg13g2_fill_1 FILLER_51_206 ();
 sg13g2_fill_1 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_220 ();
 sg13g2_fill_1 FILLER_51_231 ();
 sg13g2_decap_4 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_298 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_329 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_4 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_415 ();
 sg13g2_decap_8 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_fill_1 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_148 ();
 sg13g2_fill_1 FILLER_52_153 ();
 sg13g2_fill_2 FILLER_52_160 ();
 sg13g2_fill_1 FILLER_52_162 ();
 sg13g2_fill_2 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_186 ();
 sg13g2_decap_4 FILLER_52_192 ();
 sg13g2_decap_4 FILLER_52_219 ();
 sg13g2_fill_2 FILLER_52_258 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_decap_4 FILLER_52_296 ();
 sg13g2_fill_2 FILLER_52_300 ();
 sg13g2_decap_8 FILLER_52_307 ();
 sg13g2_decap_4 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_318 ();
 sg13g2_decap_4 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_338 ();
 sg13g2_decap_8 FILLER_52_345 ();
 sg13g2_decap_8 FILLER_52_352 ();
 sg13g2_decap_8 FILLER_52_359 ();
 sg13g2_decap_8 FILLER_52_366 ();
 sg13g2_fill_2 FILLER_52_391 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_418 ();
 sg13g2_decap_4 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_4 FILLER_53_112 ();
 sg13g2_fill_2 FILLER_53_116 ();
 sg13g2_decap_8 FILLER_53_123 ();
 sg13g2_decap_4 FILLER_53_130 ();
 sg13g2_decap_4 FILLER_53_139 ();
 sg13g2_decap_8 FILLER_53_178 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_2 FILLER_53_227 ();
 sg13g2_decap_8 FILLER_53_250 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_fill_2 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_312 ();
 sg13g2_fill_1 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_343 ();
 sg13g2_fill_1 FILLER_53_349 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_1 FILLER_53_366 ();
 sg13g2_fill_2 FILLER_53_397 ();
 sg13g2_fill_1 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_fill_2 FILLER_54_119 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_143 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_fill_2 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_decap_4 FILLER_54_164 ();
 sg13g2_fill_2 FILLER_54_168 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_180 ();
 sg13g2_fill_1 FILLER_54_187 ();
 sg13g2_fill_1 FILLER_54_198 ();
 sg13g2_fill_1 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_fill_1 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_fill_1 FILLER_54_232 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_1 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_295 ();
 sg13g2_fill_2 FILLER_54_302 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_fill_1 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_348 ();
 sg13g2_fill_1 FILLER_54_380 ();
 sg13g2_decap_4 FILLER_54_389 ();
 sg13g2_decap_4 FILLER_54_398 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_fill_2 FILLER_54_427 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_4 FILLER_55_119 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_133 ();
 sg13g2_fill_1 FILLER_55_135 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_decap_4 FILLER_55_153 ();
 sg13g2_fill_2 FILLER_55_157 ();
 sg13g2_decap_4 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_223 ();
 sg13g2_fill_1 FILLER_55_230 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_decap_4 FILLER_55_248 ();
 sg13g2_decap_4 FILLER_55_257 ();
 sg13g2_fill_2 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_272 ();
 sg13g2_fill_2 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_297 ();
 sg13g2_decap_4 FILLER_55_304 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_314 ();
 sg13g2_decap_4 FILLER_55_321 ();
 sg13g2_fill_2 FILLER_55_348 ();
 sg13g2_fill_1 FILLER_55_350 ();
 sg13g2_fill_1 FILLER_55_360 ();
 sg13g2_decap_4 FILLER_55_370 ();
 sg13g2_fill_2 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_fill_1 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_181 ();
 sg13g2_decap_8 FILLER_56_188 ();
 sg13g2_decap_8 FILLER_56_195 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_215 ();
 sg13g2_decap_4 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_249 ();
 sg13g2_fill_2 FILLER_56_258 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_fill_2 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_267 ();
 sg13g2_fill_2 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_275 ();
 sg13g2_fill_2 FILLER_56_281 ();
 sg13g2_decap_8 FILLER_56_299 ();
 sg13g2_decap_8 FILLER_56_306 ();
 sg13g2_decap_8 FILLER_56_313 ();
 sg13g2_decap_8 FILLER_56_320 ();
 sg13g2_fill_2 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_345 ();
 sg13g2_decap_4 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_decap_4 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_379 ();
 sg13g2_decap_8 FILLER_56_386 ();
 sg13g2_decap_8 FILLER_56_393 ();
 sg13g2_decap_4 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_176 ();
 sg13g2_fill_2 FILLER_57_183 ();
 sg13g2_decap_8 FILLER_57_211 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_fill_2 FILLER_57_225 ();
 sg13g2_fill_2 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_decap_4 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_277 ();
 sg13g2_decap_8 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_333 ();
 sg13g2_fill_2 FILLER_57_354 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_fill_1 FILLER_57_398 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_4 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_199 ();
 sg13g2_fill_2 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_decap_8 FILLER_58_269 ();
 sg13g2_decap_8 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_fill_2 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_decap_8 FILLER_58_351 ();
 sg13g2_fill_2 FILLER_58_358 ();
 sg13g2_fill_1 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_4 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_410 ();
 sg13g2_decap_8 FILLER_58_419 ();
 sg13g2_decap_4 FILLER_58_426 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_160 ();
 sg13g2_fill_1 FILLER_59_165 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_decap_4 FILLER_59_216 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_240 ();
 sg13g2_fill_1 FILLER_59_242 ();
 sg13g2_decap_8 FILLER_59_247 ();
 sg13g2_decap_8 FILLER_59_254 ();
 sg13g2_decap_4 FILLER_59_261 ();
 sg13g2_fill_1 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_decap_4 FILLER_59_277 ();
 sg13g2_decap_4 FILLER_59_285 ();
 sg13g2_decap_4 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_302 ();
 sg13g2_decap_4 FILLER_59_309 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_fill_1 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_388 ();
 sg13g2_decap_4 FILLER_59_395 ();
 sg13g2_fill_1 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_4 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_141 ();
 sg13g2_decap_4 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_157 ();
 sg13g2_decap_8 FILLER_60_164 ();
 sg13g2_decap_8 FILLER_60_171 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_204 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_decap_8 FILLER_60_218 ();
 sg13g2_decap_8 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_decap_8 FILLER_60_242 ();
 sg13g2_decap_4 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_309 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_decap_4 FILLER_60_320 ();
 sg13g2_decap_4 FILLER_60_328 ();
 sg13g2_fill_2 FILLER_60_332 ();
 sg13g2_decap_4 FILLER_60_347 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_4 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_fill_1 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_419 ();
 sg13g2_decap_4 FILLER_60_426 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_4 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_158 ();
 sg13g2_decap_8 FILLER_61_164 ();
 sg13g2_decap_8 FILLER_61_171 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_decap_8 FILLER_61_185 ();
 sg13g2_fill_2 FILLER_61_192 ();
 sg13g2_fill_2 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_205 ();
 sg13g2_decap_8 FILLER_61_209 ();
 sg13g2_decap_8 FILLER_61_216 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_230 ();
 sg13g2_decap_8 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_fill_2 FILLER_61_261 ();
 sg13g2_fill_2 FILLER_61_272 ();
 sg13g2_decap_4 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_324 ();
 sg13g2_decap_8 FILLER_61_331 ();
 sg13g2_decap_8 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_decap_4 FILLER_61_352 ();
 sg13g2_fill_2 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_362 ();
 sg13g2_fill_2 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_61_420 ();
 sg13g2_fill_2 FILLER_61_427 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_189 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_222 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_234 ();
 sg13g2_fill_2 FILLER_62_252 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_decap_8 FILLER_62_269 ();
 sg13g2_decap_4 FILLER_62_276 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_2 FILLER_62_297 ();
 sg13g2_fill_1 FILLER_62_299 ();
 sg13g2_decap_8 FILLER_62_326 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_decap_8 FILLER_62_347 ();
 sg13g2_decap_8 FILLER_62_354 ();
 sg13g2_decap_8 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_376 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_fill_1 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_167 ();
 sg13g2_fill_1 FILLER_63_172 ();
 sg13g2_fill_1 FILLER_63_183 ();
 sg13g2_fill_2 FILLER_63_189 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_fill_1 FILLER_63_213 ();
 sg13g2_fill_1 FILLER_63_219 ();
 sg13g2_fill_2 FILLER_63_229 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_decap_8 FILLER_63_251 ();
 sg13g2_decap_4 FILLER_63_258 ();
 sg13g2_decap_4 FILLER_63_298 ();
 sg13g2_decap_4 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_decap_8 FILLER_63_321 ();
 sg13g2_decap_8 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_335 ();
 sg13g2_fill_1 FILLER_63_337 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_4 FILLER_64_133 ();
 sg13g2_fill_1 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_181 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_2 FILLER_64_245 ();
 sg13g2_fill_2 FILLER_64_254 ();
 sg13g2_decap_8 FILLER_64_261 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_270 ();
 sg13g2_fill_2 FILLER_64_276 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_fill_2 FILLER_64_283 ();
 sg13g2_fill_1 FILLER_64_285 ();
 sg13g2_decap_8 FILLER_64_297 ();
 sg13g2_fill_2 FILLER_64_304 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_312 ();
 sg13g2_fill_1 FILLER_64_319 ();
 sg13g2_fill_2 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_147 ();
 sg13g2_decap_4 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_fill_2 FILLER_65_185 ();
 sg13g2_fill_1 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_193 ();
 sg13g2_fill_1 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_206 ();
 sg13g2_fill_2 FILLER_65_217 ();
 sg13g2_fill_1 FILLER_65_219 ();
 sg13g2_fill_1 FILLER_65_235 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_251 ();
 sg13g2_decap_4 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_fill_1 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_278 ();
 sg13g2_decap_8 FILLER_65_285 ();
 sg13g2_decap_8 FILLER_65_292 ();
 sg13g2_decap_8 FILLER_65_299 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_fill_2 FILLER_65_332 ();
 sg13g2_decap_8 FILLER_65_354 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_fill_1 FILLER_65_368 ();
 sg13g2_fill_1 FILLER_65_377 ();
 sg13g2_decap_4 FILLER_65_382 ();
 sg13g2_fill_1 FILLER_65_400 ();
 sg13g2_decap_8 FILLER_65_415 ();
 sg13g2_decap_8 FILLER_65_422 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_decap_8 FILLER_66_180 ();
 sg13g2_decap_4 FILLER_66_191 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_fill_1 FILLER_66_213 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_265 ();
 sg13g2_fill_2 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_284 ();
 sg13g2_decap_8 FILLER_66_291 ();
 sg13g2_decap_4 FILLER_66_298 ();
 sg13g2_fill_1 FILLER_66_314 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_343 ();
 sg13g2_fill_1 FILLER_66_345 ();
 sg13g2_decap_4 FILLER_66_350 ();
 sg13g2_decap_4 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_fill_1 FILLER_66_425 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_156 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_190 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_209 ();
 sg13g2_decap_8 FILLER_67_216 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_decap_4 FILLER_67_251 ();
 sg13g2_fill_2 FILLER_67_262 ();
 sg13g2_fill_2 FILLER_67_269 ();
 sg13g2_decap_8 FILLER_67_291 ();
 sg13g2_fill_2 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_300 ();
 sg13g2_decap_4 FILLER_67_311 ();
 sg13g2_decap_8 FILLER_67_335 ();
 sg13g2_decap_4 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_346 ();
 sg13g2_decap_8 FILLER_67_351 ();
 sg13g2_decap_8 FILLER_67_358 ();
 sg13g2_fill_1 FILLER_67_365 ();
 sg13g2_fill_1 FILLER_67_382 ();
 sg13g2_decap_8 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_67_414 ();
 sg13g2_decap_8 FILLER_67_421 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_156 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_212 ();
 sg13g2_fill_2 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_257 ();
 sg13g2_decap_4 FILLER_68_271 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_decap_4 FILLER_68_337 ();
 sg13g2_decap_4 FILLER_68_362 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_fill_1 FILLER_68_377 ();
 sg13g2_fill_2 FILLER_68_382 ();
 sg13g2_decap_4 FILLER_68_389 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_fill_2 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_156 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_decap_4 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_189 ();
 sg13g2_fill_2 FILLER_69_194 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_212 ();
 sg13g2_fill_2 FILLER_69_226 ();
 sg13g2_fill_2 FILLER_69_277 ();
 sg13g2_fill_1 FILLER_69_279 ();
 sg13g2_decap_4 FILLER_69_297 ();
 sg13g2_fill_2 FILLER_69_317 ();
 sg13g2_fill_2 FILLER_69_335 ();
 sg13g2_fill_1 FILLER_69_373 ();
 sg13g2_fill_2 FILLER_69_394 ();
 sg13g2_fill_1 FILLER_69_401 ();
 sg13g2_decap_4 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_decap_8 FILLER_69_415 ();
 sg13g2_decap_8 FILLER_69_422 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_fill_1 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_173 ();
 sg13g2_decap_8 FILLER_70_180 ();
 sg13g2_decap_8 FILLER_70_187 ();
 sg13g2_decap_8 FILLER_70_207 ();
 sg13g2_fill_2 FILLER_70_214 ();
 sg13g2_fill_1 FILLER_70_216 ();
 sg13g2_decap_4 FILLER_70_229 ();
 sg13g2_fill_2 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_262 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_decap_8 FILLER_70_274 ();
 sg13g2_decap_4 FILLER_70_281 ();
 sg13g2_decap_8 FILLER_70_289 ();
 sg13g2_decap_4 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_decap_4 FILLER_70_333 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_373 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_fill_2 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_409 ();
 sg13g2_fill_2 FILLER_70_416 ();
 sg13g2_decap_8 FILLER_70_423 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_decap_4 FILLER_71_180 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_decap_8 FILLER_71_220 ();
 sg13g2_fill_2 FILLER_71_227 ();
 sg13g2_decap_4 FILLER_71_234 ();
 sg13g2_fill_1 FILLER_71_238 ();
 sg13g2_fill_2 FILLER_71_244 ();
 sg13g2_fill_1 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_decap_8 FILLER_71_289 ();
 sg13g2_decap_8 FILLER_71_296 ();
 sg13g2_decap_8 FILLER_71_303 ();
 sg13g2_decap_8 FILLER_71_310 ();
 sg13g2_decap_8 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_338 ();
 sg13g2_decap_8 FILLER_71_345 ();
 sg13g2_decap_4 FILLER_71_352 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_381 ();
 sg13g2_fill_2 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_4 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_178 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_2 FILLER_72_190 ();
 sg13g2_decap_4 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_fill_1 FILLER_72_239 ();
 sg13g2_decap_4 FILLER_72_246 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_1 FILLER_72_261 ();
 sg13g2_fill_1 FILLER_72_281 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_299 ();
 sg13g2_decap_8 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_313 ();
 sg13g2_fill_2 FILLER_72_351 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_368 ();
 sg13g2_fill_1 FILLER_72_375 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_4 FILLER_73_168 ();
 sg13g2_fill_1 FILLER_73_172 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_2 FILLER_73_187 ();
 sg13g2_fill_1 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_2 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_251 ();
 sg13g2_fill_1 FILLER_73_258 ();
 sg13g2_decap_4 FILLER_73_264 ();
 sg13g2_decap_8 FILLER_73_297 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_fill_1 FILLER_73_345 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_368 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_fill_1 FILLER_73_379 ();
 sg13g2_fill_1 FILLER_73_398 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_4 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_2 FILLER_74_183 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_1 FILLER_74_197 ();
 sg13g2_fill_2 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_fill_1 FILLER_74_224 ();
 sg13g2_fill_1 FILLER_74_231 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_309 ();
 sg13g2_fill_2 FILLER_74_313 ();
 sg13g2_decap_4 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_fill_2 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_74_376 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_decap_4 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_404 ();
 sg13g2_fill_2 FILLER_74_410 ();
 sg13g2_fill_2 FILLER_74_416 ();
 sg13g2_fill_1 FILLER_74_418 ();
 sg13g2_decap_8 FILLER_74_423 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_fill_1 FILLER_75_168 ();
 sg13g2_decap_4 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_206 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_fill_2 FILLER_75_227 ();
 sg13g2_decap_4 FILLER_75_239 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_fill_2 FILLER_75_254 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_decap_4 FILLER_75_262 ();
 sg13g2_fill_1 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_300 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_fill_2 FILLER_75_314 ();
 sg13g2_fill_1 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_321 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_4 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_394 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_417 ();
 sg13g2_decap_4 FILLER_75_424 ();
 sg13g2_fill_2 FILLER_75_428 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_4 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_186 ();
 sg13g2_decap_8 FILLER_76_211 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_decap_4 FILLER_76_225 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_271 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_fill_1 FILLER_76_280 ();
 sg13g2_decap_4 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_353 ();
 sg13g2_fill_2 FILLER_76_360 ();
 sg13g2_fill_1 FILLER_76_362 ();
 sg13g2_decap_8 FILLER_76_367 ();
 sg13g2_fill_2 FILLER_76_374 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_1 FILLER_76_396 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_208 ();
 sg13g2_decap_8 FILLER_77_215 ();
 sg13g2_decap_8 FILLER_77_222 ();
 sg13g2_decap_8 FILLER_77_229 ();
 sg13g2_decap_8 FILLER_77_240 ();
 sg13g2_decap_8 FILLER_77_247 ();
 sg13g2_decap_4 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_decap_8 FILLER_77_299 ();
 sg13g2_decap_8 FILLER_77_306 ();
 sg13g2_fill_1 FILLER_77_313 ();
 sg13g2_decap_8 FILLER_77_318 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_334 ();
 sg13g2_fill_2 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_77_366 ();
 sg13g2_decap_4 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_2 FILLER_77_387 ();
 sg13g2_fill_1 FILLER_77_389 ();
 sg13g2_fill_2 FILLER_77_393 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_4 FILLER_78_137 ();
 sg13g2_fill_1 FILLER_78_141 ();
 sg13g2_decap_8 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_fill_2 FILLER_78_160 ();
 sg13g2_fill_1 FILLER_78_162 ();
 sg13g2_fill_1 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_181 ();
 sg13g2_fill_1 FILLER_78_188 ();
 sg13g2_decap_4 FILLER_78_193 ();
 sg13g2_fill_1 FILLER_78_202 ();
 sg13g2_decap_4 FILLER_78_237 ();
 sg13g2_fill_2 FILLER_78_267 ();
 sg13g2_fill_1 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_296 ();
 sg13g2_fill_1 FILLER_78_303 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_423 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_4 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_4 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_128 ();
 sg13g2_decap_8 FILLER_79_135 ();
 sg13g2_decap_8 FILLER_79_146 ();
 sg13g2_fill_1 FILLER_79_153 ();
 sg13g2_decap_4 FILLER_79_166 ();
 sg13g2_fill_2 FILLER_79_170 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_183 ();
 sg13g2_decap_8 FILLER_79_190 ();
 sg13g2_decap_4 FILLER_79_197 ();
 sg13g2_fill_1 FILLER_79_201 ();
 sg13g2_decap_4 FILLER_79_222 ();
 sg13g2_fill_1 FILLER_79_226 ();
 sg13g2_fill_1 FILLER_79_257 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_283 ();
 sg13g2_decap_4 FILLER_79_290 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_361 ();
 sg13g2_fill_1 FILLER_79_363 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_412 ();
 sg13g2_decap_8 FILLER_79_419 ();
 sg13g2_decap_4 FILLER_79_426 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_4 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_74 ();
 sg13g2_decap_8 FILLER_80_103 ();
 sg13g2_decap_4 FILLER_80_114 ();
 sg13g2_decap_8 FILLER_80_134 ();
 sg13g2_decap_4 FILLER_80_141 ();
 sg13g2_fill_2 FILLER_80_145 ();
 sg13g2_decap_4 FILLER_80_151 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_179 ();
 sg13g2_fill_2 FILLER_80_199 ();
 sg13g2_fill_1 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_224 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_241 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_258 ();
 sg13g2_decap_4 FILLER_80_269 ();
 sg13g2_fill_2 FILLER_80_281 ();
 sg13g2_decap_4 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_291 ();
 sg13g2_decap_4 FILLER_80_301 ();
 sg13g2_fill_2 FILLER_80_305 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_fill_2 FILLER_80_316 ();
 sg13g2_fill_1 FILLER_80_326 ();
 sg13g2_fill_2 FILLER_80_347 ();
 sg13g2_decap_4 FILLER_80_403 ();
 sg13g2_fill_1 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
endmodule
