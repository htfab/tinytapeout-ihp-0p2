module tt_um_vga_clock (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire clknet_0_clk;
 wire net63;
 wire \vga_clock.col_index[0] ;
 wire \vga_clock.col_index[1] ;
 wire \vga_clock.col_index_q[0] ;
 wire \vga_clock.col_index_q[1] ;
 wire \vga_clock.color[0] ;
 wire \vga_clock.color[1] ;
 wire \vga_clock.color[2] ;
 wire \vga_clock.color[3] ;
 wire \vga_clock.color[4] ;
 wire \vga_clock.color[5] ;
 wire \vga_clock.color_offset[0] ;
 wire \vga_clock.color_offset[1] ;
 wire \vga_clock.color_offset[2] ;
 wire \vga_clock.digit_0.char[0] ;
 wire \vga_clock.digit_0.char[1] ;
 wire \vga_clock.digit_0.char[2] ;
 wire \vga_clock.digit_0.char[3] ;
 wire \vga_clock.digit_0.digit_index[0] ;
 wire \vga_clock.digit_0.digit_index[1] ;
 wire \vga_clock.digit_0.digit_index[2] ;
 wire \vga_clock.digit_0.digit_index[3] ;
 wire \vga_clock.digit_0.digit_index[4] ;
 wire \vga_clock.digit_0.digit_index[5] ;
 wire \vga_clock.digit_0.number[0] ;
 wire \vga_clock.digit_0.number[1] ;
 wire \vga_clock.digit_0.x_block[0] ;
 wire \vga_clock.digit_0.x_block[1] ;
 wire \vga_clock.draw ;
 wire \vga_clock.font_0.dout[1] ;
 wire \vga_clock.font_0.dout[2] ;
 wire \vga_clock.font_0.dout[3] ;
 wire \vga_clock.hrs_d[0] ;
 wire \vga_clock.hrs_d[1] ;
 wire \vga_clock.hrs_u[0] ;
 wire \vga_clock.hrs_u[1] ;
 wire \vga_clock.hrs_u[2] ;
 wire \vga_clock.hrs_u[3] ;
 wire \vga_clock.min_d[0] ;
 wire \vga_clock.min_d[1] ;
 wire \vga_clock.min_d[2] ;
 wire \vga_clock.min_u[0] ;
 wire \vga_clock.min_u[1] ;
 wire \vga_clock.min_u[2] ;
 wire \vga_clock.min_u[3] ;
 wire \vga_clock.pulse_hrs.comp[0] ;
 wire \vga_clock.pulse_hrs.comp[1] ;
 wire \vga_clock.pulse_hrs.comp[2] ;
 wire \vga_clock.pulse_hrs.comp[3] ;
 wire \vga_clock.pulse_hrs.comp[4] ;
 wire \vga_clock.pulse_hrs.count[0] ;
 wire \vga_clock.pulse_hrs.count[1] ;
 wire \vga_clock.pulse_hrs.count[2] ;
 wire \vga_clock.pulse_hrs.count[3] ;
 wire \vga_clock.pulse_hrs.count[4] ;
 wire \vga_clock.pulse_min.comp[0] ;
 wire \vga_clock.pulse_min.comp[1] ;
 wire \vga_clock.pulse_min.comp[2] ;
 wire \vga_clock.pulse_min.comp[3] ;
 wire \vga_clock.pulse_min.comp[4] ;
 wire \vga_clock.pulse_min.count[0] ;
 wire \vga_clock.pulse_min.count[1] ;
 wire \vga_clock.pulse_min.count[2] ;
 wire \vga_clock.pulse_min.count[3] ;
 wire \vga_clock.pulse_min.count[4] ;
 wire \vga_clock.pulse_sec.comp[0] ;
 wire \vga_clock.pulse_sec.comp[1] ;
 wire \vga_clock.pulse_sec.comp[2] ;
 wire \vga_clock.pulse_sec.comp[3] ;
 wire \vga_clock.pulse_sec.comp[4] ;
 wire \vga_clock.pulse_sec.count[0] ;
 wire \vga_clock.pulse_sec.count[1] ;
 wire \vga_clock.pulse_sec.count[2] ;
 wire \vga_clock.pulse_sec.count[3] ;
 wire \vga_clock.pulse_sec.count[4] ;
 wire \vga_clock.sec_counter[0] ;
 wire \vga_clock.sec_counter[10] ;
 wire \vga_clock.sec_counter[11] ;
 wire \vga_clock.sec_counter[12] ;
 wire \vga_clock.sec_counter[13] ;
 wire \vga_clock.sec_counter[14] ;
 wire \vga_clock.sec_counter[15] ;
 wire \vga_clock.sec_counter[16] ;
 wire \vga_clock.sec_counter[17] ;
 wire \vga_clock.sec_counter[18] ;
 wire \vga_clock.sec_counter[19] ;
 wire \vga_clock.sec_counter[1] ;
 wire \vga_clock.sec_counter[20] ;
 wire \vga_clock.sec_counter[21] ;
 wire \vga_clock.sec_counter[22] ;
 wire \vga_clock.sec_counter[23] ;
 wire \vga_clock.sec_counter[24] ;
 wire \vga_clock.sec_counter[25] ;
 wire \vga_clock.sec_counter[2] ;
 wire \vga_clock.sec_counter[3] ;
 wire \vga_clock.sec_counter[4] ;
 wire \vga_clock.sec_counter[5] ;
 wire \vga_clock.sec_counter[6] ;
 wire \vga_clock.sec_counter[7] ;
 wire \vga_clock.sec_counter[8] ;
 wire \vga_clock.sec_counter[9] ;
 wire \vga_clock.sec_d[0] ;
 wire \vga_clock.sec_d[1] ;
 wire \vga_clock.sec_d[2] ;
 wire \vga_clock.sec_u[0] ;
 wire \vga_clock.sec_u[1] ;
 wire \vga_clock.sec_u[2] ;
 wire \vga_clock.sec_u[3] ;
 wire \vga_clock.vga_0.hc[0] ;
 wire \vga_clock.vga_0.hc[1] ;
 wire \vga_clock.vga_0.hc[2] ;
 wire \vga_clock.vga_0.hc[3] ;
 wire \vga_clock.vga_0.hc[4] ;
 wire \vga_clock.vga_0.hc[5] ;
 wire \vga_clock.vga_0.hc[6] ;
 wire \vga_clock.vga_0.hc[7] ;
 wire \vga_clock.vga_0.hc[8] ;
 wire \vga_clock.vga_0.hc[9] ;
 wire \vga_clock.vga_0.vc[0] ;
 wire \vga_clock.vga_0.vc[1] ;
 wire \vga_clock.vga_0.vc[2] ;
 wire \vga_clock.vga_0.vc[3] ;
 wire \vga_clock.vga_0.vc[4] ;
 wire \vga_clock.vga_0.vc[5] ;
 wire \vga_clock.vga_0.vc[6] ;
 wire \vga_clock.vga_0.vc[7] ;
 wire \vga_clock.vga_0.vc[8] ;
 wire \vga_clock.vga_0.vc[9] ;
 wire \vga_clock.vga_0.x_px[0] ;
 wire \vga_clock.vga_0.x_px[1] ;
 wire \vga_clock.vga_0.x_px[2] ;
 wire \vga_clock.vga_0.x_px[3] ;
 wire \vga_clock.vga_0.x_px[6] ;
 wire \vga_clock.vga_0.x_px[7] ;
 wire \vga_clock.vga_0.x_px[8] ;
 wire \vga_clock.vga_0.x_px[9] ;
 wire \vga_clock.vga_0.y_px[0] ;
 wire \vga_clock.vga_0.y_px[1] ;
 wire \vga_clock.vga_0.y_px[2] ;
 wire \vga_clock.vga_0.y_px[3] ;
 wire \vga_clock.vga_0.y_px[4] ;
 wire \vga_clock.vga_0.y_px[5] ;
 wire \vga_clock.vga_0.y_px[6] ;
 wire \vga_clock.vga_0.y_px[7] ;
 wire \vga_clock.vga_0.y_px[8] ;
 wire \vga_clock.vga_0.y_px[9] ;
 wire \vga_clock.x_block_q[5] ;
 wire \vga_clock.y_block[0] ;
 wire \vga_clock.y_block[1] ;
 wire \vga_clock.y_block[2] ;
 wire \vga_clock.y_block[3] ;
 wire \vga_clock.y_block[4] ;
 wire \vga_clock.y_block[5] ;
 wire \vga_clock.y_block_q[0] ;
 wire \vga_clock.y_block_q[1] ;
 wire \vga_clock.y_block_q[2] ;
 wire \vga_clock.y_block_q[3] ;
 wire \vga_clock.y_block_q[4] ;
 wire \vga_clock.y_block_q[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_2 _1070_ (.A(\vga_clock.vga_0.x_px[8] ),
    .X(_0365_));
 sg13g2_buf_1 _1071_ (.A(_0365_),
    .X(_0366_));
 sg13g2_xor2_1 _1072_ (.B(\vga_clock.color_offset[2] ),
    .A(net29),
    .X(_0367_));
 sg13g2_buf_1 _1073_ (.A(\vga_clock.vga_0.x_px[7] ),
    .X(_0368_));
 sg13g2_buf_1 _1074_ (.A(net43),
    .X(_0369_));
 sg13g2_buf_2 _1075_ (.A(\vga_clock.color_offset[1] ),
    .X(_0370_));
 sg13g2_nor2_1 _1076_ (.A(net28),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_buf_1 _1077_ (.A(\vga_clock.vga_0.x_px[6] ),
    .X(_0372_));
 sg13g2_buf_1 _1078_ (.A(net42),
    .X(_0373_));
 sg13g2_buf_2 _1079_ (.A(\vga_clock.color_offset[0] ),
    .X(_0374_));
 sg13g2_nand2_1 _1080_ (.Y(_0375_),
    .A(net27),
    .B(_0374_));
 sg13g2_nand2_2 _1081_ (.Y(_0376_),
    .A(net28),
    .B(_0370_));
 sg13g2_o21ai_1 _1082_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0371_),
    .A2(_0375_));
 sg13g2_nor2_1 _1083_ (.A(net27),
    .B(_0374_),
    .Y(_0378_));
 sg13g2_a21oi_1 _1084_ (.A1(_0376_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(_0371_));
 sg13g2_nand2_1 _1085_ (.Y(_0380_),
    .A(_0379_),
    .B(_0367_));
 sg13g2_o21ai_1 _1086_ (.B1(_0380_),
    .Y(_0000_),
    .A1(_0367_),
    .A2(_0377_));
 sg13g2_xnor2_1 _1087_ (.Y(_0381_),
    .A(net29),
    .B(\vga_clock.color_offset[2] ));
 sg13g2_xnor2_1 _1088_ (.Y(_0382_),
    .A(net27),
    .B(_0374_));
 sg13g2_a21oi_1 _1089_ (.A1(net28),
    .A2(_0370_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_nor3_1 _1090_ (.A(net27),
    .B(net28),
    .C(_0370_),
    .Y(_0384_));
 sg13g2_nor3_1 _1091_ (.A(_0381_),
    .B(_0383_),
    .C(_0384_),
    .Y(_0385_));
 sg13g2_xor2_1 _1092_ (.B(_0370_),
    .A(net28),
    .X(_0386_));
 sg13g2_nor2b_1 _1093_ (.A(_0375_),
    .B_N(_0386_),
    .Y(_0387_));
 sg13g2_nor2b_1 _1094_ (.A(_0376_),
    .B_N(_0375_),
    .Y(_0388_));
 sg13g2_nor3_1 _1095_ (.A(_0367_),
    .B(_0387_),
    .C(_0388_),
    .Y(_0389_));
 sg13g2_or2_1 _1096_ (.X(_0001_),
    .B(_0389_),
    .A(_0385_));
 sg13g2_inv_1 _1097_ (.Y(_0390_),
    .A(\vga_clock.digit_0.digit_index[4] ));
 sg13g2_buf_1 _1098_ (.A(\vga_clock.vga_0.y_px[4] ),
    .X(_0391_));
 sg13g2_or2_1 _1099_ (.X(_0392_),
    .B(\vga_clock.digit_0.digit_index[0] ),
    .A(net41));
 sg13g2_buf_8 _1100_ (.A(\vga_clock.vga_0.y_px[5] ),
    .X(_0393_));
 sg13g2_buf_2 _1101_ (.A(\vga_clock.digit_0.digit_index[1] ),
    .X(_0394_));
 sg13g2_and2_1 _1102_ (.A(_0393_),
    .B(_0394_),
    .X(_0395_));
 sg13g2_buf_8 _1103_ (.A(\vga_clock.vga_0.y_px[3] ),
    .X(_0396_));
 sg13g2_and2_1 _1104_ (.A(_0396_),
    .B(_0393_),
    .X(_0397_));
 sg13g2_a21o_1 _1105_ (.A2(\vga_clock.digit_0.digit_index[0] ),
    .A1(_0391_),
    .B1(_0394_),
    .X(_0398_));
 sg13g2_and4_1 _1106_ (.A(_0396_),
    .B(net41),
    .C(_0394_),
    .D(\vga_clock.digit_0.digit_index[0] ),
    .X(_0399_));
 sg13g2_a221oi_1 _1107_ (.B2(_0398_),
    .C1(_0399_),
    .B1(_0397_),
    .A1(_0392_),
    .Y(_0400_),
    .A2(_0395_));
 sg13g2_buf_1 _1108_ (.A(_0400_),
    .X(_0401_));
 sg13g2_nor3_2 _1109_ (.A(_0396_),
    .B(_0393_),
    .C(net41),
    .Y(_0402_));
 sg13g2_or2_1 _1110_ (.X(_0403_),
    .B(\vga_clock.digit_0.digit_index[0] ),
    .A(_0394_));
 sg13g2_buf_1 _1111_ (.A(_0403_),
    .X(_0404_));
 sg13g2_nand2_1 _1112_ (.Y(_0405_),
    .A(_0402_),
    .B(_0404_));
 sg13g2_buf_1 _1113_ (.A(\vga_clock.digit_0.digit_index[2] ),
    .X(_0406_));
 sg13g2_inv_1 _1114_ (.Y(_0407_),
    .A(net40));
 sg13g2_a21o_1 _1115_ (.A2(_0405_),
    .A1(net19),
    .B1(_0407_),
    .X(_0408_));
 sg13g2_buf_1 _1116_ (.A(\vga_clock.vga_0.y_px[6] ),
    .X(_0409_));
 sg13g2_or3_1 _1117_ (.A(_0396_),
    .B(_0393_),
    .C(net41),
    .X(_0410_));
 sg13g2_buf_8 _1118_ (.A(_0410_),
    .X(_0411_));
 sg13g2_xnor2_1 _1119_ (.Y(_0412_),
    .A(net39),
    .B(net21));
 sg13g2_a21o_1 _1120_ (.A2(_0405_),
    .A1(net19),
    .B1(_0412_),
    .X(_0413_));
 sg13g2_buf_1 _1121_ (.A(\vga_clock.digit_0.digit_index[3] ),
    .X(_0414_));
 sg13g2_buf_8 _1122_ (.A(\vga_clock.vga_0.y_px[7] ),
    .X(_0415_));
 sg13g2_a21o_1 _1123_ (.A2(net21),
    .A1(_0409_),
    .B1(net37),
    .X(_0416_));
 sg13g2_inv_1 _1124_ (.Y(\vga_clock.y_block[2] ),
    .A(_0412_));
 sg13g2_a22oi_1 _1125_ (.Y(_0417_),
    .B1(\vga_clock.y_block[2] ),
    .B2(net40),
    .A2(_0416_),
    .A1(net38));
 sg13g2_nand4_1 _1126_ (.B(_0408_),
    .C(_0413_),
    .A(_0390_),
    .Y(_0418_),
    .D(_0417_));
 sg13g2_nand2_1 _1127_ (.Y(_0419_),
    .A(_0409_),
    .B(net21));
 sg13g2_nor2_1 _1128_ (.A(net37),
    .B(net38),
    .Y(_0420_));
 sg13g2_buf_8 _1129_ (.A(_0016_),
    .X(_0421_));
 sg13g2_and4_1 _1130_ (.A(\vga_clock.vga_0.y_px[7] ),
    .B(net39),
    .C(_0421_),
    .D(net21),
    .X(_0422_));
 sg13g2_a21oi_1 _1131_ (.A1(_0419_),
    .A2(_0420_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_or2_1 _1132_ (.X(_0424_),
    .B(_0423_),
    .A(\vga_clock.digit_0.digit_index[4] ));
 sg13g2_nand2_1 _1133_ (.Y(_0425_),
    .A(net40),
    .B(net38));
 sg13g2_o21ai_1 _1134_ (.B1(_0422_),
    .Y(_0426_),
    .A1(net19),
    .A2(_0425_));
 sg13g2_nor2_2 _1135_ (.A(\vga_clock.vga_0.y_px[6] ),
    .B(net40),
    .Y(_0427_));
 sg13g2_or4_1 _1136_ (.A(_0396_),
    .B(_0393_),
    .C(net41),
    .D(net40),
    .X(_0428_));
 sg13g2_or4_1 _1137_ (.A(_0396_),
    .B(_0393_),
    .C(net41),
    .D(\vga_clock.vga_0.y_px[6] ),
    .X(_0429_));
 sg13g2_a22oi_1 _1138_ (.Y(_0430_),
    .B1(_0428_),
    .B2(_0429_),
    .A2(_0404_),
    .A1(_0402_));
 sg13g2_a21o_1 _1139_ (.A2(_0427_),
    .A1(net19),
    .B1(_0430_),
    .X(_0431_));
 sg13g2_a21oi_1 _1140_ (.A1(_0415_),
    .A2(net38),
    .Y(_0432_),
    .B1(_0421_));
 sg13g2_nand2_1 _1141_ (.Y(_0433_),
    .A(net39),
    .B(_0406_));
 sg13g2_a22oi_1 _1142_ (.Y(_0434_),
    .B1(\vga_clock.digit_0.digit_index[4] ),
    .B2(net21),
    .A2(net38),
    .A1(net37));
 sg13g2_or3_1 _1143_ (.A(net19),
    .B(_0433_),
    .C(_0434_),
    .X(_0435_));
 sg13g2_nor2_1 _1144_ (.A(_0390_),
    .B(_0420_),
    .Y(_0436_));
 sg13g2_nor2_1 _1145_ (.A(_0421_),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_a22oi_1 _1146_ (.Y(_0438_),
    .B1(_0435_),
    .B2(_0437_),
    .A2(_0432_),
    .A1(_0431_));
 sg13g2_nand4_1 _1147_ (.B(_0424_),
    .C(_0426_),
    .A(_0418_),
    .Y(_0439_),
    .D(_0438_));
 sg13g2_buf_2 _1148_ (.A(_0439_),
    .X(_0440_));
 sg13g2_and3_1 _1149_ (.X(_0441_),
    .A(net37),
    .B(net39),
    .C(_0411_));
 sg13g2_nor2b_1 _1150_ (.A(\vga_clock.vga_0.y_px[8] ),
    .B_N(\vga_clock.vga_0.y_px[9] ),
    .Y(_0442_));
 sg13g2_nor2b_1 _1151_ (.A(\vga_clock.vga_0.y_px[9] ),
    .B_N(_0421_),
    .Y(_0443_));
 sg13g2_inv_1 _1152_ (.Y(_0444_),
    .A(\vga_clock.vga_0.y_px[8] ));
 sg13g2_nand4_1 _1153_ (.B(net39),
    .C(_0444_),
    .A(net37),
    .Y(_0445_),
    .D(_0411_));
 sg13g2_nor2b_1 _1154_ (.A(_0421_),
    .B_N(\vga_clock.vga_0.y_px[9] ),
    .Y(_0446_));
 sg13g2_a221oi_1 _1155_ (.B2(_0445_),
    .C1(_0446_),
    .B1(_0443_),
    .A1(_0441_),
    .Y(_0447_),
    .A2(_0442_));
 sg13g2_xnor2_1 _1156_ (.Y(_0448_),
    .A(\vga_clock.digit_0.digit_index[5] ),
    .B(_0447_));
 sg13g2_xor2_1 _1157_ (.B(_0448_),
    .A(_0440_),
    .X(_0449_));
 sg13g2_o21ai_1 _1158_ (.B1(_0393_),
    .Y(_0450_),
    .A1(_0396_),
    .A2(net41));
 sg13g2_and2_1 _1159_ (.A(net21),
    .B(_0450_),
    .X(_0451_));
 sg13g2_xnor2_1 _1160_ (.Y(_0452_),
    .A(_0394_),
    .B(_0451_));
 sg13g2_buf_1 _1161_ (.A(_0452_),
    .X(_0453_));
 sg13g2_xor2_1 _1162_ (.B(net41),
    .A(_0396_),
    .X(_0454_));
 sg13g2_inv_1 _1163_ (.Y(\vga_clock.y_block[0] ),
    .A(_0454_));
 sg13g2_nor2_1 _1164_ (.A(net16),
    .B(net20),
    .Y(_0455_));
 sg13g2_xnor2_1 _1165_ (.Y(_0456_),
    .A(\vga_clock.vga_0.y_px[7] ),
    .B(net38));
 sg13g2_nand2_1 _1166_ (.Y(_0457_),
    .A(_0402_),
    .B(_0456_));
 sg13g2_a221oi_1 _1167_ (.B2(_0404_),
    .C1(_0457_),
    .B1(_0402_),
    .A1(net39),
    .Y(_0458_),
    .A2(net40));
 sg13g2_and4_1 _1168_ (.A(net19),
    .B(_0405_),
    .C(_0427_),
    .D(_0456_),
    .X(_0459_));
 sg13g2_xor2_1 _1169_ (.B(net38),
    .A(\vga_clock.vga_0.y_px[7] ),
    .X(_0460_));
 sg13g2_nor4_1 _1170_ (.A(_0402_),
    .B(net19),
    .C(_0433_),
    .D(_0460_),
    .Y(_0461_));
 sg13g2_nor4_1 _1171_ (.A(net39),
    .B(net40),
    .C(net21),
    .D(_0460_),
    .Y(_0462_));
 sg13g2_nor4_2 _1172_ (.A(_0458_),
    .B(_0459_),
    .C(_0461_),
    .Y(_0463_),
    .D(_0462_));
 sg13g2_nor2_1 _1173_ (.A(_0400_),
    .B(_0433_),
    .Y(_0464_));
 sg13g2_and3_1 _1174_ (.X(_0465_),
    .A(_0400_),
    .B(_0405_),
    .C(_0427_));
 sg13g2_a21o_1 _1175_ (.A2(_0427_),
    .A1(_0402_),
    .B1(_0456_),
    .X(_0466_));
 sg13g2_or4_1 _1176_ (.A(_0430_),
    .B(_0464_),
    .C(_0465_),
    .D(_0466_),
    .X(_0467_));
 sg13g2_buf_2 _1177_ (.A(_0467_),
    .X(_0468_));
 sg13g2_nand2_1 _1178_ (.Y(_0469_),
    .A(_0463_),
    .B(_0468_));
 sg13g2_nand2_1 _1179_ (.Y(_0470_),
    .A(_0401_),
    .B(_0405_));
 sg13g2_xnor2_1 _1180_ (.Y(_0471_),
    .A(net40),
    .B(_0412_));
 sg13g2_xor2_1 _1181_ (.B(_0471_),
    .A(_0470_),
    .X(_0472_));
 sg13g2_buf_1 _1182_ (.A(_0472_),
    .X(_0473_));
 sg13g2_nor2_1 _1183_ (.A(_0469_),
    .B(net13),
    .Y(_0474_));
 sg13g2_nand3_1 _1184_ (.B(_0455_),
    .C(_0474_),
    .A(_0449_),
    .Y(_0475_));
 sg13g2_buf_1 _1185_ (.A(_0469_),
    .X(_0476_));
 sg13g2_xor2_1 _1186_ (.B(_0451_),
    .A(_0394_),
    .X(_0477_));
 sg13g2_xnor2_1 _1187_ (.Y(_0478_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_nor2_1 _1188_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_nand2_1 _1189_ (.Y(_0480_),
    .A(_0476_),
    .B(_0479_));
 sg13g2_buf_1 _1190_ (.A(\vga_clock.digit_0.digit_index[0] ),
    .X(_0481_));
 sg13g2_a21o_1 _1191_ (.A2(_0480_),
    .A1(_0475_),
    .B1(_0481_),
    .X(_0482_));
 sg13g2_xnor2_1 _1192_ (.Y(_0483_),
    .A(_0440_),
    .B(_0448_));
 sg13g2_and2_1 _1193_ (.A(_0463_),
    .B(_0468_),
    .X(_0484_));
 sg13g2_buf_2 _1194_ (.A(_0484_),
    .X(_0485_));
 sg13g2_o21ai_1 _1195_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net16),
    .A2(_0483_));
 sg13g2_nor2_1 _1196_ (.A(net36),
    .B(\vga_clock.y_block[0] ),
    .Y(_0487_));
 sg13g2_buf_1 _1197_ (.A(_0477_),
    .X(_0488_));
 sg13g2_nand2_1 _1198_ (.Y(_0489_),
    .A(net36),
    .B(net20));
 sg13g2_a21oi_1 _1199_ (.A1(_0476_),
    .A2(net15),
    .Y(_0490_),
    .B1(_0489_));
 sg13g2_nor3_1 _1200_ (.A(_0487_),
    .B(_0478_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_nor4_1 _1201_ (.A(net12),
    .B(net15),
    .C(_0483_),
    .D(net13),
    .Y(_0492_));
 sg13g2_and2_1 _1202_ (.A(net36),
    .B(net20),
    .X(_0493_));
 sg13g2_buf_1 _1203_ (.A(_0493_),
    .X(_0494_));
 sg13g2_inv_1 _1204_ (.Y(_0495_),
    .A(net38));
 sg13g2_nand2_1 _1205_ (.Y(_0496_),
    .A(net37),
    .B(_0414_));
 sg13g2_nor3_1 _1206_ (.A(net19),
    .B(_0433_),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_a21o_1 _1207_ (.A2(_0431_),
    .A1(_0495_),
    .B1(_0497_),
    .X(_0498_));
 sg13g2_o21ai_1 _1208_ (.B1(_0401_),
    .Y(_0499_),
    .A1(_0495_),
    .A2(_0427_));
 sg13g2_o21ai_1 _1209_ (.B1(_0414_),
    .Y(_0500_),
    .A1(net21),
    .A2(_0404_));
 sg13g2_nand2_1 _1210_ (.Y(_0501_),
    .A(_0433_),
    .B(_0500_));
 sg13g2_a21oi_1 _1211_ (.A1(_0499_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(_0415_));
 sg13g2_xnor2_1 _1212_ (.Y(_0503_),
    .A(_0421_),
    .B(\vga_clock.digit_0.digit_index[4] ));
 sg13g2_o21ai_1 _1213_ (.B1(_0503_),
    .Y(_0504_),
    .A1(_0498_),
    .A2(_0502_));
 sg13g2_or3_1 _1214_ (.A(_0498_),
    .B(_0502_),
    .C(_0503_),
    .X(_0505_));
 sg13g2_and2_1 _1215_ (.A(_0504_),
    .B(_0505_),
    .X(_0506_));
 sg13g2_buf_1 _1216_ (.A(_0506_),
    .X(_0507_));
 sg13g2_a221oi_1 _1217_ (.B2(_0494_),
    .C1(_0507_),
    .B1(_0492_),
    .A1(_0486_),
    .Y(_0508_),
    .A2(_0491_));
 sg13g2_nand2_1 _1218_ (.Y(_0509_),
    .A(net12),
    .B(_0478_));
 sg13g2_nor2_1 _1219_ (.A(net15),
    .B(net13),
    .Y(_0510_));
 sg13g2_o21ai_1 _1220_ (.B1(_0449_),
    .Y(_0511_),
    .A1(net12),
    .A2(_0510_));
 sg13g2_xnor2_1 _1221_ (.Y(_0512_),
    .A(_0488_),
    .B(_0494_));
 sg13g2_nand2_1 _1222_ (.Y(_0513_),
    .A(net16),
    .B(_0487_));
 sg13g2_o21ai_1 _1223_ (.B1(_0507_),
    .Y(_0514_),
    .A1(net12),
    .A2(_0513_));
 sg13g2_a221oi_1 _1224_ (.B2(_0512_),
    .C1(_0514_),
    .B1(_0511_),
    .A1(_0483_),
    .Y(_0515_),
    .A2(_0509_));
 sg13g2_a21o_1 _1225_ (.A2(_0508_),
    .A1(_0482_),
    .B1(_0515_),
    .X(_0005_));
 sg13g2_nand2_1 _1226_ (.Y(_0516_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_nand2_1 _1227_ (.Y(_0517_),
    .A(net12),
    .B(net16));
 sg13g2_a221oi_1 _1228_ (.B2(_0487_),
    .C1(_0490_),
    .B1(_0517_),
    .A1(_0488_),
    .Y(_0518_),
    .A2(_0474_));
 sg13g2_nand3_1 _1229_ (.B(_0468_),
    .C(net15),
    .A(_0463_),
    .Y(_0519_));
 sg13g2_xnor2_1 _1230_ (.Y(_0520_),
    .A(net36),
    .B(net20));
 sg13g2_a21oi_1 _1231_ (.A1(net13),
    .A2(_0519_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_nor2_1 _1232_ (.A(_0516_),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_a21o_1 _1233_ (.A2(_0518_),
    .A1(_0516_),
    .B1(_0522_),
    .X(_0523_));
 sg13g2_nor2_1 _1234_ (.A(net12),
    .B(net16),
    .Y(_0524_));
 sg13g2_nand2_1 _1235_ (.Y(_0525_),
    .A(net15),
    .B(_0494_));
 sg13g2_a21o_1 _1236_ (.A2(_0525_),
    .A1(_0513_),
    .B1(_0485_),
    .X(_0526_));
 sg13g2_o21ai_1 _1237_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0507_),
    .A2(_0524_));
 sg13g2_a21oi_1 _1238_ (.A1(net13),
    .A2(_0527_),
    .Y(_0528_),
    .B1(_0483_));
 sg13g2_nand3_1 _1239_ (.B(_0468_),
    .C(net13),
    .A(_0463_),
    .Y(_0529_));
 sg13g2_nor2_1 _1240_ (.A(_0454_),
    .B(_0478_),
    .Y(_0530_));
 sg13g2_nand3_1 _1241_ (.B(_0468_),
    .C(net16),
    .A(_0463_),
    .Y(_0531_));
 sg13g2_a22oi_1 _1242_ (.Y(_0532_),
    .B1(_0530_),
    .B2(_0531_),
    .A2(_0529_),
    .A1(_0454_));
 sg13g2_nor2_1 _1243_ (.A(_0453_),
    .B(_0473_),
    .Y(_0533_));
 sg13g2_nor3_1 _1244_ (.A(_0485_),
    .B(_0479_),
    .C(_0533_),
    .Y(_0534_));
 sg13g2_a22oi_1 _1245_ (.Y(_0535_),
    .B1(_0534_),
    .B2(_0454_),
    .A2(_0532_),
    .A1(_0516_));
 sg13g2_nor2_1 _1246_ (.A(net20),
    .B(_0478_),
    .Y(_0536_));
 sg13g2_a22oi_1 _1247_ (.Y(_0537_),
    .B1(_0519_),
    .B2(_0536_),
    .A2(_0529_),
    .A1(net20));
 sg13g2_a221oi_1 _1248_ (.B2(_0516_),
    .C1(net36),
    .B1(_0537_),
    .A1(net20),
    .Y(_0538_),
    .A2(_0534_));
 sg13g2_a21o_1 _1249_ (.A2(_0535_),
    .A1(net36),
    .B1(_0538_),
    .X(_0539_));
 sg13g2_a22oi_1 _1250_ (.Y(_0006_),
    .B1(_0539_),
    .B2(_0483_),
    .A2(_0528_),
    .A1(_0523_));
 sg13g2_nor2_1 _1251_ (.A(net16),
    .B(_0448_),
    .Y(_0540_));
 sg13g2_nand2_1 _1252_ (.Y(_0541_),
    .A(_0440_),
    .B(_0540_));
 sg13g2_or3_1 _1253_ (.A(net15),
    .B(_0440_),
    .C(_0448_),
    .X(_0542_));
 sg13g2_nand2_1 _1254_ (.Y(_0543_),
    .A(net15),
    .B(_0448_));
 sg13g2_nand2_1 _1255_ (.Y(_0544_),
    .A(net16),
    .B(_0448_));
 sg13g2_mux2_1 _1256_ (.A0(_0543_),
    .A1(_0544_),
    .S(_0440_),
    .X(_0545_));
 sg13g2_o21ai_1 _1257_ (.B1(net36),
    .Y(_0546_),
    .A1(net15),
    .A2(net20));
 sg13g2_nand4_1 _1258_ (.B(_0542_),
    .C(_0545_),
    .A(_0541_),
    .Y(_0547_),
    .D(_0546_));
 sg13g2_nand2_1 _1259_ (.Y(_0548_),
    .A(_0452_),
    .B(_0494_));
 sg13g2_mux2_1 _1260_ (.A0(_0548_),
    .A1(_0525_),
    .S(_0449_),
    .X(_0549_));
 sg13g2_a221oi_1 _1261_ (.B2(_0549_),
    .C1(_0478_),
    .B1(_0547_),
    .A1(_0463_),
    .Y(_0550_),
    .A2(_0468_));
 sg13g2_nor2_1 _1262_ (.A(_0477_),
    .B(_0520_),
    .Y(_0551_));
 sg13g2_mux2_1 _1263_ (.A0(_0520_),
    .A1(_0551_),
    .S(net13),
    .X(_0552_));
 sg13g2_nand2_1 _1264_ (.Y(_0553_),
    .A(_0477_),
    .B(_0454_));
 sg13g2_o21ai_1 _1265_ (.B1(_0548_),
    .Y(_0554_),
    .A1(_0481_),
    .A2(_0553_));
 sg13g2_mux2_1 _1266_ (.A0(_0552_),
    .A1(_0554_),
    .S(_0485_),
    .X(_0555_));
 sg13g2_a21oi_1 _1267_ (.A1(_0504_),
    .A2(_0505_),
    .Y(_0556_),
    .B1(net36));
 sg13g2_a221oi_1 _1268_ (.B2(_0474_),
    .C1(_0483_),
    .B1(_0556_),
    .A1(_0507_),
    .Y(_0557_),
    .A2(_0555_));
 sg13g2_nor2_1 _1269_ (.A(_0478_),
    .B(_0553_),
    .Y(_0558_));
 sg13g2_a221oi_1 _1270_ (.B2(net12),
    .C1(_0507_),
    .B1(_0558_),
    .A1(_0449_),
    .Y(_0559_),
    .A2(_0455_));
 sg13g2_nor3_1 _1271_ (.A(net12),
    .B(_0487_),
    .C(net13),
    .Y(_0560_));
 sg13g2_nand3_1 _1272_ (.B(_0449_),
    .C(_0560_),
    .A(_0453_),
    .Y(_0561_));
 sg13g2_o21ai_1 _1273_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0557_),
    .A2(_0559_));
 sg13g2_nand2_1 _1274_ (.Y(_0563_),
    .A(_0507_),
    .B(_0557_));
 sg13g2_o21ai_1 _1275_ (.B1(_0563_),
    .Y(_0007_),
    .A1(_0550_),
    .A2(_0562_));
 sg13g2_buf_1 _1276_ (.A(\vga_clock.vga_0.x_px[9] ),
    .X(_0564_));
 sg13g2_buf_1 _1277_ (.A(_0564_),
    .X(_0565_));
 sg13g2_nor3_2 _1278_ (.A(\vga_clock.vga_0.x_px[6] ),
    .B(\vga_clock.vga_0.x_px[7] ),
    .C(_0365_),
    .Y(_0566_));
 sg13g2_xnor2_1 _1279_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_inv_1 _1280_ (.Y(\vga_clock.digit_0.char[3] ),
    .A(_0567_));
 sg13g2_xnor2_1 _1281_ (.Y(\vga_clock.digit_0.char[1] ),
    .A(net42),
    .B(_0369_));
 sg13g2_inv_1 _1282_ (.Y(_0568_),
    .A(_0368_));
 sg13g2_inv_1 _1283_ (.Y(_0569_),
    .A(_0365_));
 sg13g2_nor2b_1 _1284_ (.A(_0564_),
    .B_N(\vga_clock.vga_0.x_px[6] ),
    .Y(_0570_));
 sg13g2_nand3_1 _1285_ (.B(_0569_),
    .C(_0570_),
    .A(_0568_),
    .Y(_0571_));
 sg13g2_buf_1 _1286_ (.A(_0571_),
    .X(_0572_));
 sg13g2_buf_2 _1287_ (.A(\vga_clock.min_u[0] ),
    .X(_0573_));
 sg13g2_nand2_1 _1288_ (.Y(_0574_),
    .A(net42),
    .B(_0573_));
 sg13g2_o21ai_1 _1289_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net42),
    .A2(net29));
 sg13g2_inv_1 _1290_ (.Y(_0576_),
    .A(_0573_));
 sg13g2_buf_1 _1291_ (.A(\vga_clock.sec_d[0] ),
    .X(_0577_));
 sg13g2_nand3_1 _1292_ (.B(net29),
    .C(_0577_),
    .A(net43),
    .Y(_0578_));
 sg13g2_o21ai_1 _1293_ (.B1(_0578_),
    .Y(_0579_),
    .A1(net29),
    .A2(_0576_));
 sg13g2_a221oi_1 _1294_ (.B2(net27),
    .C1(net26),
    .B1(_0579_),
    .A1(_0568_),
    .Y(_0580_),
    .A2(_0575_));
 sg13g2_nor2_2 _1295_ (.A(_0372_),
    .B(net43),
    .Y(_0581_));
 sg13g2_nor2b_1 _1296_ (.A(\vga_clock.sec_u[0] ),
    .B_N(_0564_),
    .Y(_0582_));
 sg13g2_a21oi_1 _1297_ (.A1(_0581_),
    .A2(_0582_),
    .Y(_0583_),
    .B1(_0570_));
 sg13g2_nor2_1 _1298_ (.A(_0366_),
    .B(_0583_),
    .Y(_0584_));
 sg13g2_nand2_1 _1299_ (.Y(_0585_),
    .A(_0365_),
    .B(\vga_clock.min_d[0] ));
 sg13g2_buf_2 _1300_ (.A(\vga_clock.hrs_u[0] ),
    .X(_0586_));
 sg13g2_nand3b_1 _1301_ (.B(_0586_),
    .C(net43),
    .Y(_0587_),
    .A_N(_0365_));
 sg13g2_o21ai_1 _1302_ (.B1(_0587_),
    .Y(_0588_),
    .A1(net43),
    .A2(_0585_));
 sg13g2_o21ai_1 _1303_ (.B1(net42),
    .Y(_0589_),
    .A1(_0368_),
    .A2(_0366_));
 sg13g2_o21ai_1 _1304_ (.B1(_0589_),
    .Y(_0590_),
    .A1(_0372_),
    .A2(_0588_));
 sg13g2_or2_1 _1305_ (.X(_0591_),
    .B(_0590_),
    .A(net26));
 sg13g2_o21ai_1 _1306_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0580_),
    .A2(_0584_));
 sg13g2_o21ai_1 _1307_ (.B1(_0592_),
    .Y(_0593_),
    .A1(\vga_clock.hrs_d[0] ),
    .A2(_0572_));
 sg13g2_inv_1 _1308_ (.Y(\vga_clock.digit_0.number[0] ),
    .A(_0593_));
 sg13g2_o21ai_1 _1309_ (.B1(net27),
    .Y(_0594_),
    .A1(net28),
    .A2(_0021_));
 sg13g2_nand2b_1 _1310_ (.Y(_0595_),
    .B(_0594_),
    .A_N(_0581_));
 sg13g2_nor2_1 _1311_ (.A(_0569_),
    .B(net26),
    .Y(_0596_));
 sg13g2_xnor2_1 _1312_ (.Y(\vga_clock.digit_0.char[2] ),
    .A(_0569_),
    .B(_0581_));
 sg13g2_nor3_1 _1313_ (.A(_0565_),
    .B(\vga_clock.digit_0.char[1] ),
    .C(\vga_clock.digit_0.char[2] ),
    .Y(_0597_));
 sg13g2_and3_1 _1314_ (.X(_0598_),
    .A(net26),
    .B(_0022_),
    .C(_0566_));
 sg13g2_a221oi_1 _1315_ (.B2(_0020_),
    .C1(_0598_),
    .B1(_0597_),
    .A1(_0595_),
    .Y(_0599_),
    .A2(_0596_));
 sg13g2_a21oi_1 _1316_ (.A1(_0369_),
    .A2(_0019_),
    .Y(_0600_),
    .B1(_0373_));
 sg13g2_nor2b_1 _1317_ (.A(net43),
    .B_N(\vga_clock.min_u[2] ),
    .Y(_0601_));
 sg13g2_o21ai_1 _1318_ (.B1(_0601_),
    .Y(_0602_),
    .A1(net42),
    .A2(net29));
 sg13g2_nand4_1 _1319_ (.B(net43),
    .C(_0365_),
    .A(net42),
    .Y(_0603_),
    .D(\vga_clock.sec_d[2] ));
 sg13g2_a21o_1 _1320_ (.A2(_0603_),
    .A1(_0602_),
    .B1(net26),
    .X(_0604_));
 sg13g2_o21ai_1 _1321_ (.B1(net26),
    .Y(_0605_),
    .A1(net27),
    .A2(\vga_clock.sec_u[2] ));
 sg13g2_nand3_1 _1322_ (.B(_0604_),
    .C(_0605_),
    .A(_0568_),
    .Y(_0606_));
 sg13g2_o21ai_1 _1323_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net26),
    .A2(_0600_));
 sg13g2_nand2_1 _1324_ (.Y(_0608_),
    .A(\vga_clock.sec_u[2] ),
    .B(_0581_));
 sg13g2_a21oi_1 _1325_ (.A1(net26),
    .A2(_0608_),
    .Y(_0609_),
    .B1(net29));
 sg13g2_nand2b_1 _1326_ (.Y(_0610_),
    .B(_0581_),
    .A_N(_0564_));
 sg13g2_nor2_1 _1327_ (.A(\vga_clock.min_d[2] ),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_a21oi_1 _1328_ (.A1(_0604_),
    .A2(_0610_),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_nor2_1 _1329_ (.A(_0609_),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_a21oi_1 _1330_ (.A1(_0569_),
    .A2(_0607_),
    .Y(_0614_),
    .B1(_0613_));
 sg13g2_nand2b_1 _1331_ (.Y(_0615_),
    .B(_0614_),
    .A_N(_0599_));
 sg13g2_xnor2_1 _1332_ (.Y(_0002_),
    .A(\vga_clock.digit_0.number[0] ),
    .B(_0615_));
 sg13g2_inv_1 _1333_ (.Y(_0616_),
    .A(\vga_clock.hrs_d[1] ));
 sg13g2_nand3b_1 _1334_ (.B(_0365_),
    .C(net43),
    .Y(_0617_),
    .A_N(\vga_clock.sec_d[1] ));
 sg13g2_o21ai_1 _1335_ (.B1(_0617_),
    .Y(_0618_),
    .A1(net28),
    .A2(\vga_clock.min_u[1] ));
 sg13g2_nor3_1 _1336_ (.A(net42),
    .B(net28),
    .C(\vga_clock.min_d[1] ),
    .Y(_0619_));
 sg13g2_a21o_1 _1337_ (.A2(_0618_),
    .A1(net27),
    .B1(_0619_),
    .X(_0620_));
 sg13g2_nand3b_1 _1338_ (.B(_0581_),
    .C(_0564_),
    .Y(_0621_),
    .A_N(\vga_clock.sec_u[1] ));
 sg13g2_o21ai_1 _1339_ (.B1(_0572_),
    .Y(_0622_),
    .A1(net29),
    .A2(_0621_));
 sg13g2_a21oi_1 _1340_ (.A1(_0596_),
    .A2(_0620_),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_inv_1 _1341_ (.Y(_0624_),
    .A(\vga_clock.hrs_u[1] ));
 sg13g2_nand2_1 _1342_ (.Y(_0625_),
    .A(_0624_),
    .B(_0597_));
 sg13g2_nand2_1 _1343_ (.Y(_0626_),
    .A(_0623_),
    .B(_0625_));
 sg13g2_o21ai_1 _1344_ (.B1(_0626_),
    .Y(\vga_clock.digit_0.number[1] ),
    .A1(_0616_),
    .A2(_0572_));
 sg13g2_nand2_1 _1345_ (.Y(_0627_),
    .A(_0018_),
    .B(_0597_));
 sg13g2_nand2_1 _1346_ (.Y(_0628_),
    .A(_0623_),
    .B(_0627_));
 sg13g2_nand2b_1 _1347_ (.Y(_0629_),
    .B(_0614_),
    .A_N(_0593_));
 sg13g2_xnor2_1 _1348_ (.Y(_0630_),
    .A(\vga_clock.digit_0.number[1] ),
    .B(_0629_));
 sg13g2_nand2_1 _1349_ (.Y(_0631_),
    .A(_0572_),
    .B(_0599_));
 sg13g2_mux2_1 _1350_ (.A0(_0628_),
    .A1(_0630_),
    .S(_0631_),
    .X(_0003_));
 sg13g2_o21ai_1 _1351_ (.B1(_0628_),
    .Y(_0632_),
    .A1(_0017_),
    .A2(_0572_));
 sg13g2_nand2b_1 _1352_ (.Y(_0633_),
    .B(_0632_),
    .A_N(_0593_));
 sg13g2_nand2_1 _1353_ (.Y(_0634_),
    .A(_0614_),
    .B(_0633_));
 sg13g2_nand3_1 _1354_ (.B(_0623_),
    .C(_0625_),
    .A(_0599_),
    .Y(_0635_));
 sg13g2_o21ai_1 _1355_ (.B1(_0635_),
    .Y(_0004_),
    .A1(_0599_),
    .A2(_0634_));
 sg13g2_nand2b_1 _1356_ (.Y(_0035_),
    .B(_0567_),
    .A_N(\vga_clock.digit_0.x_block[0] ));
 sg13g2_nand2b_1 _1357_ (.Y(_0036_),
    .B(_0567_),
    .A_N(\vga_clock.digit_0.x_block[1] ));
 sg13g2_nand2b_1 _1358_ (.Y(_0636_),
    .B(_0381_),
    .A_N(_0376_));
 sg13g2_nand2_1 _1359_ (.Y(_0637_),
    .A(_0371_),
    .B(_0367_));
 sg13g2_a21oi_1 _1360_ (.A1(_0636_),
    .A2(_0637_),
    .Y(_0037_),
    .B1(_0382_));
 sg13g2_and2_1 _1361_ (.A(_0376_),
    .B(_0381_),
    .X(_0638_));
 sg13g2_nor2_1 _1362_ (.A(_0376_),
    .B(_0381_),
    .Y(_0639_));
 sg13g2_nor3_1 _1363_ (.A(_0373_),
    .B(_0374_),
    .C(_0386_),
    .Y(_0640_));
 sg13g2_nor4_1 _1364_ (.A(_0387_),
    .B(_0638_),
    .C(_0639_),
    .D(_0640_),
    .Y(_0038_));
 sg13g2_nand2_1 _1365_ (.Y(_0641_),
    .A(_0381_),
    .B(_0386_));
 sg13g2_nor2_1 _1366_ (.A(_0382_),
    .B(_0641_),
    .Y(_0039_));
 sg13g2_o21ai_1 _1367_ (.B1(_0631_),
    .Y(_0041_),
    .A1(_0615_),
    .A2(_0633_));
 sg13g2_inv_1 _1368_ (.Y(_0642_),
    .A(\vga_clock.hrs_u[3] ));
 sg13g2_nor4_2 _1369_ (.A(_0624_),
    .B(_0586_),
    .C(\vga_clock.hrs_u[2] ),
    .Y(_0643_),
    .D(_0642_));
 sg13g2_nand2_1 _1370_ (.Y(_0644_),
    .A(_0030_),
    .B(_0643_));
 sg13g2_inv_1 _1371_ (.Y(_0645_),
    .A(_0643_));
 sg13g2_nand2_1 _1372_ (.Y(_0646_),
    .A(\vga_clock.hrs_d[0] ),
    .B(_0645_));
 sg13g2_buf_1 _1373_ (.A(rst_n),
    .X(_0647_));
 sg13g2_nor4_1 _1374_ (.A(\vga_clock.hrs_u[1] ),
    .B(_0586_),
    .C(_0616_),
    .D(\vga_clock.hrs_d[0] ),
    .Y(_0648_));
 sg13g2_nand3_1 _1375_ (.B(_0642_),
    .C(_0648_),
    .A(\vga_clock.hrs_u[2] ),
    .Y(_0649_));
 sg13g2_nand2_1 _1376_ (.Y(_0650_),
    .A(_0647_),
    .B(_0649_));
 sg13g2_a21oi_1 _1377_ (.A1(_0644_),
    .A2(_0646_),
    .Y(_0043_),
    .B1(_0650_));
 sg13g2_nand2_1 _1378_ (.Y(_0651_),
    .A(\vga_clock.hrs_d[0] ),
    .B(_0643_));
 sg13g2_xnor2_1 _1379_ (.Y(_0652_),
    .A(_0616_),
    .B(_0651_));
 sg13g2_nor2_1 _1380_ (.A(_0650_),
    .B(_0652_),
    .Y(_0044_));
 sg13g2_buf_1 _1381_ (.A(net46),
    .X(_0653_));
 sg13g2_inv_1 _1382_ (.Y(_0654_),
    .A(\vga_clock.min_u[1] ));
 sg13g2_inv_1 _1383_ (.Y(_0655_),
    .A(\vga_clock.min_u[3] ));
 sg13g2_nor4_2 _1384_ (.A(_0654_),
    .B(_0573_),
    .C(\vga_clock.min_u[2] ),
    .Y(_0656_),
    .D(_0655_));
 sg13g2_mux2_1 _1385_ (.A0(\vga_clock.min_d[0] ),
    .A1(_0029_),
    .S(_0656_),
    .X(_0657_));
 sg13g2_nand3b_1 _1386_ (.B(\vga_clock.min_d[1] ),
    .C(\vga_clock.min_d[2] ),
    .Y(_0658_),
    .A_N(\vga_clock.min_d[0] ));
 sg13g2_and3_1 _1387_ (.X(_0049_),
    .A(net35),
    .B(_0657_),
    .C(_0658_));
 sg13g2_inv_2 _1388_ (.Y(_0659_),
    .A(net46));
 sg13g2_buf_1 _1389_ (.A(_0659_),
    .X(_0660_));
 sg13g2_inv_1 _1390_ (.Y(_0661_),
    .A(\vga_clock.min_d[1] ));
 sg13g2_xnor2_1 _1391_ (.Y(_0662_),
    .A(_0661_),
    .B(_0656_));
 sg13g2_nor3_1 _1392_ (.A(\vga_clock.min_d[0] ),
    .B(_0661_),
    .C(\vga_clock.min_d[2] ),
    .Y(_0663_));
 sg13g2_a21oi_1 _1393_ (.A1(\vga_clock.min_d[0] ),
    .A2(_0662_),
    .Y(_0664_),
    .B1(_0663_));
 sg13g2_nor2_1 _1394_ (.A(net25),
    .B(_0664_),
    .Y(_0050_));
 sg13g2_nor2_1 _1395_ (.A(_0661_),
    .B(\vga_clock.min_d[2] ),
    .Y(_0665_));
 sg13g2_mux2_1 _1396_ (.A0(\vga_clock.min_d[2] ),
    .A1(_0665_),
    .S(_0656_),
    .X(_0666_));
 sg13g2_a22oi_1 _1397_ (.Y(_0667_),
    .B1(_0666_),
    .B2(\vga_clock.min_d[0] ),
    .A2(\vga_clock.min_d[2] ),
    .A1(_0661_));
 sg13g2_nor2_1 _1398_ (.A(net25),
    .B(_0667_),
    .Y(_0051_));
 sg13g2_inv_1 _1399_ (.Y(_0668_),
    .A(_0031_));
 sg13g2_buf_1 _1400_ (.A(\vga_clock.sec_counter[20] ),
    .X(_0669_));
 sg13g2_buf_2 _1401_ (.A(\vga_clock.sec_counter[19] ),
    .X(_0670_));
 sg13g2_buf_2 _1402_ (.A(\vga_clock.sec_counter[18] ),
    .X(_0671_));
 sg13g2_and2_1 _1403_ (.A(\vga_clock.sec_counter[6] ),
    .B(\vga_clock.sec_counter[7] ),
    .X(_0672_));
 sg13g2_and4_1 _1404_ (.A(\vga_clock.sec_counter[3] ),
    .B(\vga_clock.sec_counter[2] ),
    .C(\vga_clock.sec_counter[1] ),
    .D(\vga_clock.sec_counter[0] ),
    .X(_0673_));
 sg13g2_and4_1 _1405_ (.A(\vga_clock.sec_counter[4] ),
    .B(\vga_clock.sec_counter[5] ),
    .C(_0672_),
    .D(_0673_),
    .X(_0674_));
 sg13g2_buf_2 _1406_ (.A(_0674_),
    .X(_0675_));
 sg13g2_inv_1 _1407_ (.Y(_0676_),
    .A(\vga_clock.sec_counter[14] ));
 sg13g2_inv_1 _1408_ (.Y(_0677_),
    .A(\vga_clock.sec_counter[15] ));
 sg13g2_buf_1 _1409_ (.A(\vga_clock.sec_counter[8] ),
    .X(_0678_));
 sg13g2_nand3_1 _1410_ (.B(\vga_clock.sec_counter[9] ),
    .C(\vga_clock.sec_counter[10] ),
    .A(_0678_),
    .Y(_0679_));
 sg13g2_buf_1 _1411_ (.A(\vga_clock.sec_counter[11] ),
    .X(_0680_));
 sg13g2_nand3_1 _1412_ (.B(_0680_),
    .C(\vga_clock.sec_counter[13] ),
    .A(\vga_clock.sec_counter[12] ),
    .Y(_0681_));
 sg13g2_nor4_1 _1413_ (.A(_0676_),
    .B(_0677_),
    .C(_0679_),
    .D(_0681_),
    .Y(_0682_));
 sg13g2_and4_1 _1414_ (.A(\vga_clock.sec_counter[17] ),
    .B(\vga_clock.sec_counter[16] ),
    .C(_0675_),
    .D(_0682_),
    .X(_0683_));
 sg13g2_buf_2 _1415_ (.A(_0683_),
    .X(_0684_));
 sg13g2_and4_1 _1416_ (.A(_0669_),
    .B(_0670_),
    .C(_0671_),
    .D(_0684_),
    .X(_0685_));
 sg13g2_xnor2_1 _1417_ (.Y(_0686_),
    .A(\vga_clock.sec_counter[21] ),
    .B(_0685_));
 sg13g2_buf_1 _1418_ (.A(\vga_clock.sec_counter[24] ),
    .X(_0687_));
 sg13g2_nor2b_1 _1419_ (.A(_0670_),
    .B_N(_0687_),
    .Y(_0688_));
 sg13g2_nand2_1 _1420_ (.Y(_0689_),
    .A(_0671_),
    .B(_0684_));
 sg13g2_inv_1 _1421_ (.Y(_0690_),
    .A(_0671_));
 sg13g2_nand2_1 _1422_ (.Y(_0691_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_nand3_1 _1423_ (.B(\vga_clock.sec_counter[22] ),
    .C(\vga_clock.sec_counter[21] ),
    .A(\vga_clock.sec_counter[23] ),
    .Y(_0692_));
 sg13g2_nor3_2 _1424_ (.A(_0690_),
    .B(_0691_),
    .C(_0692_),
    .Y(_0693_));
 sg13g2_xor2_1 _1425_ (.B(_0693_),
    .A(_0687_),
    .X(_0694_));
 sg13g2_and4_1 _1426_ (.A(_0670_),
    .B(_0671_),
    .C(_0684_),
    .D(_0694_),
    .X(_0695_));
 sg13g2_a21oi_1 _1427_ (.A1(_0688_),
    .A2(_0689_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_and2_1 _1428_ (.A(\vga_clock.sec_counter[22] ),
    .B(\vga_clock.sec_counter[21] ),
    .X(_0697_));
 sg13g2_or2_1 _1429_ (.X(_0698_),
    .B(_0670_),
    .A(_0669_));
 sg13g2_o21ai_1 _1430_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0691_),
    .A2(_0697_));
 sg13g2_inv_1 _1431_ (.Y(_0700_),
    .A(\vga_clock.sec_counter[23] ));
 sg13g2_and3_1 _1432_ (.X(_0701_),
    .A(_0700_),
    .B(_0669_),
    .C(_0670_));
 sg13g2_a22oi_1 _1433_ (.Y(_0702_),
    .B1(_0701_),
    .B2(_0697_),
    .A2(_0699_),
    .A1(\vga_clock.sec_counter[23] ));
 sg13g2_nand2_1 _1434_ (.Y(_0703_),
    .A(_0671_),
    .B(\vga_clock.sec_counter[17] ));
 sg13g2_or4_1 _1435_ (.A(_0700_),
    .B(_0669_),
    .C(_0671_),
    .D(\vga_clock.sec_counter[17] ),
    .X(_0704_));
 sg13g2_o21ai_1 _1436_ (.B1(_0704_),
    .Y(_0705_),
    .A1(_0702_),
    .A2(_0703_));
 sg13g2_nor2_1 _1437_ (.A(_0679_),
    .B(_0681_),
    .Y(_0706_));
 sg13g2_and4_1 _1438_ (.A(\vga_clock.sec_counter[14] ),
    .B(\vga_clock.sec_counter[15] ),
    .C(_0675_),
    .D(_0706_),
    .X(_0707_));
 sg13g2_buf_1 _1439_ (.A(_0707_),
    .X(_0708_));
 sg13g2_nand2_1 _1440_ (.Y(_0709_),
    .A(_0687_),
    .B(_0693_));
 sg13g2_and4_1 _1441_ (.A(\vga_clock.sec_counter[17] ),
    .B(\vga_clock.sec_counter[16] ),
    .C(_0708_),
    .D(_0709_),
    .X(_0710_));
 sg13g2_nor3_1 _1442_ (.A(\vga_clock.sec_counter[16] ),
    .B(_0708_),
    .C(_0704_),
    .Y(_0711_));
 sg13g2_a21oi_1 _1443_ (.A1(_0705_),
    .A2(_0710_),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_nand3_1 _1444_ (.B(_0675_),
    .C(_0706_),
    .A(\vga_clock.sec_counter[14] ),
    .Y(_0713_));
 sg13g2_xnor2_1 _1445_ (.Y(_0714_),
    .A(_0677_),
    .B(_0713_));
 sg13g2_nand2_1 _1446_ (.Y(_0715_),
    .A(_0678_),
    .B(_0675_));
 sg13g2_xor2_1 _1447_ (.B(_0715_),
    .A(\vga_clock.sec_counter[9] ),
    .X(_0716_));
 sg13g2_and2_1 _1448_ (.A(\vga_clock.sec_counter[4] ),
    .B(_0673_),
    .X(_0717_));
 sg13g2_buf_1 _1449_ (.A(_0717_),
    .X(_0718_));
 sg13g2_nor2b_1 _1450_ (.A(\vga_clock.sec_counter[14] ),
    .B_N(\vga_clock.sec_counter[22] ),
    .Y(_0719_));
 sg13g2_inv_1 _1451_ (.Y(_0720_),
    .A(\vga_clock.sec_counter[10] ));
 sg13g2_nor4_1 _1452_ (.A(\vga_clock.sec_counter[5] ),
    .B(_0678_),
    .C(_0720_),
    .D(\vga_clock.sec_counter[25] ),
    .Y(_0721_));
 sg13g2_nand4_1 _1453_ (.B(_0718_),
    .C(_0719_),
    .A(_0672_),
    .Y(_0722_),
    .D(_0721_));
 sg13g2_nor2_1 _1454_ (.A(\vga_clock.sec_counter[12] ),
    .B(_0680_),
    .Y(_0723_));
 sg13g2_nand2_1 _1455_ (.Y(_0724_),
    .A(\vga_clock.sec_counter[13] ),
    .B(_0723_));
 sg13g2_nand3b_1 _1456_ (.B(_0680_),
    .C(\vga_clock.sec_counter[12] ),
    .Y(_0725_),
    .A_N(\vga_clock.sec_counter[13] ));
 sg13g2_and4_1 _1457_ (.A(_0678_),
    .B(\vga_clock.sec_counter[9] ),
    .C(\vga_clock.sec_counter[10] ),
    .D(_0675_),
    .X(_0726_));
 sg13g2_buf_1 _1458_ (.A(_0726_),
    .X(_0727_));
 sg13g2_mux2_1 _1459_ (.A0(_0724_),
    .A1(_0725_),
    .S(_0727_),
    .X(_0728_));
 sg13g2_or4_1 _1460_ (.A(_0714_),
    .B(_0716_),
    .C(_0722_),
    .D(_0728_),
    .X(_0729_));
 sg13g2_nor4_2 _1461_ (.A(_0686_),
    .B(_0696_),
    .C(_0712_),
    .Y(_0730_),
    .D(_0729_));
 sg13g2_nand2b_1 _1462_ (.Y(_0731_),
    .B(net46),
    .A_N(_0730_));
 sg13g2_buf_2 _1463_ (.A(_0731_),
    .X(_0732_));
 sg13g2_buf_1 _1464_ (.A(_0732_),
    .X(_0733_));
 sg13g2_nor2_1 _1465_ (.A(_0668_),
    .B(net10),
    .Y(_0086_));
 sg13g2_nand3_1 _1466_ (.B(\vga_clock.sec_counter[9] ),
    .C(_0675_),
    .A(_0678_),
    .Y(_0734_));
 sg13g2_xnor2_1 _1467_ (.Y(_0735_),
    .A(_0720_),
    .B(_0734_));
 sg13g2_nor2_1 _1468_ (.A(net10),
    .B(_0735_),
    .Y(_0087_));
 sg13g2_xnor2_1 _1469_ (.Y(_0736_),
    .A(_0680_),
    .B(_0727_));
 sg13g2_nor2_1 _1470_ (.A(net10),
    .B(_0736_),
    .Y(_0088_));
 sg13g2_nand2_1 _1471_ (.Y(_0737_),
    .A(_0680_),
    .B(_0727_));
 sg13g2_xor2_1 _1472_ (.B(_0737_),
    .A(\vga_clock.sec_counter[12] ),
    .X(_0738_));
 sg13g2_nor2_1 _1473_ (.A(net10),
    .B(_0738_),
    .Y(_0089_));
 sg13g2_nand3_1 _1474_ (.B(_0680_),
    .C(_0727_),
    .A(\vga_clock.sec_counter[12] ),
    .Y(_0739_));
 sg13g2_xor2_1 _1475_ (.B(_0739_),
    .A(\vga_clock.sec_counter[13] ),
    .X(_0740_));
 sg13g2_nor2_1 _1476_ (.A(_0733_),
    .B(_0740_),
    .Y(_0090_));
 sg13g2_nand2_1 _1477_ (.Y(_0741_),
    .A(_0675_),
    .B(_0706_));
 sg13g2_xnor2_1 _1478_ (.Y(_0742_),
    .A(_0676_),
    .B(_0741_));
 sg13g2_nor2_1 _1479_ (.A(net10),
    .B(_0742_),
    .Y(_0091_));
 sg13g2_nor2_1 _1480_ (.A(_0714_),
    .B(net10),
    .Y(_0092_));
 sg13g2_xnor2_1 _1481_ (.Y(_0743_),
    .A(\vga_clock.sec_counter[16] ),
    .B(_0708_));
 sg13g2_nor2_1 _1482_ (.A(net10),
    .B(_0743_),
    .Y(_0093_));
 sg13g2_buf_1 _1483_ (.A(_0732_),
    .X(_0744_));
 sg13g2_nand2_1 _1484_ (.Y(_0745_),
    .A(\vga_clock.sec_counter[16] ),
    .B(_0708_));
 sg13g2_xor2_1 _1485_ (.B(_0745_),
    .A(\vga_clock.sec_counter[17] ),
    .X(_0746_));
 sg13g2_nor2_1 _1486_ (.A(_0744_),
    .B(_0746_),
    .Y(_0094_));
 sg13g2_xnor2_1 _1487_ (.Y(_0747_),
    .A(_0671_),
    .B(_0684_));
 sg13g2_nor2_1 _1488_ (.A(net9),
    .B(_0747_),
    .Y(_0095_));
 sg13g2_xor2_1 _1489_ (.B(_0689_),
    .A(_0670_),
    .X(_0748_));
 sg13g2_nor2_1 _1490_ (.A(net25),
    .B(_0748_),
    .Y(_0096_));
 sg13g2_xnor2_1 _1491_ (.Y(_0749_),
    .A(\vga_clock.sec_counter[1] ),
    .B(\vga_clock.sec_counter[0] ));
 sg13g2_nor2_1 _1492_ (.A(net9),
    .B(_0749_),
    .Y(_0097_));
 sg13g2_buf_1 _1493_ (.A(net46),
    .X(_0750_));
 sg13g2_nand3_1 _1494_ (.B(_0671_),
    .C(_0684_),
    .A(_0670_),
    .Y(_0751_));
 sg13g2_xnor2_1 _1495_ (.Y(_0752_),
    .A(_0669_),
    .B(_0751_));
 sg13g2_and2_1 _1496_ (.A(net34),
    .B(_0752_),
    .X(_0098_));
 sg13g2_nor2_1 _1497_ (.A(_0686_),
    .B(net10),
    .Y(_0099_));
 sg13g2_nand2_1 _1498_ (.Y(_0753_),
    .A(\vga_clock.sec_counter[21] ),
    .B(_0685_));
 sg13g2_xor2_1 _1499_ (.B(_0753_),
    .A(\vga_clock.sec_counter[22] ),
    .X(_0754_));
 sg13g2_nor2_1 _1500_ (.A(net9),
    .B(_0754_),
    .Y(_0100_));
 sg13g2_nand2_1 _1501_ (.Y(_0755_),
    .A(_0685_),
    .B(_0697_));
 sg13g2_xnor2_1 _1502_ (.Y(_0756_),
    .A(_0700_),
    .B(_0755_));
 sg13g2_nor2_1 _1503_ (.A(net9),
    .B(_0756_),
    .Y(_0101_));
 sg13g2_and2_1 _1504_ (.A(_0684_),
    .B(_0693_),
    .X(_0757_));
 sg13g2_xnor2_1 _1505_ (.Y(_0758_),
    .A(_0687_),
    .B(_0757_));
 sg13g2_nor2_1 _1506_ (.A(_0744_),
    .B(_0758_),
    .Y(_0102_));
 sg13g2_nand2_1 _1507_ (.Y(_0759_),
    .A(_0687_),
    .B(_0757_));
 sg13g2_xor2_1 _1508_ (.B(_0759_),
    .A(\vga_clock.sec_counter[25] ),
    .X(_0760_));
 sg13g2_nor2_1 _1509_ (.A(net25),
    .B(_0760_),
    .Y(_0103_));
 sg13g2_nand2_1 _1510_ (.Y(_0761_),
    .A(\vga_clock.sec_counter[1] ),
    .B(\vga_clock.sec_counter[0] ));
 sg13g2_xor2_1 _1511_ (.B(_0761_),
    .A(\vga_clock.sec_counter[2] ),
    .X(_0762_));
 sg13g2_nor2_1 _1512_ (.A(net9),
    .B(_0762_),
    .Y(_0104_));
 sg13g2_nand3_1 _1513_ (.B(\vga_clock.sec_counter[1] ),
    .C(\vga_clock.sec_counter[0] ),
    .A(\vga_clock.sec_counter[2] ),
    .Y(_0763_));
 sg13g2_xor2_1 _1514_ (.B(_0763_),
    .A(\vga_clock.sec_counter[3] ),
    .X(_0764_));
 sg13g2_nor2_1 _1515_ (.A(net9),
    .B(_0764_),
    .Y(_0105_));
 sg13g2_xnor2_1 _1516_ (.Y(_0765_),
    .A(\vga_clock.sec_counter[4] ),
    .B(_0673_));
 sg13g2_nor2_1 _1517_ (.A(net9),
    .B(_0765_),
    .Y(_0106_));
 sg13g2_xnor2_1 _1518_ (.Y(_0766_),
    .A(\vga_clock.sec_counter[5] ),
    .B(_0718_));
 sg13g2_nor2_1 _1519_ (.A(net9),
    .B(_0766_),
    .Y(_0107_));
 sg13g2_nand2_1 _1520_ (.Y(_0767_),
    .A(\vga_clock.sec_counter[5] ),
    .B(_0718_));
 sg13g2_xor2_1 _1521_ (.B(_0767_),
    .A(\vga_clock.sec_counter[6] ),
    .X(_0768_));
 sg13g2_nor2_1 _1522_ (.A(_0732_),
    .B(_0768_),
    .Y(_0108_));
 sg13g2_nand3_1 _1523_ (.B(\vga_clock.sec_counter[6] ),
    .C(_0718_),
    .A(\vga_clock.sec_counter[5] ),
    .Y(_0769_));
 sg13g2_xor2_1 _1524_ (.B(_0769_),
    .A(\vga_clock.sec_counter[7] ),
    .X(_0770_));
 sg13g2_nor2_1 _1525_ (.A(_0732_),
    .B(_0770_),
    .Y(_0109_));
 sg13g2_xnor2_1 _1526_ (.Y(_0771_),
    .A(_0678_),
    .B(_0675_));
 sg13g2_nor2_1 _1527_ (.A(_0732_),
    .B(_0771_),
    .Y(_0110_));
 sg13g2_nor2_1 _1528_ (.A(_0716_),
    .B(_0733_),
    .Y(_0111_));
 sg13g2_nor2b_1 _1529_ (.A(\vga_clock.sec_u[2] ),
    .B_N(\vga_clock.sec_u[3] ),
    .Y(_0772_));
 sg13g2_nor2b_1 _1530_ (.A(\vga_clock.sec_u[0] ),
    .B_N(\vga_clock.sec_u[1] ),
    .Y(_0773_));
 sg13g2_nand2_1 _1531_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_o21ai_1 _1532_ (.B1(net46),
    .Y(_0775_),
    .A1(_0027_),
    .A2(_0774_));
 sg13g2_and2_1 _1533_ (.A(_0772_),
    .B(_0773_),
    .X(_0776_));
 sg13g2_nand2_1 _1534_ (.Y(_0777_),
    .A(\vga_clock.sec_d[1] ),
    .B(\vga_clock.sec_d[2] ));
 sg13g2_a21oi_1 _1535_ (.A1(_0776_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(_0577_));
 sg13g2_nor2_1 _1536_ (.A(_0775_),
    .B(_0778_),
    .Y(_0112_));
 sg13g2_inv_1 _1537_ (.Y(_0779_),
    .A(\vga_clock.sec_d[1] ));
 sg13g2_xnor2_1 _1538_ (.Y(_0780_),
    .A(_0779_),
    .B(_0776_));
 sg13g2_nor3_1 _1539_ (.A(_0577_),
    .B(_0779_),
    .C(\vga_clock.sec_d[2] ),
    .Y(_0781_));
 sg13g2_a21oi_1 _1540_ (.A1(_0577_),
    .A2(_0780_),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_nor2_1 _1541_ (.A(net25),
    .B(_0782_),
    .Y(_0113_));
 sg13g2_nor2_1 _1542_ (.A(_0779_),
    .B(\vga_clock.sec_d[2] ),
    .Y(_0783_));
 sg13g2_mux2_1 _1543_ (.A0(\vga_clock.sec_d[2] ),
    .A1(_0783_),
    .S(_0776_),
    .X(_0784_));
 sg13g2_a22oi_1 _1544_ (.Y(_0785_),
    .B1(_0784_),
    .B2(_0577_),
    .A2(\vga_clock.sec_d[2] ),
    .A1(_0779_));
 sg13g2_nor2_1 _1545_ (.A(net25),
    .B(_0785_),
    .Y(_0114_));
 sg13g2_buf_2 _1546_ (.A(ui_in[1]),
    .X(_0786_));
 sg13g2_inv_1 _1547_ (.Y(_0787_),
    .A(_0786_));
 sg13g2_inv_1 _1548_ (.Y(_0788_),
    .A(\vga_clock.pulse_min.count[2] ));
 sg13g2_buf_2 _1549_ (.A(\vga_clock.pulse_min.count[1] ),
    .X(_0789_));
 sg13g2_buf_1 _1550_ (.A(\vga_clock.pulse_min.count[0] ),
    .X(_0790_));
 sg13g2_nor3_1 _1551_ (.A(_0789_),
    .B(net33),
    .C(\vga_clock.pulse_min.count[3] ),
    .Y(_0791_));
 sg13g2_nand3_1 _1552_ (.B(_0014_),
    .C(_0791_),
    .A(_0788_),
    .Y(_0792_));
 sg13g2_nand2_1 _1553_ (.Y(_0793_),
    .A(_0402_),
    .B(_0566_));
 sg13g2_nor2_1 _1554_ (.A(\vga_clock.vga_0.y_px[2] ),
    .B(\vga_clock.vga_0.x_px[0] ),
    .Y(_0794_));
 sg13g2_nor4_1 _1555_ (.A(net37),
    .B(net39),
    .C(\vga_clock.vga_0.y_px[9] ),
    .D(\vga_clock.vga_0.y_px[8] ),
    .Y(_0795_));
 sg13g2_nand2_1 _1556_ (.Y(_0796_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nor4_1 _1557_ (.A(\vga_clock.vga_0.y_px[0] ),
    .B(\vga_clock.vga_0.x_px[1] ),
    .C(\vga_clock.vga_0.x_px[3] ),
    .D(\vga_clock.vga_0.x_px[2] ),
    .Y(_0797_));
 sg13g2_nor4_1 _1558_ (.A(\vga_clock.vga_0.y_px[1] ),
    .B(\vga_clock.digit_0.x_block[1] ),
    .C(\vga_clock.digit_0.x_block[0] ),
    .D(_0564_),
    .Y(_0798_));
 sg13g2_nand2_1 _1559_ (.Y(_0799_),
    .A(_0797_),
    .B(_0798_));
 sg13g2_or3_1 _1560_ (.A(_0793_),
    .B(_0796_),
    .C(_0799_),
    .X(_0800_));
 sg13g2_buf_1 _1561_ (.A(_0800_),
    .X(_0801_));
 sg13g2_nor3_1 _1562_ (.A(_0787_),
    .B(_0792_),
    .C(net18),
    .Y(_0802_));
 sg13g2_nor2_1 _1563_ (.A(_0577_),
    .B(_0777_),
    .Y(_0803_));
 sg13g2_or2_1 _1564_ (.X(_0804_),
    .B(_0803_),
    .A(_0802_));
 sg13g2_buf_2 _1565_ (.A(_0804_),
    .X(_0805_));
 sg13g2_mux2_1 _1566_ (.A0(_0374_),
    .A1(_0028_),
    .S(_0805_),
    .X(_0806_));
 sg13g2_and2_1 _1567_ (.A(net34),
    .B(_0806_),
    .X(_0032_));
 sg13g2_nand2_1 _1568_ (.Y(_0807_),
    .A(_0374_),
    .B(_0805_));
 sg13g2_xor2_1 _1569_ (.B(_0807_),
    .A(_0370_),
    .X(_0808_));
 sg13g2_nor2_1 _1570_ (.A(net25),
    .B(_0808_),
    .Y(_0033_));
 sg13g2_nand3_1 _1571_ (.B(_0374_),
    .C(_0805_),
    .A(_0370_),
    .Y(_0809_));
 sg13g2_xnor2_1 _1572_ (.Y(_0810_),
    .A(\vga_clock.color_offset[2] ),
    .B(_0809_));
 sg13g2_and2_1 _1573_ (.A(net34),
    .B(_0810_),
    .X(_0034_));
 sg13g2_a21oi_1 _1574_ (.A1(_0568_),
    .A2(_0381_),
    .Y(_0811_),
    .B1(_0639_));
 sg13g2_o21ai_1 _1575_ (.B1(_0637_),
    .Y(_0812_),
    .A1(_0568_),
    .A2(_0367_));
 sg13g2_a22oi_1 _1576_ (.Y(_0813_),
    .B1(_0812_),
    .B2(_0378_),
    .A2(_0386_),
    .A1(_0381_));
 sg13g2_o21ai_1 _1577_ (.B1(_0813_),
    .Y(_0040_),
    .A1(_0375_),
    .A2(_0811_));
 sg13g2_nand2b_1 _1578_ (.Y(_0814_),
    .B(\vga_clock.font_0.dout[1] ),
    .A_N(\vga_clock.col_index_q[0] ));
 sg13g2_nand2b_1 _1579_ (.Y(_0815_),
    .B(\vga_clock.col_index_q[0] ),
    .A_N(\vga_clock.font_0.dout[2] ));
 sg13g2_nor4_1 _1580_ (.A(\vga_clock.x_block_q[5] ),
    .B(\vga_clock.y_block_q[5] ),
    .C(\vga_clock.y_block_q[4] ),
    .D(\vga_clock.y_block_q[3] ),
    .Y(_0816_));
 sg13g2_o21ai_1 _1581_ (.B1(\vga_clock.y_block_q[2] ),
    .Y(_0817_),
    .A1(\vga_clock.y_block_q[1] ),
    .A2(\vga_clock.y_block_q[0] ));
 sg13g2_or3_1 _1582_ (.A(\vga_clock.font_0.dout[3] ),
    .B(\vga_clock.col_index_q[0] ),
    .C(\vga_clock.col_index_q[1] ),
    .X(_0818_));
 sg13g2_nand4_1 _1583_ (.B(_0816_),
    .C(_0817_),
    .A(_0815_),
    .Y(_0819_),
    .D(_0818_));
 sg13g2_a21oi_1 _1584_ (.A1(\vga_clock.col_index_q[1] ),
    .A2(_0814_),
    .Y(_0042_),
    .B1(_0819_));
 sg13g2_nand2_1 _1585_ (.Y(_0820_),
    .A(_0649_),
    .B(_0645_));
 sg13g2_buf_1 _1586_ (.A(ui_in[0]),
    .X(_0821_));
 sg13g2_nor3_2 _1587_ (.A(_0793_),
    .B(_0796_),
    .C(_0799_),
    .Y(_0822_));
 sg13g2_buf_2 _1588_ (.A(\vga_clock.pulse_hrs.count[1] ),
    .X(_0823_));
 sg13g2_buf_2 _1589_ (.A(\vga_clock.pulse_hrs.count[0] ),
    .X(_0824_));
 sg13g2_nor4_1 _1590_ (.A(_0823_),
    .B(_0824_),
    .C(\vga_clock.pulse_hrs.count[3] ),
    .D(\vga_clock.pulse_hrs.count[2] ),
    .Y(_0825_));
 sg13g2_and2_1 _1591_ (.A(_0013_),
    .B(_0825_),
    .X(_0826_));
 sg13g2_nand3_1 _1592_ (.B(_0822_),
    .C(_0826_),
    .A(net45),
    .Y(_0827_));
 sg13g2_o21ai_1 _1593_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_0658_),
    .A2(_0820_));
 sg13g2_nand2_1 _1594_ (.Y(_0829_),
    .A(_0658_),
    .B(_0827_));
 sg13g2_nor2_1 _1595_ (.A(_0820_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_a22oi_1 _1596_ (.Y(_0831_),
    .B1(_0830_),
    .B2(_0586_),
    .A2(_0828_),
    .A1(_0011_));
 sg13g2_nor2_1 _1597_ (.A(net25),
    .B(_0831_),
    .Y(_0045_));
 sg13g2_buf_1 _1598_ (.A(_0659_),
    .X(_0832_));
 sg13g2_nand2_1 _1599_ (.Y(_0833_),
    .A(\vga_clock.hrs_u[1] ),
    .B(_0586_));
 sg13g2_a21oi_1 _1600_ (.A1(_0658_),
    .A2(_0827_),
    .Y(_0834_),
    .B1(_0833_));
 sg13g2_a21oi_1 _1601_ (.A1(_0586_),
    .A2(_0829_),
    .Y(_0835_),
    .B1(\vga_clock.hrs_u[1] ));
 sg13g2_and2_1 _1602_ (.A(_0827_),
    .B(_0820_),
    .X(_0836_));
 sg13g2_nor4_1 _1603_ (.A(net24),
    .B(_0834_),
    .C(_0835_),
    .D(_0836_),
    .Y(_0046_));
 sg13g2_xor2_1 _1604_ (.B(_0833_),
    .A(_0019_),
    .X(_0837_));
 sg13g2_a22oi_1 _1605_ (.Y(_0838_),
    .B1(_0837_),
    .B2(_0828_),
    .A2(_0830_),
    .A1(\vga_clock.hrs_u[2] ));
 sg13g2_nor2_1 _1606_ (.A(_0660_),
    .B(_0838_),
    .Y(_0047_));
 sg13g2_nand3_1 _1607_ (.B(_0586_),
    .C(\vga_clock.hrs_u[2] ),
    .A(\vga_clock.hrs_u[1] ),
    .Y(_0839_));
 sg13g2_xor2_1 _1608_ (.B(_0839_),
    .A(_0020_),
    .X(_0840_));
 sg13g2_a22oi_1 _1609_ (.Y(_0841_),
    .B1(_0840_),
    .B2(_0828_),
    .A2(_0830_),
    .A1(\vga_clock.hrs_u[3] ));
 sg13g2_nor2_1 _1610_ (.A(_0660_),
    .B(_0841_),
    .Y(_0048_));
 sg13g2_nor2_1 _1611_ (.A(_0656_),
    .B(_0805_),
    .Y(_0842_));
 sg13g2_nand2_1 _1612_ (.Y(_0843_),
    .A(_0573_),
    .B(_0842_));
 sg13g2_o21ai_1 _1613_ (.B1(_0010_),
    .Y(_0844_),
    .A1(_0656_),
    .A2(_0805_));
 sg13g2_inv_1 _1614_ (.Y(_0845_),
    .A(_0656_));
 sg13g2_o21ai_1 _1615_ (.B1(net46),
    .Y(_0846_),
    .A1(_0845_),
    .A2(_0802_));
 sg13g2_a21oi_1 _1616_ (.A1(_0843_),
    .A2(_0844_),
    .Y(_0052_),
    .B1(_0846_));
 sg13g2_nand2_1 _1617_ (.Y(_0847_),
    .A(_0573_),
    .B(_0805_));
 sg13g2_xnor2_1 _1618_ (.Y(_0848_),
    .A(_0654_),
    .B(_0847_));
 sg13g2_nor2_1 _1619_ (.A(_0846_),
    .B(_0848_),
    .Y(_0053_));
 sg13g2_nand3_1 _1620_ (.B(_0573_),
    .C(_0805_),
    .A(\vga_clock.min_u[1] ),
    .Y(_0849_));
 sg13g2_xor2_1 _1621_ (.B(_0849_),
    .A(\vga_clock.min_u[2] ),
    .X(_0850_));
 sg13g2_nor2_1 _1622_ (.A(_0846_),
    .B(_0850_),
    .Y(_0054_));
 sg13g2_nand3_1 _1623_ (.B(_0573_),
    .C(\vga_clock.min_u[2] ),
    .A(\vga_clock.min_u[1] ),
    .Y(_0851_));
 sg13g2_xor2_1 _1624_ (.B(_0851_),
    .A(_0021_),
    .X(_0852_));
 sg13g2_nor2_1 _1625_ (.A(_0842_),
    .B(_0852_),
    .Y(_0853_));
 sg13g2_nor2_1 _1626_ (.A(\vga_clock.min_u[3] ),
    .B(_0805_),
    .Y(_0854_));
 sg13g2_nor3_1 _1627_ (.A(_0846_),
    .B(_0853_),
    .C(_0854_),
    .Y(_0055_));
 sg13g2_buf_1 _1628_ (.A(net46),
    .X(_0855_));
 sg13g2_buf_1 _1629_ (.A(\vga_clock.pulse_hrs.comp[0] ),
    .X(_0856_));
 sg13g2_nor3_1 _1630_ (.A(\vga_clock.pulse_hrs.comp[3] ),
    .B(\vga_clock.pulse_hrs.comp[4] ),
    .C(\vga_clock.pulse_hrs.comp[2] ),
    .Y(_0857_));
 sg13g2_nand2b_1 _1631_ (.Y(_0858_),
    .B(_0826_),
    .A_N(_0857_));
 sg13g2_a21oi_1 _1632_ (.A1(net45),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0801_));
 sg13g2_nand2_1 _1633_ (.Y(_0860_),
    .A(net45),
    .B(_0859_));
 sg13g2_nor2b_1 _1634_ (.A(_0856_),
    .B_N(_0859_),
    .Y(_0861_));
 sg13g2_a21oi_1 _1635_ (.A1(_0856_),
    .A2(_0860_),
    .Y(_0862_),
    .B1(_0861_));
 sg13g2_nand2_1 _1636_ (.Y(_0056_),
    .A(_0855_),
    .B(_0862_));
 sg13g2_buf_2 _1637_ (.A(\vga_clock.pulse_hrs.comp[1] ),
    .X(_0863_));
 sg13g2_buf_1 _1638_ (.A(_0822_),
    .X(_0864_));
 sg13g2_nor2_1 _1639_ (.A(_0856_),
    .B(_0858_),
    .Y(_0865_));
 sg13g2_nand3_1 _1640_ (.B(net17),
    .C(_0865_),
    .A(_0863_),
    .Y(_0866_));
 sg13g2_o21ai_1 _1641_ (.B1(_0866_),
    .Y(_0867_),
    .A1(_0863_),
    .A2(_0865_));
 sg13g2_nand2_1 _1642_ (.Y(_0868_),
    .A(net45),
    .B(_0867_));
 sg13g2_o21ai_1 _1643_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_0863_),
    .A2(net17));
 sg13g2_nand2_1 _1644_ (.Y(_0057_),
    .A(net32),
    .B(_0869_));
 sg13g2_nand2b_1 _1645_ (.Y(_0870_),
    .B(_0865_),
    .A_N(_0863_));
 sg13g2_a21oi_1 _1646_ (.A1(net45),
    .A2(_0870_),
    .Y(_0871_),
    .B1(net18));
 sg13g2_nor3_1 _1647_ (.A(_0856_),
    .B(_0863_),
    .C(_0858_),
    .Y(_0872_));
 sg13g2_nand4_1 _1648_ (.B(net45),
    .C(net17),
    .A(\vga_clock.pulse_hrs.comp[2] ),
    .Y(_0873_),
    .D(_0872_));
 sg13g2_o21ai_1 _1649_ (.B1(_0873_),
    .Y(_0874_),
    .A1(\vga_clock.pulse_hrs.comp[2] ),
    .A2(_0871_));
 sg13g2_nand2_1 _1650_ (.Y(_0058_),
    .A(_0855_),
    .B(_0874_));
 sg13g2_or3_1 _1651_ (.A(\vga_clock.pulse_hrs.comp[2] ),
    .B(_0856_),
    .C(_0863_),
    .X(_0875_));
 sg13g2_nand2_1 _1652_ (.Y(_0876_),
    .A(net45),
    .B(_0875_));
 sg13g2_a21oi_1 _1653_ (.A1(_0859_),
    .A2(_0876_),
    .Y(_0877_),
    .B1(\vga_clock.pulse_hrs.comp[3] ));
 sg13g2_inv_1 _1654_ (.Y(_0878_),
    .A(\vga_clock.pulse_hrs.comp[3] ));
 sg13g2_nor3_1 _1655_ (.A(_0878_),
    .B(_0860_),
    .C(_0875_),
    .Y(_0879_));
 sg13g2_o21ai_1 _1656_ (.B1(net32),
    .Y(_0059_),
    .A1(_0877_),
    .A2(_0879_));
 sg13g2_o21ai_1 _1657_ (.B1(_0821_),
    .Y(_0880_),
    .A1(\vga_clock.pulse_hrs.comp[3] ),
    .A2(_0875_));
 sg13g2_nand2_1 _1658_ (.Y(_0881_),
    .A(\vga_clock.pulse_hrs.comp[4] ),
    .B(net35));
 sg13g2_a21oi_1 _1659_ (.A1(_0859_),
    .A2(_0880_),
    .Y(_0060_),
    .B1(_0881_));
 sg13g2_buf_1 _1660_ (.A(_0659_),
    .X(_0882_));
 sg13g2_buf_1 _1661_ (.A(net18),
    .X(_0883_));
 sg13g2_xor2_1 _1662_ (.B(\vga_clock.pulse_hrs.comp[3] ),
    .A(\vga_clock.pulse_hrs.count[3] ),
    .X(_0884_));
 sg13g2_xor2_1 _1663_ (.B(_0863_),
    .A(_0823_),
    .X(_0885_));
 sg13g2_xor2_1 _1664_ (.B(\vga_clock.pulse_hrs.count[4] ),
    .A(\vga_clock.pulse_hrs.comp[4] ),
    .X(_0886_));
 sg13g2_nor3_1 _1665_ (.A(_0884_),
    .B(_0885_),
    .C(_0886_),
    .Y(_0887_));
 sg13g2_xnor2_1 _1666_ (.Y(_0888_),
    .A(\vga_clock.pulse_hrs.count[2] ),
    .B(\vga_clock.pulse_hrs.comp[2] ));
 sg13g2_xnor2_1 _1667_ (.Y(_0889_),
    .A(_0824_),
    .B(_0856_));
 sg13g2_nand3_1 _1668_ (.B(_0888_),
    .C(_0889_),
    .A(_0887_),
    .Y(_0890_));
 sg13g2_nand3_1 _1669_ (.B(net17),
    .C(_0890_),
    .A(net45),
    .Y(_0891_));
 sg13g2_nor2_1 _1670_ (.A(_0824_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_a21oi_1 _1671_ (.A1(_0824_),
    .A2(_0883_),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_nor2_1 _1672_ (.A(_0882_),
    .B(_0893_),
    .Y(_0061_));
 sg13g2_o21ai_1 _1673_ (.B1(_0823_),
    .Y(_0894_),
    .A1(_0883_),
    .A2(_0892_));
 sg13g2_inv_1 _1674_ (.Y(_0895_),
    .A(_0891_));
 sg13g2_nand3b_1 _1675_ (.B(_0824_),
    .C(_0895_),
    .Y(_0896_),
    .A_N(_0823_));
 sg13g2_a21oi_1 _1676_ (.A1(_0894_),
    .A2(_0896_),
    .Y(_0062_),
    .B1(net24));
 sg13g2_a21oi_1 _1677_ (.A1(_0823_),
    .A2(_0824_),
    .Y(_0897_),
    .B1(_0891_));
 sg13g2_o21ai_1 _1678_ (.B1(\vga_clock.pulse_hrs.count[2] ),
    .Y(_0898_),
    .A1(net14),
    .A2(_0897_));
 sg13g2_inv_1 _1679_ (.Y(_0899_),
    .A(\vga_clock.pulse_hrs.count[2] ));
 sg13g2_nand4_1 _1680_ (.B(_0824_),
    .C(_0899_),
    .A(_0823_),
    .Y(_0900_),
    .D(_0895_));
 sg13g2_a21oi_1 _1681_ (.A1(_0898_),
    .A2(_0900_),
    .Y(_0063_),
    .B1(net24));
 sg13g2_and3_1 _1682_ (.X(_0901_),
    .A(_0823_),
    .B(_0824_),
    .C(\vga_clock.pulse_hrs.count[2] ));
 sg13g2_o21ai_1 _1683_ (.B1(_0864_),
    .Y(_0902_),
    .A1(_0891_),
    .A2(_0901_));
 sg13g2_nor2b_1 _1684_ (.A(\vga_clock.pulse_hrs.count[3] ),
    .B_N(_0901_),
    .Y(_0903_));
 sg13g2_a22oi_1 _1685_ (.Y(_0904_),
    .B1(_0903_),
    .B2(_0895_),
    .A2(_0902_),
    .A1(\vga_clock.pulse_hrs.count[3] ));
 sg13g2_nor2_1 _1686_ (.A(net23),
    .B(_0904_),
    .Y(_0064_));
 sg13g2_nand2_1 _1687_ (.Y(_0905_),
    .A(\vga_clock.pulse_hrs.count[3] ),
    .B(_0901_));
 sg13g2_xor2_1 _1688_ (.B(_0905_),
    .A(_0013_),
    .X(_0906_));
 sg13g2_a22oi_1 _1689_ (.Y(_0907_),
    .B1(_0895_),
    .B2(_0906_),
    .A2(net14),
    .A1(\vga_clock.pulse_hrs.count[4] ));
 sg13g2_nor2_1 _1690_ (.A(net23),
    .B(_0907_),
    .Y(_0065_));
 sg13g2_buf_2 _1691_ (.A(\vga_clock.pulse_min.comp[0] ),
    .X(_0908_));
 sg13g2_nor3_1 _1692_ (.A(\vga_clock.pulse_min.comp[3] ),
    .B(\vga_clock.pulse_min.comp[4] ),
    .C(\vga_clock.pulse_min.comp[2] ),
    .Y(_0909_));
 sg13g2_or2_1 _1693_ (.X(_0910_),
    .B(_0909_),
    .A(_0792_));
 sg13g2_a21oi_2 _1694_ (.B1(net18),
    .Y(_0911_),
    .A2(_0910_),
    .A1(_0786_));
 sg13g2_nand3_1 _1695_ (.B(_0908_),
    .C(_0911_),
    .A(_0786_),
    .Y(_0912_));
 sg13g2_o21ai_1 _1696_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0908_),
    .A2(_0911_));
 sg13g2_nand2_1 _1697_ (.Y(_0066_),
    .A(net32),
    .B(_0913_));
 sg13g2_buf_1 _1698_ (.A(\vga_clock.pulse_min.comp[1] ),
    .X(_0914_));
 sg13g2_nor2b_1 _1699_ (.A(_0908_),
    .B_N(_0914_),
    .Y(_0915_));
 sg13g2_nor2b_1 _1700_ (.A(_0914_),
    .B_N(_0908_),
    .Y(_0916_));
 sg13g2_a21oi_1 _1701_ (.A1(_0911_),
    .A2(_0915_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_or2_1 _1702_ (.X(_0918_),
    .B(_0911_),
    .A(_0914_));
 sg13g2_o21ai_1 _1703_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0787_),
    .A2(_0917_));
 sg13g2_nand2_1 _1704_ (.Y(_0067_),
    .A(net32),
    .B(_0919_));
 sg13g2_nor3_1 _1705_ (.A(_0908_),
    .B(_0914_),
    .C(_0910_),
    .Y(_0920_));
 sg13g2_o21ai_1 _1706_ (.B1(net17),
    .Y(_0921_),
    .A1(_0787_),
    .A2(_0920_));
 sg13g2_nor2b_1 _1707_ (.A(\vga_clock.pulse_min.comp[2] ),
    .B_N(_0921_),
    .Y(_0922_));
 sg13g2_and4_1 _1708_ (.A(\vga_clock.pulse_min.comp[2] ),
    .B(_0786_),
    .C(net17),
    .D(_0920_),
    .X(_0923_));
 sg13g2_o21ai_1 _1709_ (.B1(net34),
    .Y(_0068_),
    .A1(_0922_),
    .A2(_0923_));
 sg13g2_or3_1 _1710_ (.A(\vga_clock.pulse_min.comp[2] ),
    .B(_0908_),
    .C(_0914_),
    .X(_0924_));
 sg13g2_nand2_1 _1711_ (.Y(_0925_),
    .A(_0786_),
    .B(_0924_));
 sg13g2_a21oi_1 _1712_ (.A1(_0911_),
    .A2(_0925_),
    .Y(_0926_),
    .B1(\vga_clock.pulse_min.comp[3] ));
 sg13g2_inv_1 _1713_ (.Y(_0927_),
    .A(\vga_clock.pulse_min.comp[3] ));
 sg13g2_nand2_1 _1714_ (.Y(_0928_),
    .A(_0786_),
    .B(_0911_));
 sg13g2_nor3_1 _1715_ (.A(_0927_),
    .B(_0928_),
    .C(_0924_),
    .Y(_0929_));
 sg13g2_o21ai_1 _1716_ (.B1(net34),
    .Y(_0069_),
    .A1(_0926_),
    .A2(_0929_));
 sg13g2_o21ai_1 _1717_ (.B1(_0786_),
    .Y(_0930_),
    .A1(\vga_clock.pulse_min.comp[3] ),
    .A2(_0924_));
 sg13g2_nand2_1 _1718_ (.Y(_0931_),
    .A(\vga_clock.pulse_min.comp[4] ),
    .B(_0653_));
 sg13g2_a21oi_1 _1719_ (.A1(_0911_),
    .A2(_0930_),
    .Y(_0070_),
    .B1(_0931_));
 sg13g2_xor2_1 _1720_ (.B(_0908_),
    .A(net33),
    .X(_0932_));
 sg13g2_xor2_1 _1721_ (.B(\vga_clock.pulse_min.comp[2] ),
    .A(\vga_clock.pulse_min.count[2] ),
    .X(_0933_));
 sg13g2_xor2_1 _1722_ (.B(\vga_clock.pulse_min.count[4] ),
    .A(\vga_clock.pulse_min.comp[4] ),
    .X(_0934_));
 sg13g2_nor3_1 _1723_ (.A(_0932_),
    .B(_0933_),
    .C(_0934_),
    .Y(_0935_));
 sg13g2_xnor2_1 _1724_ (.Y(_0936_),
    .A(\vga_clock.pulse_min.count[3] ),
    .B(\vga_clock.pulse_min.comp[3] ));
 sg13g2_xnor2_1 _1725_ (.Y(_0937_),
    .A(_0789_),
    .B(_0914_));
 sg13g2_nand3_1 _1726_ (.B(_0936_),
    .C(_0937_),
    .A(_0935_),
    .Y(_0938_));
 sg13g2_and3_1 _1727_ (.X(_0939_),
    .A(_0786_),
    .B(_0822_),
    .C(_0938_));
 sg13g2_buf_1 _1728_ (.A(_0939_),
    .X(_0940_));
 sg13g2_inv_1 _1729_ (.Y(_0941_),
    .A(_0940_));
 sg13g2_nor2_1 _1730_ (.A(net33),
    .B(_0941_),
    .Y(_0942_));
 sg13g2_a21oi_1 _1731_ (.A1(_0790_),
    .A2(net14),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_nor2_1 _1732_ (.A(net23),
    .B(_0943_),
    .Y(_0071_));
 sg13g2_o21ai_1 _1733_ (.B1(_0789_),
    .Y(_0944_),
    .A1(net18),
    .A2(_0942_));
 sg13g2_nand3b_1 _1734_ (.B(net33),
    .C(_0940_),
    .Y(_0945_),
    .A_N(_0789_));
 sg13g2_a21oi_1 _1735_ (.A1(_0944_),
    .A2(_0945_),
    .Y(_0072_),
    .B1(_0832_));
 sg13g2_a21oi_1 _1736_ (.A1(_0789_),
    .A2(net33),
    .Y(_0946_),
    .B1(_0941_));
 sg13g2_o21ai_1 _1737_ (.B1(\vga_clock.pulse_min.count[2] ),
    .Y(_0159_),
    .A1(net18),
    .A2(_0946_));
 sg13g2_nand4_1 _1738_ (.B(net33),
    .C(_0788_),
    .A(_0789_),
    .Y(_0160_),
    .D(_0940_));
 sg13g2_a21oi_1 _1739_ (.A1(_0159_),
    .A2(_0160_),
    .Y(_0073_),
    .B1(net24));
 sg13g2_nand3_1 _1740_ (.B(net33),
    .C(\vga_clock.pulse_min.count[2] ),
    .A(_0789_),
    .Y(_0161_));
 sg13g2_a21oi_1 _1741_ (.A1(_0940_),
    .A2(_0161_),
    .Y(_0162_),
    .B1(net18));
 sg13g2_nand2b_1 _1742_ (.Y(_0163_),
    .B(\vga_clock.pulse_min.count[3] ),
    .A_N(_0162_));
 sg13g2_or3_1 _1743_ (.A(\vga_clock.pulse_min.count[3] ),
    .B(_0941_),
    .C(_0161_),
    .X(_0164_));
 sg13g2_a21oi_1 _1744_ (.A1(_0163_),
    .A2(_0164_),
    .Y(_0074_),
    .B1(net24));
 sg13g2_nand4_1 _1745_ (.B(net33),
    .C(\vga_clock.pulse_min.count[3] ),
    .A(_0789_),
    .Y(_0165_),
    .D(\vga_clock.pulse_min.count[2] ));
 sg13g2_xor2_1 _1746_ (.B(_0165_),
    .A(_0014_),
    .X(_0166_));
 sg13g2_a22oi_1 _1747_ (.Y(_0167_),
    .B1(_0940_),
    .B2(_0166_),
    .A2(net14),
    .A1(\vga_clock.pulse_min.count[4] ));
 sg13g2_nor2_1 _1748_ (.A(net23),
    .B(_0167_),
    .Y(_0075_));
 sg13g2_buf_1 _1749_ (.A(\vga_clock.pulse_sec.comp[0] ),
    .X(_0168_));
 sg13g2_buf_1 _1750_ (.A(ui_in[2]),
    .X(_0169_));
 sg13g2_buf_2 _1751_ (.A(\vga_clock.pulse_sec.comp[3] ),
    .X(_0170_));
 sg13g2_buf_1 _1752_ (.A(\vga_clock.pulse_sec.comp[2] ),
    .X(_0171_));
 sg13g2_nor3_1 _1753_ (.A(_0170_),
    .B(\vga_clock.pulse_sec.comp[4] ),
    .C(_0171_),
    .Y(_0172_));
 sg13g2_buf_2 _1754_ (.A(\vga_clock.pulse_sec.count[1] ),
    .X(_0173_));
 sg13g2_buf_2 _1755_ (.A(\vga_clock.pulse_sec.count[0] ),
    .X(_0174_));
 sg13g2_buf_2 _1756_ (.A(\vga_clock.pulse_sec.count[2] ),
    .X(_0175_));
 sg13g2_nor4_1 _1757_ (.A(_0173_),
    .B(_0174_),
    .C(\vga_clock.pulse_sec.count[3] ),
    .D(_0175_),
    .Y(_0176_));
 sg13g2_and2_1 _1758_ (.A(_0015_),
    .B(_0176_),
    .X(_0177_));
 sg13g2_nand2b_1 _1759_ (.Y(_0178_),
    .B(_0177_),
    .A_N(_0172_));
 sg13g2_a21oi_2 _1760_ (.B1(net18),
    .Y(_0179_),
    .A2(_0178_),
    .A1(net44));
 sg13g2_nand3_1 _1761_ (.B(_0168_),
    .C(_0179_),
    .A(net44),
    .Y(_0180_));
 sg13g2_o21ai_1 _1762_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0168_),
    .A2(_0179_));
 sg13g2_nand2_1 _1763_ (.Y(_0076_),
    .A(net32),
    .B(_0181_));
 sg13g2_buf_2 _1764_ (.A(\vga_clock.pulse_sec.comp[1] ),
    .X(_0182_));
 sg13g2_inv_1 _1765_ (.Y(_0183_),
    .A(_0168_));
 sg13g2_nand3_1 _1766_ (.B(_0182_),
    .C(_0179_),
    .A(_0183_),
    .Y(_0184_));
 sg13g2_o21ai_1 _1767_ (.B1(_0184_),
    .Y(_0185_),
    .A1(_0183_),
    .A2(_0182_));
 sg13g2_nand2_1 _1768_ (.Y(_0186_),
    .A(net44),
    .B(_0185_));
 sg13g2_o21ai_1 _1769_ (.B1(_0186_),
    .Y(_0187_),
    .A1(_0182_),
    .A2(_0179_));
 sg13g2_nand2_1 _1770_ (.Y(_0077_),
    .A(net32),
    .B(_0187_));
 sg13g2_nor3_1 _1771_ (.A(_0168_),
    .B(_0182_),
    .C(_0178_),
    .Y(_0188_));
 sg13g2_nand3_1 _1772_ (.B(net17),
    .C(_0188_),
    .A(_0171_),
    .Y(_0189_));
 sg13g2_o21ai_1 _1773_ (.B1(_0189_),
    .Y(_0190_),
    .A1(_0171_),
    .A2(_0188_));
 sg13g2_nand2_1 _1774_ (.Y(_0191_),
    .A(net44),
    .B(_0190_));
 sg13g2_o21ai_1 _1775_ (.B1(_0191_),
    .Y(_0192_),
    .A1(_0171_),
    .A2(_0864_));
 sg13g2_nand2_1 _1776_ (.Y(_0078_),
    .A(net32),
    .B(_0192_));
 sg13g2_nor3_1 _1777_ (.A(_0171_),
    .B(_0168_),
    .C(_0182_),
    .Y(_0193_));
 sg13g2_nand3_1 _1778_ (.B(_0179_),
    .C(_0193_),
    .A(_0170_),
    .Y(_0194_));
 sg13g2_o21ai_1 _1779_ (.B1(_0194_),
    .Y(_0195_),
    .A1(_0170_),
    .A2(_0193_));
 sg13g2_nand2_1 _1780_ (.Y(_0196_),
    .A(net44),
    .B(_0195_));
 sg13g2_o21ai_1 _1781_ (.B1(_0196_),
    .Y(_0197_),
    .A1(_0170_),
    .A2(_0179_));
 sg13g2_nand2_1 _1782_ (.Y(_0079_),
    .A(net32),
    .B(_0197_));
 sg13g2_inv_1 _1783_ (.Y(_0198_),
    .A(_0193_));
 sg13g2_o21ai_1 _1784_ (.B1(_0169_),
    .Y(_0199_),
    .A1(_0170_),
    .A2(_0198_));
 sg13g2_nand2_1 _1785_ (.Y(_0200_),
    .A(_0653_),
    .B(\vga_clock.pulse_sec.comp[4] ));
 sg13g2_a21oi_1 _1786_ (.A1(_0179_),
    .A2(_0199_),
    .Y(_0080_),
    .B1(_0200_));
 sg13g2_xor2_1 _1787_ (.B(_0182_),
    .A(_0173_),
    .X(_0201_));
 sg13g2_xor2_1 _1788_ (.B(_0168_),
    .A(_0174_),
    .X(_0202_));
 sg13g2_xor2_1 _1789_ (.B(\vga_clock.pulse_sec.count[4] ),
    .A(\vga_clock.pulse_sec.comp[4] ),
    .X(_0203_));
 sg13g2_nor3_1 _1790_ (.A(_0201_),
    .B(_0202_),
    .C(_0203_),
    .Y(_0204_));
 sg13g2_xnor2_1 _1791_ (.Y(_0205_),
    .A(\vga_clock.pulse_sec.count[3] ),
    .B(_0170_));
 sg13g2_xnor2_1 _1792_ (.Y(_0206_),
    .A(_0175_),
    .B(_0171_));
 sg13g2_nand3_1 _1793_ (.B(_0205_),
    .C(_0206_),
    .A(_0204_),
    .Y(_0207_));
 sg13g2_nand3_1 _1794_ (.B(net17),
    .C(_0207_),
    .A(net44),
    .Y(_0208_));
 sg13g2_nor2_1 _1795_ (.A(_0174_),
    .B(_0208_),
    .Y(_0209_));
 sg13g2_a21oi_1 _1796_ (.A1(_0174_),
    .A2(net14),
    .Y(_0210_),
    .B1(_0209_));
 sg13g2_nor2_1 _1797_ (.A(net23),
    .B(_0210_),
    .Y(_0081_));
 sg13g2_and3_1 _1798_ (.X(_0211_),
    .A(net44),
    .B(_0822_),
    .C(_0207_));
 sg13g2_buf_1 _1799_ (.A(_0211_),
    .X(_0212_));
 sg13g2_xor2_1 _1800_ (.B(_0174_),
    .A(_0173_),
    .X(_0213_));
 sg13g2_a22oi_1 _1801_ (.Y(_0214_),
    .B1(_0212_),
    .B2(_0213_),
    .A2(net14),
    .A1(_0173_));
 sg13g2_nor2_1 _1802_ (.A(net23),
    .B(_0214_),
    .Y(_0082_));
 sg13g2_nand2_1 _1803_ (.Y(_0215_),
    .A(_0173_),
    .B(_0174_));
 sg13g2_xnor2_1 _1804_ (.Y(_0216_),
    .A(_0175_),
    .B(_0215_));
 sg13g2_a22oi_1 _1805_ (.Y(_0217_),
    .B1(_0212_),
    .B2(_0216_),
    .A2(net14),
    .A1(_0175_));
 sg13g2_nor2_1 _1806_ (.A(net23),
    .B(_0217_),
    .Y(_0083_));
 sg13g2_nand3_1 _1807_ (.B(_0174_),
    .C(_0175_),
    .A(_0173_),
    .Y(_0218_));
 sg13g2_a21oi_1 _1808_ (.A1(_0212_),
    .A2(_0218_),
    .Y(_0219_),
    .B1(_0801_));
 sg13g2_nand2b_1 _1809_ (.Y(_0220_),
    .B(\vga_clock.pulse_sec.count[3] ),
    .A_N(_0219_));
 sg13g2_or3_1 _1810_ (.A(\vga_clock.pulse_sec.count[3] ),
    .B(_0208_),
    .C(_0218_),
    .X(_0221_));
 sg13g2_a21oi_1 _1811_ (.A1(_0220_),
    .A2(_0221_),
    .Y(_0084_),
    .B1(_0832_));
 sg13g2_nand4_1 _1812_ (.B(_0174_),
    .C(\vga_clock.pulse_sec.count[3] ),
    .A(_0173_),
    .Y(_0222_),
    .D(_0175_));
 sg13g2_xor2_1 _1813_ (.B(_0222_),
    .A(_0015_),
    .X(_0223_));
 sg13g2_a22oi_1 _1814_ (.Y(_0224_),
    .B1(_0212_),
    .B2(_0223_),
    .A2(net14),
    .A1(\vga_clock.pulse_sec.count[4] ));
 sg13g2_nor2_1 _1815_ (.A(_0882_),
    .B(_0224_),
    .Y(_0085_));
 sg13g2_and3_1 _1816_ (.X(_0225_),
    .A(net44),
    .B(_0822_),
    .C(_0177_));
 sg13g2_xor2_1 _1817_ (.B(_0730_),
    .A(\vga_clock.sec_u[0] ),
    .X(_0226_));
 sg13g2_nor2_1 _1818_ (.A(_0225_),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_nor2b_1 _1819_ (.A(_0009_),
    .B_N(_0225_),
    .Y(_0228_));
 sg13g2_nor3_1 _1820_ (.A(net24),
    .B(_0227_),
    .C(_0228_),
    .Y(_0115_));
 sg13g2_nand2_1 _1821_ (.Y(_0229_),
    .A(\vga_clock.sec_u[1] ),
    .B(_0774_));
 sg13g2_xnor2_1 _1822_ (.Y(_0230_),
    .A(\vga_clock.sec_u[1] ),
    .B(\vga_clock.sec_u[0] ));
 sg13g2_or2_1 _1823_ (.X(_0231_),
    .B(_0225_),
    .A(_0730_));
 sg13g2_mux2_1 _1824_ (.A0(_0229_),
    .A1(_0230_),
    .S(_0231_),
    .X(_0232_));
 sg13g2_nor2_1 _1825_ (.A(net23),
    .B(_0232_),
    .Y(_0116_));
 sg13g2_and2_1 _1826_ (.A(\vga_clock.sec_u[1] ),
    .B(\vga_clock.sec_u[0] ),
    .X(_0233_));
 sg13g2_o21ai_1 _1827_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_0730_),
    .A2(_0225_));
 sg13g2_xnor2_1 _1828_ (.Y(_0235_),
    .A(\vga_clock.sec_u[2] ),
    .B(_0234_));
 sg13g2_and2_1 _1829_ (.A(net34),
    .B(_0235_),
    .X(_0117_));
 sg13g2_buf_1 _1830_ (.A(_0659_),
    .X(_0236_));
 sg13g2_nand2_1 _1831_ (.Y(_0237_),
    .A(\vga_clock.sec_u[3] ),
    .B(_0774_));
 sg13g2_nand2_1 _1832_ (.Y(_0238_),
    .A(\vga_clock.sec_u[2] ),
    .B(_0233_));
 sg13g2_xnor2_1 _1833_ (.Y(_0239_),
    .A(_0022_),
    .B(_0238_));
 sg13g2_mux2_1 _1834_ (.A0(_0237_),
    .A1(_0239_),
    .S(_0231_),
    .X(_0240_));
 sg13g2_nor2_1 _1835_ (.A(_0236_),
    .B(_0240_),
    .Y(_0118_));
 sg13g2_buf_1 _1836_ (.A(\vga_clock.vga_0.hc[8] ),
    .X(_0241_));
 sg13g2_buf_1 _1837_ (.A(\vga_clock.vga_0.hc[9] ),
    .X(_0242_));
 sg13g2_buf_2 _1838_ (.A(\vga_clock.vga_0.hc[7] ),
    .X(_0243_));
 sg13g2_buf_2 _1839_ (.A(\vga_clock.vga_0.hc[6] ),
    .X(_0244_));
 sg13g2_nand3_1 _1840_ (.B(\vga_clock.vga_0.hc[1] ),
    .C(\vga_clock.vga_0.hc[0] ),
    .A(\vga_clock.vga_0.hc[2] ),
    .Y(_0245_));
 sg13g2_nand2_1 _1841_ (.Y(_0246_),
    .A(\vga_clock.vga_0.hc[3] ),
    .B(\vga_clock.vga_0.hc[4] ));
 sg13g2_nor2_1 _1842_ (.A(_0245_),
    .B(_0246_),
    .Y(_0247_));
 sg13g2_and2_1 _1843_ (.A(\vga_clock.vga_0.hc[5] ),
    .B(_0247_),
    .X(_0248_));
 sg13g2_buf_1 _1844_ (.A(_0248_),
    .X(_0249_));
 sg13g2_or3_1 _1845_ (.A(_0243_),
    .B(_0244_),
    .C(_0249_),
    .X(_0250_));
 sg13g2_and3_1 _1846_ (.X(_0251_),
    .A(_0241_),
    .B(_0242_),
    .C(_0250_));
 sg13g2_buf_2 _1847_ (.A(_0251_),
    .X(_0252_));
 sg13g2_nor2_2 _1848_ (.A(_0659_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_and2_1 _1849_ (.A(_0025_),
    .B(_0253_),
    .X(_0119_));
 sg13g2_nand2b_1 _1850_ (.Y(_0254_),
    .B(net46),
    .A_N(_0252_));
 sg13g2_buf_1 _1851_ (.A(_0254_),
    .X(_0255_));
 sg13g2_xnor2_1 _1852_ (.Y(_0256_),
    .A(\vga_clock.vga_0.hc[1] ),
    .B(\vga_clock.vga_0.hc[0] ));
 sg13g2_nor2_1 _1853_ (.A(net11),
    .B(_0256_),
    .Y(_0120_));
 sg13g2_nand2_1 _1854_ (.Y(_0257_),
    .A(\vga_clock.vga_0.hc[1] ),
    .B(\vga_clock.vga_0.hc[0] ));
 sg13g2_xor2_1 _1855_ (.B(_0257_),
    .A(\vga_clock.vga_0.hc[2] ),
    .X(_0258_));
 sg13g2_nor2_1 _1856_ (.A(net11),
    .B(_0258_),
    .Y(_0121_));
 sg13g2_xor2_1 _1857_ (.B(_0245_),
    .A(\vga_clock.vga_0.hc[3] ),
    .X(_0259_));
 sg13g2_nor2_1 _1858_ (.A(_0255_),
    .B(_0259_),
    .Y(_0122_));
 sg13g2_nand4_1 _1859_ (.B(\vga_clock.vga_0.hc[2] ),
    .C(\vga_clock.vga_0.hc[1] ),
    .A(\vga_clock.vga_0.hc[3] ),
    .Y(_0260_),
    .D(\vga_clock.vga_0.hc[0] ));
 sg13g2_xor2_1 _1860_ (.B(_0260_),
    .A(\vga_clock.vga_0.hc[4] ),
    .X(_0261_));
 sg13g2_nor2_1 _1861_ (.A(_0255_),
    .B(_0261_),
    .Y(_0123_));
 sg13g2_xnor2_1 _1862_ (.Y(_0262_),
    .A(\vga_clock.vga_0.hc[5] ),
    .B(_0247_));
 sg13g2_nor2_1 _1863_ (.A(net11),
    .B(_0262_),
    .Y(_0124_));
 sg13g2_xnor2_1 _1864_ (.Y(_0263_),
    .A(_0244_),
    .B(_0249_));
 sg13g2_nor2_1 _1865_ (.A(net11),
    .B(_0263_),
    .Y(_0125_));
 sg13g2_nand2_1 _1866_ (.Y(_0264_),
    .A(_0244_),
    .B(_0249_));
 sg13g2_xor2_1 _1867_ (.B(_0264_),
    .A(_0243_),
    .X(_0265_));
 sg13g2_nor2_1 _1868_ (.A(net11),
    .B(_0265_),
    .Y(_0126_));
 sg13g2_inv_1 _1869_ (.Y(_0266_),
    .A(_0241_));
 sg13g2_nand3_1 _1870_ (.B(_0244_),
    .C(_0249_),
    .A(_0243_),
    .Y(_0267_));
 sg13g2_xnor2_1 _1871_ (.Y(_0268_),
    .A(_0266_),
    .B(_0267_));
 sg13g2_nor2_1 _1872_ (.A(net11),
    .B(_0268_),
    .Y(_0127_));
 sg13g2_nand2_1 _1873_ (.Y(_0269_),
    .A(_0241_),
    .B(_0250_));
 sg13g2_nand2_2 _1874_ (.Y(_0270_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_nor3_1 _1875_ (.A(_0266_),
    .B(_0242_),
    .C(_0270_),
    .Y(_0271_));
 sg13g2_a22oi_1 _1876_ (.Y(_0272_),
    .B1(_0271_),
    .B2(_0249_),
    .A2(_0269_),
    .A1(_0242_));
 sg13g2_nor2_1 _1877_ (.A(net22),
    .B(_0272_),
    .Y(_0128_));
 sg13g2_inv_1 _1878_ (.Y(_0273_),
    .A(\vga_clock.vga_0.vc[5] ));
 sg13g2_buf_1 _1879_ (.A(\vga_clock.vga_0.vc[2] ),
    .X(_0274_));
 sg13g2_buf_1 _1880_ (.A(\vga_clock.vga_0.vc[1] ),
    .X(_0275_));
 sg13g2_buf_2 _1881_ (.A(\vga_clock.vga_0.vc[0] ),
    .X(_0276_));
 sg13g2_nand3_1 _1882_ (.B(_0275_),
    .C(_0276_),
    .A(_0274_),
    .Y(_0277_));
 sg13g2_buf_1 _1883_ (.A(\vga_clock.vga_0.vc[4] ),
    .X(_0278_));
 sg13g2_nor2_1 _1884_ (.A(\vga_clock.vga_0.vc[3] ),
    .B(net31),
    .Y(_0279_));
 sg13g2_buf_1 _1885_ (.A(\vga_clock.vga_0.vc[7] ),
    .X(_0280_));
 sg13g2_buf_1 _1886_ (.A(\vga_clock.vga_0.vc[6] ),
    .X(_0281_));
 sg13g2_nor3_1 _1887_ (.A(_0280_),
    .B(_0281_),
    .C(\vga_clock.vga_0.vc[8] ),
    .Y(_0282_));
 sg13g2_nand4_1 _1888_ (.B(_0277_),
    .C(_0279_),
    .A(_0273_),
    .Y(_0283_),
    .D(_0282_));
 sg13g2_a21oi_2 _1889_ (.B1(_0659_),
    .Y(_0284_),
    .A2(_0283_),
    .A1(\vga_clock.vga_0.vc[9] ));
 sg13g2_nor2_1 _1890_ (.A(_0253_),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_xnor2_1 _1891_ (.Y(_0286_),
    .A(_0276_),
    .B(_0252_));
 sg13g2_nor2_1 _1892_ (.A(_0285_),
    .B(_0286_),
    .Y(_0129_));
 sg13g2_and2_1 _1893_ (.A(_0252_),
    .B(_0284_),
    .X(_0287_));
 sg13g2_nand2_1 _1894_ (.Y(_0288_),
    .A(_0276_),
    .B(_0287_));
 sg13g2_inv_1 _1895_ (.Y(_0289_),
    .A(_0284_));
 sg13g2_nor2_1 _1896_ (.A(_0276_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_o21ai_1 _1897_ (.B1(_0275_),
    .Y(_0291_),
    .A1(_0253_),
    .A2(_0290_));
 sg13g2_o21ai_1 _1898_ (.B1(_0291_),
    .Y(_0130_),
    .A1(_0275_),
    .A2(_0288_));
 sg13g2_nand3_1 _1899_ (.B(_0276_),
    .C(_0287_),
    .A(_0275_),
    .Y(_0292_));
 sg13g2_a21oi_1 _1900_ (.A1(_0275_),
    .A2(_0276_),
    .Y(_0293_),
    .B1(_0289_));
 sg13g2_o21ai_1 _1901_ (.B1(_0274_),
    .Y(_0294_),
    .A1(_0253_),
    .A2(_0293_));
 sg13g2_o21ai_1 _1902_ (.B1(_0294_),
    .Y(_0131_),
    .A1(_0274_),
    .A2(_0292_));
 sg13g2_inv_1 _1903_ (.Y(_0295_),
    .A(_0024_));
 sg13g2_xnor2_1 _1904_ (.Y(_0296_),
    .A(_0295_),
    .B(_0277_));
 sg13g2_nand2_1 _1905_ (.Y(_0297_),
    .A(_0284_),
    .B(_0296_));
 sg13g2_nor2_1 _1906_ (.A(\vga_clock.vga_0.vc[3] ),
    .B(_0252_),
    .Y(_0298_));
 sg13g2_a21oi_1 _1907_ (.A1(net11),
    .A2(_0297_),
    .Y(_0132_),
    .B1(_0298_));
 sg13g2_inv_1 _1908_ (.Y(_0299_),
    .A(\vga_clock.vga_0.vc[3] ));
 sg13g2_nor2_1 _1909_ (.A(_0299_),
    .B(_0277_),
    .Y(_0300_));
 sg13g2_nand2_1 _1910_ (.Y(_0301_),
    .A(_0287_),
    .B(_0300_));
 sg13g2_nor2_1 _1911_ (.A(_0289_),
    .B(_0300_),
    .Y(_0302_));
 sg13g2_o21ai_1 _1912_ (.B1(net31),
    .Y(_0303_),
    .A1(_0253_),
    .A2(_0302_));
 sg13g2_o21ai_1 _1913_ (.B1(_0303_),
    .Y(_0133_),
    .A1(net31),
    .A2(_0301_));
 sg13g2_nand2_1 _1914_ (.Y(_0304_),
    .A(net31),
    .B(_0300_));
 sg13g2_xor2_1 _1915_ (.B(_0304_),
    .A(_0023_),
    .X(_0305_));
 sg13g2_nand2_1 _1916_ (.Y(_0306_),
    .A(_0284_),
    .B(_0305_));
 sg13g2_nor2_1 _1917_ (.A(\vga_clock.vga_0.vc[5] ),
    .B(_0252_),
    .Y(_0307_));
 sg13g2_a21oi_1 _1918_ (.A1(net11),
    .A2(_0306_),
    .Y(_0134_),
    .B1(_0307_));
 sg13g2_nand3_1 _1919_ (.B(\vga_clock.vga_0.vc[5] ),
    .C(_0300_),
    .A(net31),
    .Y(_0308_));
 sg13g2_xor2_1 _1920_ (.B(_0308_),
    .A(_0008_),
    .X(_0309_));
 sg13g2_nand2_1 _1921_ (.Y(_0310_),
    .A(_0284_),
    .B(_0309_));
 sg13g2_nor2_1 _1922_ (.A(_0281_),
    .B(_0252_),
    .Y(_0311_));
 sg13g2_a21oi_1 _1923_ (.A1(_0254_),
    .A2(_0310_),
    .Y(_0135_),
    .B1(_0311_));
 sg13g2_inv_1 _1924_ (.Y(_0312_),
    .A(_0308_));
 sg13g2_and3_1 _1925_ (.X(_0313_),
    .A(_0281_),
    .B(_0252_),
    .C(_0312_));
 sg13g2_xnor2_1 _1926_ (.Y(_0314_),
    .A(_0280_),
    .B(_0313_));
 sg13g2_nor2_1 _1927_ (.A(_0285_),
    .B(_0314_),
    .Y(_0136_));
 sg13g2_and2_1 _1928_ (.A(_0280_),
    .B(_0313_),
    .X(_0315_));
 sg13g2_xnor2_1 _1929_ (.Y(_0316_),
    .A(\vga_clock.vga_0.vc[8] ),
    .B(_0315_));
 sg13g2_nor2_1 _1930_ (.A(_0285_),
    .B(_0316_),
    .Y(_0137_));
 sg13g2_a21oi_1 _1931_ (.A1(\vga_clock.vga_0.vc[8] ),
    .A2(_0315_),
    .Y(_0317_),
    .B1(\vga_clock.vga_0.vc[9] ));
 sg13g2_nor2_1 _1932_ (.A(_0285_),
    .B(_0317_),
    .Y(_0138_));
 sg13g2_and2_1 _1933_ (.A(\vga_clock.vga_0.hc[0] ),
    .B(net35),
    .X(_0139_));
 sg13g2_and2_1 _1934_ (.A(\vga_clock.vga_0.hc[1] ),
    .B(net35),
    .X(_0140_));
 sg13g2_and2_1 _1935_ (.A(\vga_clock.vga_0.hc[2] ),
    .B(net35),
    .X(_0141_));
 sg13g2_and2_1 _1936_ (.A(\vga_clock.vga_0.hc[3] ),
    .B(net35),
    .X(_0142_));
 sg13g2_and2_1 _1937_ (.A(\vga_clock.vga_0.hc[4] ),
    .B(net35),
    .X(_0143_));
 sg13g2_and2_1 _1938_ (.A(\vga_clock.vga_0.hc[5] ),
    .B(net35),
    .X(_0144_));
 sg13g2_and2_1 _1939_ (.A(net34),
    .B(_0026_),
    .X(_0145_));
 sg13g2_xnor2_1 _1940_ (.Y(_0318_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_nor2_1 _1941_ (.A(net22),
    .B(_0318_),
    .Y(_0146_));
 sg13g2_xor2_1 _1942_ (.B(_0270_),
    .A(_0012_),
    .X(_0319_));
 sg13g2_nor2_1 _1943_ (.A(net22),
    .B(_0319_),
    .Y(_0147_));
 sg13g2_o21ai_1 _1944_ (.B1(_0012_),
    .Y(_0320_),
    .A1(_0241_),
    .A2(_0270_));
 sg13g2_xor2_1 _1945_ (.B(_0320_),
    .A(_0242_),
    .X(_0321_));
 sg13g2_nor2_1 _1946_ (.A(net22),
    .B(_0321_),
    .Y(_0148_));
 sg13g2_and2_1 _1947_ (.A(net34),
    .B(_0276_),
    .X(_0149_));
 sg13g2_and2_1 _1948_ (.A(_0750_),
    .B(_0275_),
    .X(_0150_));
 sg13g2_and2_1 _1949_ (.A(_0750_),
    .B(_0274_),
    .X(_0151_));
 sg13g2_nor2_1 _1950_ (.A(net22),
    .B(_0295_),
    .Y(_0152_));
 sg13g2_xor2_1 _1951_ (.B(net31),
    .A(\vga_clock.vga_0.vc[3] ),
    .X(_0322_));
 sg13g2_nor2_1 _1952_ (.A(net22),
    .B(_0322_),
    .Y(_0153_));
 sg13g2_xnor2_1 _1953_ (.Y(_0323_),
    .A(_0023_),
    .B(_0279_));
 sg13g2_nor2_1 _1954_ (.A(net22),
    .B(_0323_),
    .Y(_0154_));
 sg13g2_o21ai_1 _1955_ (.B1(\vga_clock.vga_0.vc[5] ),
    .Y(_0324_),
    .A1(\vga_clock.vga_0.vc[3] ),
    .A2(net31));
 sg13g2_xnor2_1 _1956_ (.Y(_0325_),
    .A(_0281_),
    .B(_0324_));
 sg13g2_nor2_1 _1957_ (.A(net22),
    .B(_0325_),
    .Y(_0155_));
 sg13g2_o21ai_1 _1958_ (.B1(_0008_),
    .Y(_0326_),
    .A1(_0281_),
    .A2(_0324_));
 sg13g2_xor2_1 _1959_ (.B(_0326_),
    .A(_0280_),
    .X(_0327_));
 sg13g2_nor2_1 _1960_ (.A(_0236_),
    .B(_0327_),
    .Y(_0156_));
 sg13g2_nor2_1 _1961_ (.A(_0280_),
    .B(_0281_),
    .Y(_0328_));
 sg13g2_nand2_1 _1962_ (.Y(_0329_),
    .A(_0328_),
    .B(_0324_));
 sg13g2_nand2_1 _1963_ (.Y(_0330_),
    .A(\vga_clock.vga_0.vc[8] ),
    .B(_0329_));
 sg13g2_nand2_1 _1964_ (.Y(_0331_),
    .A(_0282_),
    .B(_0324_));
 sg13g2_a21oi_1 _1965_ (.A1(_0330_),
    .A2(_0331_),
    .Y(_0157_),
    .B1(net24));
 sg13g2_xor2_1 _1966_ (.B(_0331_),
    .A(\vga_clock.vga_0.vc[9] ),
    .X(_0332_));
 sg13g2_nor2_1 _1967_ (.A(net24),
    .B(_0332_),
    .Y(_0158_));
 sg13g2_buf_1 _1968_ (.A(ui_in[3]),
    .X(_0333_));
 sg13g2_buf_1 _1969_ (.A(_0333_),
    .X(_0334_));
 sg13g2_or2_1 _1970_ (.X(_0335_),
    .B(_0276_),
    .A(_0275_));
 sg13g2_nor3_1 _1971_ (.A(_0274_),
    .B(_0299_),
    .C(_0335_),
    .Y(_0336_));
 sg13g2_nor3_1 _1972_ (.A(net31),
    .B(_0295_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_nor2b_1 _1973_ (.A(\vga_clock.vga_0.vc[9] ),
    .B_N(_0282_),
    .Y(_0338_));
 sg13g2_o21ai_1 _1974_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0273_),
    .A2(_0337_));
 sg13g2_nor2_1 _1975_ (.A(_0241_),
    .B(_0242_),
    .Y(_0340_));
 sg13g2_nand2_1 _1976_ (.Y(_0341_),
    .A(_0270_),
    .B(_0340_));
 sg13g2_nand3_1 _1977_ (.B(_0339_),
    .C(_0341_),
    .A(\vga_clock.draw ),
    .Y(_0342_));
 sg13g2_buf_1 _1978_ (.A(_0342_),
    .X(_0343_));
 sg13g2_inv_1 _1979_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_nand2_1 _1980_ (.Y(_0345_),
    .A(\vga_clock.color[5] ),
    .B(_0344_));
 sg13g2_a21oi_1 _1981_ (.A1(\vga_clock.vga_0.hc[3] ),
    .A2(\vga_clock.vga_0.hc[4] ),
    .Y(_0346_),
    .B1(\vga_clock.vga_0.hc[5] ));
 sg13g2_nor4_1 _1982_ (.A(_0241_),
    .B(_0242_),
    .C(_0243_),
    .D(_0244_),
    .Y(_0347_));
 sg13g2_nand2b_1 _1983_ (.Y(_0348_),
    .B(_0347_),
    .A_N(_0346_));
 sg13g2_nand2_1 _1984_ (.Y(_0349_),
    .A(net30),
    .B(_0348_));
 sg13g2_o21ai_1 _1985_ (.B1(_0349_),
    .Y(net1),
    .A1(net30),
    .A2(_0345_));
 sg13g2_nand2_1 _1986_ (.Y(_0350_),
    .A(\vga_clock.color[3] ),
    .B(_0344_));
 sg13g2_nor4_1 _1987_ (.A(_0274_),
    .B(_0299_),
    .C(_0278_),
    .D(\vga_clock.vga_0.vc[5] ),
    .Y(_0351_));
 sg13g2_nand3_1 _1988_ (.B(_0335_),
    .C(_0351_),
    .A(_0338_),
    .Y(_0352_));
 sg13g2_nand2_1 _1989_ (.Y(_0353_),
    .A(net30),
    .B(_0352_));
 sg13g2_o21ai_1 _1990_ (.B1(_0353_),
    .Y(net2),
    .A1(net30),
    .A2(_0350_));
 sg13g2_nor2b_1 _1991_ (.A(_0333_),
    .B_N(\vga_clock.color[1] ),
    .Y(_0354_));
 sg13g2_a21oi_1 _1992_ (.A1(\vga_clock.color[0] ),
    .A2(_0334_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_nor2_1 _1993_ (.A(_0343_),
    .B(_0355_),
    .Y(net3));
 sg13g2_nand2_1 _1994_ (.Y(_0356_),
    .A(\vga_clock.color[1] ),
    .B(_0344_));
 sg13g2_nor2_1 _1995_ (.A(net30),
    .B(_0352_),
    .Y(_0357_));
 sg13g2_a21oi_1 _1996_ (.A1(_0334_),
    .A2(_0356_),
    .Y(net4),
    .B1(_0357_));
 sg13g2_nor2b_1 _1997_ (.A(_0333_),
    .B_N(\vga_clock.color[4] ),
    .Y(_0358_));
 sg13g2_a21oi_1 _1998_ (.A1(\vga_clock.color[2] ),
    .A2(net30),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_nor2_1 _1999_ (.A(_0343_),
    .B(_0359_),
    .Y(net5));
 sg13g2_nor2b_1 _2000_ (.A(_0333_),
    .B_N(\vga_clock.color[2] ),
    .Y(_0360_));
 sg13g2_a21oi_1 _2001_ (.A1(\vga_clock.color[3] ),
    .A2(_0333_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_nor2_1 _2002_ (.A(_0343_),
    .B(_0361_),
    .Y(net6));
 sg13g2_nor2b_1 _2003_ (.A(_0333_),
    .B_N(\vga_clock.color[0] ),
    .Y(_0362_));
 sg13g2_a21oi_1 _2004_ (.A1(\vga_clock.color[4] ),
    .A2(_0333_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nor2_1 _2005_ (.A(_0343_),
    .B(_0363_),
    .Y(net7));
 sg13g2_nor2_1 _2006_ (.A(net30),
    .B(_0348_),
    .Y(_0364_));
 sg13g2_a21oi_1 _2007_ (.A1(net30),
    .A2(_0345_),
    .Y(net8),
    .B1(_0364_));
 sg13g2_inv_1 _2008_ (.Y(\vga_clock.y_block[1] ),
    .A(_0451_));
 sg13g2_xnor2_1 _2009_ (.Y(\vga_clock.y_block[3] ),
    .A(net37),
    .B(_0419_));
 sg13g2_xor2_1 _2010_ (.B(_0441_),
    .A(_0421_),
    .X(\vga_clock.y_block[4] ));
 sg13g2_inv_1 _2011_ (.Y(\vga_clock.y_block[5] ),
    .A(_0447_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \vga_clock.col_index_q[0]$_DFF_P__63  (.L_HI(net63));
 sg13g2_buf_1 _2014_ (.A(net47),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2015_ (.A(net48),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2016_ (.A(net49),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2017_ (.A(net50),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2018_ (.A(net51),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2019_ (.A(net52),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2020_ (.A(net53),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2021_ (.A(net54),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2022_ (.A(net55),
    .X(uio_out[0]));
 sg13g2_buf_1 _2023_ (.A(net56),
    .X(uio_out[1]));
 sg13g2_buf_1 _2024_ (.A(net57),
    .X(uio_out[2]));
 sg13g2_buf_1 _2025_ (.A(net58),
    .X(uio_out[3]));
 sg13g2_buf_1 _2026_ (.A(net59),
    .X(uio_out[4]));
 sg13g2_buf_1 _2027_ (.A(net60),
    .X(uio_out[5]));
 sg13g2_buf_1 _2028_ (.A(net61),
    .X(uio_out[6]));
 sg13g2_buf_1 _2029_ (.A(net62),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \vga_clock.col_index_q[0]$_DFF_P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net63),
    .D(\vga_clock.col_index[0] ),
    .Q_N(_1050_),
    .Q(\vga_clock.col_index_q[0] ));
 sg13g2_dfrbp_1 \vga_clock.col_index_q[1]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net64),
    .D(\vga_clock.col_index[1] ),
    .Q_N(_1049_),
    .Q(\vga_clock.col_index_q[1] ));
 sg13g2_dfrbp_1 \vga_clock.color_offset[0]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net65),
    .D(_0032_),
    .Q_N(_0028_),
    .Q(\vga_clock.color_offset[0] ));
 sg13g2_dfrbp_1 \vga_clock.color_offset[1]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net66),
    .D(_0033_),
    .Q_N(_1048_),
    .Q(\vga_clock.color_offset[1] ));
 sg13g2_dfrbp_1 \vga_clock.color_offset[2]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net67),
    .D(_0034_),
    .Q_N(_1047_),
    .Q(\vga_clock.color_offset[2] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.col_index[0]$_SDFF_PP1_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net68),
    .D(_0035_),
    .Q_N(_1046_),
    .Q(\vga_clock.col_index[0] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.col_index[1]$_SDFF_PP1_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net69),
    .D(_0036_),
    .Q_N(_1045_),
    .Q(\vga_clock.col_index[1] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[0]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net70),
    .D(_0037_),
    .Q_N(_1044_),
    .Q(\vga_clock.color[0] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[1]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net71),
    .D(_0038_),
    .Q_N(_1043_),
    .Q(\vga_clock.color[1] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[2]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net72),
    .D(_0039_),
    .Q_N(_1042_),
    .Q(\vga_clock.color[2] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[3]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net73),
    .D(_0040_),
    .Q_N(_1051_),
    .Q(\vga_clock.color[3] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[4]$_DFF_P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net74),
    .D(_0000_),
    .Q_N(_1052_),
    .Q(\vga_clock.color[4] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.color[5]$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net75),
    .D(_0001_),
    .Q_N(_1053_),
    .Q(\vga_clock.color[5] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[0]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net76),
    .D(\vga_clock.digit_0.number[0] ),
    .Q_N(_1054_),
    .Q(\vga_clock.digit_0.digit_index[0] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[1]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net77),
    .D(\vga_clock.digit_0.number[1] ),
    .Q_N(_1055_),
    .Q(\vga_clock.digit_0.digit_index[1] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[2]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net78),
    .D(_0002_),
    .Q_N(_1056_),
    .Q(\vga_clock.digit_0.digit_index[2] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[3]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net79),
    .D(_0003_),
    .Q_N(_1057_),
    .Q(\vga_clock.digit_0.digit_index[3] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[4]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net80),
    .D(_0004_),
    .Q_N(_1041_),
    .Q(\vga_clock.digit_0.digit_index[4] ));
 sg13g2_dfrbp_1 \vga_clock.digit_0.digit_index[5]$_SDFF_PP1_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net81),
    .D(_0041_),
    .Q_N(_1040_),
    .Q(\vga_clock.digit_0.digit_index[5] ));
 sg13g2_dfrbp_1 \vga_clock.draw$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net82),
    .D(_0042_),
    .Q_N(_1058_),
    .Q(\vga_clock.draw ));
 sg13g2_dfrbp_1 \vga_clock.font_0.dout[1]$_DFF_P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net83),
    .D(_0005_),
    .Q_N(_1059_),
    .Q(\vga_clock.font_0.dout[1] ));
 sg13g2_dfrbp_1 \vga_clock.font_0.dout[2]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net84),
    .D(_0006_),
    .Q_N(_1060_),
    .Q(\vga_clock.font_0.dout[2] ));
 sg13g2_dfrbp_1 \vga_clock.font_0.dout[3]$_DFF_P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net85),
    .D(_0007_),
    .Q_N(_1039_),
    .Q(\vga_clock.font_0.dout[3] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_d[0]$_SDFFE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net86),
    .D(_0043_),
    .Q_N(_0030_),
    .Q(\vga_clock.hrs_d[0] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_d[1]$_SDFFE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net87),
    .D(_0044_),
    .Q_N(_0017_),
    .Q(\vga_clock.hrs_d[1] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_u[0]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net88),
    .D(_0045_),
    .Q_N(_0011_),
    .Q(\vga_clock.hrs_u[0] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_u[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net89),
    .D(_0046_),
    .Q_N(_0018_),
    .Q(\vga_clock.hrs_u[1] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_u[2]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net90),
    .D(_0047_),
    .Q_N(_0019_),
    .Q(\vga_clock.hrs_u[2] ));
 sg13g2_dfrbp_1 \vga_clock.hrs_u[3]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net91),
    .D(_0048_),
    .Q_N(_0020_),
    .Q(\vga_clock.hrs_u[3] ));
 sg13g2_dfrbp_1 \vga_clock.min_d[0]$_SDFFE_PP0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net92),
    .D(_0049_),
    .Q_N(_0029_),
    .Q(\vga_clock.min_d[0] ));
 sg13g2_dfrbp_1 \vga_clock.min_d[1]$_SDFFE_PP0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net93),
    .D(_0050_),
    .Q_N(_1038_),
    .Q(\vga_clock.min_d[1] ));
 sg13g2_dfrbp_1 \vga_clock.min_d[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net94),
    .D(_0051_),
    .Q_N(_1037_),
    .Q(\vga_clock.min_d[2] ));
 sg13g2_dfrbp_1 \vga_clock.min_u[0]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net95),
    .D(_0052_),
    .Q_N(_0010_),
    .Q(\vga_clock.min_u[0] ));
 sg13g2_dfrbp_1 \vga_clock.min_u[1]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net96),
    .D(_0053_),
    .Q_N(_1036_),
    .Q(\vga_clock.min_u[1] ));
 sg13g2_dfrbp_1 \vga_clock.min_u[2]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net97),
    .D(_0054_),
    .Q_N(_1035_),
    .Q(\vga_clock.min_u[2] ));
 sg13g2_dfrbp_1 \vga_clock.min_u[3]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net98),
    .D(_0055_),
    .Q_N(_0021_),
    .Q(\vga_clock.min_u[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.comp[0]$_SDFFE_PN1P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net99),
    .D(_0056_),
    .Q_N(_1034_),
    .Q(\vga_clock.pulse_hrs.comp[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.comp[1]$_SDFFE_PN1P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net100),
    .D(_0057_),
    .Q_N(_1033_),
    .Q(\vga_clock.pulse_hrs.comp[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.comp[2]$_SDFFE_PN1P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net101),
    .D(_0058_),
    .Q_N(_1032_),
    .Q(\vga_clock.pulse_hrs.comp[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.comp[3]$_SDFFE_PN1P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net102),
    .D(_0059_),
    .Q_N(_1031_),
    .Q(\vga_clock.pulse_hrs.comp[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.comp[4]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net103),
    .D(_0060_),
    .Q_N(_1030_),
    .Q(\vga_clock.pulse_hrs.comp[4] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.count[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net104),
    .D(_0061_),
    .Q_N(_1029_),
    .Q(\vga_clock.pulse_hrs.count[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.count[1]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net105),
    .D(_0062_),
    .Q_N(_1028_),
    .Q(\vga_clock.pulse_hrs.count[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.count[2]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net106),
    .D(_0063_),
    .Q_N(_1027_),
    .Q(\vga_clock.pulse_hrs.count[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.count[3]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net107),
    .D(_0064_),
    .Q_N(_1026_),
    .Q(\vga_clock.pulse_hrs.count[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_hrs.count[4]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net108),
    .D(_0065_),
    .Q_N(_0013_),
    .Q(\vga_clock.pulse_hrs.count[4] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.comp[0]$_SDFFE_PN1P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net109),
    .D(_0066_),
    .Q_N(_1025_),
    .Q(\vga_clock.pulse_min.comp[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.comp[1]$_SDFFE_PN1P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net110),
    .D(_0067_),
    .Q_N(_1024_),
    .Q(\vga_clock.pulse_min.comp[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.comp[2]$_SDFFE_PN1P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net111),
    .D(_0068_),
    .Q_N(_1023_),
    .Q(\vga_clock.pulse_min.comp[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.comp[3]$_SDFFE_PN1P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net112),
    .D(_0069_),
    .Q_N(_1022_),
    .Q(\vga_clock.pulse_min.comp[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.comp[4]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net113),
    .D(_0070_),
    .Q_N(_1021_),
    .Q(\vga_clock.pulse_min.comp[4] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.count[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net114),
    .D(_0071_),
    .Q_N(_1020_),
    .Q(\vga_clock.pulse_min.count[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.count[1]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net115),
    .D(_0072_),
    .Q_N(_1019_),
    .Q(\vga_clock.pulse_min.count[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.count[2]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net116),
    .D(_0073_),
    .Q_N(_1018_),
    .Q(\vga_clock.pulse_min.count[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.count[3]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net117),
    .D(_0074_),
    .Q_N(_1017_),
    .Q(\vga_clock.pulse_min.count[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_min.count[4]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net118),
    .D(_0075_),
    .Q_N(_0014_),
    .Q(\vga_clock.pulse_min.count[4] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.comp[0]$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net119),
    .D(_0076_),
    .Q_N(_1016_),
    .Q(\vga_clock.pulse_sec.comp[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.comp[1]$_SDFFE_PN1P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net120),
    .D(_0077_),
    .Q_N(_1015_),
    .Q(\vga_clock.pulse_sec.comp[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.comp[2]$_SDFFE_PN1P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net121),
    .D(_0078_),
    .Q_N(_1014_),
    .Q(\vga_clock.pulse_sec.comp[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.comp[3]$_SDFFE_PN1P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net122),
    .D(_0079_),
    .Q_N(_1013_),
    .Q(\vga_clock.pulse_sec.comp[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.comp[4]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net123),
    .D(_0080_),
    .Q_N(_1012_),
    .Q(\vga_clock.pulse_sec.comp[4] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.count[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net124),
    .D(_0081_),
    .Q_N(_1011_),
    .Q(\vga_clock.pulse_sec.count[0] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.count[1]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net125),
    .D(_0082_),
    .Q_N(_1010_),
    .Q(\vga_clock.pulse_sec.count[1] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.count[2]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net126),
    .D(_0083_),
    .Q_N(_1009_),
    .Q(\vga_clock.pulse_sec.count[2] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.count[3]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net127),
    .D(_0084_),
    .Q_N(_1008_),
    .Q(\vga_clock.pulse_sec.count[3] ));
 sg13g2_dfrbp_1 \vga_clock.pulse_sec.count[4]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net128),
    .D(_0085_),
    .Q_N(_0015_),
    .Q(\vga_clock.pulse_sec.count[4] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[0]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net129),
    .D(_0086_),
    .Q_N(_0031_),
    .Q(\vga_clock.sec_counter[0] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[10]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0087_),
    .Q_N(_1007_),
    .Q(\vga_clock.sec_counter[10] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[11]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net131),
    .D(_0088_),
    .Q_N(_1006_),
    .Q(\vga_clock.sec_counter[11] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[12]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net132),
    .D(_0089_),
    .Q_N(_1005_),
    .Q(\vga_clock.sec_counter[12] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[13]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net133),
    .D(_0090_),
    .Q_N(_1004_),
    .Q(\vga_clock.sec_counter[13] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[14]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net134),
    .D(_0091_),
    .Q_N(_1003_),
    .Q(\vga_clock.sec_counter[14] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[15]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net135),
    .D(_0092_),
    .Q_N(_1002_),
    .Q(\vga_clock.sec_counter[15] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[16]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net136),
    .D(_0093_),
    .Q_N(_1001_),
    .Q(\vga_clock.sec_counter[16] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[17]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net137),
    .D(_0094_),
    .Q_N(_1000_),
    .Q(\vga_clock.sec_counter[17] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[18]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net138),
    .D(_0095_),
    .Q_N(_0999_),
    .Q(\vga_clock.sec_counter[18] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[19]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net139),
    .D(_0096_),
    .Q_N(_0998_),
    .Q(\vga_clock.sec_counter[19] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[1]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net140),
    .D(_0097_),
    .Q_N(_0997_),
    .Q(\vga_clock.sec_counter[1] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[20]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net141),
    .D(_0098_),
    .Q_N(_0996_),
    .Q(\vga_clock.sec_counter[20] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[21]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net142),
    .D(_0099_),
    .Q_N(_0995_),
    .Q(\vga_clock.sec_counter[21] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[22]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_0100_),
    .Q_N(_0994_),
    .Q(\vga_clock.sec_counter[22] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[23]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net144),
    .D(_0101_),
    .Q_N(_0993_),
    .Q(\vga_clock.sec_counter[23] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[24]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net145),
    .D(_0102_),
    .Q_N(_0992_),
    .Q(\vga_clock.sec_counter[24] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[25]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net146),
    .D(_0103_),
    .Q_N(_0991_),
    .Q(\vga_clock.sec_counter[25] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[2]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net147),
    .D(_0104_),
    .Q_N(_0990_),
    .Q(\vga_clock.sec_counter[2] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[3]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net148),
    .D(_0105_),
    .Q_N(_0989_),
    .Q(\vga_clock.sec_counter[3] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[4]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net149),
    .D(_0106_),
    .Q_N(_0988_),
    .Q(\vga_clock.sec_counter[4] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[5]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net150),
    .D(_0107_),
    .Q_N(_0987_),
    .Q(\vga_clock.sec_counter[5] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[6]$_SDFF_PP0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net151),
    .D(_0108_),
    .Q_N(_0986_),
    .Q(\vga_clock.sec_counter[6] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[7]$_SDFF_PP0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net152),
    .D(_0109_),
    .Q_N(_0985_),
    .Q(\vga_clock.sec_counter[7] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[8]$_SDFF_PP0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net153),
    .D(_0110_),
    .Q_N(_0984_),
    .Q(\vga_clock.sec_counter[8] ));
 sg13g2_dfrbp_1 \vga_clock.sec_counter[9]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net154),
    .D(_0111_),
    .Q_N(_0983_),
    .Q(\vga_clock.sec_counter[9] ));
 sg13g2_dfrbp_1 \vga_clock.sec_d[0]$_SDFFE_PP0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net155),
    .D(_0112_),
    .Q_N(_0027_),
    .Q(\vga_clock.sec_d[0] ));
 sg13g2_dfrbp_1 \vga_clock.sec_d[1]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net156),
    .D(_0113_),
    .Q_N(_0982_),
    .Q(\vga_clock.sec_d[1] ));
 sg13g2_dfrbp_1 \vga_clock.sec_d[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net157),
    .D(_0114_),
    .Q_N(_0981_),
    .Q(\vga_clock.sec_d[2] ));
 sg13g2_dfrbp_1 \vga_clock.sec_u[0]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net158),
    .D(_0115_),
    .Q_N(_0009_),
    .Q(\vga_clock.sec_u[0] ));
 sg13g2_dfrbp_1 \vga_clock.sec_u[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net159),
    .D(_0116_),
    .Q_N(_0980_),
    .Q(\vga_clock.sec_u[1] ));
 sg13g2_dfrbp_1 \vga_clock.sec_u[2]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net160),
    .D(_0117_),
    .Q_N(_0979_),
    .Q(\vga_clock.sec_u[2] ));
 sg13g2_dfrbp_1 \vga_clock.sec_u[3]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net161),
    .D(_0118_),
    .Q_N(_0022_),
    .Q(\vga_clock.sec_u[3] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[0]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net162),
    .D(_0119_),
    .Q_N(_0025_),
    .Q(\vga_clock.vga_0.hc[0] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[1]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net163),
    .D(_0120_),
    .Q_N(_0978_),
    .Q(\vga_clock.vga_0.hc[1] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[2]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net164),
    .D(_0121_),
    .Q_N(_0977_),
    .Q(\vga_clock.vga_0.hc[2] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[3]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net165),
    .D(_0122_),
    .Q_N(_0976_),
    .Q(\vga_clock.vga_0.hc[3] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[4]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net166),
    .D(_0123_),
    .Q_N(_0975_),
    .Q(\vga_clock.vga_0.hc[4] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[5]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net167),
    .D(_0124_),
    .Q_N(_0974_),
    .Q(\vga_clock.vga_0.hc[5] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[6]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net168),
    .D(_0125_),
    .Q_N(_0026_),
    .Q(\vga_clock.vga_0.hc[6] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[7]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net169),
    .D(_0126_),
    .Q_N(_0973_),
    .Q(\vga_clock.vga_0.hc[7] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[8]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net170),
    .D(_0127_),
    .Q_N(_0012_),
    .Q(\vga_clock.vga_0.hc[8] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.hc[9]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net171),
    .D(_0128_),
    .Q_N(_0972_),
    .Q(\vga_clock.vga_0.hc[9] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[0]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net172),
    .D(_0129_),
    .Q_N(_0971_),
    .Q(\vga_clock.vga_0.vc[0] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[1]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net173),
    .D(_0130_),
    .Q_N(_0970_),
    .Q(\vga_clock.vga_0.vc[1] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[2]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net174),
    .D(_0131_),
    .Q_N(_0969_),
    .Q(\vga_clock.vga_0.vc[2] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[3]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net175),
    .D(_0132_),
    .Q_N(_0024_),
    .Q(\vga_clock.vga_0.vc[3] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[4]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net176),
    .D(_0133_),
    .Q_N(_0968_),
    .Q(\vga_clock.vga_0.vc[4] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[5]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net177),
    .D(_0134_),
    .Q_N(_0023_),
    .Q(\vga_clock.vga_0.vc[5] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[6]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net178),
    .D(_0135_),
    .Q_N(_0008_),
    .Q(\vga_clock.vga_0.vc[6] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[7]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net179),
    .D(_0136_),
    .Q_N(_0967_),
    .Q(\vga_clock.vga_0.vc[7] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[8]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net180),
    .D(_0137_),
    .Q_N(_0966_),
    .Q(\vga_clock.vga_0.vc[8] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.vc[9]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net181),
    .D(_0138_),
    .Q_N(_0965_),
    .Q(\vga_clock.vga_0.vc[9] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[0]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net182),
    .D(_0139_),
    .Q_N(_0964_),
    .Q(\vga_clock.vga_0.x_px[0] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[1]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net183),
    .D(_0140_),
    .Q_N(_0963_),
    .Q(\vga_clock.vga_0.x_px[1] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[2]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net184),
    .D(_0141_),
    .Q_N(_0962_),
    .Q(\vga_clock.vga_0.x_px[2] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[3]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net185),
    .D(_0142_),
    .Q_N(_0961_),
    .Q(\vga_clock.vga_0.x_px[3] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[4]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net186),
    .D(_0143_),
    .Q_N(_0960_),
    .Q(\vga_clock.digit_0.x_block[0] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[5]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net187),
    .D(_0144_),
    .Q_N(_0959_),
    .Q(\vga_clock.digit_0.x_block[1] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[6]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net188),
    .D(_0145_),
    .Q_N(\vga_clock.digit_0.char[0] ),
    .Q(\vga_clock.vga_0.x_px[6] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[7]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net189),
    .D(_0146_),
    .Q_N(_0958_),
    .Q(\vga_clock.vga_0.x_px[7] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[8]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net190),
    .D(_0147_),
    .Q_N(_0957_),
    .Q(\vga_clock.vga_0.x_px[8] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.x_px[9]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net191),
    .D(_0148_),
    .Q_N(_0956_),
    .Q(\vga_clock.vga_0.x_px[9] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[0]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net192),
    .D(_0149_),
    .Q_N(_0955_),
    .Q(\vga_clock.vga_0.y_px[0] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[1]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net193),
    .D(_0150_),
    .Q_N(_0954_),
    .Q(\vga_clock.vga_0.y_px[1] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[2]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net194),
    .D(_0151_),
    .Q_N(_0953_),
    .Q(\vga_clock.vga_0.y_px[2] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[3]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net195),
    .D(_0152_),
    .Q_N(_0952_),
    .Q(\vga_clock.vga_0.y_px[3] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[4]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net196),
    .D(_0153_),
    .Q_N(_0951_),
    .Q(\vga_clock.vga_0.y_px[4] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[5]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net197),
    .D(_0154_),
    .Q_N(_0950_),
    .Q(\vga_clock.vga_0.y_px[5] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[6]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net198),
    .D(_0155_),
    .Q_N(_0949_),
    .Q(\vga_clock.vga_0.y_px[6] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[7]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net199),
    .D(_0156_),
    .Q_N(_0948_),
    .Q(\vga_clock.vga_0.y_px[7] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[8]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net200),
    .D(_0157_),
    .Q_N(_0016_),
    .Q(\vga_clock.vga_0.y_px[8] ));
 sg13g2_dfrbp_1 \vga_clock.vga_0.y_px[9]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net201),
    .D(_0158_),
    .Q_N(_1061_),
    .Q(\vga_clock.vga_0.y_px[9] ));
 sg13g2_dfrbp_1 \vga_clock.x_block_q[5]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net202),
    .D(\vga_clock.digit_0.char[3] ),
    .Q_N(_1062_),
    .Q(\vga_clock.x_block_q[5] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[0]$_DFF_P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net203),
    .D(\vga_clock.y_block[0] ),
    .Q_N(_1063_),
    .Q(\vga_clock.y_block_q[0] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[1]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net204),
    .D(\vga_clock.y_block[1] ),
    .Q_N(_1064_),
    .Q(\vga_clock.y_block_q[1] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[2]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net205),
    .D(\vga_clock.y_block[2] ),
    .Q_N(_1065_),
    .Q(\vga_clock.y_block_q[2] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[3]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net206),
    .D(\vga_clock.y_block[3] ),
    .Q_N(_1066_),
    .Q(\vga_clock.y_block_q[3] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[4]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net207),
    .D(\vga_clock.y_block[4] ),
    .Q_N(_1067_),
    .Q(\vga_clock.y_block_q[4] ));
 sg13g2_dfrbp_1 \vga_clock.y_block_q[5]$_DFF_P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net208),
    .D(\vga_clock.y_block[5] ),
    .Q_N(_0947_),
    .Q(\vga_clock.y_block_q[5] ));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uo_out[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[1]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[2]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[3]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[4]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[5]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[6]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout9 (.A(_0744_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_0733_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0255_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0476_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0473_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0883_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0488_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0453_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0864_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0801_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0401_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(\vga_clock.y_block[0] ),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0411_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0236_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0882_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0832_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0660_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0565_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0373_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0369_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0366_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0334_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0278_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0855_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0790_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0750_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0653_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0481_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0415_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0414_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0409_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0406_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0391_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0372_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0368_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0169_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0821_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0647_),
    .X(net46));
 sg13g2_tielo _2014__47 (.L_LO(net47));
 sg13g2_tielo _2015__48 (.L_LO(net48));
 sg13g2_tielo _2016__49 (.L_LO(net49));
 sg13g2_tielo _2017__50 (.L_LO(net50));
 sg13g2_tielo _2018__51 (.L_LO(net51));
 sg13g2_tielo _2019__52 (.L_LO(net52));
 sg13g2_tielo _2020__53 (.L_LO(net53));
 sg13g2_tielo _2021__54 (.L_LO(net54));
 sg13g2_tielo _2022__55 (.L_LO(net55));
 sg13g2_tielo _2023__56 (.L_LO(net56));
 sg13g2_tielo _2024__57 (.L_LO(net57));
 sg13g2_tielo _2025__58 (.L_LO(net58));
 sg13g2_tielo _2026__59 (.L_LO(net59));
 sg13g2_tielo _2027__60 (.L_LO(net60));
 sg13g2_tielo _2028__61 (.L_LO(net61));
 sg13g2_tielo _2029__62 (.L_LO(net62));
 sg13g2_tiehi \vga_clock.col_index_q[1]$_DFF_P__64  (.L_HI(net64));
 sg13g2_tiehi \vga_clock.color_offset[0]$_SDFFE_PN0P__65  (.L_HI(net65));
 sg13g2_tiehi \vga_clock.color_offset[1]$_SDFFE_PN0P__66  (.L_HI(net66));
 sg13g2_tiehi \vga_clock.color_offset[2]$_SDFFE_PN0P__67  (.L_HI(net67));
 sg13g2_tiehi \vga_clock.digit_0.col_index[0]$_SDFF_PP1__68  (.L_HI(net68));
 sg13g2_tiehi \vga_clock.digit_0.col_index[1]$_SDFF_PP1__69  (.L_HI(net69));
 sg13g2_tiehi \vga_clock.digit_0.color[0]$_SDFF_PP0__70  (.L_HI(net70));
 sg13g2_tiehi \vga_clock.digit_0.color[1]$_SDFF_PP0__71  (.L_HI(net71));
 sg13g2_tiehi \vga_clock.digit_0.color[2]$_SDFF_PP0__72  (.L_HI(net72));
 sg13g2_tiehi \vga_clock.digit_0.color[3]$_SDFF_PN0__73  (.L_HI(net73));
 sg13g2_tiehi \vga_clock.digit_0.color[4]$_DFF_P__74  (.L_HI(net74));
 sg13g2_tiehi \vga_clock.digit_0.color[5]$_DFF_P__75  (.L_HI(net75));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[0]$_DFF_P__76  (.L_HI(net76));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[1]$_DFF_P__77  (.L_HI(net77));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[2]$_DFF_P__78  (.L_HI(net78));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[3]$_DFF_P__79  (.L_HI(net79));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[4]$_DFF_P__80  (.L_HI(net80));
 sg13g2_tiehi \vga_clock.digit_0.digit_index[5]$_SDFF_PP1__81  (.L_HI(net81));
 sg13g2_tiehi \vga_clock.draw$_SDFF_PN0__82  (.L_HI(net82));
 sg13g2_tiehi \vga_clock.font_0.dout[1]$_DFF_P__83  (.L_HI(net83));
 sg13g2_tiehi \vga_clock.font_0.dout[2]$_DFF_P__84  (.L_HI(net84));
 sg13g2_tiehi \vga_clock.font_0.dout[3]$_DFF_P__85  (.L_HI(net85));
 sg13g2_tiehi \vga_clock.hrs_d[0]$_SDFFE_PP0P__86  (.L_HI(net86));
 sg13g2_tiehi \vga_clock.hrs_d[1]$_SDFFE_PP0P__87  (.L_HI(net87));
 sg13g2_tiehi \vga_clock.hrs_u[0]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \vga_clock.hrs_u[1]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \vga_clock.hrs_u[2]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \vga_clock.hrs_u[3]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \vga_clock.min_d[0]$_SDFFE_PP0P__92  (.L_HI(net92));
 sg13g2_tiehi \vga_clock.min_d[1]$_SDFFE_PP0P__93  (.L_HI(net93));
 sg13g2_tiehi \vga_clock.min_d[2]$_SDFFE_PP0P__94  (.L_HI(net94));
 sg13g2_tiehi \vga_clock.min_u[0]$_SDFFE_PN0P__95  (.L_HI(net95));
 sg13g2_tiehi \vga_clock.min_u[1]$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \vga_clock.min_u[2]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \vga_clock.min_u[3]$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \vga_clock.pulse_hrs.comp[0]$_SDFFE_PN1P__99  (.L_HI(net99));
 sg13g2_tiehi \vga_clock.pulse_hrs.comp[1]$_SDFFE_PN1P__100  (.L_HI(net100));
 sg13g2_tiehi \vga_clock.pulse_hrs.comp[2]$_SDFFE_PN1P__101  (.L_HI(net101));
 sg13g2_tiehi \vga_clock.pulse_hrs.comp[3]$_SDFFE_PN1P__102  (.L_HI(net102));
 sg13g2_tiehi \vga_clock.pulse_hrs.comp[4]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \vga_clock.pulse_hrs.count[0]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \vga_clock.pulse_hrs.count[1]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \vga_clock.pulse_hrs.count[2]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \vga_clock.pulse_hrs.count[3]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \vga_clock.pulse_hrs.count[4]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \vga_clock.pulse_min.comp[0]$_SDFFE_PN1P__109  (.L_HI(net109));
 sg13g2_tiehi \vga_clock.pulse_min.comp[1]$_SDFFE_PN1P__110  (.L_HI(net110));
 sg13g2_tiehi \vga_clock.pulse_min.comp[2]$_SDFFE_PN1P__111  (.L_HI(net111));
 sg13g2_tiehi \vga_clock.pulse_min.comp[3]$_SDFFE_PN1P__112  (.L_HI(net112));
 sg13g2_tiehi \vga_clock.pulse_min.comp[4]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \vga_clock.pulse_min.count[0]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \vga_clock.pulse_min.count[1]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \vga_clock.pulse_min.count[2]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \vga_clock.pulse_min.count[3]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \vga_clock.pulse_min.count[4]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \vga_clock.pulse_sec.comp[0]$_SDFFE_PN1P__119  (.L_HI(net119));
 sg13g2_tiehi \vga_clock.pulse_sec.comp[1]$_SDFFE_PN1P__120  (.L_HI(net120));
 sg13g2_tiehi \vga_clock.pulse_sec.comp[2]$_SDFFE_PN1P__121  (.L_HI(net121));
 sg13g2_tiehi \vga_clock.pulse_sec.comp[3]$_SDFFE_PN1P__122  (.L_HI(net122));
 sg13g2_tiehi \vga_clock.pulse_sec.comp[4]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \vga_clock.pulse_sec.count[0]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \vga_clock.pulse_sec.count[1]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \vga_clock.pulse_sec.count[2]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \vga_clock.pulse_sec.count[3]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \vga_clock.pulse_sec.count[4]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \vga_clock.sec_counter[0]$_SDFF_PP0__129  (.L_HI(net129));
 sg13g2_tiehi \vga_clock.sec_counter[10]$_SDFF_PP0__130  (.L_HI(net130));
 sg13g2_tiehi \vga_clock.sec_counter[11]$_SDFF_PP0__131  (.L_HI(net131));
 sg13g2_tiehi \vga_clock.sec_counter[12]$_SDFF_PP0__132  (.L_HI(net132));
 sg13g2_tiehi \vga_clock.sec_counter[13]$_SDFF_PP0__133  (.L_HI(net133));
 sg13g2_tiehi \vga_clock.sec_counter[14]$_SDFF_PP0__134  (.L_HI(net134));
 sg13g2_tiehi \vga_clock.sec_counter[15]$_SDFF_PP0__135  (.L_HI(net135));
 sg13g2_tiehi \vga_clock.sec_counter[16]$_SDFF_PP0__136  (.L_HI(net136));
 sg13g2_tiehi \vga_clock.sec_counter[17]$_SDFF_PP0__137  (.L_HI(net137));
 sg13g2_tiehi \vga_clock.sec_counter[18]$_SDFF_PP0__138  (.L_HI(net138));
 sg13g2_tiehi \vga_clock.sec_counter[19]$_SDFF_PP0__139  (.L_HI(net139));
 sg13g2_tiehi \vga_clock.sec_counter[1]$_SDFF_PP0__140  (.L_HI(net140));
 sg13g2_tiehi \vga_clock.sec_counter[20]$_SDFF_PP0__141  (.L_HI(net141));
 sg13g2_tiehi \vga_clock.sec_counter[21]$_SDFF_PP0__142  (.L_HI(net142));
 sg13g2_tiehi \vga_clock.sec_counter[22]$_SDFF_PP0__143  (.L_HI(net143));
 sg13g2_tiehi \vga_clock.sec_counter[23]$_SDFF_PP0__144  (.L_HI(net144));
 sg13g2_tiehi \vga_clock.sec_counter[24]$_SDFF_PP0__145  (.L_HI(net145));
 sg13g2_tiehi \vga_clock.sec_counter[25]$_SDFF_PP0__146  (.L_HI(net146));
 sg13g2_tiehi \vga_clock.sec_counter[2]$_SDFF_PP0__147  (.L_HI(net147));
 sg13g2_tiehi \vga_clock.sec_counter[3]$_SDFF_PP0__148  (.L_HI(net148));
 sg13g2_tiehi \vga_clock.sec_counter[4]$_SDFF_PP0__149  (.L_HI(net149));
 sg13g2_tiehi \vga_clock.sec_counter[5]$_SDFF_PP0__150  (.L_HI(net150));
 sg13g2_tiehi \vga_clock.sec_counter[6]$_SDFF_PP0__151  (.L_HI(net151));
 sg13g2_tiehi \vga_clock.sec_counter[7]$_SDFF_PP0__152  (.L_HI(net152));
 sg13g2_tiehi \vga_clock.sec_counter[8]$_SDFF_PP0__153  (.L_HI(net153));
 sg13g2_tiehi \vga_clock.sec_counter[9]$_SDFF_PP0__154  (.L_HI(net154));
 sg13g2_tiehi \vga_clock.sec_d[0]$_SDFFE_PP0P__155  (.L_HI(net155));
 sg13g2_tiehi \vga_clock.sec_d[1]$_SDFFE_PP0P__156  (.L_HI(net156));
 sg13g2_tiehi \vga_clock.sec_d[2]$_SDFFE_PP0P__157  (.L_HI(net157));
 sg13g2_tiehi \vga_clock.sec_u[0]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \vga_clock.sec_u[1]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \vga_clock.sec_u[2]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \vga_clock.sec_u[3]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \vga_clock.vga_0.hc[0]$_SDFF_PN0__162  (.L_HI(net162));
 sg13g2_tiehi \vga_clock.vga_0.hc[1]$_SDFF_PN0__163  (.L_HI(net163));
 sg13g2_tiehi \vga_clock.vga_0.hc[2]$_SDFF_PN0__164  (.L_HI(net164));
 sg13g2_tiehi \vga_clock.vga_0.hc[3]$_SDFF_PN0__165  (.L_HI(net165));
 sg13g2_tiehi \vga_clock.vga_0.hc[4]$_SDFF_PN0__166  (.L_HI(net166));
 sg13g2_tiehi \vga_clock.vga_0.hc[5]$_SDFF_PN0__167  (.L_HI(net167));
 sg13g2_tiehi \vga_clock.vga_0.hc[6]$_SDFF_PN0__168  (.L_HI(net168));
 sg13g2_tiehi \vga_clock.vga_0.hc[7]$_SDFF_PN0__169  (.L_HI(net169));
 sg13g2_tiehi \vga_clock.vga_0.hc[8]$_SDFF_PN0__170  (.L_HI(net170));
 sg13g2_tiehi \vga_clock.vga_0.hc[9]$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_tiehi \vga_clock.vga_0.vc[0]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \vga_clock.vga_0.vc[1]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \vga_clock.vga_0.vc[2]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \vga_clock.vga_0.vc[3]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \vga_clock.vga_0.vc[4]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \vga_clock.vga_0.vc[5]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \vga_clock.vga_0.vc[6]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \vga_clock.vga_0.vc[7]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \vga_clock.vga_0.vc[8]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \vga_clock.vga_0.vc[9]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \vga_clock.vga_0.x_px[0]$_SDFF_PN0__182  (.L_HI(net182));
 sg13g2_tiehi \vga_clock.vga_0.x_px[1]$_SDFF_PN0__183  (.L_HI(net183));
 sg13g2_tiehi \vga_clock.vga_0.x_px[2]$_SDFF_PN0__184  (.L_HI(net184));
 sg13g2_tiehi \vga_clock.vga_0.x_px[3]$_SDFF_PN0__185  (.L_HI(net185));
 sg13g2_tiehi \vga_clock.vga_0.x_px[4]$_SDFF_PN0__186  (.L_HI(net186));
 sg13g2_tiehi \vga_clock.vga_0.x_px[5]$_SDFF_PN0__187  (.L_HI(net187));
 sg13g2_tiehi \vga_clock.vga_0.x_px[6]$_SDFF_PN0__188  (.L_HI(net188));
 sg13g2_tiehi \vga_clock.vga_0.x_px[7]$_SDFF_PN0__189  (.L_HI(net189));
 sg13g2_tiehi \vga_clock.vga_0.x_px[8]$_SDFF_PN0__190  (.L_HI(net190));
 sg13g2_tiehi \vga_clock.vga_0.x_px[9]$_SDFF_PN0__191  (.L_HI(net191));
 sg13g2_tiehi \vga_clock.vga_0.y_px[0]$_SDFF_PN0__192  (.L_HI(net192));
 sg13g2_tiehi \vga_clock.vga_0.y_px[1]$_SDFF_PN0__193  (.L_HI(net193));
 sg13g2_tiehi \vga_clock.vga_0.y_px[2]$_SDFF_PN0__194  (.L_HI(net194));
 sg13g2_tiehi \vga_clock.vga_0.y_px[3]$_SDFF_PN0__195  (.L_HI(net195));
 sg13g2_tiehi \vga_clock.vga_0.y_px[4]$_SDFF_PN0__196  (.L_HI(net196));
 sg13g2_tiehi \vga_clock.vga_0.y_px[5]$_SDFF_PN0__197  (.L_HI(net197));
 sg13g2_tiehi \vga_clock.vga_0.y_px[6]$_SDFF_PN0__198  (.L_HI(net198));
 sg13g2_tiehi \vga_clock.vga_0.y_px[7]$_SDFF_PN0__199  (.L_HI(net199));
 sg13g2_tiehi \vga_clock.vga_0.y_px[8]$_SDFF_PN0__200  (.L_HI(net200));
 sg13g2_tiehi \vga_clock.vga_0.y_px[9]$_SDFF_PN0__201  (.L_HI(net201));
 sg13g2_tiehi \vga_clock.x_block_q[5]$_DFF_P__202  (.L_HI(net202));
 sg13g2_tiehi \vga_clock.y_block_q[0]$_DFF_P__203  (.L_HI(net203));
 sg13g2_tiehi \vga_clock.y_block_q[1]$_DFF_P__204  (.L_HI(net204));
 sg13g2_tiehi \vga_clock.y_block_q[2]$_DFF_P__205  (.L_HI(net205));
 sg13g2_tiehi \vga_clock.y_block_q[3]$_DFF_P__206  (.L_HI(net206));
 sg13g2_tiehi \vga_clock.y_block_q[4]$_DFF_P__207  (.L_HI(net207));
 sg13g2_tiehi \vga_clock.y_block_q[5]$_DFF_P__208  (.L_HI(net208));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_fill_1 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_33 ();
 sg13g2_decap_8 FILLER_0_40 ();
 sg13g2_decap_8 FILLER_0_47 ();
 sg13g2_decap_4 FILLER_0_54 ();
 sg13g2_fill_2 FILLER_0_58 ();
 sg13g2_decap_8 FILLER_0_64 ();
 sg13g2_decap_8 FILLER_0_71 ();
 sg13g2_decap_8 FILLER_0_78 ();
 sg13g2_decap_4 FILLER_0_85 ();
 sg13g2_fill_1 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_94 ();
 sg13g2_decap_8 FILLER_0_101 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_decap_8 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_122 ();
 sg13g2_decap_8 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_136 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_15 ();
 sg13g2_fill_1 FILLER_1_52 ();
 sg13g2_fill_1 FILLER_1_79 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_fill_1 FILLER_1_117 ();
 sg13g2_decap_8 FILLER_1_122 ();
 sg13g2_decap_8 FILLER_1_129 ();
 sg13g2_decap_4 FILLER_1_136 ();
 sg13g2_fill_2 FILLER_1_140 ();
 sg13g2_decap_4 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_176 ();
 sg13g2_decap_8 FILLER_1_183 ();
 sg13g2_decap_8 FILLER_1_190 ();
 sg13g2_decap_8 FILLER_1_197 ();
 sg13g2_decap_8 FILLER_1_204 ();
 sg13g2_decap_8 FILLER_1_211 ();
 sg13g2_decap_8 FILLER_1_218 ();
 sg13g2_decap_8 FILLER_1_225 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_decap_8 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_246 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_4 FILLER_2_38 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_60 ();
 sg13g2_fill_2 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_92 ();
 sg13g2_decap_8 FILLER_2_99 ();
 sg13g2_fill_1 FILLER_2_106 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_4 FILLER_2_144 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_fill_1 FILLER_2_153 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_18 ();
 sg13g2_fill_2 FILLER_3_23 ();
 sg13g2_fill_1 FILLER_3_25 ();
 sg13g2_fill_2 FILLER_3_38 ();
 sg13g2_fill_2 FILLER_3_66 ();
 sg13g2_fill_1 FILLER_3_68 ();
 sg13g2_decap_8 FILLER_3_94 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_4 FILLER_3_130 ();
 sg13g2_fill_1 FILLER_3_142 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_177 ();
 sg13g2_decap_8 FILLER_3_188 ();
 sg13g2_decap_8 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_202 ();
 sg13g2_decap_8 FILLER_3_209 ();
 sg13g2_decap_8 FILLER_3_216 ();
 sg13g2_decap_8 FILLER_3_223 ();
 sg13g2_decap_8 FILLER_3_230 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_251 ();
 sg13g2_decap_8 FILLER_3_258 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_300 ();
 sg13g2_decap_8 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_328 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_27 ();
 sg13g2_fill_1 FILLER_4_33 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_fill_2 FILLER_4_46 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_87 ();
 sg13g2_fill_2 FILLER_4_94 ();
 sg13g2_decap_8 FILLER_4_145 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_206 ();
 sg13g2_decap_8 FILLER_4_213 ();
 sg13g2_decap_8 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_227 ();
 sg13g2_decap_8 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_241 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_255 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_9 ();
 sg13g2_decap_8 FILLER_5_16 ();
 sg13g2_fill_2 FILLER_5_23 ();
 sg13g2_decap_8 FILLER_5_33 ();
 sg13g2_decap_8 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_decap_4 FILLER_5_54 ();
 sg13g2_fill_2 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_77 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_fill_2 FILLER_5_101 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_4 FILLER_5_116 ();
 sg13g2_fill_2 FILLER_5_120 ();
 sg13g2_decap_4 FILLER_5_131 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_decap_4 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_90 ();
 sg13g2_decap_4 FILLER_6_97 ();
 sg13g2_fill_2 FILLER_6_101 ();
 sg13g2_fill_1 FILLER_6_107 ();
 sg13g2_decap_4 FILLER_6_113 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_132 ();
 sg13g2_decap_8 FILLER_6_173 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_fill_2 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_8 FILLER_6_250 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_fill_1 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_4 FILLER_6_424 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_11 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_decap_4 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_61 ();
 sg13g2_decap_4 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_111 ();
 sg13g2_decap_8 FILLER_7_146 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_fill_2 FILLER_7_167 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_fill_1 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_decap_4 FILLER_7_265 ();
 sg13g2_fill_2 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_4 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_335 ();
 sg13g2_decap_4 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_4 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_fill_1 FILLER_7_389 ();
 sg13g2_fill_2 FILLER_7_394 ();
 sg13g2_fill_1 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_fill_2 FILLER_8_18 ();
 sg13g2_fill_1 FILLER_8_20 ();
 sg13g2_decap_8 FILLER_8_37 ();
 sg13g2_decap_4 FILLER_8_44 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_decap_8 FILLER_8_79 ();
 sg13g2_decap_8 FILLER_8_86 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_decap_8 FILLER_8_110 ();
 sg13g2_decap_8 FILLER_8_117 ();
 sg13g2_decap_8 FILLER_8_124 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_fill_2 FILLER_8_166 ();
 sg13g2_fill_1 FILLER_8_168 ();
 sg13g2_decap_4 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_222 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_241 ();
 sg13g2_decap_4 FILLER_8_264 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_decap_4 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_4 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_345 ();
 sg13g2_fill_1 FILLER_8_352 ();
 sg13g2_decap_4 FILLER_8_363 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_381 ();
 sg13g2_fill_2 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_4 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_41 ();
 sg13g2_fill_1 FILLER_9_43 ();
 sg13g2_decap_8 FILLER_9_48 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_fill_2 FILLER_9_137 ();
 sg13g2_fill_2 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_decap_4 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_257 ();
 sg13g2_fill_1 FILLER_9_259 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_318 ();
 sg13g2_decap_4 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_fill_1 FILLER_9_345 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_fill_2 FILLER_9_382 ();
 sg13g2_fill_1 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_decap_4 FILLER_10_54 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_4 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_4 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_120 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_180 ();
 sg13g2_decap_4 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_fill_1 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_4 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_decap_4 FILLER_11_75 ();
 sg13g2_fill_2 FILLER_11_79 ();
 sg13g2_decap_8 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_decap_4 FILLER_11_111 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_155 ();
 sg13g2_decap_8 FILLER_11_183 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_4 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_4 FILLER_11_328 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_342 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_decap_4 FILLER_11_356 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_375 ();
 sg13g2_fill_2 FILLER_11_388 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_410 ();
 sg13g2_fill_1 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_418 ();
 sg13g2_decap_4 FILLER_11_425 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_decap_4 FILLER_12_115 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_decap_8 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_285 ();
 sg13g2_fill_1 FILLER_12_290 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_328 ();
 sg13g2_decap_4 FILLER_12_334 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_decap_4 FILLER_12_374 ();
 sg13g2_fill_2 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_12_398 ();
 sg13g2_fill_1 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_13_31 ();
 sg13g2_decap_8 FILLER_13_41 ();
 sg13g2_decap_4 FILLER_13_48 ();
 sg13g2_decap_4 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_79 ();
 sg13g2_fill_1 FILLER_13_90 ();
 sg13g2_fill_1 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_decap_4 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_4 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_344 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_378 ();
 sg13g2_fill_1 FILLER_13_384 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_395 ();
 sg13g2_fill_1 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_25 ();
 sg13g2_fill_2 FILLER_14_36 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_64 ();
 sg13g2_decap_4 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_fill_1 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_decap_4 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_fill_2 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_4 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_decap_4 FILLER_14_337 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_4 FILLER_14_395 ();
 sg13g2_fill_1 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_4 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_87 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_140 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_decap_4 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_289 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_4 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_decap_4 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_16_31 ();
 sg13g2_decap_8 FILLER_16_38 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_decap_4 FILLER_16_110 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_fill_2 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_11 ();
 sg13g2_decap_8 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_32 ();
 sg13g2_decap_8 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_decap_4 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_decap_4 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_4 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_decap_4 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_375 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_4 FILLER_18_30 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_decap_4 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_decap_4 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_decap_4 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_fill_2 FILLER_18_405 ();
 sg13g2_fill_1 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_8 FILLER_19_15 ();
 sg13g2_decap_4 FILLER_19_22 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_decap_4 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_65 ();
 sg13g2_fill_1 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_decap_4 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_decap_4 FILLER_20_44 ();
 sg13g2_decap_4 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_58 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_decap_8 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_4 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_52 ();
 sg13g2_decap_4 FILLER_21_59 ();
 sg13g2_decap_4 FILLER_21_72 ();
 sg13g2_decap_4 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_142 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_4 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_decap_4 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_decap_4 FILLER_21_372 ();
 sg13g2_decap_4 FILLER_21_389 ();
 sg13g2_fill_2 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_20 ();
 sg13g2_decap_8 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_decap_8 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_decap_4 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_4 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_404 ();
 sg13g2_fill_2 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_decap_4 FILLER_23_48 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_decap_4 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_79 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_decap_8 FILLER_23_99 ();
 sg13g2_decap_8 FILLER_23_106 ();
 sg13g2_decap_8 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_decap_4 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_decap_4 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_4 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_4 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_decap_4 FILLER_23_415 ();
 sg13g2_decap_4 FILLER_23_424 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_33 ();
 sg13g2_decap_4 FILLER_24_40 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_decap_4 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_146 ();
 sg13g2_decap_8 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_4 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_4 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_decap_4 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_decap_4 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_decap_4 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_decap_4 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_decap_4 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_4 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_13 ();
 sg13g2_fill_2 FILLER_26_20 ();
 sg13g2_fill_1 FILLER_26_22 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_decap_8 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_4 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_4 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_52 ();
 sg13g2_decap_4 FILLER_27_59 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_4 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_299 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_27_409 ();
 sg13g2_decap_4 FILLER_27_415 ();
 sg13g2_fill_1 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_17 ();
 sg13g2_decap_8 FILLER_28_24 ();
 sg13g2_decap_4 FILLER_28_31 ();
 sg13g2_decap_8 FILLER_28_48 ();
 sg13g2_decap_8 FILLER_28_55 ();
 sg13g2_decap_4 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_decap_4 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_decap_4 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_29 ();
 sg13g2_decap_8 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_decap_4 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_decap_4 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_decap_4 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_10 ();
 sg13g2_fill_2 FILLER_30_41 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_decap_4 FILLER_30_374 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_2 FILLER_31_29 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_37 ();
 sg13g2_decap_8 FILLER_31_54 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_decap_4 FILLER_31_149 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_decap_4 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_decap_4 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_decap_4 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_4 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_31_401 ();
 sg13g2_fill_2 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_15 ();
 sg13g2_fill_2 FILLER_32_22 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_2 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_289 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_412 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_4 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_decap_8 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_decap_4 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_decap_4 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_245 ();
 sg13g2_decap_4 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_61 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_82 ();
 sg13g2_decap_8 FILLER_34_101 ();
 sg13g2_decap_4 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_44 ();
 sg13g2_decap_4 FILLER_35_51 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_decap_8 FILLER_35_80 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_113 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_215 ();
 sg13g2_decap_4 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_decap_4 FILLER_35_318 ();
 sg13g2_decap_4 FILLER_35_356 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_35_413 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_decap_4 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_16 ();
 sg13g2_decap_8 FILLER_36_23 ();
 sg13g2_decap_8 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_decap_4 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_48 ();
 sg13g2_decap_4 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_decap_4 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_decap_4 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_decap_4 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_decap_4 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_4 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_397 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_decap_4 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_decap_4 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_1 FILLER_37_407 ();
 sg13g2_decap_4 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_decap_4 FILLER_38_366 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_decap_4 FILLER_38_376 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_1 FILLER_38_394 ();
 sg13g2_fill_2 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
