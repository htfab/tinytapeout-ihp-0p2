module tt_um_tomkeddie_a (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire clknet_0_clk;
 wire net93;
 wire b0;
 wire g0;
 wire hs;
 wire \vga.ball_angle[0] ;
 wire \vga.ball_angle[1] ;
 wire \vga.ball_angle[2] ;
 wire \vga.ball_angle[3] ;
 wire \vga.ball_motion_l ;
 wire \vga.ball_pos_h[0] ;
 wire \vga.ball_pos_h[1] ;
 wire \vga.ball_pos_h[2] ;
 wire \vga.ball_pos_h[3] ;
 wire \vga.ball_pos_h[4] ;
 wire \vga.ball_pos_h[5] ;
 wire \vga.ball_pos_h[6] ;
 wire \vga.ball_pos_h[7] ;
 wire \vga.ball_pos_h[8] ;
 wire \vga.ball_pos_h[9] ;
 wire \vga.ball_pos_v[0] ;
 wire \vga.ball_pos_v[1] ;
 wire \vga.ball_pos_v[2] ;
 wire \vga.ball_pos_v[3] ;
 wire \vga.ball_pos_v[4] ;
 wire \vga.ball_pos_v[5] ;
 wire \vga.ball_pos_v[6] ;
 wire \vga.ball_pos_v[7] ;
 wire \vga.ball_pos_v[8] ;
 wire \vga.ball_ratio[0] ;
 wire \vga.ball_ratio[1] ;
 wire \vga.ball_ratio[2] ;
 wire \vga.blank_h ;
 wire \vga.blank_v ;
 wire \vga.count_h[0] ;
 wire \vga.count_h[1] ;
 wire \vga.count_h[2] ;
 wire \vga.count_h[3] ;
 wire \vga.count_h[4] ;
 wire \vga.count_h[5] ;
 wire \vga.count_h[6] ;
 wire \vga.count_h[7] ;
 wire \vga.count_h[8] ;
 wire \vga.count_h[9] ;
 wire \vga.count_v[0] ;
 wire \vga.count_v[1] ;
 wire \vga.count_v[2] ;
 wire \vga.count_v[3] ;
 wire \vga.count_v[4] ;
 wire \vga.count_v[5] ;
 wire \vga.count_v[6] ;
 wire \vga.count_v[7] ;
 wire \vga.count_v[8] ;
 wire \vga.count_v[9] ;
 wire \vga.hs_out ;
 wire \vga.interval_counter[0] ;
 wire \vga.interval_counter[10] ;
 wire \vga.interval_counter[11] ;
 wire \vga.interval_counter[12] ;
 wire \vga.interval_counter[13] ;
 wire \vga.interval_counter[14] ;
 wire \vga.interval_counter[15] ;
 wire \vga.interval_counter[16] ;
 wire \vga.interval_counter[17] ;
 wire \vga.interval_counter[18] ;
 wire \vga.interval_counter[19] ;
 wire \vga.interval_counter[1] ;
 wire \vga.interval_counter[20] ;
 wire \vga.interval_counter[21] ;
 wire \vga.interval_counter[22] ;
 wire \vga.interval_counter[23] ;
 wire \vga.interval_counter[24] ;
 wire \vga.interval_counter[2] ;
 wire \vga.interval_counter[3] ;
 wire \vga.interval_counter[4] ;
 wire \vga.interval_counter[5] ;
 wire \vga.interval_counter[6] ;
 wire \vga.interval_counter[7] ;
 wire \vga.interval_counter[8] ;
 wire \vga.interval_counter[9] ;
 wire \vga.left_down_1d ;
 wire \vga.left_down_pressed ;
 wire \vga.left_up_1d ;
 wire \vga.left_up_pressed ;
 wire \vga.paddle_l_pos_v[0] ;
 wire \vga.paddle_l_pos_v[1] ;
 wire \vga.paddle_l_pos_v[2] ;
 wire \vga.paddle_l_pos_v[3] ;
 wire \vga.paddle_l_pos_v[4] ;
 wire \vga.paddle_l_pos_v[5] ;
 wire \vga.paddle_l_pos_v[6] ;
 wire \vga.paddle_l_pos_v[7] ;
 wire \vga.paddle_l_pos_v[8] ;
 wire \vga.paddle_r_pos_v[0] ;
 wire \vga.paddle_r_pos_v[1] ;
 wire \vga.paddle_r_pos_v[2] ;
 wire \vga.paddle_r_pos_v[3] ;
 wire \vga.paddle_r_pos_v[4] ;
 wire \vga.paddle_r_pos_v[5] ;
 wire \vga.paddle_r_pos_v[6] ;
 wire \vga.paddle_r_pos_v[7] ;
 wire \vga.paddle_r_pos_v[8] ;
 wire \vga.right_down_1d ;
 wire \vga.right_down_pressed ;
 wire \vga.right_up_1d ;
 wire \vga.right_up_pressed ;
 wire \vga.score_l[0] ;
 wire \vga.score_l[1] ;
 wire \vga.score_l[2] ;
 wire \vga.score_l[3] ;
 wire \vga.score_l[4] ;
 wire \vga.score_l_ten_enable ;
 wire \vga.score_l_unit_pixels[0] ;
 wire \vga.score_l_unit_pixels[1] ;
 wire \vga.score_l_unit_pixels[2] ;
 wire \vga.score_r[0] ;
 wire \vga.score_r[1] ;
 wire \vga.score_r[2] ;
 wire \vga.score_r[3] ;
 wire \vga.score_r[4] ;
 wire \vga.score_r_ten_enable ;
 wire \vga.score_r_unit_pixels[0] ;
 wire \vga.score_r_unit_pixels[1] ;
 wire \vga.score_r_unit_pixels[2] ;
 wire \vga.speed_lsb_1d ;
 wire \vga.speed_msb_1d ;
 wire \vga.vs ;
 wire \vga.vs_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_1 _2120_ (.Y(_1404_),
    .A(\vga.score_l[4] ));
 sg13g2_buf_1 _2121_ (.A(\vga.score_l[1] ),
    .X(_1405_));
 sg13g2_buf_1 _2122_ (.A(\vga.score_l[0] ),
    .X(_1406_));
 sg13g2_nand2_1 _2123_ (.Y(_1407_),
    .A(_1405_),
    .B(_1406_));
 sg13g2_nor4_1 _2124_ (.A(\vga.score_l[3] ),
    .B(\vga.score_l[2] ),
    .C(_1404_),
    .D(_1407_),
    .Y(_1408_));
 sg13g2_inv_1 _2125_ (.Y(_1409_),
    .A(\vga.score_l[2] ));
 sg13g2_nand2_1 _2126_ (.Y(_1410_),
    .A(_1407_),
    .B(_1409_));
 sg13g2_nand3_1 _2127_ (.B(_1406_),
    .C(\vga.score_l[2] ),
    .A(_1405_),
    .Y(_1411_));
 sg13g2_nand2_1 _2128_ (.Y(_1412_),
    .A(_1410_),
    .B(_1411_));
 sg13g2_buf_2 _2129_ (.A(\vga.ball_pos_v[7] ),
    .X(_1413_));
 sg13g2_buf_2 _2130_ (.A(\vga.paddle_r_pos_v[7] ),
    .X(_1414_));
 sg13g2_inv_1 _2131_ (.Y(_1415_),
    .A(_1414_));
 sg13g2_buf_8 _2132_ (.A(\vga.paddle_r_pos_v[3] ),
    .X(_1416_));
 sg13g2_buf_8 _2133_ (.A(\vga.paddle_r_pos_v[2] ),
    .X(_1417_));
 sg13g2_nand2_2 _2134_ (.Y(_1418_),
    .A(_1416_),
    .B(_1417_));
 sg13g2_inv_4 _2135_ (.A(_1418_),
    .Y(_1419_));
 sg13g2_buf_2 _2136_ (.A(\vga.paddle_r_pos_v[4] ),
    .X(_1420_));
 sg13g2_inv_2 _2137_ (.Y(_1421_),
    .A(_1420_));
 sg13g2_nand2_1 _2138_ (.Y(_1422_),
    .A(_1419_),
    .B(_1421_));
 sg13g2_nand2_1 _2139_ (.Y(_1423_),
    .A(_1422_),
    .B(_0061_));
 sg13g2_buf_8 _2140_ (.A(\vga.paddle_r_pos_v[5] ),
    .X(_1424_));
 sg13g2_buf_8 _2141_ (.A(\vga.paddle_r_pos_v[6] ),
    .X(_1425_));
 sg13g2_nand2_1 _2142_ (.Y(_1426_),
    .A(_1424_),
    .B(_1425_));
 sg13g2_inv_2 _2143_ (.Y(_1427_),
    .A(_1426_));
 sg13g2_nand2_1 _2144_ (.Y(_1428_),
    .A(_1423_),
    .B(_1427_));
 sg13g2_xnor2_1 _2145_ (.Y(_1429_),
    .A(_1415_),
    .B(_1428_));
 sg13g2_buf_1 _2146_ (.A(_0067_),
    .X(_1430_));
 sg13g2_inv_2 _2147_ (.Y(_1431_),
    .A(_1430_));
 sg13g2_buf_2 _2148_ (.A(\vga.paddle_r_pos_v[8] ),
    .X(_1432_));
 sg13g2_o21ai_1 _2149_ (.B1(_1427_),
    .Y(_1433_),
    .A1(_1420_),
    .A2(_1419_));
 sg13g2_nor2_1 _2150_ (.A(_1415_),
    .B(_1433_),
    .Y(_1434_));
 sg13g2_xor2_1 _2151_ (.B(_1434_),
    .A(_1432_),
    .X(_1435_));
 sg13g2_xnor2_1 _2152_ (.Y(_1436_),
    .A(_1431_),
    .B(_1435_));
 sg13g2_o21ai_1 _2153_ (.B1(_1436_),
    .Y(_1437_),
    .A1(_1413_),
    .A2(_1429_));
 sg13g2_buf_1 _2154_ (.A(\vga.ball_pos_v[4] ),
    .X(_1438_));
 sg13g2_buf_1 _2155_ (.A(_1438_),
    .X(_1439_));
 sg13g2_xnor2_1 _2156_ (.Y(_1440_),
    .A(_1421_),
    .B(_1418_));
 sg13g2_inv_1 _2157_ (.Y(_1441_),
    .A(_1440_));
 sg13g2_nor2_1 _2158_ (.A(net70),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_buf_1 _2159_ (.A(\vga.ball_pos_v[1] ),
    .X(_1443_));
 sg13g2_inv_1 _2160_ (.Y(_1444_),
    .A(net88));
 sg13g2_buf_2 _2161_ (.A(\vga.paddle_r_pos_v[1] ),
    .X(_1445_));
 sg13g2_nand2_1 _2162_ (.Y(_1446_),
    .A(_1444_),
    .B(_1445_));
 sg13g2_buf_1 _2163_ (.A(\vga.ball_pos_v[0] ),
    .X(_1447_));
 sg13g2_inv_2 _2164_ (.Y(_1448_),
    .A(net87));
 sg13g2_buf_2 _2165_ (.A(\vga.paddle_r_pos_v[0] ),
    .X(_1449_));
 sg13g2_nand2_1 _2166_ (.Y(_1450_),
    .A(net69),
    .B(_1449_));
 sg13g2_nor2_1 _2167_ (.A(_1445_),
    .B(_1444_),
    .Y(_1451_));
 sg13g2_a21oi_1 _2168_ (.A1(_1446_),
    .A2(_1450_),
    .Y(_1452_),
    .B1(_1451_));
 sg13g2_buf_1 _2169_ (.A(\vga.ball_pos_v[2] ),
    .X(_1453_));
 sg13g2_nand2_1 _2170_ (.Y(_1454_),
    .A(_1417_),
    .B(net86));
 sg13g2_inv_1 _2171_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_buf_1 _2172_ (.A(_1417_),
    .X(_1456_));
 sg13g2_nor2_1 _2173_ (.A(_1456_),
    .B(net86),
    .Y(_1457_));
 sg13g2_inv_1 _2174_ (.Y(_1458_),
    .A(_0075_));
 sg13g2_nor2_2 _2175_ (.A(_1416_),
    .B(_1417_),
    .Y(_1459_));
 sg13g2_inv_1 _2176_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_nand2_2 _2177_ (.Y(_1461_),
    .A(_1460_),
    .B(_1418_));
 sg13g2_xnor2_1 _2178_ (.Y(_1462_),
    .A(_1458_),
    .B(_1461_));
 sg13g2_nor3_1 _2179_ (.A(_1455_),
    .B(_1457_),
    .C(_1462_),
    .Y(_1463_));
 sg13g2_nand2b_1 _2180_ (.Y(_1464_),
    .B(_1463_),
    .A_N(_1452_));
 sg13g2_buf_1 _2181_ (.A(\vga.ball_pos_v[3] ),
    .X(_1465_));
 sg13g2_nor2_1 _2182_ (.A(_1454_),
    .B(_1462_),
    .Y(_1466_));
 sg13g2_a21oi_1 _2183_ (.A1(net85),
    .A2(_1461_),
    .Y(_1467_),
    .B1(_1466_));
 sg13g2_nand2_1 _2184_ (.Y(_1468_),
    .A(_1464_),
    .B(_1467_));
 sg13g2_nand2b_1 _2185_ (.Y(_1469_),
    .B(_1468_),
    .A_N(_1442_));
 sg13g2_buf_1 _2186_ (.A(\vga.ball_pos_v[5] ),
    .X(_1470_));
 sg13g2_buf_1 _2187_ (.A(_1470_),
    .X(_1471_));
 sg13g2_inv_2 _2188_ (.Y(_1472_),
    .A(_1424_));
 sg13g2_xnor2_1 _2189_ (.Y(_1473_),
    .A(_1472_),
    .B(_1423_));
 sg13g2_inv_1 _2190_ (.Y(_1474_),
    .A(_1473_));
 sg13g2_a22oi_1 _2191_ (.Y(_1475_),
    .B1(net67),
    .B2(_1474_),
    .A2(_1441_),
    .A1(net70));
 sg13g2_nand2_1 _2192_ (.Y(_1476_),
    .A(_1469_),
    .B(_1475_));
 sg13g2_buf_2 _2193_ (.A(_0071_),
    .X(_1477_));
 sg13g2_o21ai_1 _2194_ (.B1(_1424_),
    .Y(_1478_),
    .A1(_1420_),
    .A2(_1419_));
 sg13g2_inv_2 _2195_ (.Y(_1479_),
    .A(_1425_));
 sg13g2_nand2_1 _2196_ (.Y(_1480_),
    .A(_1478_),
    .B(_1479_));
 sg13g2_nand2_1 _2197_ (.Y(_1481_),
    .A(_1480_),
    .B(_1433_));
 sg13g2_xnor2_1 _2198_ (.Y(_1482_),
    .A(_1477_),
    .B(_1481_));
 sg13g2_nand2_1 _2199_ (.Y(_1483_),
    .A(_1429_),
    .B(_1413_));
 sg13g2_nand2_1 _2200_ (.Y(_1484_),
    .A(_1482_),
    .B(_1483_));
 sg13g2_inv_1 _2201_ (.Y(_1485_),
    .A(net67));
 sg13g2_nand2_1 _2202_ (.Y(_1486_),
    .A(_1473_),
    .B(_1485_));
 sg13g2_nor2b_1 _2203_ (.A(_1484_),
    .B_N(_1486_),
    .Y(_1487_));
 sg13g2_nand2_1 _2204_ (.Y(_1488_),
    .A(_1476_),
    .B(_1487_));
 sg13g2_buf_1 _2205_ (.A(\vga.ball_pos_v[6] ),
    .X(_1489_));
 sg13g2_a22oi_1 _2206_ (.Y(_1490_),
    .B1(_1413_),
    .B2(_1429_),
    .A2(_1481_),
    .A1(_1489_));
 sg13g2_nand2_1 _2207_ (.Y(_1491_),
    .A(_1488_),
    .B(_1490_));
 sg13g2_nand2b_1 _2208_ (.Y(_1492_),
    .B(_1491_),
    .A_N(_1437_));
 sg13g2_buf_1 _2209_ (.A(\vga.ball_pos_v[8] ),
    .X(_1493_));
 sg13g2_nand2b_1 _2210_ (.Y(_1494_),
    .B(net83),
    .A_N(_1435_));
 sg13g2_nand2_1 _2211_ (.Y(_1495_),
    .A(_1492_),
    .B(_1494_));
 sg13g2_nand2_1 _2212_ (.Y(_1496_),
    .A(_1414_),
    .B(_1432_));
 sg13g2_nor2_1 _2213_ (.A(_1496_),
    .B(_1428_),
    .Y(_1497_));
 sg13g2_inv_1 _2214_ (.Y(_1498_),
    .A(_1449_));
 sg13g2_inv_2 _2215_ (.Y(_1499_),
    .A(_1438_));
 sg13g2_nand3b_1 _2216_ (.B(_1446_),
    .C(_1450_),
    .Y(_1500_),
    .A_N(_1451_));
 sg13g2_a221oi_1 _2217_ (.B2(_1499_),
    .C1(_1500_),
    .B1(_1440_),
    .A1(_1498_),
    .Y(_1501_),
    .A2(net87));
 sg13g2_nand4_1 _2218_ (.B(_1501_),
    .C(_1463_),
    .A(_1475_),
    .Y(_1502_),
    .D(_1486_));
 sg13g2_nor3_1 _2219_ (.A(_1484_),
    .B(_1502_),
    .C(_1437_),
    .Y(_1503_));
 sg13g2_nor2_1 _2220_ (.A(_1497_),
    .B(_1503_),
    .Y(_1504_));
 sg13g2_nand2_1 _2221_ (.Y(_1505_),
    .A(_1495_),
    .B(_1504_));
 sg13g2_inv_1 _2222_ (.Y(_1506_),
    .A(_0073_));
 sg13g2_nand2_1 _2223_ (.Y(_1507_),
    .A(_1472_),
    .B(_1479_));
 sg13g2_nor2_2 _2224_ (.A(_1421_),
    .B(_1459_),
    .Y(_1508_));
 sg13g2_nor2_1 _2225_ (.A(_1507_),
    .B(_1508_),
    .Y(_1509_));
 sg13g2_xnor2_1 _2226_ (.Y(_1510_),
    .A(_1414_),
    .B(_1509_));
 sg13g2_inv_1 _2227_ (.Y(_1511_),
    .A(_0069_));
 sg13g2_a21oi_2 _2228_ (.B1(_1511_),
    .Y(_1512_),
    .A2(_1472_),
    .A1(_1508_));
 sg13g2_nand3_1 _2229_ (.B(_1415_),
    .C(_1479_),
    .A(_1512_),
    .Y(_1513_));
 sg13g2_xnor2_1 _2230_ (.Y(_1514_),
    .A(_0068_),
    .B(_1513_));
 sg13g2_xnor2_1 _2231_ (.Y(_1515_),
    .A(_1479_),
    .B(_1512_));
 sg13g2_inv_2 _2232_ (.Y(_1516_),
    .A(_1413_));
 sg13g2_xnor2_1 _2233_ (.Y(_1517_),
    .A(_0070_),
    .B(_1509_));
 sg13g2_xnor2_1 _2234_ (.Y(_1518_),
    .A(net66),
    .B(_1517_));
 sg13g2_nor3_1 _2235_ (.A(_1477_),
    .B(_1515_),
    .C(_1518_),
    .Y(_1519_));
 sg13g2_a221oi_1 _2236_ (.B2(_1514_),
    .C1(_1519_),
    .B1(net83),
    .A1(_1506_),
    .Y(_1520_),
    .A2(_1510_));
 sg13g2_inv_1 _2237_ (.Y(_1521_),
    .A(net85));
 sg13g2_a21o_1 _2238_ (.A2(_1454_),
    .A1(_1452_),
    .B1(_1457_),
    .X(_1522_));
 sg13g2_o21ai_1 _2239_ (.B1(_1522_),
    .Y(_1523_),
    .A1(_1521_),
    .A2(_1461_));
 sg13g2_xnor2_1 _2240_ (.Y(_1524_),
    .A(_1511_),
    .B(_1508_));
 sg13g2_xnor2_1 _2241_ (.Y(_1525_),
    .A(net67),
    .B(_1524_));
 sg13g2_xnor2_1 _2242_ (.Y(_1526_),
    .A(_1421_),
    .B(_1459_));
 sg13g2_inv_1 _2243_ (.Y(_1527_),
    .A(_1526_));
 sg13g2_inv_1 _2244_ (.Y(_1528_),
    .A(_1461_));
 sg13g2_nand2_1 _2245_ (.Y(_1529_),
    .A(_1526_),
    .B(_1438_));
 sg13g2_o21ai_1 _2246_ (.B1(_1529_),
    .Y(_1530_),
    .A1(net85),
    .A2(_1528_));
 sg13g2_a21oi_1 _2247_ (.A1(_1499_),
    .A2(_1527_),
    .Y(_1531_),
    .B1(_1530_));
 sg13g2_nand3_1 _2248_ (.B(_1525_),
    .C(_1531_),
    .A(_1523_),
    .Y(_1532_));
 sg13g2_inv_1 _2249_ (.Y(_1533_),
    .A(_0074_));
 sg13g2_xnor2_1 _2250_ (.Y(_1534_),
    .A(_1472_),
    .B(_1508_));
 sg13g2_inv_1 _2251_ (.Y(_1535_),
    .A(_1529_));
 sg13g2_a22oi_1 _2252_ (.Y(_1536_),
    .B1(_1535_),
    .B2(_1525_),
    .A2(_1534_),
    .A1(_1533_));
 sg13g2_nand2_1 _2253_ (.Y(_1537_),
    .A(_1532_),
    .B(_1536_));
 sg13g2_xnor2_1 _2254_ (.Y(_1538_),
    .A(_0072_),
    .B(_1512_));
 sg13g2_inv_2 _2255_ (.Y(_1539_),
    .A(_1477_));
 sg13g2_nand2b_1 _2256_ (.Y(_1540_),
    .B(_1539_),
    .A_N(_1538_));
 sg13g2_a21oi_1 _2257_ (.A1(_1477_),
    .A2(_1538_),
    .Y(_1541_),
    .B1(_1518_));
 sg13g2_nand3_1 _2258_ (.B(_1540_),
    .C(_1541_),
    .A(_1537_),
    .Y(_1542_));
 sg13g2_nand2_1 _2259_ (.Y(_1543_),
    .A(_1520_),
    .B(_1542_));
 sg13g2_o21ai_1 _2260_ (.B1(_1514_),
    .Y(_1544_),
    .A1(_1430_),
    .A2(net83));
 sg13g2_inv_1 _2261_ (.Y(_1545_),
    .A(_1514_));
 sg13g2_nand2_1 _2262_ (.Y(_1546_),
    .A(_1545_),
    .B(_1431_));
 sg13g2_nor2_1 _2263_ (.A(_1414_),
    .B(_1432_),
    .Y(_1547_));
 sg13g2_nand2_1 _2264_ (.Y(_1548_),
    .A(_1509_),
    .B(_1547_));
 sg13g2_inv_1 _2265_ (.Y(_1549_),
    .A(_1548_));
 sg13g2_a21oi_1 _2266_ (.A1(_1544_),
    .A2(_1546_),
    .Y(_1550_),
    .B1(_1549_));
 sg13g2_nand2_1 _2267_ (.Y(_1551_),
    .A(_1543_),
    .B(_1550_));
 sg13g2_inv_1 _2268_ (.Y(_1552_),
    .A(_1551_));
 sg13g2_nand2_1 _2269_ (.Y(_1553_),
    .A(_1505_),
    .B(_1552_));
 sg13g2_buf_8 _2270_ (.A(_1553_),
    .X(_1554_));
 sg13g2_o21ai_1 _2271_ (.B1(_1554_),
    .Y(_1555_),
    .A1(_1408_),
    .A2(_1412_));
 sg13g2_a21oi_1 _2272_ (.A1(_1495_),
    .A2(_1504_),
    .Y(_1556_),
    .B1(_1551_));
 sg13g2_buf_2 _2273_ (.A(ui_in[4]),
    .X(_1557_));
 sg13g2_nor2_1 _2274_ (.A(_1557_),
    .B(_1409_),
    .Y(_1558_));
 sg13g2_inv_1 _2275_ (.Y(_1559_),
    .A(_1558_));
 sg13g2_nand2_1 _2276_ (.Y(_1560_),
    .A(_1556_),
    .B(_1559_));
 sg13g2_buf_1 _2277_ (.A(\vga.ball_motion_l ),
    .X(_1561_));
 sg13g2_buf_2 _2278_ (.A(\vga.ball_pos_h[3] ),
    .X(_1562_));
 sg13g2_buf_2 _2279_ (.A(\vga.ball_pos_h[2] ),
    .X(_1563_));
 sg13g2_nand2_2 _2280_ (.Y(_1564_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_buf_8 _2281_ (.A(\vga.ball_pos_h[0] ),
    .X(_1565_));
 sg13g2_buf_1 _2282_ (.A(\vga.ball_pos_h[1] ),
    .X(_1566_));
 sg13g2_nand2_1 _2283_ (.Y(_1567_),
    .A(_1565_),
    .B(_1566_));
 sg13g2_nor2_1 _2284_ (.A(_1564_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_buf_2 _2285_ (.A(\vga.ball_pos_h[7] ),
    .X(_1569_));
 sg13g2_buf_1 _2286_ (.A(\vga.ball_pos_h[8] ),
    .X(_1570_));
 sg13g2_buf_1 _2287_ (.A(\vga.ball_pos_h[9] ),
    .X(_1571_));
 sg13g2_inv_1 _2288_ (.Y(_1572_),
    .A(_1571_));
 sg13g2_nor3_1 _2289_ (.A(_1569_),
    .B(net81),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_buf_1 _2290_ (.A(\vga.ball_pos_h[4] ),
    .X(_1574_));
 sg13g2_inv_1 _2291_ (.Y(_1575_),
    .A(net80));
 sg13g2_buf_2 _2292_ (.A(\vga.ball_pos_h[5] ),
    .X(_1576_));
 sg13g2_buf_2 _2293_ (.A(\vga.ball_pos_h[6] ),
    .X(_1577_));
 sg13g2_nand2_1 _2294_ (.Y(_1578_),
    .A(_1576_),
    .B(_1577_));
 sg13g2_inv_1 _2295_ (.Y(_1579_),
    .A(_1578_));
 sg13g2_nand4_1 _2296_ (.B(_1573_),
    .C(_1575_),
    .A(_1568_),
    .Y(_1580_),
    .D(_1579_));
 sg13g2_nor2_1 _2297_ (.A(net82),
    .B(_1580_),
    .Y(_1581_));
 sg13g2_buf_2 _2298_ (.A(_1581_),
    .X(_1582_));
 sg13g2_nand3_1 _2299_ (.B(_1560_),
    .C(_1582_),
    .A(_1555_),
    .Y(_1583_));
 sg13g2_inv_4 _2300_ (.A(_1582_),
    .Y(_1584_));
 sg13g2_inv_1 _2301_ (.Y(_1585_),
    .A(\vga.interval_counter[23] ));
 sg13g2_inv_1 _2302_ (.Y(_1586_),
    .A(\vga.interval_counter[22] ));
 sg13g2_inv_1 _2303_ (.Y(_1587_),
    .A(\vga.interval_counter[24] ));
 sg13g2_nand3_1 _2304_ (.B(_1586_),
    .C(_1587_),
    .A(_1585_),
    .Y(_1588_));
 sg13g2_nor3_1 _2305_ (.A(\vga.interval_counter[21] ),
    .B(\vga.interval_counter[20] ),
    .C(_1588_),
    .Y(_1589_));
 sg13g2_buf_1 _2306_ (.A(\vga.interval_counter[7] ),
    .X(_1590_));
 sg13g2_buf_1 _2307_ (.A(\vga.interval_counter[6] ),
    .X(_1591_));
 sg13g2_nor2_1 _2308_ (.A(_1590_),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_buf_1 _2309_ (.A(\vga.interval_counter[3] ),
    .X(_1593_));
 sg13g2_buf_8 _2310_ (.A(\vga.interval_counter[2] ),
    .X(_1594_));
 sg13g2_nor2_1 _2311_ (.A(\vga.interval_counter[19] ),
    .B(\vga.interval_counter[18] ),
    .Y(_1595_));
 sg13g2_inv_1 _2312_ (.Y(_1596_),
    .A(_1595_));
 sg13g2_nor3_1 _2313_ (.A(_1593_),
    .B(_1594_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_nand3_1 _2314_ (.B(_1592_),
    .C(_1597_),
    .A(_1589_),
    .Y(_1598_));
 sg13g2_buf_8 _2315_ (.A(\vga.interval_counter[0] ),
    .X(_1599_));
 sg13g2_buf_1 _2316_ (.A(\vga.interval_counter[15] ),
    .X(_1600_));
 sg13g2_buf_2 _2317_ (.A(\vga.interval_counter[13] ),
    .X(_1601_));
 sg13g2_nor2_1 _2318_ (.A(_1601_),
    .B(\vga.interval_counter[12] ),
    .Y(_1602_));
 sg13g2_inv_1 _2319_ (.Y(_1603_),
    .A(\vga.interval_counter[4] ));
 sg13g2_buf_1 _2320_ (.A(\vga.interval_counter[5] ),
    .X(_1604_));
 sg13g2_inv_1 _2321_ (.Y(_1605_),
    .A(_1604_));
 sg13g2_nand3_1 _2322_ (.B(_1603_),
    .C(_1605_),
    .A(_1602_),
    .Y(_1606_));
 sg13g2_nor4_1 _2323_ (.A(\vga.interval_counter[1] ),
    .B(_1599_),
    .C(_1600_),
    .D(_1606_),
    .Y(_1607_));
 sg13g2_buf_1 _2324_ (.A(\vga.interval_counter[8] ),
    .X(_1608_));
 sg13g2_nor4_1 _2325_ (.A(_1608_),
    .B(\vga.interval_counter[9] ),
    .C(\vga.interval_counter[11] ),
    .D(\vga.interval_counter[10] ),
    .Y(_1609_));
 sg13g2_buf_2 _2326_ (.A(\vga.interval_counter[14] ),
    .X(_1610_));
 sg13g2_nor3_1 _2327_ (.A(_1610_),
    .B(\vga.interval_counter[16] ),
    .C(\vga.interval_counter[17] ),
    .Y(_1611_));
 sg13g2_nand3_1 _2328_ (.B(_1609_),
    .C(_1611_),
    .A(_1607_),
    .Y(_1612_));
 sg13g2_nor2_1 _2329_ (.A(_1598_),
    .B(_1612_),
    .Y(_1613_));
 sg13g2_inv_1 _2330_ (.Y(_1614_),
    .A(_1613_));
 sg13g2_buf_1 _2331_ (.A(_1614_),
    .X(_1615_));
 sg13g2_a21oi_1 _2332_ (.A1(net51),
    .A2(_1558_),
    .Y(_1616_),
    .B1(net48));
 sg13g2_nand2_1 _2333_ (.Y(_1617_),
    .A(_1583_),
    .B(_1616_));
 sg13g2_buf_1 _2334_ (.A(rst_n),
    .X(_1618_));
 sg13g2_inv_1 _2335_ (.Y(_1619_),
    .A(_1618_));
 sg13g2_buf_1 _2336_ (.A(_1619_),
    .X(_1620_));
 sg13g2_a21oi_1 _2337_ (.A1(net48),
    .A2(_1559_),
    .Y(_1621_),
    .B1(net65));
 sg13g2_nand2_1 _2338_ (.Y(_1622_),
    .A(_1617_),
    .B(_1621_));
 sg13g2_buf_8 _2339_ (.A(_1622_),
    .X(_1623_));
 sg13g2_inv_1 _2340_ (.Y(_1624_),
    .A(_1408_));
 sg13g2_nor2_1 _2341_ (.A(net51),
    .B(net48),
    .Y(_1625_));
 sg13g2_nand3_1 _2342_ (.B(_1624_),
    .C(_1625_),
    .A(_1554_),
    .Y(_1626_));
 sg13g2_nor2b_1 _2343_ (.A(_1557_),
    .B_N(_1405_),
    .Y(_1627_));
 sg13g2_inv_1 _2344_ (.Y(_1628_),
    .A(_1625_));
 sg13g2_xor2_1 _2345_ (.B(_1406_),
    .A(_1405_),
    .X(_1629_));
 sg13g2_inv_1 _2346_ (.Y(_1630_),
    .A(_1629_));
 sg13g2_nor3_1 _2347_ (.A(_1628_),
    .B(_1630_),
    .C(_1556_),
    .Y(_1631_));
 sg13g2_a21oi_2 _2348_ (.B1(_1631_),
    .Y(_1632_),
    .A2(_1627_),
    .A1(_1626_));
 sg13g2_nor2_1 _2349_ (.A(net65),
    .B(_1632_),
    .Y(_0197_));
 sg13g2_inv_1 _2350_ (.Y(_1633_),
    .A(_1557_));
 sg13g2_nand2_1 _2351_ (.Y(_1634_),
    .A(_1633_),
    .B(_1406_));
 sg13g2_nand2_1 _2352_ (.Y(_1635_),
    .A(_1626_),
    .B(_1634_));
 sg13g2_nand4_1 _2353_ (.B(_1406_),
    .C(_1624_),
    .A(_1554_),
    .Y(_1636_),
    .D(_1625_));
 sg13g2_nand3_1 _2354_ (.B(_1636_),
    .C(_1618_),
    .A(_1635_),
    .Y(_1637_));
 sg13g2_buf_2 _2355_ (.A(_1637_),
    .X(_1638_));
 sg13g2_nand2_1 _2356_ (.Y(_1639_),
    .A(_0197_),
    .B(_1638_));
 sg13g2_nor2_1 _2357_ (.A(_1623_),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_nand2_1 _2358_ (.Y(_1641_),
    .A(_1554_),
    .B(_1624_));
 sg13g2_inv_1 _2359_ (.Y(_1642_),
    .A(\vga.score_l[3] ));
 sg13g2_nor2_1 _2360_ (.A(_1557_),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_inv_1 _2361_ (.Y(_1644_),
    .A(_1643_));
 sg13g2_nand2_1 _2362_ (.Y(_1645_),
    .A(_1641_),
    .B(_1644_));
 sg13g2_xnor2_1 _2363_ (.Y(_1646_),
    .A(_1642_),
    .B(_1411_));
 sg13g2_nand3_1 _2364_ (.B(_1646_),
    .C(_1624_),
    .A(_1554_),
    .Y(_1647_));
 sg13g2_nand3_1 _2365_ (.B(_1647_),
    .C(_1582_),
    .A(_1645_),
    .Y(_1648_));
 sg13g2_a21oi_1 _2366_ (.A1(net51),
    .A2(_1643_),
    .Y(_1649_),
    .B1(net48));
 sg13g2_buf_1 _2367_ (.A(_1613_),
    .X(_1650_));
 sg13g2_o21ai_1 _2368_ (.B1(_1618_),
    .Y(_1651_),
    .A1(_1643_),
    .A2(net50));
 sg13g2_a21oi_1 _2369_ (.A1(_1648_),
    .A2(_1649_),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_buf_2 _2370_ (.A(_1652_),
    .X(_0199_));
 sg13g2_inv_2 _2371_ (.Y(_1653_),
    .A(_0199_));
 sg13g2_buf_1 _2372_ (.A(_1653_),
    .X(_1654_));
 sg13g2_nand2_1 _2373_ (.Y(_1655_),
    .A(_1623_),
    .B(_1638_));
 sg13g2_inv_2 _2374_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_a21oi_1 _2375_ (.A1(_1640_),
    .A2(net29),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_nand2_1 _2376_ (.Y(_1658_),
    .A(_1626_),
    .B(_1627_));
 sg13g2_nand2b_1 _2377_ (.Y(_1659_),
    .B(_1658_),
    .A_N(_1631_));
 sg13g2_buf_1 _2378_ (.A(_1618_),
    .X(_1660_));
 sg13g2_nand2_1 _2379_ (.Y(_1661_),
    .A(_1659_),
    .B(net79));
 sg13g2_nand2_1 _2380_ (.Y(_1662_),
    .A(_1661_),
    .B(_1638_));
 sg13g2_inv_1 _2381_ (.Y(_1663_),
    .A(_1662_));
 sg13g2_inv_1 _2382_ (.Y(_1664_),
    .A(_1621_));
 sg13g2_a21oi_1 _2383_ (.A1(_1583_),
    .A2(_1616_),
    .Y(_1665_),
    .B1(_1664_));
 sg13g2_buf_2 _2384_ (.A(_1665_),
    .X(_0198_));
 sg13g2_nand3_1 _2385_ (.B(_0199_),
    .C(_0198_),
    .A(_1663_),
    .Y(_1666_));
 sg13g2_nor2_1 _2386_ (.A(_1628_),
    .B(_1556_),
    .Y(_1667_));
 sg13g2_a22oi_1 _2387_ (.Y(_1668_),
    .B1(_1624_),
    .B2(_1667_),
    .A2(_1633_),
    .A1(\vga.score_l[4] ));
 sg13g2_nor2_1 _2388_ (.A(_1642_),
    .B(_1411_),
    .Y(_1669_));
 sg13g2_xnor2_1 _2389_ (.Y(_1670_),
    .A(\vga.score_l[4] ),
    .B(_1669_));
 sg13g2_a21oi_1 _2390_ (.A1(_1667_),
    .A2(_1670_),
    .Y(_1671_),
    .B1(net65));
 sg13g2_nor2b_1 _2391_ (.A(_1668_),
    .B_N(_1671_),
    .Y(_1672_));
 sg13g2_buf_1 _2392_ (.A(_1672_),
    .X(_0200_));
 sg13g2_inv_2 _2393_ (.Y(_1673_),
    .A(net38));
 sg13g2_a21oi_1 _2394_ (.A1(_1656_),
    .A2(net29),
    .Y(_1674_),
    .B1(_1673_));
 sg13g2_a21oi_1 _2395_ (.A1(_1657_),
    .A2(_1666_),
    .Y(_0008_),
    .B1(_1674_));
 sg13g2_buf_8 _2396_ (.A(\vga.paddle_l_pos_v[4] ),
    .X(_1675_));
 sg13g2_inv_8 _2397_ (.Y(_1676_),
    .A(_1675_));
 sg13g2_buf_8 _2398_ (.A(\vga.paddle_l_pos_v[3] ),
    .X(_1677_));
 sg13g2_buf_8 _2399_ (.A(\vga.paddle_l_pos_v[2] ),
    .X(_1678_));
 sg13g2_nand3_1 _2400_ (.B(_1677_),
    .C(_1678_),
    .A(_1676_),
    .Y(_1679_));
 sg13g2_buf_1 _2401_ (.A(_1679_),
    .X(_1680_));
 sg13g2_nand2_1 _2402_ (.Y(_1681_),
    .A(_1680_),
    .B(_0059_));
 sg13g2_buf_2 _2403_ (.A(\vga.paddle_l_pos_v[6] ),
    .X(_1682_));
 sg13g2_buf_2 _2404_ (.A(\vga.paddle_l_pos_v[5] ),
    .X(_1683_));
 sg13g2_nand2_1 _2405_ (.Y(_1684_),
    .A(_1682_),
    .B(_1683_));
 sg13g2_inv_1 _2406_ (.Y(_1685_),
    .A(_1684_));
 sg13g2_nand2_1 _2407_ (.Y(_1686_),
    .A(_1681_),
    .B(_1685_));
 sg13g2_buf_1 _2408_ (.A(\vga.paddle_l_pos_v[7] ),
    .X(_1687_));
 sg13g2_inv_2 _2409_ (.Y(_1688_),
    .A(_1687_));
 sg13g2_nand2_1 _2410_ (.Y(_1689_),
    .A(_1686_),
    .B(net64));
 sg13g2_nand3_1 _2411_ (.B(_1687_),
    .C(_1685_),
    .A(_1681_),
    .Y(_1690_));
 sg13g2_nand2_1 _2412_ (.Y(_1691_),
    .A(_1689_),
    .B(_1690_));
 sg13g2_nand2_1 _2413_ (.Y(_1692_),
    .A(_1691_),
    .B(_1413_));
 sg13g2_nand3_1 _2414_ (.B(_1690_),
    .C(_1516_),
    .A(_1689_),
    .Y(_1693_));
 sg13g2_nand2_1 _2415_ (.Y(_1694_),
    .A(_1692_),
    .B(_1693_));
 sg13g2_nand2_1 _2416_ (.Y(_1695_),
    .A(_1677_),
    .B(_1678_));
 sg13g2_nand2_1 _2417_ (.Y(_1696_),
    .A(_1695_),
    .B(_1676_));
 sg13g2_nand2_1 _2418_ (.Y(_1697_),
    .A(_1696_),
    .B(_1683_));
 sg13g2_inv_1 _2419_ (.Y(_1698_),
    .A(_1682_));
 sg13g2_nand2_1 _2420_ (.Y(_1699_),
    .A(_1697_),
    .B(_1698_));
 sg13g2_nand2_1 _2421_ (.Y(_1700_),
    .A(_1696_),
    .B(_1685_));
 sg13g2_nand2_1 _2422_ (.Y(_1701_),
    .A(_1699_),
    .B(_1700_));
 sg13g2_xnor2_1 _2423_ (.Y(_1702_),
    .A(_1477_),
    .B(_1701_));
 sg13g2_nor2b_1 _2424_ (.A(_1694_),
    .B_N(_1702_),
    .Y(_1703_));
 sg13g2_nand2_1 _2425_ (.Y(_1704_),
    .A(_1681_),
    .B(_1683_));
 sg13g2_inv_1 _2426_ (.Y(_1705_),
    .A(_1683_));
 sg13g2_nand3_1 _2427_ (.B(_1705_),
    .C(_0059_),
    .A(_1680_),
    .Y(_1706_));
 sg13g2_nand2_1 _2428_ (.Y(_1707_),
    .A(_1704_),
    .B(_1706_));
 sg13g2_nand2_1 _2429_ (.Y(_1708_),
    .A(_1707_),
    .B(_1470_));
 sg13g2_nand2_1 _2430_ (.Y(_1709_),
    .A(_1695_),
    .B(_1675_));
 sg13g2_nand2_1 _2431_ (.Y(_1710_),
    .A(_1680_),
    .B(_1709_));
 sg13g2_nand2_1 _2432_ (.Y(_1711_),
    .A(_1710_),
    .B(_1438_));
 sg13g2_nor2_1 _2433_ (.A(_1470_),
    .B(_1707_),
    .Y(_1712_));
 sg13g2_a21oi_1 _2434_ (.A1(_1708_),
    .A2(_1711_),
    .Y(_1713_),
    .B1(_1712_));
 sg13g2_inv_1 _2435_ (.Y(_1714_),
    .A(net84));
 sg13g2_a21oi_1 _2436_ (.A1(_1699_),
    .A2(_1700_),
    .Y(_1715_),
    .B1(_1714_));
 sg13g2_nand2_1 _2437_ (.Y(_1716_),
    .A(_1693_),
    .B(_1715_));
 sg13g2_nand2_1 _2438_ (.Y(_1717_),
    .A(_1716_),
    .B(_1692_));
 sg13g2_a21oi_1 _2439_ (.A1(_1703_),
    .A2(_1713_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_nor2_1 _2440_ (.A(_1439_),
    .B(_1710_),
    .Y(_1719_));
 sg13g2_nand2_1 _2441_ (.Y(_1720_),
    .A(_1708_),
    .B(_1711_));
 sg13g2_nor3_1 _2442_ (.A(_1712_),
    .B(_1719_),
    .C(_1720_),
    .Y(_1721_));
 sg13g2_nor2_2 _2443_ (.A(_1677_),
    .B(_1678_),
    .Y(_1722_));
 sg13g2_inv_1 _2444_ (.Y(_1723_),
    .A(_1722_));
 sg13g2_nand2_2 _2445_ (.Y(_1724_),
    .A(_1723_),
    .B(_1695_));
 sg13g2_buf_2 _2446_ (.A(\vga.paddle_l_pos_v[1] ),
    .X(_1725_));
 sg13g2_nand2_1 _2447_ (.Y(_1726_),
    .A(_1444_),
    .B(_1725_));
 sg13g2_buf_1 _2448_ (.A(\vga.paddle_l_pos_v[0] ),
    .X(_1727_));
 sg13g2_nand2_1 _2449_ (.Y(_1728_),
    .A(_1448_),
    .B(_1727_));
 sg13g2_nor2_1 _2450_ (.A(_1725_),
    .B(_1444_),
    .Y(_1729_));
 sg13g2_a21oi_1 _2451_ (.A1(_1726_),
    .A2(_1728_),
    .Y(_1730_),
    .B1(_1729_));
 sg13g2_buf_1 _2452_ (.A(_1678_),
    .X(_1731_));
 sg13g2_xor2_1 _2453_ (.B(net86),
    .A(net63),
    .X(_1732_));
 sg13g2_nor2b_1 _2454_ (.A(_1730_),
    .B_N(_1732_),
    .Y(_1733_));
 sg13g2_xnor2_1 _2455_ (.Y(_1734_),
    .A(_0075_),
    .B(_1724_));
 sg13g2_a22oi_1 _2456_ (.Y(_1735_),
    .B1(_1733_),
    .B2(_1734_),
    .A2(_1724_),
    .A1(net85));
 sg13g2_nand3_1 _2457_ (.B(net63),
    .C(net86),
    .A(_1734_),
    .Y(_1736_));
 sg13g2_nand2_1 _2458_ (.Y(_1737_),
    .A(_1735_),
    .B(_1736_));
 sg13g2_nand3_1 _2459_ (.B(_1721_),
    .C(_1737_),
    .A(_1703_),
    .Y(_1738_));
 sg13g2_nand2_1 _2460_ (.Y(_1739_),
    .A(_1718_),
    .B(_1738_));
 sg13g2_nand2_1 _2461_ (.Y(_1740_),
    .A(\vga.paddle_l_pos_v[8] ),
    .B(_1687_));
 sg13g2_nor2_1 _2462_ (.A(_1740_),
    .B(_1686_),
    .Y(_1741_));
 sg13g2_nor2_1 _2463_ (.A(net64),
    .B(_1700_),
    .Y(_1742_));
 sg13g2_xnor2_1 _2464_ (.Y(_1743_),
    .A(\vga.paddle_l_pos_v[8] ),
    .B(_1742_));
 sg13g2_xnor2_1 _2465_ (.Y(_1744_),
    .A(_1431_),
    .B(_1743_));
 sg13g2_nor2_1 _2466_ (.A(_1741_),
    .B(_1744_),
    .Y(_1745_));
 sg13g2_nand2_1 _2467_ (.Y(_1746_),
    .A(_1739_),
    .B(_1745_));
 sg13g2_nand3b_1 _2468_ (.B(_1743_),
    .C(net83),
    .Y(_1747_),
    .A_N(_1741_));
 sg13g2_nand2_1 _2469_ (.Y(_1748_),
    .A(_1746_),
    .B(_1747_));
 sg13g2_inv_1 _2470_ (.Y(_1749_),
    .A(_1727_));
 sg13g2_nand3b_1 _2471_ (.B(_1726_),
    .C(_1728_),
    .Y(_1750_),
    .A_N(_1729_));
 sg13g2_a21oi_1 _2472_ (.A1(_1749_),
    .A2(net87),
    .Y(_1751_),
    .B1(_1750_));
 sg13g2_and3_1 _2473_ (.X(_1752_),
    .A(_1751_),
    .B(_1732_),
    .C(_1734_));
 sg13g2_nand4_1 _2474_ (.B(_1703_),
    .C(_1721_),
    .A(_1745_),
    .Y(_1753_),
    .D(_1752_));
 sg13g2_nand2_1 _2475_ (.Y(_1754_),
    .A(_1748_),
    .B(_1753_));
 sg13g2_nor2_2 _2476_ (.A(_1676_),
    .B(_1722_),
    .Y(_1755_));
 sg13g2_nand2_1 _2477_ (.Y(_1756_),
    .A(_1755_),
    .B(_1705_));
 sg13g2_nand2_1 _2478_ (.Y(_1757_),
    .A(_1756_),
    .B(_0077_));
 sg13g2_xnor2_1 _2479_ (.Y(_1758_),
    .A(_1698_),
    .B(_1757_));
 sg13g2_nand2_1 _2480_ (.Y(_1759_),
    .A(_1758_),
    .B(_1539_));
 sg13g2_inv_1 _2481_ (.Y(_1760_),
    .A(_0078_));
 sg13g2_inv_1 _2482_ (.Y(_1761_),
    .A(_1755_));
 sg13g2_nor2_1 _2483_ (.A(_1682_),
    .B(_1683_),
    .Y(_1762_));
 sg13g2_nand2_1 _2484_ (.Y(_1763_),
    .A(_1761_),
    .B(_1762_));
 sg13g2_xnor2_1 _2485_ (.Y(_1764_),
    .A(_1760_),
    .B(_1763_));
 sg13g2_xnor2_1 _2486_ (.Y(_1765_),
    .A(net66),
    .B(_1764_));
 sg13g2_xnor2_1 _2487_ (.Y(_1766_),
    .A(net64),
    .B(_1763_));
 sg13g2_nand2_1 _2488_ (.Y(_1767_),
    .A(_1766_),
    .B(_1506_));
 sg13g2_o21ai_1 _2489_ (.B1(_1767_),
    .Y(_1768_),
    .A1(_1759_),
    .A2(_1765_));
 sg13g2_xnor2_1 _2490_ (.Y(_1769_),
    .A(_1683_),
    .B(_1755_));
 sg13g2_inv_1 _2491_ (.Y(_1770_),
    .A(_1769_));
 sg13g2_xnor2_1 _2492_ (.Y(_1771_),
    .A(_1675_),
    .B(_1722_));
 sg13g2_nor2_1 _2493_ (.A(_1499_),
    .B(_1771_),
    .Y(_1772_));
 sg13g2_inv_1 _2494_ (.Y(_1773_),
    .A(_0077_));
 sg13g2_xnor2_1 _2495_ (.Y(_1774_),
    .A(_1773_),
    .B(_1755_));
 sg13g2_xnor2_1 _2496_ (.Y(_1775_),
    .A(_1470_),
    .B(_1774_));
 sg13g2_a22oi_1 _2497_ (.Y(_1776_),
    .B1(_1772_),
    .B2(_1775_),
    .A2(_1770_),
    .A1(_1533_));
 sg13g2_inv_1 _2498_ (.Y(_1777_),
    .A(_0079_));
 sg13g2_xnor2_1 _2499_ (.Y(_1778_),
    .A(_1777_),
    .B(_1757_));
 sg13g2_xnor2_1 _2500_ (.Y(_1779_),
    .A(_1539_),
    .B(_1778_));
 sg13g2_nand2b_1 _2501_ (.Y(_1780_),
    .B(_1779_),
    .A_N(_1765_));
 sg13g2_nor2_1 _2502_ (.A(_1776_),
    .B(_1780_),
    .Y(_1781_));
 sg13g2_nor2_1 _2503_ (.A(_1768_),
    .B(_1781_),
    .Y(_1782_));
 sg13g2_xnor2_1 _2504_ (.Y(_1783_),
    .A(_1499_),
    .B(_1771_));
 sg13g2_nand2b_1 _2505_ (.Y(_1784_),
    .B(_1775_),
    .A_N(_1783_));
 sg13g2_nor2_1 _2506_ (.A(_1784_),
    .B(_1780_),
    .Y(_1785_));
 sg13g2_inv_1 _2507_ (.Y(_1786_),
    .A(_1724_));
 sg13g2_a221oi_1 _2508_ (.B2(_1786_),
    .C1(_1733_),
    .B1(net85),
    .A1(net63),
    .Y(_1787_),
    .A2(net86));
 sg13g2_a21oi_1 _2509_ (.A1(_1521_),
    .A2(_1724_),
    .Y(_1788_),
    .B1(_1787_));
 sg13g2_nand2_1 _2510_ (.Y(_1789_),
    .A(_1785_),
    .B(_1788_));
 sg13g2_nand2_1 _2511_ (.Y(_1790_),
    .A(_1782_),
    .B(_1789_));
 sg13g2_inv_1 _2512_ (.Y(_1791_),
    .A(\vga.paddle_l_pos_v[8] ));
 sg13g2_nand3_1 _2513_ (.B(_1791_),
    .C(net64),
    .A(_1762_),
    .Y(_1792_));
 sg13g2_nor2_1 _2514_ (.A(_1755_),
    .B(_1792_),
    .Y(_1793_));
 sg13g2_nand4_1 _2515_ (.B(_1688_),
    .C(_1698_),
    .A(_1756_),
    .Y(_1794_),
    .D(_0077_));
 sg13g2_xnor2_1 _2516_ (.Y(_1795_),
    .A(_0076_),
    .B(_1794_));
 sg13g2_xnor2_1 _2517_ (.Y(_1796_),
    .A(_1431_),
    .B(_1795_));
 sg13g2_nor2_1 _2518_ (.A(_1793_),
    .B(_1796_),
    .Y(_1797_));
 sg13g2_nand2_1 _2519_ (.Y(_1798_),
    .A(_1790_),
    .B(_1797_));
 sg13g2_inv_1 _2520_ (.Y(_1799_),
    .A(_1793_));
 sg13g2_nand3_1 _2521_ (.B(net83),
    .C(_1799_),
    .A(_1795_),
    .Y(_1800_));
 sg13g2_nand2_1 _2522_ (.Y(_1801_),
    .A(_1798_),
    .B(_1800_));
 sg13g2_nand2_1 _2523_ (.Y(_1802_),
    .A(_1754_),
    .B(_1801_));
 sg13g2_buf_8 _2524_ (.A(_1802_),
    .X(_1803_));
 sg13g2_nor2_1 _2525_ (.A(_1569_),
    .B(_1577_),
    .Y(_1804_));
 sg13g2_inv_1 _2526_ (.Y(_1805_),
    .A(_1804_));
 sg13g2_nor2_1 _2527_ (.A(net80),
    .B(_1576_),
    .Y(_1806_));
 sg13g2_inv_1 _2528_ (.Y(_1807_),
    .A(_1806_));
 sg13g2_nor4_1 _2529_ (.A(net81),
    .B(_1571_),
    .C(_1805_),
    .D(_1807_),
    .Y(_1808_));
 sg13g2_inv_1 _2530_ (.Y(_1809_),
    .A(_1565_));
 sg13g2_buf_1 _2531_ (.A(_1566_),
    .X(_1810_));
 sg13g2_nor3_1 _2532_ (.A(net62),
    .B(net61),
    .C(_1564_),
    .Y(_1811_));
 sg13g2_nand2_1 _2533_ (.Y(_1812_),
    .A(_1808_),
    .B(_1811_));
 sg13g2_inv_1 _2534_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_nand2_1 _2535_ (.Y(_1814_),
    .A(_1803_),
    .B(_1813_));
 sg13g2_buf_1 _2536_ (.A(\vga.score_r[1] ),
    .X(_1815_));
 sg13g2_nand2_1 _2537_ (.Y(_1816_),
    .A(_1633_),
    .B(_1815_));
 sg13g2_inv_1 _2538_ (.Y(_1817_),
    .A(_1816_));
 sg13g2_nand2_1 _2539_ (.Y(_1818_),
    .A(_1814_),
    .B(_1817_));
 sg13g2_buf_1 _2540_ (.A(\vga.score_r[3] ),
    .X(_1819_));
 sg13g2_buf_1 _2541_ (.A(\vga.score_r[2] ),
    .X(_1820_));
 sg13g2_inv_1 _2542_ (.Y(_1821_),
    .A(\vga.score_r[4] ));
 sg13g2_nand2_1 _2543_ (.Y(_1822_),
    .A(_1815_),
    .B(\vga.score_r[0] ));
 sg13g2_nor4_2 _2544_ (.A(_1819_),
    .B(_1820_),
    .C(_1821_),
    .Y(_1823_),
    .D(_1822_));
 sg13g2_xor2_1 _2545_ (.B(\vga.score_r[0] ),
    .A(_1815_),
    .X(_1824_));
 sg13g2_a21oi_1 _2546_ (.A1(_1823_),
    .A2(_1817_),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_inv_1 _2547_ (.Y(_1826_),
    .A(_1825_));
 sg13g2_nand3_1 _2548_ (.B(_1813_),
    .C(_1826_),
    .A(_1803_),
    .Y(_1827_));
 sg13g2_inv_2 _2549_ (.Y(_1828_),
    .A(net82));
 sg13g2_nor2_1 _2550_ (.A(_1828_),
    .B(net48),
    .Y(_1829_));
 sg13g2_nand3_1 _2551_ (.B(_1827_),
    .C(_1829_),
    .A(_1818_),
    .Y(_1830_));
 sg13g2_inv_1 _2552_ (.Y(_1831_),
    .A(_1823_));
 sg13g2_nor2_1 _2553_ (.A(net81),
    .B(_1571_),
    .Y(_1832_));
 sg13g2_nand2b_1 _2554_ (.Y(_1833_),
    .B(_1832_),
    .A_N(net61));
 sg13g2_nor2_1 _2555_ (.A(_1805_),
    .B(_1807_),
    .Y(_1834_));
 sg13g2_inv_1 _2556_ (.Y(_1835_),
    .A(_1834_));
 sg13g2_nor4_2 _2557_ (.A(net62),
    .B(_1564_),
    .C(_1833_),
    .Y(_1836_),
    .D(_1835_));
 sg13g2_nand2_2 _2558_ (.Y(_1837_),
    .A(_1836_),
    .B(net82));
 sg13g2_nor2_1 _2559_ (.A(_1837_),
    .B(_1614_),
    .Y(_1838_));
 sg13g2_nand3_1 _2560_ (.B(_1831_),
    .C(_1838_),
    .A(_1803_),
    .Y(_1839_));
 sg13g2_nor2b_1 _2561_ (.A(_1557_),
    .B_N(\vga.score_r[0] ),
    .Y(_1840_));
 sg13g2_inv_1 _2562_ (.Y(_1841_),
    .A(_1840_));
 sg13g2_nand2_1 _2563_ (.Y(_1842_),
    .A(_1839_),
    .B(_1841_));
 sg13g2_nand4_1 _2564_ (.B(\vga.score_r[0] ),
    .C(_1831_),
    .A(_1803_),
    .Y(_1843_),
    .D(_1838_));
 sg13g2_nand2_1 _2565_ (.Y(_1844_),
    .A(_1842_),
    .B(_1843_));
 sg13g2_inv_1 _2566_ (.Y(_1845_),
    .A(_1829_));
 sg13g2_a21oi_1 _2567_ (.A1(_1845_),
    .A2(_1816_),
    .Y(_1846_),
    .B1(net65));
 sg13g2_nand3_1 _2568_ (.B(_1844_),
    .C(_1846_),
    .A(_1830_),
    .Y(_1847_));
 sg13g2_inv_2 _2569_ (.Y(_1848_),
    .A(_1847_));
 sg13g2_nor2_1 _2570_ (.A(_1828_),
    .B(_1812_),
    .Y(_1849_));
 sg13g2_inv_1 _2571_ (.Y(_1850_),
    .A(_1822_));
 sg13g2_nand2_1 _2572_ (.Y(_1851_),
    .A(_1850_),
    .B(_1820_));
 sg13g2_nand2b_1 _2573_ (.Y(_1852_),
    .B(_1822_),
    .A_N(_1820_));
 sg13g2_nand3_1 _2574_ (.B(_1851_),
    .C(_1852_),
    .A(_1849_),
    .Y(_1853_));
 sg13g2_nand3b_1 _2575_ (.B(_1803_),
    .C(_1831_),
    .Y(_1854_),
    .A_N(_1853_));
 sg13g2_nor2b_1 _2576_ (.A(_1557_),
    .B_N(_1820_),
    .Y(_1855_));
 sg13g2_a21oi_1 _2577_ (.A1(_1855_),
    .A2(_1837_),
    .Y(_1856_),
    .B1(net48));
 sg13g2_nand2_1 _2578_ (.Y(_1857_),
    .A(_1854_),
    .B(_1856_));
 sg13g2_buf_1 _2579_ (.A(_1849_),
    .X(_1858_));
 sg13g2_nand4_1 _2580_ (.B(_1801_),
    .C(_1855_),
    .A(_1754_),
    .Y(_1859_),
    .D(_1858_));
 sg13g2_nor2b_1 _2581_ (.A(_1857_),
    .B_N(_1859_),
    .Y(_1860_));
 sg13g2_nor2_1 _2582_ (.A(_1855_),
    .B(_1613_),
    .Y(_1861_));
 sg13g2_nor2_1 _2583_ (.A(_1620_),
    .B(_1861_),
    .Y(_1862_));
 sg13g2_nor2b_1 _2584_ (.A(_1860_),
    .B_N(_1862_),
    .Y(_1863_));
 sg13g2_buf_1 _2585_ (.A(_1863_),
    .X(_0207_));
 sg13g2_inv_1 _2586_ (.Y(_1864_),
    .A(net35));
 sg13g2_inv_1 _2587_ (.Y(_1865_),
    .A(_1819_));
 sg13g2_nor2_1 _2588_ (.A(_1865_),
    .B(_1851_),
    .Y(_1866_));
 sg13g2_a21oi_1 _2589_ (.A1(_1850_),
    .A2(_1820_),
    .Y(_1867_),
    .B1(_1819_));
 sg13g2_o21ai_1 _2590_ (.B1(_1803_),
    .Y(_1868_),
    .A1(_1866_),
    .A2(_1867_));
 sg13g2_nor2_1 _2591_ (.A(_1557_),
    .B(_1865_),
    .Y(_1869_));
 sg13g2_inv_1 _2592_ (.Y(_1870_),
    .A(_1869_));
 sg13g2_nand3_1 _2593_ (.B(_1801_),
    .C(_1870_),
    .A(_1754_),
    .Y(_1871_));
 sg13g2_nand3_1 _2594_ (.B(_1858_),
    .C(_1871_),
    .A(_1868_),
    .Y(_1872_));
 sg13g2_a21oi_1 _2595_ (.A1(_1837_),
    .A2(_1869_),
    .Y(_1873_),
    .B1(_1615_));
 sg13g2_o21ai_1 _2596_ (.B1(_1618_),
    .Y(_1874_),
    .A1(_1869_),
    .A2(_1613_));
 sg13g2_a21oi_1 _2597_ (.A1(_1872_),
    .A2(_1873_),
    .Y(_1875_),
    .B1(_1874_));
 sg13g2_buf_1 _2598_ (.A(_1875_),
    .X(_0208_));
 sg13g2_nand3_1 _2599_ (.B(_1864_),
    .C(net37),
    .A(_1848_),
    .Y(_1876_));
 sg13g2_nor2_2 _2600_ (.A(net65),
    .B(_1844_),
    .Y(_0205_));
 sg13g2_nor2_1 _2601_ (.A(_0205_),
    .B(net35),
    .Y(_1877_));
 sg13g2_inv_4 _2602_ (.A(net37),
    .Y(_1878_));
 sg13g2_nand2_1 _2603_ (.Y(_1879_),
    .A(_1830_),
    .B(_1846_));
 sg13g2_buf_1 _2604_ (.A(_1879_),
    .X(_1880_));
 sg13g2_nand3_1 _2605_ (.B(net34),
    .C(net33),
    .A(_1877_),
    .Y(_1881_));
 sg13g2_nor2_1 _2606_ (.A(_1844_),
    .B(net33),
    .Y(_1882_));
 sg13g2_nand3_1 _2607_ (.B(_1882_),
    .C(net35),
    .A(net34),
    .Y(_1883_));
 sg13g2_nand3_1 _2608_ (.B(_1881_),
    .C(_1883_),
    .A(_1876_),
    .Y(_1884_));
 sg13g2_nor2_1 _2609_ (.A(_1557_),
    .B(_1821_),
    .Y(_1885_));
 sg13g2_inv_1 _2610_ (.Y(_1886_),
    .A(_1885_));
 sg13g2_nand2_1 _2611_ (.Y(_1887_),
    .A(_1803_),
    .B(_1836_));
 sg13g2_inv_1 _2612_ (.Y(_1888_),
    .A(_1866_));
 sg13g2_nand2_1 _2613_ (.Y(_1889_),
    .A(_1866_),
    .B(\vga.score_r[4] ));
 sg13g2_o21ai_1 _2614_ (.B1(_1889_),
    .Y(_1890_),
    .A1(_1885_),
    .A2(_1831_));
 sg13g2_a21oi_1 _2615_ (.A1(_1821_),
    .A2(_1888_),
    .Y(_1891_),
    .B1(_1890_));
 sg13g2_nor2_1 _2616_ (.A(_1891_),
    .B(_1887_),
    .Y(_1892_));
 sg13g2_a21oi_1 _2617_ (.A1(_1886_),
    .A2(_1887_),
    .Y(_1893_),
    .B1(_1892_));
 sg13g2_a21oi_1 _2618_ (.A1(_1845_),
    .A2(_1886_),
    .Y(_1894_),
    .B1(_1620_));
 sg13g2_o21ai_1 _2619_ (.B1(_1894_),
    .Y(_1895_),
    .A1(_1845_),
    .A2(_1893_));
 sg13g2_buf_2 _2620_ (.A(_1895_),
    .X(_1896_));
 sg13g2_nand2_1 _2621_ (.Y(_1897_),
    .A(_0205_),
    .B(net33));
 sg13g2_nor2_1 _2622_ (.A(_1863_),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_inv_2 _2623_ (.Y(_1899_),
    .A(_1898_));
 sg13g2_nor3_1 _2624_ (.A(_1896_),
    .B(net37),
    .C(_1899_),
    .Y(_1900_));
 sg13g2_a21oi_1 _2625_ (.A1(_1884_),
    .A2(_1896_),
    .Y(_0006_),
    .B1(_1900_));
 sg13g2_inv_2 _2626_ (.Y(_0209_),
    .A(_1896_));
 sg13g2_nor2_1 _2627_ (.A(_0209_),
    .B(_1883_),
    .Y(_1901_));
 sg13g2_nor2_1 _2628_ (.A(net37),
    .B(_1898_),
    .Y(_1902_));
 sg13g2_nand3_1 _2629_ (.B(_1843_),
    .C(_1618_),
    .A(_1842_),
    .Y(_1903_));
 sg13g2_nor3_1 _2630_ (.A(_1903_),
    .B(net33),
    .C(_1863_),
    .Y(_1904_));
 sg13g2_o21ai_1 _2631_ (.B1(_1896_),
    .Y(_1905_),
    .A1(net34),
    .A2(_1904_));
 sg13g2_nor2_1 _2632_ (.A(_1902_),
    .B(_1905_),
    .Y(_0086_));
 sg13g2_nor3_1 _2633_ (.A(_1900_),
    .B(_1901_),
    .C(_0086_),
    .Y(_0007_));
 sg13g2_nor2_1 _2634_ (.A(_0198_),
    .B(_1639_),
    .Y(_1906_));
 sg13g2_a21oi_1 _2635_ (.A1(_1906_),
    .A2(_0199_),
    .Y(_1907_),
    .B1(net38));
 sg13g2_nor2_2 _2636_ (.A(_1632_),
    .B(_1638_),
    .Y(_1908_));
 sg13g2_inv_2 _2637_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_nand2_1 _2638_ (.Y(_1910_),
    .A(_1909_),
    .B(_0198_));
 sg13g2_nand2_1 _2639_ (.Y(_1911_),
    .A(_1662_),
    .B(_1623_));
 sg13g2_nand3_1 _2640_ (.B(net29),
    .C(_1911_),
    .A(_1910_),
    .Y(_1912_));
 sg13g2_nand2_1 _2641_ (.Y(_1913_),
    .A(_1907_),
    .B(_1912_));
 sg13g2_nor2_1 _2642_ (.A(_1659_),
    .B(_1638_),
    .Y(_1914_));
 sg13g2_nand3_1 _2643_ (.B(_1623_),
    .C(_1914_),
    .A(_1654_),
    .Y(_1915_));
 sg13g2_nand2_1 _2644_ (.Y(_1916_),
    .A(_1915_),
    .B(net38));
 sg13g2_nand2_1 _2645_ (.Y(_0004_),
    .A(_1913_),
    .B(_1916_));
 sg13g2_a21oi_1 _2646_ (.A1(_1908_),
    .A2(_1623_),
    .Y(_1917_),
    .B1(_1653_));
 sg13g2_nor2_1 _2647_ (.A(net38),
    .B(_1917_),
    .Y(_1918_));
 sg13g2_a21oi_1 _2648_ (.A1(_1914_),
    .A2(_1623_),
    .Y(_1919_),
    .B1(_0199_));
 sg13g2_nand2_1 _2649_ (.Y(_1920_),
    .A(_1908_),
    .B(_0198_));
 sg13g2_nand2_1 _2650_ (.Y(_1921_),
    .A(_1919_),
    .B(_1920_));
 sg13g2_nor2_1 _2651_ (.A(_1673_),
    .B(_1915_),
    .Y(_1922_));
 sg13g2_a21oi_1 _2652_ (.A1(_1918_),
    .A2(_1921_),
    .Y(_0005_),
    .B1(_1922_));
 sg13g2_nand2_1 _2653_ (.Y(_1923_),
    .A(_1848_),
    .B(net35));
 sg13g2_nand2_1 _2654_ (.Y(_1924_),
    .A(_1923_),
    .B(net37));
 sg13g2_nand3_1 _2655_ (.B(_1847_),
    .C(_0207_),
    .A(_1897_),
    .Y(_1925_));
 sg13g2_nand2_1 _2656_ (.Y(_1926_),
    .A(_1925_),
    .B(net34));
 sg13g2_o21ai_1 _2657_ (.B1(_1926_),
    .Y(_1927_),
    .A1(_1898_),
    .A2(_1924_));
 sg13g2_nand2_1 _2658_ (.Y(_1928_),
    .A(_1927_),
    .B(_1896_));
 sg13g2_nand3_1 _2659_ (.B(_1877_),
    .C(net34),
    .A(_0209_),
    .Y(_1929_));
 sg13g2_nand2_1 _2660_ (.Y(_0012_),
    .A(_1928_),
    .B(_1929_));
 sg13g2_nand3_1 _2661_ (.B(_1899_),
    .C(_1878_),
    .A(_1925_),
    .Y(_1930_));
 sg13g2_nand2_1 _2662_ (.Y(_1931_),
    .A(_1864_),
    .B(_0205_));
 sg13g2_nand3_1 _2663_ (.B(net37),
    .C(_1931_),
    .A(_1923_),
    .Y(_1932_));
 sg13g2_nand2_1 _2664_ (.Y(_1933_),
    .A(_1930_),
    .B(_1932_));
 sg13g2_nand2_1 _2665_ (.Y(_1934_),
    .A(_1933_),
    .B(_1896_));
 sg13g2_nand2_1 _2666_ (.Y(_0013_),
    .A(_1934_),
    .B(_1929_));
 sg13g2_a21oi_1 _2667_ (.A1(_0205_),
    .A2(net33),
    .Y(_1935_),
    .B1(net35));
 sg13g2_a21oi_1 _2668_ (.A1(_1882_),
    .A2(_0208_),
    .Y(_1936_),
    .B1(_0209_));
 sg13g2_o21ai_1 _2669_ (.B1(_1936_),
    .Y(_1937_),
    .A1(_1935_),
    .A2(_1926_));
 sg13g2_nand2_1 _2670_ (.Y(_1938_),
    .A(_1881_),
    .B(_0209_));
 sg13g2_nand2_1 _2671_ (.Y(_0002_),
    .A(_1937_),
    .B(_1938_));
 sg13g2_nand3_1 _2672_ (.B(net35),
    .C(net33),
    .A(_1896_),
    .Y(_1939_));
 sg13g2_nand2_1 _2673_ (.Y(_1940_),
    .A(_1905_),
    .B(_1939_));
 sg13g2_nand2_1 _2674_ (.Y(_1941_),
    .A(net33),
    .B(_1903_));
 sg13g2_o21ai_1 _2675_ (.B1(_1941_),
    .Y(_1942_),
    .A1(_1864_),
    .A2(_1882_));
 sg13g2_nand2_1 _2676_ (.Y(_1943_),
    .A(_1942_),
    .B(net34));
 sg13g2_a21oi_1 _2677_ (.A1(_1940_),
    .A2(_1943_),
    .Y(_0003_),
    .B1(_1900_));
 sg13g2_nand2_1 _2678_ (.Y(_1944_),
    .A(_1639_),
    .B(_0198_));
 sg13g2_nand2_1 _2679_ (.Y(_1945_),
    .A(net29),
    .B(_1914_));
 sg13g2_nand2_1 _2680_ (.Y(_1946_),
    .A(_1945_),
    .B(_1673_));
 sg13g2_a21oi_1 _2681_ (.A1(net29),
    .A2(_1944_),
    .Y(_1947_),
    .B1(_1946_));
 sg13g2_nor2_1 _2682_ (.A(net29),
    .B(_1640_),
    .Y(_1948_));
 sg13g2_nand2_1 _2683_ (.Y(_1949_),
    .A(_1914_),
    .B(_1623_));
 sg13g2_nand2_1 _2684_ (.Y(_1950_),
    .A(_1948_),
    .B(_1949_));
 sg13g2_a21oi_1 _2685_ (.A1(_1947_),
    .A2(_1950_),
    .Y(_0010_),
    .B1(_1674_));
 sg13g2_nand2_1 _2686_ (.Y(_1951_),
    .A(_1944_),
    .B(_1655_));
 sg13g2_a21oi_1 _2687_ (.A1(_1951_),
    .A2(_0199_),
    .Y(_1952_),
    .B1(net38));
 sg13g2_nand2_1 _2688_ (.Y(_1953_),
    .A(_1663_),
    .B(_0198_));
 sg13g2_nand3_1 _2689_ (.B(_1953_),
    .C(_1920_),
    .A(_1919_),
    .Y(_1954_));
 sg13g2_a21oi_1 _2690_ (.A1(_1952_),
    .A2(_1954_),
    .Y(_0011_),
    .B1(_1674_));
 sg13g2_a21oi_1 _2691_ (.A1(_1659_),
    .A2(net38),
    .Y(_1955_),
    .B1(_1674_));
 sg13g2_a21oi_1 _2692_ (.A1(_0199_),
    .A2(_1908_),
    .Y(_1956_),
    .B1(net38));
 sg13g2_nand2_1 _2693_ (.Y(_1957_),
    .A(_1640_),
    .B(net29));
 sg13g2_nand3_1 _2694_ (.B(_1957_),
    .C(_1945_),
    .A(_1956_),
    .Y(_1958_));
 sg13g2_nand2_1 _2695_ (.Y(_0000_),
    .A(_1955_),
    .B(_1958_));
 sg13g2_nand3_1 _2696_ (.B(net29),
    .C(_1909_),
    .A(_1911_),
    .Y(_1959_));
 sg13g2_nand2_1 _2697_ (.Y(_1960_),
    .A(_1908_),
    .B(_1623_));
 sg13g2_nand2_1 _2698_ (.Y(_1961_),
    .A(_0198_),
    .B(_1632_));
 sg13g2_nand3_1 _2699_ (.B(_1961_),
    .C(_0199_),
    .A(_1960_),
    .Y(_1962_));
 sg13g2_nand2_1 _2700_ (.Y(_1963_),
    .A(_1959_),
    .B(_1962_));
 sg13g2_nand2_1 _2701_ (.Y(_1964_),
    .A(_1963_),
    .B(_1673_));
 sg13g2_nand2_1 _2702_ (.Y(_0001_),
    .A(_1964_),
    .B(_1916_));
 sg13g2_nand3_1 _2703_ (.B(_1880_),
    .C(_1903_),
    .A(net35),
    .Y(_1965_));
 sg13g2_inv_1 _2704_ (.Y(_1966_),
    .A(_1877_));
 sg13g2_a21oi_1 _2705_ (.A1(_1965_),
    .A2(_1966_),
    .Y(_1967_),
    .B1(net34));
 sg13g2_a21oi_1 _2706_ (.A1(_1923_),
    .A2(_1966_),
    .Y(_1968_),
    .B1(net37));
 sg13g2_o21ai_1 _2707_ (.B1(_1896_),
    .Y(_1969_),
    .A1(_1967_),
    .A2(_1968_));
 sg13g2_nand2_1 _2708_ (.Y(_0009_),
    .A(_1969_),
    .B(_1929_));
 sg13g2_buf_1 _2709_ (.A(\vga.count_v[1] ),
    .X(_1970_));
 sg13g2_buf_1 _2710_ (.A(\vga.count_v[0] ),
    .X(_1971_));
 sg13g2_nor2_1 _2711_ (.A(net78),
    .B(net77),
    .Y(_1972_));
 sg13g2_inv_1 _2712_ (.Y(_1973_),
    .A(_1972_));
 sg13g2_buf_2 _2713_ (.A(\vga.count_v[9] ),
    .X(_1974_));
 sg13g2_nor2_1 _2714_ (.A(_1974_),
    .B(\vga.count_v[8] ),
    .Y(_1975_));
 sg13g2_inv_1 _2715_ (.Y(_1976_),
    .A(_1975_));
 sg13g2_buf_1 _2716_ (.A(\vga.count_v[2] ),
    .X(_1977_));
 sg13g2_buf_1 _2717_ (.A(\vga.count_v[3] ),
    .X(_1978_));
 sg13g2_nand2_1 _2718_ (.Y(_1979_),
    .A(net76),
    .B(net75));
 sg13g2_buf_1 _2719_ (.A(\vga.count_v[5] ),
    .X(_1980_));
 sg13g2_buf_1 _2720_ (.A(\vga.count_v[4] ),
    .X(_1981_));
 sg13g2_inv_1 _2721_ (.Y(_1982_),
    .A(net73));
 sg13g2_buf_2 _2722_ (.A(\vga.count_v[7] ),
    .X(_1983_));
 sg13g2_buf_1 _2723_ (.A(\vga.count_v[6] ),
    .X(_1984_));
 sg13g2_nor2_1 _2724_ (.A(_1983_),
    .B(_1984_),
    .Y(_1985_));
 sg13g2_inv_1 _2725_ (.Y(_1986_),
    .A(_1985_));
 sg13g2_nor3_1 _2726_ (.A(net74),
    .B(_1982_),
    .C(_1986_),
    .Y(_1987_));
 sg13g2_inv_1 _2727_ (.Y(_1988_),
    .A(_1987_));
 sg13g2_nor4_1 _2728_ (.A(_1973_),
    .B(net56),
    .C(_1979_),
    .D(_1988_),
    .Y(_1989_));
 sg13g2_buf_2 _2729_ (.A(_1989_),
    .X(_1990_));
 sg13g2_nor2_1 _2730_ (.A(net76),
    .B(net75),
    .Y(_1991_));
 sg13g2_inv_1 _2731_ (.Y(_1992_),
    .A(_1991_));
 sg13g2_nand2_1 _2732_ (.Y(_1993_),
    .A(net74),
    .B(net73));
 sg13g2_nor2_1 _2733_ (.A(_1993_),
    .B(_1986_),
    .Y(_1994_));
 sg13g2_inv_1 _2734_ (.Y(_1995_),
    .A(_1994_));
 sg13g2_nor4_1 _2735_ (.A(_1973_),
    .B(net56),
    .C(_1992_),
    .D(_1995_),
    .Y(_1996_));
 sg13g2_buf_2 _2736_ (.A(_1996_),
    .X(_1997_));
 sg13g2_nor2b_1 _2737_ (.A(_1997_),
    .B_N(_0015_),
    .Y(_1998_));
 sg13g2_a21oi_1 _2738_ (.A1(_0028_),
    .A2(_1997_),
    .Y(_1999_),
    .B1(_1998_));
 sg13g2_nand2_1 _2739_ (.Y(_2000_),
    .A(_1990_),
    .B(_0018_));
 sg13g2_o21ai_1 _2740_ (.B1(_2000_),
    .Y(_2001_),
    .A1(_1990_),
    .A2(_1999_));
 sg13g2_inv_1 _2741_ (.Y(_2002_),
    .A(net78));
 sg13g2_nor2_1 _2742_ (.A(net77),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_inv_1 _2743_ (.Y(_2004_),
    .A(net76));
 sg13g2_nand3_1 _2744_ (.B(_2004_),
    .C(net75),
    .A(_2003_),
    .Y(_2005_));
 sg13g2_nor3_1 _2745_ (.A(net56),
    .B(_1995_),
    .C(_2005_),
    .Y(_2006_));
 sg13g2_nor3_1 _2746_ (.A(_1997_),
    .B(_2006_),
    .C(_1990_),
    .Y(_2007_));
 sg13g2_inv_2 _2747_ (.Y(_2008_),
    .A(_2003_));
 sg13g2_nor2_1 _2748_ (.A(net75),
    .B(_2004_),
    .Y(_2009_));
 sg13g2_inv_1 _2749_ (.Y(_2010_),
    .A(_2009_));
 sg13g2_inv_2 _2750_ (.Y(_2011_),
    .A(net74));
 sg13g2_nor2_1 _2751_ (.A(net73),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_inv_1 _2752_ (.Y(_2013_),
    .A(_2012_));
 sg13g2_nor2_1 _2753_ (.A(_1986_),
    .B(_1976_),
    .Y(_2014_));
 sg13g2_inv_1 _2754_ (.Y(_2015_),
    .A(_2014_));
 sg13g2_nor4_2 _2755_ (.A(_2008_),
    .B(_2010_),
    .C(_2013_),
    .Y(_2016_),
    .D(_2015_));
 sg13g2_nor4_2 _2756_ (.A(net56),
    .B(_2008_),
    .C(_1992_),
    .Y(_2017_),
    .D(_1988_));
 sg13g2_nor2_1 _2757_ (.A(_2016_),
    .B(_2017_),
    .Y(_2018_));
 sg13g2_nand2_1 _2758_ (.Y(_2019_),
    .A(_2007_),
    .B(_2018_));
 sg13g2_buf_2 _2759_ (.A(_2019_),
    .X(_2020_));
 sg13g2_mux2_1 _2760_ (.A0(\vga.score_l_unit_pixels[0] ),
    .A1(_2001_),
    .S(_2020_),
    .X(_0202_));
 sg13g2_inv_1 _2761_ (.Y(_2021_),
    .A(\vga.score_l_unit_pixels[1] ));
 sg13g2_inv_1 _2762_ (.Y(_2022_),
    .A(_2020_));
 sg13g2_a21oi_1 _2763_ (.A1(_0014_),
    .A2(_2017_),
    .Y(_0217_),
    .B1(_2022_));
 sg13g2_inv_1 _2764_ (.Y(_0218_),
    .A(_0019_));
 sg13g2_nor4_2 _2765_ (.A(_1973_),
    .B(net56),
    .C(_1992_),
    .Y(_0219_),
    .D(_1995_));
 sg13g2_nor4_2 _2766_ (.A(_1973_),
    .B(net56),
    .C(_1979_),
    .Y(_0220_),
    .D(_1988_));
 sg13g2_or2_1 _2767_ (.X(_0221_),
    .B(_0220_),
    .A(_0219_));
 sg13g2_inv_1 _2768_ (.Y(_0222_),
    .A(_1990_));
 sg13g2_nor4_2 _2769_ (.A(_2008_),
    .B(_2010_),
    .C(_2013_),
    .Y(_0223_),
    .D(_2015_));
 sg13g2_inv_1 _2770_ (.Y(_0224_),
    .A(_0223_));
 sg13g2_nor2_2 _2771_ (.A(_0219_),
    .B(_0223_),
    .Y(_0225_));
 sg13g2_nand2b_1 _2772_ (.Y(_0226_),
    .B(_0225_),
    .A_N(_0032_));
 sg13g2_o21ai_1 _2773_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0024_),
    .A2(_0224_));
 sg13g2_a22oi_1 _2774_ (.Y(_0228_),
    .B1(_0222_),
    .B2(_0227_),
    .A2(_0221_),
    .A1(_0218_));
 sg13g2_inv_1 _2775_ (.Y(_0229_),
    .A(_2017_));
 sg13g2_nand2_1 _2776_ (.Y(_0230_),
    .A(_0228_),
    .B(_0229_));
 sg13g2_a22oi_1 _2777_ (.Y(_0203_),
    .B1(_0217_),
    .B2(_0230_),
    .A2(_2022_),
    .A1(_2021_));
 sg13g2_inv_1 _2778_ (.Y(_0231_),
    .A(_0020_));
 sg13g2_nor4_1 _2779_ (.A(net56),
    .B(_2008_),
    .C(_1992_),
    .D(_1988_),
    .Y(_0232_));
 sg13g2_a21oi_1 _2780_ (.A1(_0220_),
    .A2(_0231_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_a22oi_1 _2781_ (.Y(_0234_),
    .B1(_0033_),
    .B2(_0225_),
    .A2(_1997_),
    .A1(_0029_));
 sg13g2_a21oi_1 _2782_ (.A1(_0025_),
    .A2(_2016_),
    .Y(_0235_),
    .B1(_1990_));
 sg13g2_nand2_1 _2783_ (.Y(_0236_),
    .A(_0234_),
    .B(_0235_));
 sg13g2_a22oi_1 _2784_ (.Y(_0237_),
    .B1(_0233_),
    .B2(_0236_),
    .A2(_2017_),
    .A1(_0015_));
 sg13g2_nor2_1 _2785_ (.A(\vga.score_l_unit_pixels[2] ),
    .B(_2020_),
    .Y(_0238_));
 sg13g2_a21oi_1 _2786_ (.A1(_0237_),
    .A2(_2020_),
    .Y(_0204_),
    .B1(_0238_));
 sg13g2_inv_1 _2787_ (.Y(_0239_),
    .A(\vga.score_r_unit_pixels[0] ));
 sg13g2_nor2b_1 _2788_ (.A(_1997_),
    .B_N(_0017_),
    .Y(_0240_));
 sg13g2_a21oi_1 _2789_ (.A1(_0030_),
    .A2(_1997_),
    .Y(_0241_),
    .B1(_0240_));
 sg13g2_nand2_1 _2790_ (.Y(_0242_),
    .A(_1990_),
    .B(_0021_));
 sg13g2_o21ai_1 _2791_ (.B1(_0242_),
    .Y(_0243_),
    .A1(_1990_),
    .A2(_0241_));
 sg13g2_nand2_1 _2792_ (.Y(_0244_),
    .A(_0243_),
    .B(_2020_));
 sg13g2_o21ai_1 _2793_ (.B1(_0244_),
    .Y(_0211_),
    .A1(_0239_),
    .A2(_2020_));
 sg13g2_inv_1 _2794_ (.Y(_0245_),
    .A(\vga.score_r_unit_pixels[1] ));
 sg13g2_a21oi_1 _2795_ (.A1(_0016_),
    .A2(_2017_),
    .Y(_0246_),
    .B1(_2022_));
 sg13g2_inv_1 _2796_ (.Y(_0247_),
    .A(_0022_));
 sg13g2_nand2b_1 _2797_ (.Y(_0248_),
    .B(_0225_),
    .A_N(_0034_));
 sg13g2_o21ai_1 _2798_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0026_),
    .A2(_0224_));
 sg13g2_a22oi_1 _2799_ (.Y(_0250_),
    .B1(_0222_),
    .B2(_0249_),
    .A2(_0221_),
    .A1(_0247_));
 sg13g2_nand2_1 _2800_ (.Y(_0251_),
    .A(_0250_),
    .B(_0229_));
 sg13g2_a22oi_1 _2801_ (.Y(_0212_),
    .B1(_0246_),
    .B2(_0251_),
    .A2(_2022_),
    .A1(_0245_));
 sg13g2_inv_1 _2802_ (.Y(_0252_),
    .A(_0023_));
 sg13g2_a21oi_1 _2803_ (.A1(_0220_),
    .A2(_0252_),
    .Y(_0253_),
    .B1(_0232_));
 sg13g2_a21oi_1 _2804_ (.A1(_0225_),
    .A2(_0035_),
    .Y(_0254_),
    .B1(_1990_));
 sg13g2_a22oi_1 _2805_ (.Y(_0255_),
    .B1(_0027_),
    .B2(_2016_),
    .A2(_0031_),
    .A1(_1997_));
 sg13g2_nand2_1 _2806_ (.Y(_0256_),
    .A(_0254_),
    .B(_0255_));
 sg13g2_a22oi_1 _2807_ (.Y(_0257_),
    .B1(_0253_),
    .B2(_0256_),
    .A2(_2017_),
    .A1(_0017_));
 sg13g2_nor2_1 _2808_ (.A(\vga.score_r_unit_pixels[2] ),
    .B(_2020_),
    .Y(_0258_));
 sg13g2_a21oi_1 _2809_ (.A1(_0257_),
    .A2(_2020_),
    .Y(_0213_),
    .B1(_0258_));
 sg13g2_inv_1 _2810_ (.Y(_0259_),
    .A(\vga.left_down_1d ));
 sg13g2_nand2_1 _2811_ (.Y(_0260_),
    .A(net50),
    .B(net2));
 sg13g2_o21ai_1 _2812_ (.B1(_0260_),
    .Y(_0169_),
    .A1(_0259_),
    .A2(net50));
 sg13g2_inv_1 _2813_ (.Y(_0261_),
    .A(\vga.left_up_1d ));
 sg13g2_nand2_1 _2814_ (.Y(_0262_),
    .A(net50),
    .B(net1));
 sg13g2_o21ai_1 _2815_ (.B1(_0262_),
    .Y(_0171_),
    .A1(_0261_),
    .A2(net50));
 sg13g2_inv_1 _2816_ (.Y(_0263_),
    .A(\vga.right_down_1d ));
 sg13g2_nand2_1 _2817_ (.Y(_0264_),
    .A(_1650_),
    .B(net4));
 sg13g2_o21ai_1 _2818_ (.B1(_0264_),
    .Y(_0192_),
    .A1(_0263_),
    .A2(_1650_));
 sg13g2_inv_1 _2819_ (.Y(_0265_),
    .A(\vga.right_up_1d ));
 sg13g2_nand2_1 _2820_ (.Y(_0266_),
    .A(net50),
    .B(net3));
 sg13g2_o21ai_1 _2821_ (.B1(_0266_),
    .Y(_0194_),
    .A1(_0265_),
    .A2(net50));
 sg13g2_o21ai_1 _2822_ (.B1(_1905_),
    .Y(_0267_),
    .A1(_0209_),
    .A2(_1965_));
 sg13g2_o21ai_1 _2823_ (.B1(_1902_),
    .Y(_0268_),
    .A1(net35),
    .A2(_1847_));
 sg13g2_nand2_1 _2824_ (.Y(_0085_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_inv_1 _2825_ (.Y(_0087_),
    .A(_0086_));
 sg13g2_inv_1 _2826_ (.Y(_0269_),
    .A(_1919_));
 sg13g2_nand2_1 _2827_ (.Y(_0088_),
    .A(_1918_),
    .B(_0269_));
 sg13g2_a21oi_1 _2828_ (.A1(_1917_),
    .A2(_1953_),
    .Y(_0270_),
    .B1(_0200_));
 sg13g2_o21ai_1 _2829_ (.B1(_0270_),
    .Y(_0089_),
    .A1(_1906_),
    .A2(_0269_));
 sg13g2_inv_2 _2830_ (.Y(_0090_),
    .A(_0088_));
 sg13g2_a21oi_1 _2831_ (.A1(_1953_),
    .A2(_1654_),
    .Y(_0271_),
    .B1(_1948_));
 sg13g2_nand2_1 _2832_ (.Y(_0091_),
    .A(_0271_),
    .B(_1673_));
 sg13g2_a21oi_1 _2833_ (.A1(_1965_),
    .A2(net34),
    .Y(_0272_),
    .B1(_0209_));
 sg13g2_nand2_1 _2834_ (.Y(_0092_),
    .A(_0272_),
    .B(_1924_));
 sg13g2_buf_1 _2835_ (.A(net65),
    .X(_0273_));
 sg13g2_buf_1 _2836_ (.A(net55),
    .X(_0274_));
 sg13g2_buf_1 _2837_ (.A(\vga.count_h[5] ),
    .X(_0275_));
 sg13g2_buf_2 _2838_ (.A(\vga.count_h[4] ),
    .X(_0276_));
 sg13g2_nand2_2 _2839_ (.Y(_0277_),
    .A(net72),
    .B(_0276_));
 sg13g2_buf_1 _2840_ (.A(\vga.count_h[7] ),
    .X(_0278_));
 sg13g2_buf_2 _2841_ (.A(\vga.count_h[6] ),
    .X(_0279_));
 sg13g2_inv_1 _2842_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nor2_1 _2843_ (.A(_0278_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_inv_1 _2844_ (.Y(_0282_),
    .A(_0281_));
 sg13g2_nor2_1 _2845_ (.A(_0277_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_buf_2 _2846_ (.A(\vga.count_h[8] ),
    .X(_0284_));
 sg13g2_buf_2 _2847_ (.A(\vga.count_h[9] ),
    .X(_0285_));
 sg13g2_inv_1 _2848_ (.Y(_0286_),
    .A(_0285_));
 sg13g2_nor2_2 _2849_ (.A(_0284_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nand2_1 _2850_ (.Y(_0288_),
    .A(_0283_),
    .B(_0287_));
 sg13g2_inv_1 _2851_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_buf_1 _2852_ (.A(\vga.count_h[0] ),
    .X(_0290_));
 sg13g2_buf_2 _2853_ (.A(\vga.count_h[1] ),
    .X(_0291_));
 sg13g2_nand2_1 _2854_ (.Y(_0292_),
    .A(_0290_),
    .B(_0291_));
 sg13g2_buf_2 _2855_ (.A(_0292_),
    .X(_0293_));
 sg13g2_buf_1 _2856_ (.A(\vga.count_h[2] ),
    .X(_0294_));
 sg13g2_buf_2 _2857_ (.A(\vga.count_h[3] ),
    .X(_0295_));
 sg13g2_nand2_2 _2858_ (.Y(_0296_),
    .A(_0294_),
    .B(_0295_));
 sg13g2_nor2_2 _2859_ (.A(_0293_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_inv_1 _2860_ (.Y(_0298_),
    .A(_0278_));
 sg13g2_a21oi_1 _2861_ (.A1(_0287_),
    .A2(_0298_),
    .Y(_0299_),
    .B1(_0066_));
 sg13g2_a21oi_1 _2862_ (.A1(_0289_),
    .A2(_0297_),
    .Y(_0300_),
    .B1(_0299_));
 sg13g2_inv_1 _2863_ (.Y(_0301_),
    .A(_0277_));
 sg13g2_nand2_1 _2864_ (.Y(_0302_),
    .A(_0278_),
    .B(_0279_));
 sg13g2_inv_1 _2865_ (.Y(_0303_),
    .A(_0302_));
 sg13g2_inv_1 _2866_ (.Y(_0304_),
    .A(_0287_));
 sg13g2_a21oi_1 _2867_ (.A1(_0301_),
    .A2(_0303_),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_inv_1 _2868_ (.Y(_0306_),
    .A(_0275_));
 sg13g2_nor2_1 _2869_ (.A(_0276_),
    .B(_0306_),
    .Y(_0307_));
 sg13g2_nand4_1 _2870_ (.B(_0287_),
    .C(_0303_),
    .A(_0297_),
    .Y(_0308_),
    .D(_0307_));
 sg13g2_o21ai_1 _2871_ (.B1(_0308_),
    .Y(_0309_),
    .A1(_0066_),
    .A2(_0305_));
 sg13g2_nor2_1 _2872_ (.A(\vga.count_h[5] ),
    .B(_0276_),
    .Y(_0310_));
 sg13g2_inv_1 _2873_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_nor3_1 _2874_ (.A(_0298_),
    .B(_0279_),
    .C(_0311_),
    .Y(_0312_));
 sg13g2_nand2_1 _2875_ (.Y(_0313_),
    .A(_0312_),
    .B(_0287_));
 sg13g2_nand2b_1 _2876_ (.Y(_0314_),
    .B(_0313_),
    .A_N(_0299_));
 sg13g2_o21ai_1 _2877_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0297_),
    .A2(_0313_));
 sg13g2_nor4_1 _2878_ (.A(net52),
    .B(_0300_),
    .C(_0309_),
    .D(_0315_),
    .Y(_0143_));
 sg13g2_buf_1 _2879_ (.A(ui_in[6]),
    .X(_0316_));
 sg13g2_inv_1 _2880_ (.Y(_0317_),
    .A(net5));
 sg13g2_inv_1 _2881_ (.Y(_0318_),
    .A(_1591_));
 sg13g2_inv_1 _2882_ (.Y(_0319_),
    .A(\vga.interval_counter[16] ));
 sg13g2_nand4_1 _2883_ (.B(_0319_),
    .C(_1590_),
    .A(_0318_),
    .Y(_0320_),
    .D(\vga.interval_counter[17] ));
 sg13g2_nand2_1 _2884_ (.Y(_0321_),
    .A(_1608_),
    .B(\vga.interval_counter[9] ));
 sg13g2_nand2_1 _2885_ (.Y(_0322_),
    .A(\vga.interval_counter[11] ),
    .B(\vga.interval_counter[10] ));
 sg13g2_nor2_1 _2886_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_inv_2 _2887_ (.Y(_0324_),
    .A(_1594_));
 sg13g2_nand4_1 _2888_ (.B(_1593_),
    .C(_0324_),
    .A(_0323_),
    .Y(_0325_),
    .D(_1595_));
 sg13g2_inv_1 _2889_ (.Y(_0326_),
    .A(_1600_));
 sg13g2_nor4_1 _2890_ (.A(_1604_),
    .B(_1610_),
    .C(_1603_),
    .D(_0326_),
    .Y(_0327_));
 sg13g2_inv_1 _2891_ (.Y(_0328_),
    .A(\vga.interval_counter[1] ));
 sg13g2_nand4_1 _2892_ (.B(_0328_),
    .C(_1599_),
    .A(_0327_),
    .Y(_0329_),
    .D(_1602_));
 sg13g2_nor4_1 _2893_ (.A(_0317_),
    .B(_0320_),
    .C(_0325_),
    .D(_0329_),
    .Y(_0330_));
 sg13g2_inv_1 _2894_ (.Y(_0331_),
    .A(\vga.interval_counter[17] ));
 sg13g2_nand2_1 _2895_ (.Y(_0332_),
    .A(_1604_),
    .B(_1591_));
 sg13g2_nand2_1 _2896_ (.Y(_0333_),
    .A(_1600_),
    .B(_1610_));
 sg13g2_nor4_1 _2897_ (.A(_0319_),
    .B(_0331_),
    .C(_0332_),
    .D(_0333_),
    .Y(_0334_));
 sg13g2_inv_1 _2898_ (.Y(_0335_),
    .A(\vga.interval_counter[10] ));
 sg13g2_nor2_1 _2899_ (.A(\vga.interval_counter[11] ),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_inv_1 _2900_ (.Y(_0337_),
    .A(_0336_));
 sg13g2_nor2_1 _2901_ (.A(_0321_),
    .B(_0337_),
    .Y(_0338_));
 sg13g2_nor3_1 _2902_ (.A(_1593_),
    .B(_0324_),
    .C(_1596_),
    .Y(_0339_));
 sg13g2_inv_1 _2903_ (.Y(_0340_),
    .A(\vga.interval_counter[12] ));
 sg13g2_nor4_1 _2904_ (.A(\vga.interval_counter[4] ),
    .B(_1590_),
    .C(_1601_),
    .D(_0340_),
    .Y(_0341_));
 sg13g2_nand4_1 _2905_ (.B(_0338_),
    .C(_0339_),
    .A(_0334_),
    .Y(_0342_),
    .D(_0341_));
 sg13g2_nor4_1 _2906_ (.A(net5),
    .B(_0328_),
    .C(_1599_),
    .D(_0342_),
    .Y(_0343_));
 sg13g2_nor3_1 _2907_ (.A(_0316_),
    .B(_0330_),
    .C(_0343_),
    .Y(_0344_));
 sg13g2_inv_1 _2908_ (.Y(_0345_),
    .A(_1593_));
 sg13g2_nand4_1 _2909_ (.B(_1592_),
    .C(_0345_),
    .A(_0336_),
    .Y(_0346_),
    .D(_0324_));
 sg13g2_inv_1 _2910_ (.Y(_0347_),
    .A(_1601_));
 sg13g2_nor2_1 _2911_ (.A(\vga.interval_counter[1] ),
    .B(_1599_),
    .Y(_0348_));
 sg13g2_nand3_1 _2912_ (.B(_0317_),
    .C(_1608_),
    .A(_0348_),
    .Y(_0349_));
 sg13g2_nor4_1 _2913_ (.A(\vga.interval_counter[9] ),
    .B(_0347_),
    .C(_0340_),
    .D(_0349_),
    .Y(_0350_));
 sg13g2_nand2_1 _2914_ (.Y(_0351_),
    .A(_0350_),
    .B(_0327_));
 sg13g2_nand4_1 _2915_ (.B(_1590_),
    .C(_1591_),
    .A(_1594_),
    .Y(_0352_),
    .D(_1610_));
 sg13g2_nor3_1 _2916_ (.A(_0317_),
    .B(_0345_),
    .C(_0352_),
    .Y(_0353_));
 sg13g2_nand3_1 _2917_ (.B(_0353_),
    .C(_0338_),
    .A(_1607_),
    .Y(_0354_));
 sg13g2_o21ai_1 _2918_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_0346_),
    .A2(_0351_));
 sg13g2_nor3_1 _2919_ (.A(_0319_),
    .B(\vga.interval_counter[17] ),
    .C(_1596_),
    .Y(_0356_));
 sg13g2_nand2_1 _2920_ (.Y(_0357_),
    .A(_0355_),
    .B(_0356_));
 sg13g2_nand2_1 _2921_ (.Y(_0358_),
    .A(_0357_),
    .B(_0316_));
 sg13g2_nand3b_1 _2922_ (.B(_1589_),
    .C(_0358_),
    .Y(_0359_),
    .A_N(_0344_));
 sg13g2_xnor2_1 _2923_ (.Y(_0360_),
    .A(_0316_),
    .B(\vga.speed_msb_1d ));
 sg13g2_o21ai_1 _2924_ (.B1(_1660_),
    .Y(_0361_),
    .A1(\vga.speed_lsb_1d ),
    .A2(_0317_));
 sg13g2_a21oi_1 _2925_ (.A1(_0317_),
    .A2(\vga.speed_lsb_1d ),
    .Y(_0362_),
    .B1(_0361_));
 sg13g2_nand3_1 _2926_ (.B(_0360_),
    .C(_0362_),
    .A(_0359_),
    .Y(_0363_));
 sg13g2_buf_1 _2927_ (.A(_0363_),
    .X(_0364_));
 sg13g2_buf_1 _2928_ (.A(_0364_),
    .X(_0365_));
 sg13g2_nor2b_1 _2929_ (.A(_0365_),
    .B_N(_0083_),
    .Y(_0144_));
 sg13g2_nand2_1 _2930_ (.Y(_0366_),
    .A(\vga.interval_counter[1] ),
    .B(_1599_));
 sg13g2_nor2_1 _2931_ (.A(_0324_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nand2_1 _2932_ (.Y(_0368_),
    .A(_0367_),
    .B(_1593_));
 sg13g2_nor2_1 _2933_ (.A(_1603_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_nand2_1 _2934_ (.Y(_0370_),
    .A(_0369_),
    .B(_1604_));
 sg13g2_nor2_1 _2935_ (.A(_0318_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nand2_1 _2936_ (.Y(_0372_),
    .A(_0371_),
    .B(_1590_));
 sg13g2_nor2_2 _2937_ (.A(_0321_),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nor2_1 _2938_ (.A(\vga.interval_counter[10] ),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_inv_4 _2939_ (.A(_0373_),
    .Y(_0375_));
 sg13g2_nor2_1 _2940_ (.A(_0335_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_nor3_1 _2941_ (.A(_0374_),
    .B(_0376_),
    .C(net42),
    .Y(_0145_));
 sg13g2_nor2_1 _2942_ (.A(\vga.interval_counter[11] ),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nor2_1 _2943_ (.A(_0322_),
    .B(_0375_),
    .Y(_0378_));
 sg13g2_nor3_1 _2944_ (.A(_0377_),
    .B(_0378_),
    .C(net42),
    .Y(_0146_));
 sg13g2_nor3_1 _2945_ (.A(_0340_),
    .B(_0322_),
    .C(_0375_),
    .Y(_0379_));
 sg13g2_nor2_1 _2946_ (.A(\vga.interval_counter[12] ),
    .B(_0378_),
    .Y(_0380_));
 sg13g2_nor3_1 _2947_ (.A(_0379_),
    .B(_0380_),
    .C(net42),
    .Y(_0147_));
 sg13g2_nor2_1 _2948_ (.A(_1601_),
    .B(_0379_),
    .Y(_0381_));
 sg13g2_nand2_1 _2949_ (.Y(_0382_),
    .A(_0379_),
    .B(_1601_));
 sg13g2_inv_2 _2950_ (.Y(_0383_),
    .A(_0382_));
 sg13g2_nor3_1 _2951_ (.A(_0381_),
    .B(_0383_),
    .C(_0365_),
    .Y(_0148_));
 sg13g2_nor2_1 _2952_ (.A(_1610_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_nand2_2 _2953_ (.Y(_0385_),
    .A(_0383_),
    .B(_1610_));
 sg13g2_inv_4 _2954_ (.A(_0385_),
    .Y(_0386_));
 sg13g2_nor3_1 _2955_ (.A(_0384_),
    .B(_0386_),
    .C(net42),
    .Y(_0149_));
 sg13g2_nand2_1 _2956_ (.Y(_0387_),
    .A(_0386_),
    .B(_0326_));
 sg13g2_nand2_1 _2957_ (.Y(_0388_),
    .A(_0385_),
    .B(_1600_));
 sg13g2_a21oi_1 _2958_ (.A1(_0387_),
    .A2(_0388_),
    .Y(_0150_),
    .B1(net42));
 sg13g2_nor2_1 _2959_ (.A(_0326_),
    .B(_0385_),
    .Y(_0389_));
 sg13g2_inv_1 _2960_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_nand2_1 _2961_ (.Y(_0391_),
    .A(_1600_),
    .B(\vga.interval_counter[16] ));
 sg13g2_nand2b_1 _2962_ (.Y(_0392_),
    .B(_0386_),
    .A_N(_0391_));
 sg13g2_nand2b_1 _2963_ (.Y(_0393_),
    .B(_0392_),
    .A_N(_0364_));
 sg13g2_a21oi_1 _2964_ (.A1(_0319_),
    .A2(_0390_),
    .Y(_0151_),
    .B1(_0393_));
 sg13g2_nor2_1 _2965_ (.A(_0331_),
    .B(_0391_),
    .Y(_0394_));
 sg13g2_buf_1 _2966_ (.A(_0364_),
    .X(_0395_));
 sg13g2_a221oi_1 _2967_ (.B2(_0386_),
    .C1(net41),
    .B1(_0394_),
    .A1(_0331_),
    .Y(_0152_),
    .A2(_0392_));
 sg13g2_a21oi_1 _2968_ (.A1(_0386_),
    .A2(_0394_),
    .Y(_0396_),
    .B1(\vga.interval_counter[18] ));
 sg13g2_and3_1 _2969_ (.X(_0397_),
    .A(_0386_),
    .B(\vga.interval_counter[18] ),
    .C(_0394_));
 sg13g2_buf_1 _2970_ (.A(_0397_),
    .X(_0398_));
 sg13g2_nor3_1 _2971_ (.A(_0396_),
    .B(_0398_),
    .C(net42),
    .Y(_0153_));
 sg13g2_nor2_1 _2972_ (.A(\vga.interval_counter[19] ),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_nand2_1 _2973_ (.Y(_0400_),
    .A(_0398_),
    .B(\vga.interval_counter[19] ));
 sg13g2_inv_2 _2974_ (.Y(_0401_),
    .A(_0400_));
 sg13g2_nor3_1 _2975_ (.A(net41),
    .B(_0399_),
    .C(_0401_),
    .Y(_0154_));
 sg13g2_inv_1 _2976_ (.Y(_0402_),
    .A(_0366_));
 sg13g2_nor3_1 _2977_ (.A(_0348_),
    .B(_0402_),
    .C(net42),
    .Y(_0155_));
 sg13g2_nor2_1 _2978_ (.A(\vga.interval_counter[20] ),
    .B(_0401_),
    .Y(_0403_));
 sg13g2_nand2_1 _2979_ (.Y(_0404_),
    .A(_0401_),
    .B(\vga.interval_counter[20] ));
 sg13g2_inv_2 _2980_ (.Y(_0405_),
    .A(_0404_));
 sg13g2_nor3_1 _2981_ (.A(net41),
    .B(_0403_),
    .C(_0405_),
    .Y(_0156_));
 sg13g2_nor2_1 _2982_ (.A(\vga.interval_counter[21] ),
    .B(_0405_),
    .Y(_0406_));
 sg13g2_nand2_1 _2983_ (.Y(_0407_),
    .A(_0405_),
    .B(\vga.interval_counter[21] ));
 sg13g2_inv_1 _2984_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nor3_1 _2985_ (.A(_0364_),
    .B(_0406_),
    .C(_0408_),
    .Y(_0157_));
 sg13g2_nor2_1 _2986_ (.A(_1586_),
    .B(_0407_),
    .Y(_0409_));
 sg13g2_nor2_1 _2987_ (.A(\vga.interval_counter[22] ),
    .B(_0408_),
    .Y(_0410_));
 sg13g2_nor3_1 _2988_ (.A(_0364_),
    .B(_0409_),
    .C(_0410_),
    .Y(_0158_));
 sg13g2_nor3_1 _2989_ (.A(_1585_),
    .B(_1586_),
    .C(_0407_),
    .Y(_0411_));
 sg13g2_nor2_1 _2990_ (.A(\vga.interval_counter[23] ),
    .B(_0409_),
    .Y(_0412_));
 sg13g2_nor3_1 _2991_ (.A(_0364_),
    .B(_0411_),
    .C(_0412_),
    .Y(_0159_));
 sg13g2_nor2_1 _2992_ (.A(\vga.interval_counter[24] ),
    .B(_0411_),
    .Y(_0413_));
 sg13g2_nor2b_1 _2993_ (.A(_1587_),
    .B_N(_0411_),
    .Y(_0414_));
 sg13g2_nor3_1 _2994_ (.A(_0364_),
    .B(_0413_),
    .C(_0414_),
    .Y(_0160_));
 sg13g2_nor2_1 _2995_ (.A(_1594_),
    .B(_0402_),
    .Y(_0415_));
 sg13g2_nor3_1 _2996_ (.A(_0367_),
    .B(_0415_),
    .C(net42),
    .Y(_0161_));
 sg13g2_inv_1 _2997_ (.Y(_0416_),
    .A(_0368_));
 sg13g2_nor2_1 _2998_ (.A(_1593_),
    .B(_0367_),
    .Y(_0417_));
 sg13g2_nor3_1 _2999_ (.A(_0416_),
    .B(_0417_),
    .C(net41),
    .Y(_0162_));
 sg13g2_nor2_1 _3000_ (.A(\vga.interval_counter[4] ),
    .B(_0416_),
    .Y(_0418_));
 sg13g2_nor3_1 _3001_ (.A(_0369_),
    .B(_0418_),
    .C(net41),
    .Y(_0163_));
 sg13g2_inv_1 _3002_ (.Y(_0419_),
    .A(_0370_));
 sg13g2_nor2_1 _3003_ (.A(_1604_),
    .B(_0369_),
    .Y(_0420_));
 sg13g2_nor3_1 _3004_ (.A(_0419_),
    .B(_0420_),
    .C(net41),
    .Y(_0164_));
 sg13g2_nor2_1 _3005_ (.A(_1591_),
    .B(_0419_),
    .Y(_0421_));
 sg13g2_nor3_1 _3006_ (.A(_0371_),
    .B(_0421_),
    .C(net41),
    .Y(_0165_));
 sg13g2_inv_1 _3007_ (.Y(_0422_),
    .A(_0372_));
 sg13g2_nor2_1 _3008_ (.A(_1590_),
    .B(_0371_),
    .Y(_0423_));
 sg13g2_nor3_1 _3009_ (.A(_0422_),
    .B(_0423_),
    .C(net41),
    .Y(_0166_));
 sg13g2_nor2b_1 _3010_ (.A(_0372_),
    .B_N(_1608_),
    .Y(_0424_));
 sg13g2_nor2_1 _3011_ (.A(_1608_),
    .B(_0422_),
    .Y(_0425_));
 sg13g2_nor3_1 _3012_ (.A(_0424_),
    .B(_0425_),
    .C(_0395_),
    .Y(_0167_));
 sg13g2_nor2_1 _3013_ (.A(\vga.interval_counter[9] ),
    .B(_0424_),
    .Y(_0426_));
 sg13g2_nor3_1 _3014_ (.A(_0373_),
    .B(_0426_),
    .C(_0395_),
    .Y(_0168_));
 sg13g2_nor2_1 _3015_ (.A(_0259_),
    .B(_0260_),
    .Y(_0170_));
 sg13g2_nor2_1 _3016_ (.A(_0261_),
    .B(_0262_),
    .Y(_0172_));
 sg13g2_nor2_2 _3017_ (.A(_1725_),
    .B(_1727_),
    .Y(_0427_));
 sg13g2_inv_1 _3018_ (.Y(_0428_),
    .A(_0427_));
 sg13g2_nor3_1 _3019_ (.A(_1705_),
    .B(_0428_),
    .C(_1680_),
    .Y(_0429_));
 sg13g2_nand2_1 _3020_ (.Y(_0430_),
    .A(_1701_),
    .B(_0429_));
 sg13g2_a21oi_1 _3021_ (.A1(_1689_),
    .A2(_1690_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_nand2_1 _3022_ (.Y(_0432_),
    .A(_0431_),
    .B(_1743_));
 sg13g2_inv_2 _3023_ (.Y(_0433_),
    .A(_1974_));
 sg13g2_a21oi_1 _3024_ (.A1(_0432_),
    .A2(_1741_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_inv_1 _3025_ (.Y(_0435_),
    .A(_0295_));
 sg13g2_nor2_1 _3026_ (.A(_0278_),
    .B(_0279_),
    .Y(_0436_));
 sg13g2_inv_1 _3027_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_nor2_1 _3028_ (.A(_0284_),
    .B(_0285_),
    .Y(_0438_));
 sg13g2_inv_1 _3029_ (.Y(_0439_),
    .A(_0438_));
 sg13g2_nor4_1 _3030_ (.A(_0435_),
    .B(_0311_),
    .C(_0437_),
    .D(_0439_),
    .Y(_0440_));
 sg13g2_inv_1 _3031_ (.Y(_0441_),
    .A(_0296_));
 sg13g2_inv_1 _3032_ (.Y(_0442_),
    .A(_0291_));
 sg13g2_nor2_1 _3033_ (.A(_0290_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_inv_1 _3034_ (.Y(_0444_),
    .A(_0294_));
 sg13g2_nor2_1 _3035_ (.A(_0444_),
    .B(_0293_),
    .Y(_0445_));
 sg13g2_a21oi_1 _3036_ (.A1(_0441_),
    .A2(_0443_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_nand3_1 _3037_ (.B(_1799_),
    .C(_0446_),
    .A(_0440_),
    .Y(_0447_));
 sg13g2_buf_1 _3038_ (.A(_0065_),
    .X(_0448_));
 sg13g2_inv_1 _3039_ (.Y(_0449_),
    .A(_0448_));
 sg13g2_nand2_1 _3040_ (.Y(_0450_),
    .A(_0432_),
    .B(_1741_));
 sg13g2_xnor2_1 _3041_ (.Y(_0451_),
    .A(_0449_),
    .B(_0450_));
 sg13g2_nor2_1 _3042_ (.A(_0428_),
    .B(_1680_),
    .Y(_0452_));
 sg13g2_xnor2_1 _3043_ (.Y(_0453_),
    .A(_0452_),
    .B(_1707_));
 sg13g2_nor2_1 _3044_ (.A(_2011_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_buf_2 _3045_ (.A(_0041_),
    .X(_0455_));
 sg13g2_xnor2_1 _3046_ (.Y(_0456_),
    .A(_0455_),
    .B(_0453_));
 sg13g2_buf_2 _3047_ (.A(_0040_),
    .X(_0457_));
 sg13g2_inv_2 _3048_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_inv_1 _3049_ (.Y(_0459_),
    .A(_1710_));
 sg13g2_nand2_1 _3050_ (.Y(_0460_),
    .A(_0427_),
    .B(_1675_));
 sg13g2_a21oi_1 _3051_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(_0452_));
 sg13g2_inv_1 _3052_ (.Y(_0462_),
    .A(_1677_));
 sg13g2_inv_1 _3053_ (.Y(_0463_),
    .A(net63));
 sg13g2_nor2_1 _3054_ (.A(_0463_),
    .B(_0427_),
    .Y(_0464_));
 sg13g2_xnor2_1 _3055_ (.Y(_0465_),
    .A(_0462_),
    .B(_0464_));
 sg13g2_inv_2 _3056_ (.Y(_0466_),
    .A(\vga.count_v[3] ));
 sg13g2_nand2_1 _3057_ (.Y(_0467_),
    .A(_0465_),
    .B(_0466_));
 sg13g2_o21ai_1 _3058_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0458_),
    .A2(_0461_));
 sg13g2_xnor2_1 _3059_ (.Y(_0469_),
    .A(net63),
    .B(_0427_));
 sg13g2_inv_1 _3060_ (.Y(_0470_),
    .A(_0469_));
 sg13g2_inv_2 _3061_ (.Y(_0471_),
    .A(_0038_));
 sg13g2_xnor2_1 _3062_ (.Y(_0472_),
    .A(_0471_),
    .B(_0469_));
 sg13g2_inv_1 _3063_ (.Y(_0473_),
    .A(_1725_));
 sg13g2_nor2_1 _3064_ (.A(net78),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_nand2_1 _3065_ (.Y(_0475_),
    .A(_1749_),
    .B(net77));
 sg13g2_a21oi_1 _3066_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0476_),
    .B1(_0427_));
 sg13g2_nand2_2 _3067_ (.Y(_0477_),
    .A(net78),
    .B(_1971_));
 sg13g2_nand2b_1 _3068_ (.Y(_0478_),
    .B(_0477_),
    .A_N(_0476_));
 sg13g2_nor2_1 _3069_ (.A(_0466_),
    .B(_0465_),
    .Y(_0479_));
 sg13g2_a221oi_1 _3070_ (.B2(_0478_),
    .C1(_0479_),
    .B1(_0472_),
    .A1(net76),
    .Y(_0480_),
    .A2(_0470_));
 sg13g2_nor2_1 _3071_ (.A(_0468_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_a21oi_1 _3072_ (.A1(_0458_),
    .A2(_0461_),
    .Y(_0482_),
    .B1(_0481_));
 sg13g2_nor2_1 _3073_ (.A(_0456_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_buf_2 _3074_ (.A(_0042_),
    .X(_0484_));
 sg13g2_inv_1 _3075_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_xnor2_1 _3076_ (.Y(_0486_),
    .A(_0429_),
    .B(_1701_));
 sg13g2_xnor2_1 _3077_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_o21ai_1 _3078_ (.B1(_0487_),
    .Y(_0488_),
    .A1(_0454_),
    .A2(_0483_));
 sg13g2_inv_1 _3079_ (.Y(_0489_),
    .A(_1984_));
 sg13g2_nor2_1 _3080_ (.A(_0489_),
    .B(_0486_),
    .Y(_0490_));
 sg13g2_inv_2 _3081_ (.Y(_0491_),
    .A(_1983_));
 sg13g2_xor2_1 _3082_ (.B(_1691_),
    .A(_0430_),
    .X(_0492_));
 sg13g2_nor2_1 _3083_ (.A(_0491_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nor2_1 _3084_ (.A(_0490_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_nand2_1 _3085_ (.Y(_0495_),
    .A(_0488_),
    .B(_0494_));
 sg13g2_buf_1 _3086_ (.A(_0044_),
    .X(_0496_));
 sg13g2_xnor2_1 _3087_ (.Y(_0497_),
    .A(_1743_),
    .B(_0431_));
 sg13g2_a22oi_1 _3088_ (.Y(_0498_),
    .B1(net71),
    .B2(_0497_),
    .A2(_0492_),
    .A1(_0491_));
 sg13g2_nor2_1 _3089_ (.A(net71),
    .B(_0497_),
    .Y(_0499_));
 sg13g2_a21oi_1 _3090_ (.A1(_0495_),
    .A2(_0498_),
    .Y(_0500_),
    .B1(_0499_));
 sg13g2_nor2_1 _3091_ (.A(_0451_),
    .B(_0500_),
    .Y(_0501_));
 sg13g2_xnor2_1 _3092_ (.Y(_0502_),
    .A(_0491_),
    .B(_1764_));
 sg13g2_xnor2_1 _3093_ (.Y(_0503_),
    .A(_0485_),
    .B(_1778_));
 sg13g2_inv_1 _3094_ (.Y(_0504_),
    .A(_0455_));
 sg13g2_nor2_1 _3095_ (.A(net77),
    .B(_1749_),
    .Y(_0505_));
 sg13g2_nand2_1 _3096_ (.Y(_0506_),
    .A(_0473_),
    .B(net78));
 sg13g2_a21oi_1 _3097_ (.A1(_0505_),
    .A2(_0506_),
    .Y(_0507_),
    .B1(_0474_));
 sg13g2_nand2_1 _3098_ (.Y(_0508_),
    .A(net76),
    .B(net63));
 sg13g2_inv_1 _3099_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_a22oi_1 _3100_ (.Y(_0510_),
    .B1(_0466_),
    .B2(_1724_),
    .A2(_0463_),
    .A1(_2004_));
 sg13g2_o21ai_1 _3101_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_0507_),
    .A2(_0509_));
 sg13g2_inv_1 _3102_ (.Y(_0512_),
    .A(_1771_));
 sg13g2_a22oi_1 _3103_ (.Y(_0513_),
    .B1(_0458_),
    .B2(_0512_),
    .A2(_1786_),
    .A1(net75));
 sg13g2_nand2_1 _3104_ (.Y(_0514_),
    .A(_1771_),
    .B(_0457_));
 sg13g2_o21ai_1 _3105_ (.B1(_0514_),
    .Y(_0515_),
    .A1(_0455_),
    .A2(_1774_));
 sg13g2_a221oi_1 _3106_ (.B2(_0513_),
    .C1(_0515_),
    .B1(_0511_),
    .A1(_0455_),
    .Y(_0516_),
    .A2(_1774_));
 sg13g2_a21o_1 _3107_ (.A2(_1770_),
    .A1(_0504_),
    .B1(_0516_),
    .X(_0517_));
 sg13g2_a22oi_1 _3108_ (.Y(_0518_),
    .B1(_0503_),
    .B2(_0517_),
    .A2(_1758_),
    .A1(_0485_));
 sg13g2_inv_1 _3109_ (.Y(_0519_),
    .A(_0043_));
 sg13g2_inv_1 _3110_ (.Y(_0520_),
    .A(net71));
 sg13g2_a22oi_1 _3111_ (.Y(_0521_),
    .B1(_0520_),
    .B2(_1795_),
    .A2(_1766_),
    .A1(_0519_));
 sg13g2_o21ai_1 _3112_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0502_),
    .A2(_0518_));
 sg13g2_inv_1 _3113_ (.Y(_0523_),
    .A(_1795_));
 sg13g2_xnor2_1 _3114_ (.Y(_0524_),
    .A(_0433_),
    .B(_1793_));
 sg13g2_a21oi_1 _3115_ (.A1(_0523_),
    .A2(net71),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_a21oi_1 _3116_ (.A1(_0522_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0449_));
 sg13g2_nor4_1 _3117_ (.A(_0434_),
    .B(_0447_),
    .C(_0501_),
    .D(_0526_),
    .Y(_0527_));
 sg13g2_nor2_2 _3118_ (.A(_1445_),
    .B(_1449_),
    .Y(_0528_));
 sg13g2_inv_1 _3119_ (.Y(_0529_),
    .A(_0528_));
 sg13g2_nor2_1 _3120_ (.A(_0529_),
    .B(_1422_),
    .Y(_0530_));
 sg13g2_nand2_1 _3121_ (.Y(_0531_),
    .A(_0530_),
    .B(_1424_));
 sg13g2_a21oi_1 _3122_ (.A1(_1480_),
    .A2(_1433_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_nand2_1 _3123_ (.Y(_0533_),
    .A(_0532_),
    .B(_1429_));
 sg13g2_o21ai_1 _3124_ (.B1(_1497_),
    .Y(_0534_),
    .A1(_1435_),
    .A2(_0533_));
 sg13g2_xnor2_1 _3125_ (.Y(_0535_),
    .A(_0448_),
    .B(_0534_));
 sg13g2_xnor2_1 _3126_ (.Y(_0536_),
    .A(_1435_),
    .B(_0533_));
 sg13g2_nor2_1 _3127_ (.A(_0530_),
    .B(_1474_),
    .Y(_0537_));
 sg13g2_nor2b_1 _3128_ (.A(_0537_),
    .B_N(_0531_),
    .Y(_0538_));
 sg13g2_inv_1 _3129_ (.Y(_0539_),
    .A(_0538_));
 sg13g2_nor2_1 _3130_ (.A(_1418_),
    .B(_0528_),
    .Y(_0540_));
 sg13g2_xnor2_1 _3131_ (.Y(_0541_),
    .A(_1420_),
    .B(_0540_));
 sg13g2_inv_1 _3132_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_a21oi_1 _3133_ (.A1(_0529_),
    .A2(net68),
    .Y(_0543_),
    .B1(_1416_));
 sg13g2_nor2_1 _3134_ (.A(_0540_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a22oi_1 _3135_ (.Y(_0545_),
    .B1(_0466_),
    .B2(_0544_),
    .A2(_1982_),
    .A1(_0541_));
 sg13g2_inv_1 _3136_ (.Y(_0546_),
    .A(_0477_));
 sg13g2_inv_1 _3137_ (.Y(_0547_),
    .A(_1445_));
 sg13g2_nor2_1 _3138_ (.A(net78),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_nand2_1 _3139_ (.Y(_0549_),
    .A(_1498_),
    .B(net77));
 sg13g2_a21oi_1 _3140_ (.A1(_0548_),
    .A2(_0549_),
    .Y(_0550_),
    .B1(_0528_));
 sg13g2_xnor2_1 _3141_ (.Y(_0551_),
    .A(net68),
    .B(_0528_));
 sg13g2_xnor2_1 _3142_ (.Y(_0552_),
    .A(_0471_),
    .B(_0551_));
 sg13g2_o21ai_1 _3143_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0546_),
    .A2(_0550_));
 sg13g2_o21ai_1 _3144_ (.B1(net75),
    .Y(_0554_),
    .A1(_0540_),
    .A2(_0543_));
 sg13g2_nand2b_1 _3145_ (.Y(_0555_),
    .B(net76),
    .A_N(_0551_));
 sg13g2_nand3_1 _3146_ (.B(_0554_),
    .C(_0555_),
    .A(_0553_),
    .Y(_0556_));
 sg13g2_a22oi_1 _3147_ (.Y(_0557_),
    .B1(_0545_),
    .B2(_0556_),
    .A2(_0542_),
    .A1(net73));
 sg13g2_o21ai_1 _3148_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_2011_),
    .A2(_0539_));
 sg13g2_xnor2_1 _3149_ (.Y(_0559_),
    .A(_0531_),
    .B(_1481_));
 sg13g2_xnor2_1 _3150_ (.Y(_0560_),
    .A(_0484_),
    .B(_0559_));
 sg13g2_nand2_1 _3151_ (.Y(_0561_),
    .A(_0539_),
    .B(_2011_));
 sg13g2_nand3_1 _3152_ (.B(_0560_),
    .C(_0561_),
    .A(_0558_),
    .Y(_0562_));
 sg13g2_xor2_1 _3153_ (.B(_0532_),
    .A(_1429_),
    .X(_0563_));
 sg13g2_a22oi_1 _3154_ (.Y(_0564_),
    .B1(_1983_),
    .B2(_0563_),
    .A2(_0559_),
    .A1(_1984_));
 sg13g2_nand2_1 _3155_ (.Y(_0565_),
    .A(_0536_),
    .B(net71));
 sg13g2_o21ai_1 _3156_ (.B1(_0565_),
    .Y(_0566_),
    .A1(_1983_),
    .A2(_0563_));
 sg13g2_a21o_1 _3157_ (.A2(_0564_),
    .A1(_0562_),
    .B1(_0566_),
    .X(_0567_));
 sg13g2_o21ai_1 _3158_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net71),
    .A2(_0536_));
 sg13g2_a22oi_1 _3159_ (.Y(_0569_),
    .B1(_0535_),
    .B2(_0568_),
    .A2(_0534_),
    .A1(_1974_));
 sg13g2_xnor2_1 _3160_ (.Y(_0570_),
    .A(_0491_),
    .B(_1517_));
 sg13g2_nor2_1 _3161_ (.A(_0466_),
    .B(_1461_),
    .Y(_0571_));
 sg13g2_inv_1 _3162_ (.Y(_0572_),
    .A(net68));
 sg13g2_nor2_1 _3163_ (.A(\vga.count_v[0] ),
    .B(_1498_),
    .Y(_0573_));
 sg13g2_nand2_1 _3164_ (.Y(_0574_),
    .A(_0547_),
    .B(net78));
 sg13g2_a21oi_1 _3165_ (.A1(_0573_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(_0548_));
 sg13g2_a21oi_1 _3166_ (.A1(net76),
    .A2(net68),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_a21oi_1 _3167_ (.A1(_2004_),
    .A2(_0572_),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_a22oi_1 _3168_ (.Y(_0578_),
    .B1(_0457_),
    .B2(_1527_),
    .A2(_1461_),
    .A1(_0466_));
 sg13g2_o21ai_1 _3169_ (.B1(_0578_),
    .Y(_0579_),
    .A1(_0571_),
    .A2(_0577_));
 sg13g2_nand2_1 _3170_ (.Y(_0580_),
    .A(_1526_),
    .B(_0458_));
 sg13g2_xnor2_1 _3171_ (.Y(_0581_),
    .A(_0455_),
    .B(_1524_));
 sg13g2_a21oi_1 _3172_ (.A1(_0579_),
    .A2(_0580_),
    .Y(_0582_),
    .B1(_0581_));
 sg13g2_a21o_1 _3173_ (.A2(_1534_),
    .A1(_0504_),
    .B1(_0582_),
    .X(_0583_));
 sg13g2_xnor2_1 _3174_ (.Y(_0584_),
    .A(_0485_),
    .B(_1538_));
 sg13g2_nor2_1 _3175_ (.A(_0484_),
    .B(_1515_),
    .Y(_0585_));
 sg13g2_a21oi_1 _3176_ (.A1(_0583_),
    .A2(_0584_),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_a22oi_1 _3177_ (.Y(_0587_),
    .B1(_0520_),
    .B2(_1514_),
    .A2(_1510_),
    .A1(_0519_));
 sg13g2_o21ai_1 _3178_ (.B1(_0587_),
    .Y(_0588_),
    .A1(_0570_),
    .A2(_0586_));
 sg13g2_xnor2_1 _3179_ (.Y(_0589_),
    .A(_0433_),
    .B(_1548_));
 sg13g2_nand2_1 _3180_ (.Y(_0590_),
    .A(_1545_),
    .B(net71));
 sg13g2_nand3_1 _3181_ (.B(_0589_),
    .C(_0590_),
    .A(_0588_),
    .Y(_0591_));
 sg13g2_nand2_1 _3182_ (.Y(_0592_),
    .A(_0591_),
    .B(_0448_));
 sg13g2_nor2_1 _3183_ (.A(_0295_),
    .B(_0444_),
    .Y(_0593_));
 sg13g2_nand2_1 _3184_ (.Y(_0594_),
    .A(_0593_),
    .B(_0291_));
 sg13g2_nand3_1 _3185_ (.B(_0435_),
    .C(_0050_),
    .A(_0594_),
    .Y(_0595_));
 sg13g2_nor3_1 _3186_ (.A(_0288_),
    .B(_0595_),
    .C(_1549_),
    .Y(_0596_));
 sg13g2_nand3_1 _3187_ (.B(_0592_),
    .C(_0596_),
    .A(_0569_),
    .Y(_0597_));
 sg13g2_inv_1 _3188_ (.Y(_0598_),
    .A(_0293_));
 sg13g2_inv_1 _3189_ (.Y(_0599_),
    .A(_0284_));
 sg13g2_nor2_2 _3190_ (.A(_0285_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_inv_1 _3191_ (.Y(_0601_),
    .A(_0600_));
 sg13g2_nor2_2 _3192_ (.A(_0282_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_nor2_1 _3193_ (.A(_0294_),
    .B(_0295_),
    .Y(_0603_));
 sg13g2_nand3_1 _3194_ (.B(_0310_),
    .C(_0603_),
    .A(_0602_),
    .Y(_0604_));
 sg13g2_nor2_1 _3195_ (.A(_0437_),
    .B(_0601_),
    .Y(_0605_));
 sg13g2_nor2_2 _3196_ (.A(_0438_),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_o21ai_1 _3197_ (.B1(_0606_),
    .Y(_0607_),
    .A1(_0598_),
    .A2(_0604_));
 sg13g2_nor2_1 _3198_ (.A(_0290_),
    .B(_0291_),
    .Y(_0608_));
 sg13g2_inv_1 _3199_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_nand2_1 _3200_ (.Y(_0610_),
    .A(_0609_),
    .B(_0441_));
 sg13g2_nand2_1 _3201_ (.Y(_0611_),
    .A(_0439_),
    .B(_0301_));
 sg13g2_inv_1 _3202_ (.Y(_0612_),
    .A(_0606_));
 sg13g2_o21ai_1 _3203_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0610_),
    .A2(_0611_));
 sg13g2_inv_1 _3204_ (.Y(_0614_),
    .A(_0603_));
 sg13g2_nor2b_1 _3205_ (.A(_0614_),
    .B_N(_0443_),
    .Y(_0615_));
 sg13g2_nand3_1 _3206_ (.B(_0602_),
    .C(_0310_),
    .A(_0615_),
    .Y(_0616_));
 sg13g2_nand4_1 _3207_ (.B(_0613_),
    .C(_0457_),
    .A(_0607_),
    .Y(_0617_),
    .D(_0616_));
 sg13g2_nand2_1 _3208_ (.Y(_0618_),
    .A(_0597_),
    .B(_0617_));
 sg13g2_inv_1 _3209_ (.Y(_0619_),
    .A(_1569_));
 sg13g2_inv_2 _3210_ (.Y(_0620_),
    .A(_1577_));
 sg13g2_inv_1 _3211_ (.Y(_0621_),
    .A(_1576_));
 sg13g2_nor3_1 _3212_ (.A(_1575_),
    .B(_0621_),
    .C(_1564_),
    .Y(_0622_));
 sg13g2_nand2_1 _3213_ (.Y(_0623_),
    .A(_0622_),
    .B(net61));
 sg13g2_nor3_2 _3214_ (.A(_0619_),
    .B(_0620_),
    .C(_0623_),
    .Y(_0624_));
 sg13g2_xor2_1 _3215_ (.B(_0624_),
    .A(_0047_),
    .X(_0625_));
 sg13g2_xnor2_1 _3216_ (.Y(_0626_),
    .A(_1577_),
    .B(_0623_));
 sg13g2_nor2_1 _3217_ (.A(_0620_),
    .B(_0623_),
    .Y(_0627_));
 sg13g2_xnor2_1 _3218_ (.Y(_0628_),
    .A(_0046_),
    .B(_0627_));
 sg13g2_nand2_1 _3219_ (.Y(_0629_),
    .A(_1566_),
    .B(_1563_));
 sg13g2_inv_1 _3220_ (.Y(_0630_),
    .A(_0629_));
 sg13g2_nand2_1 _3221_ (.Y(_0631_),
    .A(_0630_),
    .B(_1562_));
 sg13g2_nor2_2 _3222_ (.A(_1575_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_xnor2_1 _3223_ (.Y(_0633_),
    .A(_0621_),
    .B(_0632_));
 sg13g2_nor2_1 _3224_ (.A(_1565_),
    .B(_0631_),
    .Y(_0634_));
 sg13g2_xnor2_1 _3225_ (.Y(_0635_),
    .A(net80),
    .B(_0631_));
 sg13g2_xnor2_1 _3226_ (.Y(_0636_),
    .A(_0052_),
    .B(_0632_));
 sg13g2_nor2_1 _3227_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_o21ai_1 _3228_ (.B1(_0637_),
    .Y(_0638_),
    .A1(_0633_),
    .A2(_0634_));
 sg13g2_nor3_1 _3229_ (.A(_0626_),
    .B(_0628_),
    .C(_0638_),
    .Y(_0639_));
 sg13g2_xnor2_1 _3230_ (.Y(_0640_),
    .A(_0625_),
    .B(_0639_));
 sg13g2_nor2_1 _3231_ (.A(_0054_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_inv_1 _3232_ (.Y(_0642_),
    .A(_0641_));
 sg13g2_nand4_1 _3233_ (.B(_1569_),
    .C(net81),
    .A(_0632_),
    .Y(_0643_),
    .D(_1579_));
 sg13g2_xnor2_1 _3234_ (.Y(_0644_),
    .A(_1571_),
    .B(_0643_));
 sg13g2_inv_1 _3235_ (.Y(_0645_),
    .A(net81));
 sg13g2_xnor2_1 _3236_ (.Y(_0646_),
    .A(_0645_),
    .B(_0624_));
 sg13g2_inv_1 _3237_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_nand4_1 _3238_ (.B(net62),
    .C(_1576_),
    .A(_0632_),
    .Y(_0648_),
    .D(_1577_));
 sg13g2_nor2_1 _3239_ (.A(_1569_),
    .B(_0627_),
    .Y(_0649_));
 sg13g2_nor2_1 _3240_ (.A(_0624_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_nor2b_1 _3241_ (.A(_0650_),
    .B_N(_0625_),
    .Y(_0651_));
 sg13g2_inv_1 _3242_ (.Y(_0652_),
    .A(_0651_));
 sg13g2_a21o_1 _3243_ (.A2(_0648_),
    .A1(_0647_),
    .B1(_0652_),
    .X(_0653_));
 sg13g2_xnor2_1 _3244_ (.Y(_0654_),
    .A(_0644_),
    .B(_0653_));
 sg13g2_xnor2_1 _3245_ (.Y(_0655_),
    .A(_0066_),
    .B(_0654_));
 sg13g2_nand2b_1 _3246_ (.Y(_0656_),
    .B(_0285_),
    .A_N(_0654_));
 sg13g2_o21ai_1 _3247_ (.B1(_0656_),
    .Y(_0657_),
    .A1(_0642_),
    .A2(_0655_));
 sg13g2_nand3b_1 _3248_ (.B(_0622_),
    .C(_1570_),
    .Y(_0658_),
    .A_N(_0057_));
 sg13g2_nor4_2 _3249_ (.A(_0619_),
    .B(_0620_),
    .C(_1572_),
    .Y(_0659_),
    .D(_0658_));
 sg13g2_nand3b_1 _3250_ (.B(_0639_),
    .C(_0647_),
    .Y(_0660_),
    .A_N(_0644_));
 sg13g2_xnor2_1 _3251_ (.Y(_0661_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_or3_1 _3252_ (.A(_0659_),
    .B(_0644_),
    .C(_0653_),
    .X(_0662_));
 sg13g2_nand2b_1 _3253_ (.Y(_0663_),
    .B(_0662_),
    .A_N(_0661_));
 sg13g2_inv_1 _3254_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_xnor2_1 _3255_ (.Y(_0665_),
    .A(_0626_),
    .B(_0638_));
 sg13g2_nor2_1 _3256_ (.A(_0280_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_xnor2_1 _3257_ (.Y(_0667_),
    .A(_0648_),
    .B(_0628_));
 sg13g2_xnor2_1 _3258_ (.Y(_0668_),
    .A(_0278_),
    .B(_0667_));
 sg13g2_nor2_1 _3259_ (.A(net62),
    .B(_0636_),
    .Y(_0669_));
 sg13g2_a21oi_1 _3260_ (.A1(net62),
    .A2(_0052_),
    .Y(_0670_),
    .B1(_0669_));
 sg13g2_xnor2_1 _3261_ (.Y(_0671_),
    .A(_0058_),
    .B(_0670_));
 sg13g2_xnor2_1 _3262_ (.Y(_0672_),
    .A(net80),
    .B(_1568_));
 sg13g2_inv_1 _3263_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_nor2_1 _3264_ (.A(_0056_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nand2b_1 _3265_ (.Y(_0675_),
    .B(_0674_),
    .A_N(_0671_));
 sg13g2_o21ai_1 _3266_ (.B1(_0675_),
    .Y(_0676_),
    .A1(_0306_),
    .A2(_0670_));
 sg13g2_xnor2_1 _3267_ (.Y(_0677_),
    .A(_0055_),
    .B(_0665_));
 sg13g2_nor2b_1 _3268_ (.A(_0677_),
    .B_N(_0668_),
    .Y(_0678_));
 sg13g2_nor2_1 _3269_ (.A(_0298_),
    .B(_0667_),
    .Y(_0679_));
 sg13g2_a221oi_1 _3270_ (.B2(_0678_),
    .C1(_0679_),
    .B1(_0676_),
    .A1(_0666_),
    .Y(_0680_),
    .A2(_0668_));
 sg13g2_inv_1 _3271_ (.Y(_0681_),
    .A(_0056_));
 sg13g2_nor2_1 _3272_ (.A(_0681_),
    .B(_0672_),
    .Y(_0682_));
 sg13g2_nor3_1 _3273_ (.A(_0674_),
    .B(_0682_),
    .C(_0671_),
    .Y(_0683_));
 sg13g2_inv_1 _3274_ (.Y(_0684_),
    .A(_0290_));
 sg13g2_nor2_1 _3275_ (.A(_0291_),
    .B(net61),
    .Y(_0685_));
 sg13g2_o21ai_1 _3276_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_0684_),
    .A2(_1565_));
 sg13g2_nand2_1 _3277_ (.Y(_0687_),
    .A(net62),
    .B(net61));
 sg13g2_a21oi_1 _3278_ (.A1(_0686_),
    .A2(_0687_),
    .Y(_0688_),
    .B1(_0598_));
 sg13g2_a21oi_1 _3279_ (.A1(_0630_),
    .A2(_1565_),
    .Y(_0689_),
    .B1(_1562_));
 sg13g2_nor2_1 _3280_ (.A(_1568_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_xnor2_1 _3281_ (.Y(_0691_),
    .A(_0295_),
    .B(_0690_));
 sg13g2_inv_1 _3282_ (.Y(_0692_),
    .A(_0053_));
 sg13g2_xnor2_1 _3283_ (.Y(_0693_),
    .A(_1563_),
    .B(_1567_));
 sg13g2_xnor2_1 _3284_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nand2_1 _3285_ (.Y(_0695_),
    .A(_0691_),
    .B(_0694_));
 sg13g2_nor2_1 _3286_ (.A(_0444_),
    .B(_0693_),
    .Y(_0696_));
 sg13g2_nor2_1 _3287_ (.A(_0435_),
    .B(_0690_),
    .Y(_0697_));
 sg13g2_a21oi_1 _3288_ (.A1(_0691_),
    .A2(_0696_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_o21ai_1 _3289_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0688_),
    .A2(_0695_));
 sg13g2_nand3_1 _3290_ (.B(_0683_),
    .C(_0699_),
    .A(_0678_),
    .Y(_0700_));
 sg13g2_nand2_1 _3291_ (.Y(_0701_),
    .A(_0680_),
    .B(_0700_));
 sg13g2_inv_1 _3292_ (.Y(_0702_),
    .A(_0054_));
 sg13g2_nor2b_1 _3293_ (.A(_0702_),
    .B_N(_0640_),
    .Y(_0703_));
 sg13g2_nor4_1 _3294_ (.A(_0641_),
    .B(_0703_),
    .C(_0663_),
    .D(_0655_),
    .Y(_0704_));
 sg13g2_a22oi_1 _3295_ (.Y(_0705_),
    .B1(_0701_),
    .B2(_0704_),
    .A2(_0664_),
    .A1(_0657_));
 sg13g2_nor2_2 _3296_ (.A(net86),
    .B(net88),
    .Y(_0706_));
 sg13g2_inv_1 _3297_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_nor2_1 _3298_ (.A(net85),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_inv_1 _3299_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_nor2_1 _3300_ (.A(net70),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_xnor2_1 _3301_ (.Y(_0711_),
    .A(_0074_),
    .B(_0710_));
 sg13g2_nor2_1 _3302_ (.A(_2011_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nand2_1 _3303_ (.Y(_0713_),
    .A(_0711_),
    .B(_2011_));
 sg13g2_xnor2_1 _3304_ (.Y(_0714_),
    .A(net70),
    .B(_0708_));
 sg13g2_xnor2_1 _3305_ (.Y(_0715_),
    .A(_0457_),
    .B(_0714_));
 sg13g2_nand3b_1 _3306_ (.B(_0713_),
    .C(_0715_),
    .Y(_0716_),
    .A_N(_0712_));
 sg13g2_nand2_1 _3307_ (.Y(_0717_),
    .A(net78),
    .B(net88));
 sg13g2_o21ai_1 _3308_ (.B1(_0717_),
    .Y(_0718_),
    .A1(\vga.count_v[0] ),
    .A2(net69));
 sg13g2_a21oi_1 _3309_ (.A1(_2002_),
    .A2(_1444_),
    .Y(_0719_),
    .B1(_0718_));
 sg13g2_nor2b_1 _3310_ (.A(_0719_),
    .B_N(_0717_),
    .Y(_0720_));
 sg13g2_nand2_1 _3311_ (.Y(_0721_),
    .A(net86),
    .B(net88));
 sg13g2_inv_1 _3312_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_nor2_2 _3313_ (.A(_0706_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_xnor2_1 _3314_ (.Y(_0724_),
    .A(_0471_),
    .B(_0723_));
 sg13g2_xnor2_1 _3315_ (.Y(_0725_),
    .A(net85),
    .B(_0706_));
 sg13g2_nand2b_1 _3316_ (.Y(_0726_),
    .B(_0466_),
    .A_N(_0725_));
 sg13g2_nand2_1 _3317_ (.Y(_0727_),
    .A(_0725_),
    .B(net75));
 sg13g2_nand3b_1 _3318_ (.B(_0726_),
    .C(_0727_),
    .Y(_0728_),
    .A_N(_0724_));
 sg13g2_o21ai_1 _3319_ (.B1(_0727_),
    .Y(_0729_),
    .A1(_0720_),
    .A2(_0728_));
 sg13g2_nand3_1 _3320_ (.B(_1977_),
    .C(_0723_),
    .A(_0726_),
    .Y(_0730_));
 sg13g2_nor2b_1 _3321_ (.A(_0729_),
    .B_N(_0730_),
    .Y(_0731_));
 sg13g2_nand2_1 _3322_ (.Y(_0732_),
    .A(_0714_),
    .B(_0458_));
 sg13g2_inv_1 _3323_ (.Y(_0733_),
    .A(_0732_));
 sg13g2_a21oi_1 _3324_ (.A1(_0713_),
    .A2(_0733_),
    .Y(_0734_),
    .B1(_0712_));
 sg13g2_o21ai_1 _3325_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0716_),
    .A2(_0731_));
 sg13g2_nand2_1 _3326_ (.Y(_0736_),
    .A(_0710_),
    .B(_1485_));
 sg13g2_xnor2_1 _3327_ (.Y(_0737_),
    .A(_1539_),
    .B(_0736_));
 sg13g2_xnor2_1 _3328_ (.Y(_0738_),
    .A(_0484_),
    .B(_0737_));
 sg13g2_nor2_1 _3329_ (.A(net84),
    .B(_0736_),
    .Y(_0739_));
 sg13g2_xnor2_1 _3330_ (.Y(_0740_),
    .A(_0073_),
    .B(_0739_));
 sg13g2_nor2_1 _3331_ (.A(_0491_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_nand2_1 _3332_ (.Y(_0742_),
    .A(_0740_),
    .B(_0491_));
 sg13g2_nand2b_1 _3333_ (.Y(_0743_),
    .B(_0742_),
    .A_N(_0741_));
 sg13g2_nor2_1 _3334_ (.A(_0738_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand2_1 _3335_ (.Y(_0745_),
    .A(_0735_),
    .B(_0744_));
 sg13g2_nor2_1 _3336_ (.A(net67),
    .B(net70),
    .Y(_0746_));
 sg13g2_nand3_1 _3337_ (.B(net66),
    .C(_1714_),
    .A(_0746_),
    .Y(_0747_));
 sg13g2_nor2_1 _3338_ (.A(_0747_),
    .B(_0709_),
    .Y(_0748_));
 sg13g2_xnor2_1 _3339_ (.Y(_0749_),
    .A(_1431_),
    .B(_0748_));
 sg13g2_nand2_1 _3340_ (.Y(_0750_),
    .A(_0749_),
    .B(_0520_));
 sg13g2_nor2_1 _3341_ (.A(_0489_),
    .B(_0737_),
    .Y(_0751_));
 sg13g2_a21oi_1 _3342_ (.A1(_0742_),
    .A2(_0751_),
    .Y(_0752_),
    .B1(_0741_));
 sg13g2_nand3_1 _3343_ (.B(_0750_),
    .C(_0752_),
    .A(_0745_),
    .Y(_0753_));
 sg13g2_nor3_1 _3344_ (.A(net83),
    .B(_0747_),
    .C(_0709_),
    .Y(_0754_));
 sg13g2_xnor2_1 _3345_ (.Y(_0755_),
    .A(_0433_),
    .B(_0754_));
 sg13g2_nor2_1 _3346_ (.A(_0520_),
    .B(_0749_),
    .Y(_0756_));
 sg13g2_nor2_1 _3347_ (.A(_0755_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_a21oi_1 _3348_ (.A1(_0753_),
    .A2(_0757_),
    .Y(_0758_),
    .B1(_0449_));
 sg13g2_nand2_1 _3349_ (.Y(_0759_),
    .A(net67),
    .B(net84));
 sg13g2_nand2_2 _3350_ (.Y(_0760_),
    .A(_0722_),
    .B(net85));
 sg13g2_nor2_2 _3351_ (.A(_1499_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_inv_1 _3352_ (.Y(_0762_),
    .A(_0761_));
 sg13g2_nor2_1 _3353_ (.A(_0759_),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_xnor2_1 _3354_ (.Y(_0764_),
    .A(_0073_),
    .B(_0763_));
 sg13g2_nor2_1 _3355_ (.A(_0491_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_nand2_1 _3356_ (.Y(_0766_),
    .A(_0761_),
    .B(net67));
 sg13g2_xnor2_1 _3357_ (.Y(_0767_),
    .A(_1539_),
    .B(_0766_));
 sg13g2_nor2_1 _3358_ (.A(_0489_),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_nor2_1 _3359_ (.A(_0038_),
    .B(_0723_),
    .Y(_0769_));
 sg13g2_nor2b_1 _3360_ (.A(_0769_),
    .B_N(_0720_),
    .Y(_0770_));
 sg13g2_xnor2_1 _3361_ (.Y(_0771_),
    .A(_0075_),
    .B(_0721_));
 sg13g2_inv_1 _3362_ (.Y(_0772_),
    .A(_0771_));
 sg13g2_a22oi_1 _3363_ (.Y(_0773_),
    .B1(_0039_),
    .B2(_0772_),
    .A2(_0723_),
    .A1(_0038_));
 sg13g2_o21ai_1 _3364_ (.B1(_0773_),
    .Y(_0774_),
    .A1(_0039_),
    .A2(_0772_));
 sg13g2_xnor2_1 _3365_ (.Y(_0775_),
    .A(_1499_),
    .B(_0760_));
 sg13g2_a22oi_1 _3366_ (.Y(_0776_),
    .B1(_0458_),
    .B2(_0775_),
    .A2(_0771_),
    .A1(net75));
 sg13g2_o21ai_1 _3367_ (.B1(_0776_),
    .Y(_0777_),
    .A1(_0770_),
    .A2(_0774_));
 sg13g2_xnor2_1 _3368_ (.Y(_0778_),
    .A(_0074_),
    .B(_0761_));
 sg13g2_nand2b_1 _3369_ (.Y(_0779_),
    .B(_0457_),
    .A_N(_0775_));
 sg13g2_o21ai_1 _3370_ (.B1(_0779_),
    .Y(_0780_),
    .A1(_0455_),
    .A2(_0778_));
 sg13g2_a21oi_1 _3371_ (.A1(_0455_),
    .A2(_0778_),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_nand2_1 _3372_ (.Y(_0782_),
    .A(_0777_),
    .B(_0781_));
 sg13g2_nand2b_1 _3373_ (.Y(_0783_),
    .B(_1980_),
    .A_N(_0778_));
 sg13g2_xnor2_1 _3374_ (.Y(_0784_),
    .A(_0484_),
    .B(_0767_));
 sg13g2_a21oi_1 _3375_ (.A1(_0782_),
    .A2(_0783_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_nor3_1 _3376_ (.A(_0765_),
    .B(_0768_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_nand4_1 _3377_ (.B(_1413_),
    .C(net67),
    .A(_0761_),
    .Y(_0787_),
    .D(net84));
 sg13g2_xnor2_1 _3378_ (.Y(_0788_),
    .A(_1431_),
    .B(_0787_));
 sg13g2_inv_1 _3379_ (.Y(_0789_),
    .A(_0788_));
 sg13g2_nand2_1 _3380_ (.Y(_0790_),
    .A(_0788_),
    .B(_0496_));
 sg13g2_inv_1 _3381_ (.Y(_0791_),
    .A(net83));
 sg13g2_nor3_1 _3382_ (.A(net66),
    .B(_0791_),
    .C(_0759_),
    .Y(_0792_));
 sg13g2_nand2_1 _3383_ (.Y(_0793_),
    .A(_0761_),
    .B(_0792_));
 sg13g2_xnor2_1 _3384_ (.Y(_0794_),
    .A(_0448_),
    .B(_0793_));
 sg13g2_nand2_1 _3385_ (.Y(_0795_),
    .A(_0790_),
    .B(_0794_));
 sg13g2_a221oi_1 _3386_ (.B2(_0789_),
    .C1(_0795_),
    .B1(_0520_),
    .A1(_0491_),
    .Y(_0796_),
    .A2(_0764_));
 sg13g2_nor2b_1 _3387_ (.A(_0786_),
    .B_N(_0796_),
    .Y(_0797_));
 sg13g2_nor2_1 _3388_ (.A(_1562_),
    .B(_1563_),
    .Y(_0798_));
 sg13g2_inv_1 _3389_ (.Y(_0799_),
    .A(_0798_));
 sg13g2_nor2_1 _3390_ (.A(_1810_),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_inv_1 _3391_ (.Y(_0801_),
    .A(_0800_));
 sg13g2_nor2_1 _3392_ (.A(_1807_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_xnor2_1 _3393_ (.Y(_0803_),
    .A(_1577_),
    .B(_0802_));
 sg13g2_nor2_1 _3394_ (.A(_0279_),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_nor2_1 _3395_ (.A(net80),
    .B(_0801_),
    .Y(_0805_));
 sg13g2_xor2_1 _3396_ (.B(_0805_),
    .A(_0052_),
    .X(_0806_));
 sg13g2_nor2_1 _3397_ (.A(net72),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_nor2b_1 _3398_ (.A(_0280_),
    .B_N(_0803_),
    .Y(_0808_));
 sg13g2_nor2_2 _3399_ (.A(net61),
    .B(_1563_),
    .Y(_0809_));
 sg13g2_xnor2_1 _3400_ (.Y(_0810_),
    .A(_1562_),
    .B(_0809_));
 sg13g2_inv_1 _3401_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nor2_1 _3402_ (.A(_0809_),
    .B(_0630_),
    .Y(_0812_));
 sg13g2_a22oi_1 _3403_ (.Y(_0813_),
    .B1(_0295_),
    .B2(_0810_),
    .A2(_0812_),
    .A1(_0294_));
 sg13g2_o21ai_1 _3404_ (.B1(_0053_),
    .Y(_0814_),
    .A1(_0809_),
    .A2(_0630_));
 sg13g2_nor2_1 _3405_ (.A(_0290_),
    .B(net62),
    .Y(_0815_));
 sg13g2_nand2_1 _3406_ (.Y(_0816_),
    .A(_0291_),
    .B(net61));
 sg13g2_a21oi_1 _3407_ (.A1(_0815_),
    .A2(_0816_),
    .Y(_0817_),
    .B1(_0685_));
 sg13g2_nand2_1 _3408_ (.Y(_0818_),
    .A(_0812_),
    .B(_0692_));
 sg13g2_nand3_1 _3409_ (.B(_0817_),
    .C(_0818_),
    .A(_0814_),
    .Y(_0819_));
 sg13g2_xnor2_1 _3410_ (.Y(_0820_),
    .A(net80),
    .B(_0800_));
 sg13g2_xnor2_1 _3411_ (.Y(_0821_),
    .A(_0276_),
    .B(_0820_));
 sg13g2_a221oi_1 _3412_ (.B2(_0819_),
    .C1(_0821_),
    .B1(_0813_),
    .A1(_0435_),
    .Y(_0822_),
    .A2(_0811_));
 sg13g2_a22oi_1 _3413_ (.Y(_0823_),
    .B1(_0275_),
    .B2(_0806_),
    .A2(_0820_),
    .A1(_0681_));
 sg13g2_nor2b_1 _3414_ (.A(_0822_),
    .B_N(_0823_),
    .Y(_0824_));
 sg13g2_nor4_1 _3415_ (.A(_0804_),
    .B(_0807_),
    .C(_0808_),
    .D(_0824_),
    .Y(_0825_));
 sg13g2_inv_1 _3416_ (.Y(_0826_),
    .A(_0055_));
 sg13g2_inv_1 _3417_ (.Y(_0827_),
    .A(_0050_));
 sg13g2_nor2_1 _3418_ (.A(_0801_),
    .B(_1835_),
    .Y(_0828_));
 sg13g2_nand2_1 _3419_ (.Y(_0829_),
    .A(_0802_),
    .B(_0620_));
 sg13g2_nand2_1 _3420_ (.Y(_0830_),
    .A(_0829_),
    .B(_1569_));
 sg13g2_nor2b_1 _3421_ (.A(_0828_),
    .B_N(_0830_),
    .Y(_0831_));
 sg13g2_a22oi_1 _3422_ (.Y(_0832_),
    .B1(_0827_),
    .B2(_0831_),
    .A2(_0803_),
    .A1(_0826_));
 sg13g2_nand2b_1 _3423_ (.Y(_0833_),
    .B(_0832_),
    .A_N(_0825_));
 sg13g2_xnor2_1 _3424_ (.Y(_0834_),
    .A(net81),
    .B(_0828_));
 sg13g2_nand2b_1 _3425_ (.Y(_0835_),
    .B(_0599_),
    .A_N(_0834_));
 sg13g2_o21ai_1 _3426_ (.B1(_0835_),
    .Y(_0836_),
    .A1(_0827_),
    .A2(_0831_));
 sg13g2_a21oi_1 _3427_ (.A1(_0284_),
    .A2(_0834_),
    .Y(_0837_),
    .B1(_0836_));
 sg13g2_nand2_1 _3428_ (.Y(_0838_),
    .A(_0833_),
    .B(_0837_));
 sg13g2_nor3_2 _3429_ (.A(net81),
    .B(_0801_),
    .C(_1835_),
    .Y(_0839_));
 sg13g2_xnor2_1 _3430_ (.Y(_0840_),
    .A(_0048_),
    .B(_0839_));
 sg13g2_nand2b_1 _3431_ (.Y(_0841_),
    .B(_0285_),
    .A_N(_0840_));
 sg13g2_nand2_1 _3432_ (.Y(_0842_),
    .A(_0834_),
    .B(_0702_));
 sg13g2_nand3_1 _3433_ (.B(_0841_),
    .C(_0842_),
    .A(_0838_),
    .Y(_0843_));
 sg13g2_inv_1 _3434_ (.Y(_0844_),
    .A(_1971_));
 sg13g2_o21ai_1 _3435_ (.B1(_0719_),
    .Y(_0845_),
    .A1(_0844_),
    .A2(net87));
 sg13g2_nand2b_1 _3436_ (.Y(_0846_),
    .B(_0744_),
    .A_N(_0716_));
 sg13g2_nor3_1 _3437_ (.A(_0728_),
    .B(_0845_),
    .C(_0846_),
    .Y(_0847_));
 sg13g2_nand3_1 _3438_ (.B(_0757_),
    .C(_0750_),
    .A(_0847_),
    .Y(_0848_));
 sg13g2_nand3_1 _3439_ (.B(\vga.count_v[8] ),
    .C(_0794_),
    .A(_0789_),
    .Y(_0849_));
 sg13g2_o21ai_1 _3440_ (.B1(_0793_),
    .Y(_0850_),
    .A1(_1974_),
    .A2(_0754_));
 sg13g2_a22oi_1 _3441_ (.Y(_0851_),
    .B1(_0286_),
    .B2(_0840_),
    .A2(_0839_),
    .A1(_1572_));
 sg13g2_and3_1 _3442_ (.X(_0852_),
    .A(_0849_),
    .B(_0850_),
    .C(_0851_));
 sg13g2_nand3_1 _3443_ (.B(_0848_),
    .C(_0852_),
    .A(_0843_),
    .Y(_0853_));
 sg13g2_nor3_1 _3444_ (.A(_0758_),
    .B(_0797_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_nand2_1 _3445_ (.Y(_0855_),
    .A(_0705_),
    .B(_0854_));
 sg13g2_inv_1 _3446_ (.Y(_0856_),
    .A(_0276_));
 sg13g2_nor2_1 _3447_ (.A(net72),
    .B(_0856_),
    .Y(_0857_));
 sg13g2_inv_1 _3448_ (.Y(_0858_),
    .A(_0857_));
 sg13g2_nor2_1 _3449_ (.A(_0614_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_a21oi_1 _3450_ (.A1(_0606_),
    .A2(_0311_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_nand2_1 _3451_ (.Y(_0861_),
    .A(_0859_),
    .B(_0293_));
 sg13g2_nor2_1 _3452_ (.A(_0291_),
    .B(_0684_),
    .Y(_0862_));
 sg13g2_nand3_1 _3453_ (.B(_0857_),
    .C(_0862_),
    .A(_0441_),
    .Y(_0863_));
 sg13g2_nand3_1 _3454_ (.B(_0863_),
    .C(_0602_),
    .A(_0861_),
    .Y(_0864_));
 sg13g2_nor2_1 _3455_ (.A(_0856_),
    .B(_0296_),
    .Y(_0865_));
 sg13g2_inv_1 _3456_ (.Y(_0866_),
    .A(_0051_));
 sg13g2_a21oi_1 _3457_ (.A1(_0865_),
    .A2(_0866_),
    .Y(_0867_),
    .B1(net72));
 sg13g2_nor2_1 _3458_ (.A(_0867_),
    .B(_0612_),
    .Y(_0868_));
 sg13g2_nor3_1 _3459_ (.A(_0860_),
    .B(_0864_),
    .C(_0868_),
    .Y(_0869_));
 sg13g2_nor2_1 _3460_ (.A(_0295_),
    .B(_0445_),
    .Y(_0870_));
 sg13g2_o21ai_1 _3461_ (.B1(_0602_),
    .Y(_0871_),
    .A1(_0277_),
    .A2(_0870_));
 sg13g2_nand2_1 _3462_ (.Y(_0872_),
    .A(_0871_),
    .B(_0606_));
 sg13g2_nand4_1 _3463_ (.B(_0443_),
    .C(_0593_),
    .A(_0283_),
    .Y(_0873_),
    .D(_0600_));
 sg13g2_nand2_1 _3464_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_));
 sg13g2_nand3_1 _3465_ (.B(_0603_),
    .C(_0608_),
    .A(_0312_),
    .Y(_0875_));
 sg13g2_nand3_1 _3466_ (.B(_0284_),
    .C(_0827_),
    .A(_0875_),
    .Y(_0876_));
 sg13g2_nand2b_1 _3467_ (.Y(_0877_),
    .B(_0600_),
    .A_N(_0875_));
 sg13g2_nor2_1 _3468_ (.A(_0285_),
    .B(_0239_),
    .Y(_0878_));
 sg13g2_nand4_1 _3469_ (.B(_0876_),
    .C(_0877_),
    .A(_0874_),
    .Y(_0879_),
    .D(_0878_));
 sg13g2_a21oi_1 _3470_ (.A1(_0614_),
    .A2(net72),
    .Y(_0880_),
    .B1(_0301_));
 sg13g2_nand2_1 _3471_ (.Y(_0881_),
    .A(_0598_),
    .B(net72));
 sg13g2_nand3_1 _3472_ (.B(_0881_),
    .C(_0602_),
    .A(_0880_),
    .Y(_0882_));
 sg13g2_nand2_1 _3473_ (.Y(_0883_),
    .A(_0882_),
    .B(_0606_));
 sg13g2_nand4_1 _3474_ (.B(_0307_),
    .C(_0281_),
    .A(_0615_),
    .Y(_0884_),
    .D(_0600_));
 sg13g2_o21ai_1 _3475_ (.B1(net72),
    .Y(_0885_),
    .A1(_0276_),
    .A2(_0441_));
 sg13g2_a21oi_1 _3476_ (.A1(_0885_),
    .A2(_0602_),
    .Y(_0886_),
    .B1(_0612_));
 sg13g2_a21oi_1 _3477_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0887_),
    .B1(_0886_));
 sg13g2_nand2_1 _3478_ (.Y(_0888_),
    .A(_0887_),
    .B(\vga.score_r_unit_pixels[2] ));
 sg13g2_nand4_1 _3479_ (.B(\vga.score_r_unit_pixels[1] ),
    .C(_0886_),
    .A(_0872_),
    .Y(_0889_),
    .D(_0873_));
 sg13g2_nand3_1 _3480_ (.B(_0888_),
    .C(_0889_),
    .A(_0879_),
    .Y(_0890_));
 sg13g2_a21oi_1 _3481_ (.A1(\vga.score_r_ten_enable ),
    .A2(_0869_),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_and2_1 _3482_ (.A(_0307_),
    .B(_0593_),
    .X(_0892_));
 sg13g2_a21oi_1 _3483_ (.A1(_0892_),
    .A2(_0293_),
    .Y(_0893_),
    .B1(_0880_));
 sg13g2_nand2_1 _3484_ (.Y(_0894_),
    .A(_0893_),
    .B(_0439_));
 sg13g2_nand3_1 _3485_ (.B(_0443_),
    .C(_0605_),
    .A(_0892_),
    .Y(_0895_));
 sg13g2_nand3_1 _3486_ (.B(_0612_),
    .C(_0895_),
    .A(_0894_),
    .Y(_0896_));
 sg13g2_nand4_1 _3487_ (.B(\vga.score_l_unit_pixels[0] ),
    .C(_0612_),
    .A(_0896_),
    .Y(_0897_),
    .D(_0611_));
 sg13g2_nand4_1 _3488_ (.B(_0436_),
    .C(_0857_),
    .A(_0615_),
    .Y(_0898_),
    .D(_0600_));
 sg13g2_nor2b_1 _3489_ (.A(_0606_),
    .B_N(_0898_),
    .Y(_0899_));
 sg13g2_nand3_1 _3490_ (.B(_0311_),
    .C(_0439_),
    .A(_0861_),
    .Y(_0900_));
 sg13g2_inv_1 _3491_ (.Y(_0901_),
    .A(_0605_));
 sg13g2_o21ai_1 _3492_ (.B1(_0306_),
    .Y(_0902_),
    .A1(_0856_),
    .A2(_0296_));
 sg13g2_o21ai_1 _3493_ (.B1(_0439_),
    .Y(_0903_),
    .A1(_0901_),
    .A2(_0902_));
 sg13g2_inv_1 _3494_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_a21oi_1 _3495_ (.A1(_0899_),
    .A2(_0900_),
    .Y(_0905_),
    .B1(_0904_));
 sg13g2_nor3_1 _3496_ (.A(_2021_),
    .B(_0903_),
    .C(_0896_),
    .Y(_0906_));
 sg13g2_nor2_1 _3497_ (.A(_0905_),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_nand3_1 _3498_ (.B(_0897_),
    .C(_0907_),
    .A(_0891_),
    .Y(_0908_));
 sg13g2_nor3_1 _3499_ (.A(_1983_),
    .B(_0489_),
    .C(net56),
    .Y(_0909_));
 sg13g2_nand2_1 _3500_ (.Y(_0910_),
    .A(_2002_),
    .B(net77));
 sg13g2_nor4_1 _3501_ (.A(net74),
    .B(net73),
    .C(_0910_),
    .D(_2010_),
    .Y(_0911_));
 sg13g2_nand2b_1 _3502_ (.Y(_0912_),
    .B(_1977_),
    .A_N(_0080_));
 sg13g2_nor2_1 _3503_ (.A(net74),
    .B(net73),
    .Y(_0913_));
 sg13g2_nand4_1 _3504_ (.B(_0466_),
    .C(_0912_),
    .A(_0909_),
    .Y(_0914_),
    .D(_0913_));
 sg13g2_a22oi_1 _3505_ (.Y(_0915_),
    .B1(_2015_),
    .B2(_0914_),
    .A2(_0911_),
    .A1(_0909_));
 sg13g2_inv_1 _3506_ (.Y(_0916_),
    .A(_0915_));
 sg13g2_nand4_1 _3507_ (.B(_1991_),
    .C(_2011_),
    .A(_0546_),
    .Y(_0917_),
    .D(net73));
 sg13g2_a21oi_1 _3508_ (.A1(_1992_),
    .A2(net73),
    .Y(_0918_),
    .B1(net74));
 sg13g2_nand3_1 _3509_ (.B(_2014_),
    .C(_0918_),
    .A(_0917_),
    .Y(_0919_));
 sg13g2_inv_1 _3510_ (.Y(_0920_),
    .A(_0919_));
 sg13g2_nor2_1 _3511_ (.A(_0290_),
    .B(_0614_),
    .Y(_0921_));
 sg13g2_a22oi_1 _3512_ (.Y(_0922_),
    .B1(_0862_),
    .B2(_0441_),
    .A2(_0442_),
    .A1(_0603_));
 sg13g2_o21ai_1 _3513_ (.B1(_0922_),
    .Y(_0923_),
    .A1(_0051_),
    .A2(_0296_));
 sg13g2_nor4_1 _3514_ (.A(_0311_),
    .B(_0901_),
    .C(_0921_),
    .D(_0923_),
    .Y(_0924_));
 sg13g2_nor2b_1 _3515_ (.A(\vga.score_l_unit_pixels[2] ),
    .B_N(_0905_),
    .Y(_0925_));
 sg13g2_nor4_1 _3516_ (.A(_0916_),
    .B(_0920_),
    .C(_0924_),
    .D(_0925_),
    .Y(_0926_));
 sg13g2_nand2_1 _3517_ (.Y(_0927_),
    .A(_0908_),
    .B(_0926_));
 sg13g2_nand4_1 _3518_ (.B(_0915_),
    .C(\vga.score_l_ten_enable ),
    .A(_0924_),
    .Y(_0928_),
    .D(_0919_));
 sg13g2_nand3_1 _3519_ (.B(_0927_),
    .C(_0928_),
    .A(_0855_),
    .Y(_0929_));
 sg13g2_nor3_1 _3520_ (.A(_0527_),
    .B(_0618_),
    .C(_0929_),
    .Y(_0930_));
 sg13g2_nor3_1 _3521_ (.A(\vga.blank_h ),
    .B(\vga.blank_v ),
    .C(net55),
    .Y(_0122_));
 sg13g2_nor2b_1 _3522_ (.A(_0930_),
    .B_N(_0122_),
    .Y(_0191_));
 sg13g2_nor2_1 _3523_ (.A(_0263_),
    .B(_0264_),
    .Y(_0193_));
 sg13g2_nor2_1 _3524_ (.A(_0265_),
    .B(_0266_),
    .Y(_0195_));
 sg13g2_buf_1 _3525_ (.A(\vga.ball_angle[0] ),
    .X(_0931_));
 sg13g2_inv_1 _3526_ (.Y(_0932_),
    .A(_0931_));
 sg13g2_nand2_1 _3527_ (.Y(_0933_),
    .A(_1580_),
    .B(_1828_));
 sg13g2_inv_1 _3528_ (.Y(_0934_),
    .A(_0933_));
 sg13g2_nor2_1 _3529_ (.A(_1828_),
    .B(_1836_),
    .Y(_0935_));
 sg13g2_nor2_1 _3530_ (.A(_0934_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_buf_2 _3531_ (.A(_0936_),
    .X(_0937_));
 sg13g2_inv_2 _3532_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_inv_1 _3533_ (.Y(_0939_),
    .A(_0064_));
 sg13g2_nand2_1 _3534_ (.Y(_0940_),
    .A(_1823_),
    .B(_0939_));
 sg13g2_inv_1 _3535_ (.Y(_0941_),
    .A(_1837_));
 sg13g2_nand3_1 _3536_ (.B(_1801_),
    .C(_0941_),
    .A(_1754_),
    .Y(_0942_));
 sg13g2_o21ai_1 _3537_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0940_),
    .A2(_1887_));
 sg13g2_nor2_1 _3538_ (.A(_1580_),
    .B(_1554_),
    .Y(_0944_));
 sg13g2_inv_1 _3539_ (.Y(_0945_),
    .A(_0944_));
 sg13g2_nor2_1 _3540_ (.A(_1624_),
    .B(net51),
    .Y(_0946_));
 sg13g2_a21oi_1 _3541_ (.A1(_1554_),
    .A2(_0946_),
    .Y(_0947_),
    .B1(net48));
 sg13g2_o21ai_1 _3542_ (.B1(_0947_),
    .Y(_0948_),
    .A1(_0939_),
    .A2(_0945_));
 sg13g2_nor2_1 _3543_ (.A(_0943_),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_inv_2 _3544_ (.Y(_0950_),
    .A(_0949_));
 sg13g2_nor2_2 _3545_ (.A(_0938_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_buf_1 _3546_ (.A(net65),
    .X(_0952_));
 sg13g2_a21oi_1 _3547_ (.A1(_0951_),
    .A2(_0084_),
    .Y(_0953_),
    .B1(net54));
 sg13g2_o21ai_1 _3548_ (.B1(_0953_),
    .Y(_0093_),
    .A1(_0932_),
    .A2(_0951_));
 sg13g2_inv_1 _3549_ (.Y(_0954_),
    .A(\vga.ball_angle[1] ));
 sg13g2_buf_1 _3550_ (.A(_0949_),
    .X(_0955_));
 sg13g2_nand2_1 _3551_ (.Y(_0956_),
    .A(_1837_),
    .B(_1584_));
 sg13g2_nand2_1 _3552_ (.Y(_0957_),
    .A(_0955_),
    .B(_0956_));
 sg13g2_nor3_1 _3553_ (.A(_0954_),
    .B(_0931_),
    .C(_0957_),
    .Y(_0958_));
 sg13g2_a21oi_1 _3554_ (.A1(_0951_),
    .A2(_0932_),
    .Y(_0959_),
    .B1(\vga.ball_angle[1] ));
 sg13g2_nor3_1 _3555_ (.A(net52),
    .B(_0958_),
    .C(_0959_),
    .Y(_0094_));
 sg13g2_nor2_1 _3556_ (.A(\vga.ball_angle[1] ),
    .B(_0931_),
    .Y(_0960_));
 sg13g2_xnor2_1 _3557_ (.Y(_0961_),
    .A(_0063_),
    .B(_0960_));
 sg13g2_buf_1 _3558_ (.A(net79),
    .X(_0962_));
 sg13g2_o21ai_1 _3559_ (.B1(net60),
    .Y(_0963_),
    .A1(\vga.ball_angle[2] ),
    .A2(_0951_));
 sg13g2_a21oi_1 _3560_ (.A1(_0951_),
    .A2(_0961_),
    .Y(_0095_),
    .B1(_0963_));
 sg13g2_buf_1 _3561_ (.A(_0950_),
    .X(_0964_));
 sg13g2_inv_1 _3562_ (.Y(_0965_),
    .A(_0960_));
 sg13g2_nand2_1 _3563_ (.Y(_0966_),
    .A(_0965_),
    .B(\vga.ball_angle[2] ));
 sg13g2_xor2_1 _3564_ (.B(_0966_),
    .A(_0049_),
    .X(_0967_));
 sg13g2_buf_1 _3565_ (.A(\vga.ball_angle[3] ),
    .X(_0968_));
 sg13g2_inv_2 _3566_ (.Y(_0969_),
    .A(_0968_));
 sg13g2_nor2b_1 _3567_ (.A(_0965_),
    .B_N(_0063_),
    .Y(_0970_));
 sg13g2_xnor2_1 _3568_ (.Y(_0971_),
    .A(\vga.ball_ratio[2] ),
    .B(\vga.ball_angle[2] ));
 sg13g2_xnor2_1 _3569_ (.Y(_0972_),
    .A(\vga.ball_angle[1] ),
    .B(\vga.ball_ratio[1] ));
 sg13g2_buf_1 _3570_ (.A(\vga.ball_ratio[0] ),
    .X(_0973_));
 sg13g2_xnor2_1 _3571_ (.Y(_0974_),
    .A(_0931_),
    .B(_0973_));
 sg13g2_nand3_1 _3572_ (.B(_0972_),
    .C(_0974_),
    .A(_0971_),
    .Y(_0975_));
 sg13g2_buf_1 _3573_ (.A(_0975_),
    .X(_0976_));
 sg13g2_nor2_2 _3574_ (.A(_0970_),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_inv_1 _3575_ (.Y(_0978_),
    .A(_0977_));
 sg13g2_a21oi_1 _3576_ (.A1(_0969_),
    .A2(_0978_),
    .Y(_0979_),
    .B1(_0937_));
 sg13g2_nand4_1 _3577_ (.B(_1485_),
    .C(_1714_),
    .A(net66),
    .Y(_0980_),
    .D(_1430_));
 sg13g2_nand2_1 _3578_ (.Y(_0981_),
    .A(_0708_),
    .B(net69));
 sg13g2_nor3_1 _3579_ (.A(net70),
    .B(_0980_),
    .C(_0981_),
    .Y(_0982_));
 sg13g2_inv_1 _3580_ (.Y(_0983_),
    .A(_0982_));
 sg13g2_nor2_1 _3581_ (.A(_0968_),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_nor4_1 _3582_ (.A(net66),
    .B(_0791_),
    .C(_1714_),
    .D(_0762_),
    .Y(_0985_));
 sg13g2_nor2_1 _3583_ (.A(_0792_),
    .B(_0985_),
    .Y(_0986_));
 sg13g2_nand2_1 _3584_ (.Y(_0987_),
    .A(_0986_),
    .B(_0968_));
 sg13g2_nand3b_1 _3585_ (.B(_0987_),
    .C(_0977_),
    .Y(_0988_),
    .A_N(_0984_));
 sg13g2_a22oi_1 _3586_ (.Y(_0989_),
    .B1(_0979_),
    .B2(_0988_),
    .A2(_0967_),
    .A1(_0937_));
 sg13g2_buf_1 _3587_ (.A(_0950_),
    .X(_0990_));
 sg13g2_buf_1 _3588_ (.A(_0968_),
    .X(_0991_));
 sg13g2_buf_1 _3589_ (.A(net65),
    .X(_0992_));
 sg13g2_a21oi_1 _3590_ (.A1(net31),
    .A2(net59),
    .Y(_0993_),
    .B1(net53));
 sg13g2_o21ai_1 _3591_ (.B1(_0993_),
    .Y(_0096_),
    .A1(net32),
    .A2(_0989_));
 sg13g2_nor2_1 _3592_ (.A(_1615_),
    .B(_0942_),
    .Y(_0994_));
 sg13g2_a21oi_1 _3593_ (.A1(_0944_),
    .A2(net50),
    .Y(_0995_),
    .B1(net82));
 sg13g2_buf_1 _3594_ (.A(net79),
    .X(_0996_));
 sg13g2_o21ai_1 _3595_ (.B1(net58),
    .Y(_0097_),
    .A1(_0994_),
    .A2(_0995_));
 sg13g2_nand2_1 _3596_ (.Y(_0997_),
    .A(net31),
    .B(_1565_));
 sg13g2_buf_1 _3597_ (.A(_0045_),
    .X(_0998_));
 sg13g2_nand2_1 _3598_ (.Y(_0999_),
    .A(net36),
    .B(_0998_));
 sg13g2_nand4_1 _3599_ (.B(_0957_),
    .C(_0999_),
    .A(_0997_),
    .Y(_0098_),
    .D(net60));
 sg13g2_a21oi_1 _3600_ (.A1(net32),
    .A2(net61),
    .Y(_1000_),
    .B1(net52));
 sg13g2_nor2_1 _3601_ (.A(_1565_),
    .B(_1810_),
    .Y(_1001_));
 sg13g2_inv_1 _3602_ (.Y(_1002_),
    .A(_1567_));
 sg13g2_nor3_1 _3603_ (.A(net82),
    .B(_1001_),
    .C(_1002_),
    .Y(_1003_));
 sg13g2_nand3_1 _3604_ (.B(_1834_),
    .C(_1832_),
    .A(_1811_),
    .Y(_1004_));
 sg13g2_buf_1 _3605_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nor2_1 _3606_ (.A(_1001_),
    .B(_1002_),
    .Y(_1006_));
 sg13g2_a21oi_1 _3607_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1007_),
    .B1(_1828_));
 sg13g2_buf_1 _3608_ (.A(net36),
    .X(_1008_));
 sg13g2_o21ai_1 _3609_ (.B1(net30),
    .Y(_1009_),
    .A1(_1003_),
    .A2(_1007_));
 sg13g2_nand2_1 _3610_ (.Y(_0099_),
    .A(_1000_),
    .B(_1009_));
 sg13g2_nor2_1 _3611_ (.A(net82),
    .B(_1567_),
    .Y(_1010_));
 sg13g2_a21oi_1 _3612_ (.A1(net82),
    .A2(_1001_),
    .Y(_1011_),
    .B1(_1010_));
 sg13g2_nor3_1 _3613_ (.A(_1563_),
    .B(_1011_),
    .C(_0950_),
    .Y(_1012_));
 sg13g2_nor3_1 _3614_ (.A(net55),
    .B(_0951_),
    .C(_1012_),
    .Y(_1013_));
 sg13g2_o21ai_1 _3615_ (.B1(_1563_),
    .Y(_1014_),
    .A1(_1011_),
    .A2(net31));
 sg13g2_nand2_1 _3616_ (.Y(_0100_),
    .A(_1013_),
    .B(_1014_));
 sg13g2_a21oi_1 _3617_ (.A1(net32),
    .A2(_1562_),
    .Y(_1015_),
    .B1(net54));
 sg13g2_inv_1 _3618_ (.Y(_1016_),
    .A(_1562_));
 sg13g2_a21oi_1 _3619_ (.A1(_0809_),
    .A2(_0998_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_a21oi_1 _3620_ (.A1(_0800_),
    .A2(_0998_),
    .Y(_1018_),
    .B1(_1017_));
 sg13g2_nand2_1 _3621_ (.Y(_1019_),
    .A(_1018_),
    .B(net82));
 sg13g2_nor2_1 _3622_ (.A(_0998_),
    .B(_0629_),
    .Y(_1020_));
 sg13g2_xnor2_1 _3623_ (.Y(_1021_),
    .A(_1562_),
    .B(_1020_));
 sg13g2_nand2_1 _3624_ (.Y(_1022_),
    .A(_0934_),
    .B(_1021_));
 sg13g2_nand3_1 _3625_ (.B(_1019_),
    .C(_1022_),
    .A(net36),
    .Y(_1023_));
 sg13g2_nand2_1 _3626_ (.Y(_0101_),
    .A(_1015_),
    .B(_1023_));
 sg13g2_nand2_1 _3627_ (.Y(_1024_),
    .A(_1001_),
    .B(_0798_));
 sg13g2_xnor2_1 _3628_ (.Y(_1025_),
    .A(net80),
    .B(_1024_));
 sg13g2_a22oi_1 _3629_ (.Y(_1026_),
    .B1(_0673_),
    .B2(_0934_),
    .A2(_1025_),
    .A1(_1561_));
 sg13g2_o21ai_1 _3630_ (.B1(_0962_),
    .Y(_1027_),
    .A1(net80),
    .A2(net36));
 sg13g2_a21oi_1 _3631_ (.A1(net30),
    .A2(_1026_),
    .Y(_0102_),
    .B1(_1027_));
 sg13g2_inv_1 _3632_ (.Y(_1028_),
    .A(_0998_));
 sg13g2_nand2_1 _3633_ (.Y(_1029_),
    .A(_0632_),
    .B(_1028_));
 sg13g2_xnor2_1 _3634_ (.Y(_1030_),
    .A(_1576_),
    .B(_1029_));
 sg13g2_nand2_1 _3635_ (.Y(_1031_),
    .A(_0802_),
    .B(_1809_));
 sg13g2_o21ai_1 _3636_ (.B1(_1576_),
    .Y(_1032_),
    .A1(_1574_),
    .A2(_1024_));
 sg13g2_nand3_1 _3637_ (.B(_1005_),
    .C(_1032_),
    .A(_1031_),
    .Y(_1033_));
 sg13g2_a22oi_1 _3638_ (.Y(_1034_),
    .B1(_1561_),
    .B2(_1033_),
    .A2(_0934_),
    .A1(_1030_));
 sg13g2_a21oi_1 _3639_ (.A1(net31),
    .A2(_1576_),
    .Y(_1035_),
    .B1(_0992_));
 sg13g2_o21ai_1 _3640_ (.B1(_1035_),
    .Y(_0103_),
    .A1(net32),
    .A2(_1034_));
 sg13g2_a21oi_1 _3641_ (.A1(_0964_),
    .A2(_1577_),
    .Y(_1036_),
    .B1(net54));
 sg13g2_nand2_1 _3642_ (.Y(_1037_),
    .A(_0622_),
    .B(_1002_));
 sg13g2_xnor2_1 _3643_ (.Y(_1038_),
    .A(_0620_),
    .B(_1037_));
 sg13g2_nor2_1 _3644_ (.A(_1038_),
    .B(_0933_),
    .Y(_1039_));
 sg13g2_xnor2_1 _3645_ (.Y(_1040_),
    .A(_0620_),
    .B(_1031_));
 sg13g2_a21oi_1 _3646_ (.A1(_1040_),
    .A2(_1005_),
    .Y(_1041_),
    .B1(_1828_));
 sg13g2_o21ai_1 _3647_ (.B1(net30),
    .Y(_1042_),
    .A1(_1039_),
    .A2(_1041_));
 sg13g2_nand2_1 _3648_ (.Y(_0104_),
    .A(_1036_),
    .B(_1042_));
 sg13g2_nor2_1 _3649_ (.A(_1028_),
    .B(_0829_),
    .Y(_1043_));
 sg13g2_xnor2_1 _3650_ (.Y(_1044_),
    .A(_0046_),
    .B(_1043_));
 sg13g2_a21oi_1 _3651_ (.A1(_0627_),
    .A2(_1028_),
    .Y(_1045_),
    .B1(_1569_));
 sg13g2_a21oi_1 _3652_ (.A1(_0624_),
    .A2(_1028_),
    .Y(_1046_),
    .B1(_1045_));
 sg13g2_a22oi_1 _3653_ (.Y(_1047_),
    .B1(_1828_),
    .B2(_1046_),
    .A2(_0935_),
    .A1(_1044_));
 sg13g2_o21ai_1 _3654_ (.B1(net79),
    .Y(_1048_),
    .A1(_1569_),
    .A2(_0955_));
 sg13g2_a21oi_1 _3655_ (.A1(net30),
    .A2(_1047_),
    .Y(_0105_),
    .B1(_1048_));
 sg13g2_nor2_1 _3656_ (.A(_1024_),
    .B(_1835_),
    .Y(_1049_));
 sg13g2_xnor2_1 _3657_ (.Y(_1050_),
    .A(_0047_),
    .B(_1049_));
 sg13g2_a21oi_1 _3658_ (.A1(net62),
    .A2(_0645_),
    .Y(_1051_),
    .B1(_0933_));
 sg13g2_nand2_1 _3659_ (.Y(_1052_),
    .A(_0647_),
    .B(_1565_));
 sg13g2_a22oi_1 _3660_ (.Y(_1053_),
    .B1(_1051_),
    .B2(_1052_),
    .A2(_1050_),
    .A1(_0935_));
 sg13g2_o21ai_1 _3661_ (.B1(net79),
    .Y(_1054_),
    .A1(net81),
    .A2(net36));
 sg13g2_a21oi_1 _3662_ (.A1(_1008_),
    .A2(_1053_),
    .Y(_0106_),
    .B1(_1054_));
 sg13g2_a21oi_1 _3663_ (.A1(_0964_),
    .A2(_1571_),
    .Y(_1055_),
    .B1(net54));
 sg13g2_a21oi_1 _3664_ (.A1(_0839_),
    .A2(_1809_),
    .Y(_1056_),
    .B1(_1572_));
 sg13g2_a21oi_1 _3665_ (.A1(_1832_),
    .A2(_1049_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_a21oi_1 _3666_ (.A1(_1057_),
    .A2(_1005_),
    .Y(_1058_),
    .B1(_1828_));
 sg13g2_nor2_1 _3667_ (.A(_0998_),
    .B(_0643_),
    .Y(_1059_));
 sg13g2_xor2_1 _3668_ (.B(_1059_),
    .A(_0048_),
    .X(_1060_));
 sg13g2_nor2_1 _3669_ (.A(_0933_),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_o21ai_1 _3670_ (.B1(_1008_),
    .Y(_1062_),
    .A1(_1058_),
    .A2(_1061_));
 sg13g2_nand2_1 _3671_ (.Y(_0107_),
    .A(_1055_),
    .B(_1062_));
 sg13g2_a21oi_1 _3672_ (.A1(net32),
    .A2(_1447_),
    .Y(_1063_),
    .B1(net54));
 sg13g2_inv_1 _3673_ (.Y(_1064_),
    .A(_0986_));
 sg13g2_a21oi_1 _3674_ (.A1(_1064_),
    .A2(_0968_),
    .Y(_1065_),
    .B1(_0978_));
 sg13g2_inv_1 _3675_ (.Y(_1066_),
    .A(_1065_));
 sg13g2_nor2_1 _3676_ (.A(_0984_),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_inv_1 _3677_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_o21ai_1 _3678_ (.B1(_0938_),
    .Y(_1069_),
    .A1(net69),
    .A2(_1066_));
 sg13g2_a21oi_1 _3679_ (.A1(net69),
    .A2(_1068_),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_nand2_1 _3680_ (.Y(_1071_),
    .A(net49),
    .B(_1449_));
 sg13g2_o21ai_1 _3681_ (.B1(_1071_),
    .Y(_1072_),
    .A1(_1749_),
    .A2(net51));
 sg13g2_o21ai_1 _3682_ (.B1(net30),
    .Y(_1073_),
    .A1(_1070_),
    .A2(_1072_));
 sg13g2_nand2_1 _3683_ (.Y(_0108_),
    .A(_1063_),
    .B(_1073_));
 sg13g2_nor2_1 _3684_ (.A(net88),
    .B(_1447_),
    .Y(_1074_));
 sg13g2_nand2_1 _3685_ (.Y(_1075_),
    .A(net88),
    .B(net87));
 sg13g2_nand2b_1 _3686_ (.Y(_1076_),
    .B(_1075_),
    .A_N(_1074_));
 sg13g2_nand3_1 _3687_ (.B(_0969_),
    .C(_1076_),
    .A(_0983_),
    .Y(_1077_));
 sg13g2_o21ai_1 _3688_ (.B1(_1077_),
    .Y(_1078_),
    .A1(_1076_),
    .A2(_0987_));
 sg13g2_a22oi_1 _3689_ (.Y(_1079_),
    .B1(net88),
    .B2(_1068_),
    .A2(_1078_),
    .A1(_0977_));
 sg13g2_nand2b_1 _3690_ (.Y(_1080_),
    .B(_0938_),
    .A_N(_1079_));
 sg13g2_a22oi_1 _3691_ (.Y(_1081_),
    .B1(_1445_),
    .B2(net49),
    .A2(_1725_),
    .A1(_1582_));
 sg13g2_a21oi_1 _3692_ (.A1(_1080_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(net31));
 sg13g2_a21oi_1 _3693_ (.A1(net31),
    .A2(net88),
    .Y(_1083_),
    .B1(_0952_));
 sg13g2_nand2b_1 _3694_ (.Y(_0109_),
    .B(_1083_),
    .A_N(_1082_));
 sg13g2_inv_1 _3695_ (.Y(_1084_),
    .A(_1453_));
 sg13g2_nand2_1 _3696_ (.Y(_1085_),
    .A(_0983_),
    .B(_1074_));
 sg13g2_nand2_1 _3697_ (.Y(_1086_),
    .A(_1085_),
    .B(_0969_));
 sg13g2_nand2_1 _3698_ (.Y(_1087_),
    .A(_1075_),
    .B(net59));
 sg13g2_nand3_1 _3699_ (.B(_1086_),
    .C(_1087_),
    .A(_1065_),
    .Y(_1088_));
 sg13g2_nor2_1 _3700_ (.A(_1084_),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nor2_1 _3701_ (.A(_0937_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_nand2_1 _3702_ (.Y(_1091_),
    .A(_1088_),
    .B(_1084_));
 sg13g2_nor2_1 _3703_ (.A(_0463_),
    .B(net51),
    .Y(_1092_));
 sg13g2_a221oi_1 _3704_ (.B2(_1091_),
    .C1(_1092_),
    .B1(_1090_),
    .A1(_1456_),
    .Y(_1093_),
    .A2(net49));
 sg13g2_a21oi_1 _3705_ (.A1(net31),
    .A2(_1453_),
    .Y(_1094_),
    .B1(net53));
 sg13g2_o21ai_1 _3706_ (.B1(_1094_),
    .Y(_0110_),
    .A1(net32),
    .A2(_1093_));
 sg13g2_nor2_1 _3707_ (.A(net86),
    .B(_1085_),
    .Y(_1095_));
 sg13g2_inv_1 _3708_ (.Y(_1096_),
    .A(_1095_));
 sg13g2_nand3_1 _3709_ (.B(net87),
    .C(net59),
    .A(_1443_),
    .Y(_1097_));
 sg13g2_a221oi_1 _3710_ (.B2(_1097_),
    .C1(_1066_),
    .B1(_1096_),
    .A1(_1084_),
    .Y(_1098_),
    .A2(_0991_));
 sg13g2_xnor2_1 _3711_ (.Y(_1099_),
    .A(_1521_),
    .B(_1098_));
 sg13g2_nor2_1 _3712_ (.A(_0462_),
    .B(net51),
    .Y(_1100_));
 sg13g2_a221oi_1 _3713_ (.B2(_0938_),
    .C1(_1100_),
    .B1(_1099_),
    .A1(_1416_),
    .Y(_1101_),
    .A2(net49));
 sg13g2_a21oi_1 _3714_ (.A1(net31),
    .A2(_1465_),
    .Y(_1102_),
    .B1(_0992_));
 sg13g2_o21ai_1 _3715_ (.B1(_1102_),
    .Y(_0111_),
    .A1(net32),
    .A2(_1101_));
 sg13g2_o21ai_1 _3716_ (.B1(net59),
    .Y(_1103_),
    .A1(net69),
    .A2(_0760_));
 sg13g2_nand2_1 _3717_ (.Y(_1104_),
    .A(_0981_),
    .B(_0969_));
 sg13g2_nand3_1 _3718_ (.B(_1103_),
    .C(_1104_),
    .A(_1067_),
    .Y(_1105_));
 sg13g2_xnor2_1 _3719_ (.Y(_1106_),
    .A(_1439_),
    .B(_1105_));
 sg13g2_nor2_1 _3720_ (.A(_1676_),
    .B(net51),
    .Y(_1107_));
 sg13g2_a221oi_1 _3721_ (.B2(_0938_),
    .C1(_1107_),
    .B1(_1106_),
    .A1(_1420_),
    .Y(_1108_),
    .A2(net49));
 sg13g2_o21ai_1 _3722_ (.B1(net79),
    .Y(_1109_),
    .A1(net70),
    .A2(net36));
 sg13g2_a21oi_1 _3723_ (.A1(net30),
    .A2(_1108_),
    .Y(_0112_),
    .B1(_1109_));
 sg13g2_nor2_1 _3724_ (.A(net70),
    .B(_0981_),
    .Y(_1110_));
 sg13g2_nand2_1 _3725_ (.Y(_1111_),
    .A(_1110_),
    .B(_0980_));
 sg13g2_a21oi_1 _3726_ (.A1(_1111_),
    .A2(_0969_),
    .Y(_1112_),
    .B1(_0978_));
 sg13g2_nor3_1 _3727_ (.A(_1485_),
    .B(net59),
    .C(_1111_),
    .Y(_1113_));
 sg13g2_nand2b_1 _3728_ (.Y(_1114_),
    .B(_0968_),
    .A_N(_0792_));
 sg13g2_a21oi_1 _3729_ (.A1(_0761_),
    .A2(net87),
    .Y(_1115_),
    .B1(net67));
 sg13g2_nor3_1 _3730_ (.A(_1485_),
    .B(net69),
    .C(_0762_),
    .Y(_1116_));
 sg13g2_nor3_1 _3731_ (.A(_1115_),
    .B(_1116_),
    .C(_0985_),
    .Y(_1117_));
 sg13g2_nor2_1 _3732_ (.A(_1114_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_o21ai_1 _3733_ (.B1(_0977_),
    .Y(_1119_),
    .A1(_1113_),
    .A2(_1118_));
 sg13g2_o21ai_1 _3734_ (.B1(_1119_),
    .Y(_1120_),
    .A1(_1471_),
    .A2(_1112_));
 sg13g2_nand2_1 _3735_ (.Y(_1121_),
    .A(_1120_),
    .B(_0938_));
 sg13g2_a22oi_1 _3736_ (.Y(_1122_),
    .B1(_1472_),
    .B2(_0941_),
    .A2(_1582_),
    .A1(_1705_));
 sg13g2_nand3_1 _3737_ (.B(_1121_),
    .C(_1122_),
    .A(net36),
    .Y(_1123_));
 sg13g2_nand2_1 _3738_ (.Y(_1124_),
    .A(net32),
    .B(_1471_));
 sg13g2_nand3_1 _3739_ (.B(_1124_),
    .C(net60),
    .A(_1123_),
    .Y(_0113_));
 sg13g2_nand2_1 _3740_ (.Y(_1125_),
    .A(_1116_),
    .B(net84));
 sg13g2_nand2b_1 _3741_ (.Y(_1126_),
    .B(_1714_),
    .A_N(_1116_));
 sg13g2_a21oi_1 _3742_ (.A1(_1125_),
    .A2(_1126_),
    .Y(_1127_),
    .B1(_0987_));
 sg13g2_nor2_1 _3743_ (.A(_0978_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nand2_1 _3744_ (.Y(_1129_),
    .A(_0746_),
    .B(_1521_));
 sg13g2_nor3_1 _3745_ (.A(net84),
    .B(_1129_),
    .C(_1096_),
    .Y(_1130_));
 sg13g2_o21ai_1 _3746_ (.B1(net84),
    .Y(_1131_),
    .A1(_1129_),
    .A2(_1096_));
 sg13g2_nand3b_1 _3747_ (.B(_1131_),
    .C(_0969_),
    .Y(_1132_),
    .A_N(_1130_));
 sg13g2_a22oi_1 _3748_ (.Y(_1133_),
    .B1(_1128_),
    .B2(_1132_),
    .A2(_0978_),
    .A1(_1489_));
 sg13g2_nand2b_1 _3749_ (.Y(_1134_),
    .B(_0938_),
    .A_N(_1133_));
 sg13g2_a22oi_1 _3750_ (.Y(_1135_),
    .B1(_1425_),
    .B2(net49),
    .A2(_1682_),
    .A1(_1582_));
 sg13g2_a21oi_1 _3751_ (.A1(_1134_),
    .A2(_1135_),
    .Y(_1136_),
    .B1(_0950_));
 sg13g2_a21oi_1 _3752_ (.A1(net84),
    .A2(_0990_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_buf_1 _3753_ (.A(net79),
    .X(_1138_));
 sg13g2_nand2_1 _3754_ (.Y(_0114_),
    .A(_1137_),
    .B(net57));
 sg13g2_a21oi_1 _3755_ (.A1(_0990_),
    .A2(_1413_),
    .Y(_1139_),
    .B1(net54));
 sg13g2_xnor2_1 _3756_ (.Y(_1140_),
    .A(net66),
    .B(_1130_));
 sg13g2_xnor2_1 _3757_ (.Y(_1141_),
    .A(net66),
    .B(_1125_));
 sg13g2_nand2_1 _3758_ (.Y(_1142_),
    .A(_1141_),
    .B(net59));
 sg13g2_o21ai_1 _3759_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_0991_),
    .A2(_1140_));
 sg13g2_a221oi_1 _3760_ (.B2(_1065_),
    .C1(_0956_),
    .B1(_1143_),
    .A1(_1516_),
    .Y(_1144_),
    .A2(_0978_));
 sg13g2_nand2_1 _3761_ (.Y(_1145_),
    .A(net49),
    .B(_1414_));
 sg13g2_o21ai_1 _3762_ (.B1(_1145_),
    .Y(_1146_),
    .A1(net64),
    .A2(_1584_));
 sg13g2_o21ai_1 _3763_ (.B1(net30),
    .Y(_1147_),
    .A1(_1144_),
    .A2(_1146_));
 sg13g2_nand2_1 _3764_ (.Y(_0115_),
    .A(_1139_),
    .B(_1147_));
 sg13g2_nor4_1 _3765_ (.A(_1430_),
    .B(net87),
    .C(_0747_),
    .D(_0709_),
    .Y(_1148_));
 sg13g2_o21ai_1 _3766_ (.B1(_0977_),
    .Y(_1149_),
    .A1(net59),
    .A2(_1148_));
 sg13g2_o21ai_1 _3767_ (.B1(_0791_),
    .Y(_1150_),
    .A1(net69),
    .A2(_0787_));
 sg13g2_nand2_1 _3768_ (.Y(_1151_),
    .A(_1150_),
    .B(net59));
 sg13g2_nand3_1 _3769_ (.B(_0791_),
    .C(_0969_),
    .A(_1148_),
    .Y(_1152_));
 sg13g2_nand2_1 _3770_ (.Y(_1153_),
    .A(_1151_),
    .B(_1152_));
 sg13g2_a22oi_1 _3771_ (.Y(_1154_),
    .B1(_0977_),
    .B2(_1153_),
    .A2(_1149_),
    .A1(net83));
 sg13g2_nor2_1 _3772_ (.A(_0937_),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_a221oi_1 _3773_ (.B2(net49),
    .C1(_1155_),
    .B1(_1432_),
    .A1(\vga.paddle_l_pos_v[8] ),
    .Y(_1156_),
    .A2(_1582_));
 sg13g2_o21ai_1 _3774_ (.B1(_1660_),
    .Y(_1157_),
    .A1(_1493_),
    .A2(net36));
 sg13g2_a21oi_1 _3775_ (.A1(net30),
    .A2(_1156_),
    .Y(_0116_),
    .B1(_1157_));
 sg13g2_nor3_2 _3776_ (.A(_0937_),
    .B(_0970_),
    .C(net48),
    .Y(_1158_));
 sg13g2_a21oi_1 _3777_ (.A1(_1158_),
    .A2(_0976_),
    .Y(_1159_),
    .B1(_0973_));
 sg13g2_a21oi_1 _3778_ (.A1(_1158_),
    .A2(_0973_),
    .Y(_1160_),
    .B1(_0273_));
 sg13g2_nor2b_1 _3779_ (.A(_1159_),
    .B_N(_1160_),
    .Y(_0117_));
 sg13g2_a21oi_1 _3780_ (.A1(_1158_),
    .A2(_0973_),
    .Y(_1161_),
    .B1(\vga.ball_ratio[1] ));
 sg13g2_nand2_1 _3781_ (.Y(_1162_),
    .A(_0973_),
    .B(\vga.ball_ratio[1] ));
 sg13g2_inv_1 _3782_ (.Y(_1163_),
    .A(_1158_));
 sg13g2_a21oi_1 _3783_ (.A1(_0976_),
    .A2(_1162_),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_nor3_1 _3784_ (.A(_0274_),
    .B(_1161_),
    .C(_1164_),
    .Y(_0118_));
 sg13g2_nand4_1 _3785_ (.B(_0973_),
    .C(\vga.ball_ratio[1] ),
    .A(_1158_),
    .Y(_1165_),
    .D(_0976_));
 sg13g2_nor2b_1 _3786_ (.A(\vga.ball_ratio[2] ),
    .B_N(_1165_),
    .Y(_1166_));
 sg13g2_a21oi_1 _3787_ (.A1(_1164_),
    .A2(\vga.ball_ratio[2] ),
    .Y(_1167_),
    .B1(_0273_));
 sg13g2_nor2b_1 _3788_ (.A(_1166_),
    .B_N(_1167_),
    .Y(_0119_));
 sg13g2_inv_1 _3789_ (.Y(_1168_),
    .A(\vga.blank_h ));
 sg13g2_nand2_1 _3790_ (.Y(_1169_),
    .A(_0865_),
    .B(_0598_));
 sg13g2_nor2_1 _3791_ (.A(net72),
    .B(_1169_),
    .Y(_1170_));
 sg13g2_inv_1 _3792_ (.Y(_1171_),
    .A(_1170_));
 sg13g2_nand2_1 _3793_ (.Y(_1172_),
    .A(_0436_),
    .B(_0058_));
 sg13g2_inv_1 _3794_ (.Y(_1173_),
    .A(_1172_));
 sg13g2_nand2_1 _3795_ (.Y(_1174_),
    .A(_0284_),
    .B(_0285_));
 sg13g2_a21oi_1 _3796_ (.A1(_1171_),
    .A2(_1173_),
    .Y(_1175_),
    .B1(_1174_));
 sg13g2_inv_1 _3797_ (.Y(_1176_),
    .A(_1175_));
 sg13g2_inv_1 _3798_ (.Y(_1177_),
    .A(_0300_));
 sg13g2_nand2_1 _3799_ (.Y(_1178_),
    .A(_0309_),
    .B(_1177_));
 sg13g2_nor2_1 _3800_ (.A(_1176_),
    .B(_1178_),
    .Y(_1179_));
 sg13g2_buf_1 _3801_ (.A(_1179_),
    .X(_1180_));
 sg13g2_a21oi_1 _3802_ (.A1(_0315_),
    .A2(_1177_),
    .Y(_1181_),
    .B1(net53));
 sg13g2_o21ai_1 _3803_ (.B1(_1181_),
    .Y(_0120_),
    .A1(_1168_),
    .A2(net40));
 sg13g2_inv_1 _3804_ (.Y(_1182_),
    .A(\vga.count_v[8] ));
 sg13g2_nand2_1 _3805_ (.Y(_1183_),
    .A(_1983_),
    .B(_1984_));
 sg13g2_nor2_1 _3806_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_inv_1 _3807_ (.Y(_1185_),
    .A(_1184_));
 sg13g2_nor2_1 _3808_ (.A(_1979_),
    .B(_0477_),
    .Y(_1186_));
 sg13g2_inv_1 _3809_ (.Y(_1187_),
    .A(_1186_));
 sg13g2_nor2_1 _3810_ (.A(_1982_),
    .B(_1187_),
    .Y(_1188_));
 sg13g2_nor2_1 _3811_ (.A(net74),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_o21ai_1 _3812_ (.B1(_0433_),
    .Y(_1190_),
    .A1(_1185_),
    .A2(_1189_));
 sg13g2_buf_1 _3813_ (.A(_1190_),
    .X(_1191_));
 sg13g2_inv_1 _3814_ (.Y(_1192_),
    .A(_1191_));
 sg13g2_o21ai_1 _3815_ (.B1(\vga.blank_v ),
    .Y(_1193_),
    .A1(_1176_),
    .A2(_1192_));
 sg13g2_nand4_1 _3816_ (.B(_0913_),
    .C(_1974_),
    .A(_1985_),
    .Y(_1194_),
    .D(_1182_));
 sg13g2_nor2_1 _3817_ (.A(_1186_),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_a21oi_1 _3818_ (.A1(_0448_),
    .A2(_1194_),
    .Y(_1196_),
    .B1(_1195_));
 sg13g2_nand3b_1 _3819_ (.B(_1175_),
    .C(_1191_),
    .Y(_1197_),
    .A_N(_1196_));
 sg13g2_nand3_1 _3820_ (.B(net60),
    .C(_1197_),
    .A(_1193_),
    .Y(_0121_));
 sg13g2_buf_1 _3821_ (.A(_1176_),
    .X(_1198_));
 sg13g2_nand3_1 _3822_ (.B(_0684_),
    .C(_0309_),
    .A(_1198_),
    .Y(_1199_));
 sg13g2_nand2_1 _3823_ (.Y(_1200_),
    .A(_1178_),
    .B(_0036_));
 sg13g2_nand3_1 _3824_ (.B(_1200_),
    .C(net60),
    .A(_1199_),
    .Y(_0123_));
 sg13g2_nand2_1 _3825_ (.Y(_1201_),
    .A(_0609_),
    .B(_0293_));
 sg13g2_o21ai_1 _3826_ (.B1(net58),
    .Y(_0124_),
    .A1(_1201_),
    .A2(net40));
 sg13g2_xnor2_1 _3827_ (.Y(_1202_),
    .A(_0444_),
    .B(_0293_));
 sg13g2_o21ai_1 _3828_ (.B1(net58),
    .Y(_0125_),
    .A1(_1202_),
    .A2(net40));
 sg13g2_inv_1 _3829_ (.Y(_1203_),
    .A(_0297_));
 sg13g2_nand2b_1 _3830_ (.Y(_1204_),
    .B(_1203_),
    .A_N(_0870_));
 sg13g2_o21ai_1 _3831_ (.B1(net58),
    .Y(_0126_),
    .A1(_1204_),
    .A2(net40));
 sg13g2_xnor2_1 _3832_ (.Y(_1205_),
    .A(_0276_),
    .B(_0297_));
 sg13g2_o21ai_1 _3833_ (.B1(net58),
    .Y(_0127_),
    .A1(_1205_),
    .A2(net40));
 sg13g2_xnor2_1 _3834_ (.Y(_1206_),
    .A(_0306_),
    .B(_1169_));
 sg13g2_o21ai_1 _3835_ (.B1(net58),
    .Y(_0128_),
    .A1(_1206_),
    .A2(net40));
 sg13g2_nor2_2 _3836_ (.A(_0277_),
    .B(_1203_),
    .Y(_1207_));
 sg13g2_xnor2_1 _3837_ (.Y(_1208_),
    .A(_0279_),
    .B(_1207_));
 sg13g2_o21ai_1 _3838_ (.B1(net58),
    .Y(_0129_),
    .A1(_1208_),
    .A2(net40));
 sg13g2_a21oi_1 _3839_ (.A1(_1207_),
    .A2(_0279_),
    .Y(_1209_),
    .B1(_0298_));
 sg13g2_a21oi_1 _3840_ (.A1(_0297_),
    .A2(_0283_),
    .Y(_1210_),
    .B1(_1209_));
 sg13g2_o21ai_1 _3841_ (.B1(net58),
    .Y(_0130_),
    .A1(_1210_),
    .A2(_1180_));
 sg13g2_a21oi_1 _3842_ (.A1(_1207_),
    .A2(_0303_),
    .Y(_1211_),
    .B1(_0284_));
 sg13g2_nand3_1 _3843_ (.B(_0284_),
    .C(_0303_),
    .A(_1207_),
    .Y(_1212_));
 sg13g2_nand2b_1 _3844_ (.Y(_1213_),
    .B(_1212_),
    .A_N(_1211_));
 sg13g2_o21ai_1 _3845_ (.B1(_0996_),
    .Y(_0131_),
    .A1(_1213_),
    .A2(net40));
 sg13g2_xnor2_1 _3846_ (.Y(_1214_),
    .A(_0286_),
    .B(_1212_));
 sg13g2_o21ai_1 _3847_ (.B1(net60),
    .Y(_0132_),
    .A1(_1214_),
    .A2(_1180_));
 sg13g2_a21oi_1 _3848_ (.A1(_1191_),
    .A2(_1196_),
    .Y(_1215_),
    .B1(_1176_));
 sg13g2_buf_1 _3849_ (.A(_1215_),
    .X(_1216_));
 sg13g2_nor2_1 _3850_ (.A(_0037_),
    .B(_1191_),
    .Y(_1217_));
 sg13g2_a21oi_1 _3851_ (.A1(net77),
    .A2(_1191_),
    .Y(_1218_),
    .B1(_1217_));
 sg13g2_a22oi_1 _3852_ (.Y(_1219_),
    .B1(net44),
    .B2(_1218_),
    .A2(net46),
    .A1(net77));
 sg13g2_nand2_1 _3853_ (.Y(_0133_),
    .A(_1219_),
    .B(net57));
 sg13g2_nand2_1 _3854_ (.Y(_1220_),
    .A(_2008_),
    .B(_0910_));
 sg13g2_a22oi_1 _3855_ (.Y(_1221_),
    .B1(_1220_),
    .B2(_1216_),
    .A2(_1198_),
    .A1(_1970_));
 sg13g2_nand2_1 _3856_ (.Y(_0134_),
    .A(_1221_),
    .B(net57));
 sg13g2_xnor2_1 _3857_ (.Y(_1222_),
    .A(_0471_),
    .B(_0477_));
 sg13g2_a22oi_1 _3858_ (.Y(_1223_),
    .B1(_1222_),
    .B2(net44),
    .A2(net46),
    .A1(net76));
 sg13g2_nand2_1 _3859_ (.Y(_0135_),
    .A(_1223_),
    .B(_1138_));
 sg13g2_nor2_1 _3860_ (.A(_2004_),
    .B(_0477_),
    .Y(_1224_));
 sg13g2_xnor2_1 _3861_ (.Y(_1225_),
    .A(_0039_),
    .B(_1224_));
 sg13g2_a22oi_1 _3862_ (.Y(_1226_),
    .B1(_1225_),
    .B2(_1216_),
    .A2(net46),
    .A1(_1978_));
 sg13g2_nand2_1 _3863_ (.Y(_0136_),
    .A(_1226_),
    .B(_1138_));
 sg13g2_xnor2_1 _3864_ (.Y(_1227_),
    .A(_0457_),
    .B(_1186_));
 sg13g2_a22oi_1 _3865_ (.Y(_1228_),
    .B1(_1227_),
    .B2(net44),
    .A2(net46),
    .A1(_1981_));
 sg13g2_nand2_1 _3866_ (.Y(_0137_),
    .A(_1228_),
    .B(net57));
 sg13g2_xnor2_1 _3867_ (.Y(_1229_),
    .A(_0455_),
    .B(_1188_));
 sg13g2_a22oi_1 _3868_ (.Y(_1230_),
    .B1(_1229_),
    .B2(net44),
    .A2(net46),
    .A1(net74));
 sg13g2_nand2_1 _3869_ (.Y(_0138_),
    .A(_1230_),
    .B(net57));
 sg13g2_nor2_1 _3870_ (.A(_1993_),
    .B(_1187_),
    .Y(_1231_));
 sg13g2_xnor2_1 _3871_ (.Y(_1232_),
    .A(_0484_),
    .B(_1231_));
 sg13g2_a22oi_1 _3872_ (.Y(_1233_),
    .B1(_1232_),
    .B2(net44),
    .A2(net46),
    .A1(_1984_));
 sg13g2_nand2_1 _3873_ (.Y(_0139_),
    .A(_1233_),
    .B(net57));
 sg13g2_nand2_1 _3874_ (.Y(_1234_),
    .A(_1231_),
    .B(_1984_));
 sg13g2_xnor2_1 _3875_ (.Y(_1235_),
    .A(_0519_),
    .B(_1234_));
 sg13g2_a22oi_1 _3876_ (.Y(_1236_),
    .B1(_1235_),
    .B2(net44),
    .A2(net46),
    .A1(_1983_));
 sg13g2_nand2_1 _3877_ (.Y(_0140_),
    .A(_1236_),
    .B(net57));
 sg13g2_nor3_1 _3878_ (.A(_1993_),
    .B(_1183_),
    .C(_1187_),
    .Y(_1237_));
 sg13g2_xnor2_1 _3879_ (.Y(_1238_),
    .A(net71),
    .B(_1237_));
 sg13g2_a22oi_1 _3880_ (.Y(_1239_),
    .B1(_1238_),
    .B2(net44),
    .A2(net46),
    .A1(\vga.count_v[8] ));
 sg13g2_nand2_1 _3881_ (.Y(_0141_),
    .A(_1239_),
    .B(net57));
 sg13g2_nand2_1 _3882_ (.Y(_1240_),
    .A(_1231_),
    .B(_1184_));
 sg13g2_xnor2_1 _3883_ (.Y(_1241_),
    .A(_0449_),
    .B(_1240_));
 sg13g2_a22oi_1 _3884_ (.Y(_1242_),
    .B1(_1241_),
    .B2(net44),
    .A2(_1176_),
    .A1(_1974_));
 sg13g2_nor2_1 _3885_ (.A(net52),
    .B(_1242_),
    .Y(_0142_));
 sg13g2_inv_1 _3886_ (.Y(_1243_),
    .A(_0082_));
 sg13g2_inv_1 _3887_ (.Y(_1244_),
    .A(\vga.left_up_pressed ));
 sg13g2_nand4_1 _3888_ (.B(_0473_),
    .C(net63),
    .A(_0462_),
    .Y(_1245_),
    .D(_0082_));
 sg13g2_a21oi_1 _3889_ (.A1(_0462_),
    .A2(_0060_),
    .Y(_1246_),
    .B1(_1676_));
 sg13g2_a21oi_1 _3890_ (.A1(_1245_),
    .A2(_1246_),
    .Y(_1247_),
    .B1(_1792_));
 sg13g2_nor2_1 _3891_ (.A(_1244_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_nand2_1 _3892_ (.Y(_1249_),
    .A(_1725_),
    .B(_1727_));
 sg13g2_nor4_1 _3893_ (.A(_1675_),
    .B(net63),
    .C(_0462_),
    .D(_1249_),
    .Y(_1250_));
 sg13g2_nor2_1 _3894_ (.A(_1698_),
    .B(_1740_),
    .Y(_1251_));
 sg13g2_o21ai_1 _3895_ (.B1(_1251_),
    .Y(_1252_),
    .A1(_1706_),
    .A2(_1250_));
 sg13g2_nand2_1 _3896_ (.Y(_1253_),
    .A(_1252_),
    .B(\vga.left_down_pressed ));
 sg13g2_buf_1 _3897_ (.A(_1253_),
    .X(_1254_));
 sg13g2_inv_1 _3898_ (.Y(_1255_),
    .A(_1254_));
 sg13g2_nor2_1 _3899_ (.A(_1248_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_buf_1 _3900_ (.A(_1256_),
    .X(_1257_));
 sg13g2_a21oi_1 _3901_ (.A1(net43),
    .A2(_1727_),
    .Y(_1258_),
    .B1(net53));
 sg13g2_o21ai_1 _3902_ (.B1(_1258_),
    .Y(_0173_),
    .A1(_1243_),
    .A2(net43));
 sg13g2_inv_1 _3903_ (.Y(_1259_),
    .A(_1256_));
 sg13g2_buf_1 _3904_ (.A(_1254_),
    .X(_1260_));
 sg13g2_xnor2_1 _3905_ (.Y(_1261_),
    .A(_1725_),
    .B(_1260_));
 sg13g2_xnor2_1 _3906_ (.Y(_1262_),
    .A(_1243_),
    .B(_1261_));
 sg13g2_a21oi_1 _3907_ (.A1(_1262_),
    .A2(_1259_),
    .Y(_1263_),
    .B1(net53));
 sg13g2_o21ai_1 _3908_ (.B1(_1263_),
    .Y(_0174_),
    .A1(_0473_),
    .A2(_1259_));
 sg13g2_inv_1 _3909_ (.Y(_1264_),
    .A(_1249_));
 sg13g2_a21oi_1 _3910_ (.A1(_1254_),
    .A2(_0428_),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_xnor2_1 _3911_ (.Y(_1266_),
    .A(_1731_),
    .B(_1254_));
 sg13g2_nor2_1 _3912_ (.A(_1265_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_nand2_1 _3913_ (.Y(_1268_),
    .A(_1266_),
    .B(_1265_));
 sg13g2_nand3b_1 _3914_ (.B(_1259_),
    .C(_1268_),
    .Y(_1269_),
    .A_N(_1267_));
 sg13g2_a21oi_1 _3915_ (.A1(net43),
    .A2(_1731_),
    .Y(_1270_),
    .B1(net54));
 sg13g2_nand2_1 _3916_ (.Y(_0175_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_nor2_1 _3917_ (.A(_1677_),
    .B(net47),
    .Y(_1271_));
 sg13g2_nor2_1 _3918_ (.A(_0462_),
    .B(_1255_),
    .Y(_1272_));
 sg13g2_nor2_1 _3919_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_inv_1 _3920_ (.Y(_1274_),
    .A(_0060_));
 sg13g2_a21oi_1 _3921_ (.A1(_1274_),
    .A2(_1254_),
    .Y(_1275_),
    .B1(_1267_));
 sg13g2_xor2_1 _3922_ (.B(_1275_),
    .A(_1273_),
    .X(_1276_));
 sg13g2_a21oi_1 _3923_ (.A1(net43),
    .A2(_1677_),
    .Y(_1277_),
    .B1(net53));
 sg13g2_o21ai_1 _3924_ (.B1(_1277_),
    .Y(_0176_),
    .A1(net43),
    .A2(_1276_));
 sg13g2_xnor2_1 _3925_ (.Y(_1278_),
    .A(_1675_),
    .B(net47));
 sg13g2_nor2_1 _3926_ (.A(_1271_),
    .B(_1275_),
    .Y(_1279_));
 sg13g2_nor2_1 _3927_ (.A(_1272_),
    .B(_1279_),
    .Y(_1280_));
 sg13g2_nor2_1 _3928_ (.A(_1278_),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_inv_1 _3929_ (.Y(_1282_),
    .A(_1281_));
 sg13g2_nand2_1 _3930_ (.Y(_1283_),
    .A(_1280_),
    .B(_1278_));
 sg13g2_nand3_1 _3931_ (.B(_1259_),
    .C(_1283_),
    .A(_1282_),
    .Y(_1284_));
 sg13g2_nand2_1 _3932_ (.Y(_1285_),
    .A(net43),
    .B(_1675_));
 sg13g2_a21oi_1 _3933_ (.A1(_1284_),
    .A2(_1285_),
    .Y(_0177_),
    .B1(_0274_));
 sg13g2_xnor2_1 _3934_ (.Y(_1286_),
    .A(_1705_),
    .B(net47));
 sg13g2_inv_1 _3935_ (.Y(_1287_),
    .A(_1286_));
 sg13g2_nand2b_1 _3936_ (.Y(_1288_),
    .B(net47),
    .A_N(_0059_));
 sg13g2_nand2_1 _3937_ (.Y(_1289_),
    .A(_1282_),
    .B(_1288_));
 sg13g2_inv_1 _3938_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_nor2_1 _3939_ (.A(_1287_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_inv_1 _3940_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nand2_1 _3941_ (.Y(_1293_),
    .A(_1290_),
    .B(_1287_));
 sg13g2_nand3_1 _3942_ (.B(_1259_),
    .C(_1293_),
    .A(_1292_),
    .Y(_1294_));
 sg13g2_a21oi_1 _3943_ (.A1(net43),
    .A2(_1683_),
    .Y(_1295_),
    .B1(net54));
 sg13g2_nand2_1 _3944_ (.Y(_0178_),
    .A(_1294_),
    .B(_1295_));
 sg13g2_xnor2_1 _3945_ (.Y(_1296_),
    .A(_1682_),
    .B(net47));
 sg13g2_nand2_1 _3946_ (.Y(_1297_),
    .A(net47),
    .B(_1773_));
 sg13g2_nand2_1 _3947_ (.Y(_1298_),
    .A(_1292_),
    .B(_1297_));
 sg13g2_inv_1 _3948_ (.Y(_1299_),
    .A(_1298_));
 sg13g2_nor2_1 _3949_ (.A(_1296_),
    .B(_1299_),
    .Y(_1300_));
 sg13g2_inv_1 _3950_ (.Y(_1301_),
    .A(_1300_));
 sg13g2_a21oi_1 _3951_ (.A1(_1299_),
    .A2(_1296_),
    .Y(_1302_),
    .B1(_1256_));
 sg13g2_a22oi_1 _3952_ (.Y(_1303_),
    .B1(_1301_),
    .B2(_1302_),
    .A2(net43),
    .A1(_1682_));
 sg13g2_nand2_1 _3953_ (.Y(_0179_),
    .A(_1303_),
    .B(_0996_));
 sg13g2_inv_1 _3954_ (.Y(_1304_),
    .A(\vga.left_down_pressed ));
 sg13g2_nor2_1 _3955_ (.A(net64),
    .B(net47),
    .Y(_1305_));
 sg13g2_a21oi_1 _3956_ (.A1(net64),
    .A2(_1304_),
    .Y(_1306_),
    .B1(_1305_));
 sg13g2_a21oi_1 _3957_ (.A1(_1777_),
    .A2(net47),
    .Y(_1307_),
    .B1(_1300_));
 sg13g2_xnor2_1 _3958_ (.Y(_1308_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_a21oi_1 _3959_ (.A1(_1257_),
    .A2(_1687_),
    .Y(_1309_),
    .B1(net53));
 sg13g2_o21ai_1 _3960_ (.B1(_1309_),
    .Y(_0180_),
    .A1(_1257_),
    .A2(_1308_));
 sg13g2_inv_1 _3961_ (.Y(_1310_),
    .A(_1306_));
 sg13g2_a21oi_1 _3962_ (.A1(net64),
    .A2(_1777_),
    .Y(_1311_),
    .B1(_1760_));
 sg13g2_nand3_1 _3963_ (.B(_1248_),
    .C(_1311_),
    .A(_1260_),
    .Y(_1312_));
 sg13g2_a21oi_1 _3964_ (.A1(_1300_),
    .A2(_1310_),
    .Y(_1313_),
    .B1(_1312_));
 sg13g2_a21oi_1 _3965_ (.A1(_1300_),
    .A2(_1305_),
    .Y(_1314_),
    .B1(_1313_));
 sg13g2_o21ai_1 _3966_ (.B1(_0962_),
    .Y(_1315_),
    .A1(_1791_),
    .A2(_1314_));
 sg13g2_nand2_1 _3967_ (.Y(_1316_),
    .A(_1314_),
    .B(_1791_));
 sg13g2_nor2b_1 _3968_ (.A(_1315_),
    .B_N(_1316_),
    .Y(_0181_));
 sg13g2_inv_1 _3969_ (.Y(_1317_),
    .A(_0081_));
 sg13g2_inv_1 _3970_ (.Y(_1318_),
    .A(_1416_));
 sg13g2_nand4_1 _3971_ (.B(_0547_),
    .C(net68),
    .A(_1318_),
    .Y(_1319_),
    .D(_0081_));
 sg13g2_a21oi_1 _3972_ (.A1(_1318_),
    .A2(_0062_),
    .Y(_1320_),
    .B1(_1421_));
 sg13g2_a21oi_1 _3973_ (.A1(_1319_),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1507_));
 sg13g2_inv_1 _3974_ (.Y(_1322_),
    .A(\vga.right_up_pressed ));
 sg13g2_a21oi_1 _3975_ (.A1(_1321_),
    .A2(_1547_),
    .Y(_1323_),
    .B1(_1322_));
 sg13g2_nor2_1 _3976_ (.A(_1426_),
    .B(_1496_),
    .Y(_1324_));
 sg13g2_nand2_1 _3977_ (.Y(_1325_),
    .A(_1445_),
    .B(_1449_));
 sg13g2_nor4_1 _3978_ (.A(_1420_),
    .B(net68),
    .C(_1318_),
    .D(_1325_),
    .Y(_1326_));
 sg13g2_nor3_1 _3979_ (.A(_1424_),
    .B(_1479_),
    .C(_1496_),
    .Y(_1327_));
 sg13g2_o21ai_1 _3980_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_1423_),
    .A2(_1326_));
 sg13g2_nand2_1 _3981_ (.Y(_1329_),
    .A(_1328_),
    .B(\vga.right_down_pressed ));
 sg13g2_nor2_1 _3982_ (.A(_1324_),
    .B(_1329_),
    .Y(_1330_));
 sg13g2_buf_1 _3983_ (.A(_1330_),
    .X(_1331_));
 sg13g2_buf_1 _3984_ (.A(_1331_),
    .X(_1332_));
 sg13g2_nor2_1 _3985_ (.A(_1323_),
    .B(net45),
    .Y(_1333_));
 sg13g2_buf_1 _3986_ (.A(_1333_),
    .X(_1334_));
 sg13g2_a21oi_1 _3987_ (.A1(net39),
    .A2(_1449_),
    .Y(_1335_),
    .B1(net53));
 sg13g2_o21ai_1 _3988_ (.B1(_1335_),
    .Y(_0182_),
    .A1(_1317_),
    .A2(net39));
 sg13g2_inv_2 _3989_ (.Y(_1336_),
    .A(_1333_));
 sg13g2_xnor2_1 _3990_ (.Y(_1337_),
    .A(_0547_),
    .B(net45));
 sg13g2_xnor2_1 _3991_ (.Y(_1338_),
    .A(_1317_),
    .B(_1337_));
 sg13g2_a21oi_1 _3992_ (.A1(_1338_),
    .A2(_1336_),
    .Y(_1339_),
    .B1(net55));
 sg13g2_o21ai_1 _3993_ (.B1(_1339_),
    .Y(_0183_),
    .A1(_0547_),
    .A2(_1336_));
 sg13g2_xnor2_1 _3994_ (.Y(_1340_),
    .A(net68),
    .B(_1331_));
 sg13g2_o21ai_1 _3995_ (.B1(_1325_),
    .Y(_1341_),
    .A1(_0528_),
    .A2(_1331_));
 sg13g2_nor2_1 _3996_ (.A(_1340_),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_nand2_1 _3997_ (.Y(_1343_),
    .A(_1341_),
    .B(_1340_));
 sg13g2_nand2_1 _3998_ (.Y(_1344_),
    .A(_1343_),
    .B(_1336_));
 sg13g2_a21oi_1 _3999_ (.A1(net39),
    .A2(net68),
    .Y(_1345_),
    .B1(net55));
 sg13g2_o21ai_1 _4000_ (.B1(_1345_),
    .Y(_0184_),
    .A1(_1342_),
    .A2(_1344_));
 sg13g2_nor2_1 _4001_ (.A(_1318_),
    .B(net45),
    .Y(_1346_));
 sg13g2_inv_1 _4002_ (.Y(_1347_),
    .A(_1331_));
 sg13g2_nor2_1 _4003_ (.A(_1416_),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_nor2_1 _4004_ (.A(_1346_),
    .B(_1348_),
    .Y(_1349_));
 sg13g2_o21ai_1 _4005_ (.B1(_1343_),
    .Y(_1350_),
    .A1(_0062_),
    .A2(_1331_));
 sg13g2_xnor2_1 _4006_ (.Y(_1351_),
    .A(_1349_),
    .B(_1350_));
 sg13g2_a21oi_1 _4007_ (.A1(net39),
    .A2(_1416_),
    .Y(_1352_),
    .B1(net55));
 sg13g2_o21ai_1 _4008_ (.B1(_1352_),
    .Y(_0185_),
    .A1(net39),
    .A2(_1351_));
 sg13g2_nand2b_1 _4009_ (.Y(_1353_),
    .B(_1350_),
    .A_N(_1348_));
 sg13g2_nand2b_1 _4010_ (.Y(_1354_),
    .B(_1353_),
    .A_N(_1346_));
 sg13g2_xnor2_1 _4011_ (.Y(_1355_),
    .A(_1421_),
    .B(net45));
 sg13g2_nand2b_1 _4012_ (.Y(_1356_),
    .B(_1355_),
    .A_N(_1354_));
 sg13g2_nand2b_1 _4013_ (.Y(_1357_),
    .B(_1354_),
    .A_N(_1355_));
 sg13g2_nand3_1 _4014_ (.B(_1336_),
    .C(_1357_),
    .A(_1356_),
    .Y(_1358_));
 sg13g2_nand2_1 _4015_ (.Y(_1359_),
    .A(net39),
    .B(_1420_));
 sg13g2_a21oi_1 _4016_ (.A1(_1358_),
    .A2(_1359_),
    .Y(_0186_),
    .B1(net52));
 sg13g2_nand2b_1 _4017_ (.Y(_1360_),
    .B(_1347_),
    .A_N(_0061_));
 sg13g2_nand2_1 _4018_ (.Y(_1361_),
    .A(_1357_),
    .B(_1360_));
 sg13g2_xnor2_1 _4019_ (.Y(_1362_),
    .A(_1424_),
    .B(net45));
 sg13g2_nand2_1 _4020_ (.Y(_1363_),
    .A(_1361_),
    .B(_1362_));
 sg13g2_inv_1 _4021_ (.Y(_1364_),
    .A(_1363_));
 sg13g2_o21ai_1 _4022_ (.B1(_1336_),
    .Y(_1365_),
    .A1(_1362_),
    .A2(_1361_));
 sg13g2_a21oi_1 _4023_ (.A1(net39),
    .A2(_1424_),
    .Y(_1366_),
    .B1(net55));
 sg13g2_o21ai_1 _4024_ (.B1(_1366_),
    .Y(_0187_),
    .A1(_1364_),
    .A2(_1365_));
 sg13g2_nand2_1 _4025_ (.Y(_1367_),
    .A(_1347_),
    .B(_1511_));
 sg13g2_xnor2_1 _4026_ (.Y(_1368_),
    .A(_1479_),
    .B(net45));
 sg13g2_a21o_1 _4027_ (.A2(_1367_),
    .A1(_1363_),
    .B1(_1368_),
    .X(_1369_));
 sg13g2_nand3_1 _4028_ (.B(_1367_),
    .C(_1368_),
    .A(_1363_),
    .Y(_1370_));
 sg13g2_nand3_1 _4029_ (.B(_1336_),
    .C(_1370_),
    .A(_1369_),
    .Y(_1371_));
 sg13g2_a21oi_1 _4030_ (.A1(net39),
    .A2(_1425_),
    .Y(_1372_),
    .B1(_0952_));
 sg13g2_nand2_1 _4031_ (.Y(_0188_),
    .A(_1371_),
    .B(_1372_));
 sg13g2_xnor2_1 _4032_ (.Y(_1373_),
    .A(_1415_),
    .B(_1332_));
 sg13g2_o21ai_1 _4033_ (.B1(_1369_),
    .Y(_1374_),
    .A1(_0072_),
    .A2(net45));
 sg13g2_xor2_1 _4034_ (.B(_1374_),
    .A(_1373_),
    .X(_1375_));
 sg13g2_a21oi_1 _4035_ (.A1(_1333_),
    .A2(_1414_),
    .Y(_1376_),
    .B1(net55));
 sg13g2_o21ai_1 _4036_ (.B1(_1376_),
    .Y(_0189_),
    .A1(_1334_),
    .A2(_1375_));
 sg13g2_xor2_1 _4037_ (.B(_1332_),
    .A(_1432_),
    .X(_1377_));
 sg13g2_inv_1 _4038_ (.Y(_1378_),
    .A(_0070_));
 sg13g2_inv_1 _4039_ (.Y(_1379_),
    .A(_1362_));
 sg13g2_o21ai_1 _4040_ (.B1(_1367_),
    .Y(_1380_),
    .A1(_1360_),
    .A2(_1379_));
 sg13g2_nor2_1 _4041_ (.A(_1368_),
    .B(_1373_),
    .Y(_1381_));
 sg13g2_nor3_1 _4042_ (.A(_1414_),
    .B(_0072_),
    .C(net45),
    .Y(_1382_));
 sg13g2_a221oi_1 _4043_ (.B2(_1381_),
    .C1(_1382_),
    .B1(_1380_),
    .A1(_1378_),
    .Y(_1383_),
    .A2(_1347_));
 sg13g2_nor2_1 _4044_ (.A(_1355_),
    .B(_1379_),
    .Y(_1384_));
 sg13g2_nand3_1 _4045_ (.B(_1384_),
    .C(_1381_),
    .A(_1354_),
    .Y(_1385_));
 sg13g2_nand2_1 _4046_ (.Y(_1386_),
    .A(_1383_),
    .B(_1385_));
 sg13g2_xnor2_1 _4047_ (.Y(_1387_),
    .A(_1377_),
    .B(_1386_));
 sg13g2_nand2_1 _4048_ (.Y(_1388_),
    .A(_1387_),
    .B(_1336_));
 sg13g2_nand2_1 _4049_ (.Y(_1389_),
    .A(_1334_),
    .B(_1432_));
 sg13g2_a21oi_1 _4050_ (.A1(_1388_),
    .A2(_1389_),
    .Y(_0190_),
    .B1(net52));
 sg13g2_inv_1 _4051_ (.Y(_0196_),
    .A(_1638_));
 sg13g2_o21ai_1 _4052_ (.B1(\vga.score_l[3] ),
    .Y(_1390_),
    .A1(_1405_),
    .A2(\vga.score_l[2] ));
 sg13g2_a21oi_1 _4053_ (.A1(_1390_),
    .A2(_1404_),
    .Y(_0201_),
    .B1(net52));
 sg13g2_inv_1 _4054_ (.Y(_0206_),
    .A(net33));
 sg13g2_o21ai_1 _4055_ (.B1(_1819_),
    .Y(_1391_),
    .A1(_1815_),
    .A2(_1820_));
 sg13g2_a21oi_1 _4056_ (.A1(_1391_),
    .A2(_1821_),
    .Y(_0210_),
    .B1(net52));
 sg13g2_nand2_1 _4057_ (.Y(_1392_),
    .A(net60),
    .B(net5));
 sg13g2_inv_1 _4058_ (.Y(_0214_),
    .A(_1392_));
 sg13g2_nand2_1 _4059_ (.Y(_1393_),
    .A(net60),
    .B(_0316_));
 sg13g2_inv_1 _4060_ (.Y(_0215_),
    .A(_1393_));
 sg13g2_inv_1 _4061_ (.Y(_1394_),
    .A(\vga.vs_out ));
 sg13g2_nand2_1 _4062_ (.Y(_1395_),
    .A(_0433_),
    .B(_1978_));
 sg13g2_nor4_1 _4063_ (.A(_1395_),
    .B(_0912_),
    .C(_2013_),
    .D(_1185_),
    .Y(_1396_));
 sg13g2_o21ai_1 _4064_ (.B1(net79),
    .Y(_1397_),
    .A1(_1396_),
    .A2(_1197_));
 sg13g2_a21oi_1 _4065_ (.A1(_1394_),
    .A2(_1197_),
    .Y(_0216_),
    .B1(_1397_));
 sg13g2_inv_1 _4066_ (.Y(net14),
    .A(net6));
 sg13g2_inv_1 _4067_ (.Y(_1398_),
    .A(b0));
 sg13g2_nand2_1 _4068_ (.Y(_1399_),
    .A(net90),
    .B(g0));
 sg13g2_o21ai_1 _4069_ (.B1(_1399_),
    .Y(net23),
    .A1(net90),
    .A2(_1398_));
 sg13g2_inv_1 _4070_ (.Y(_1400_),
    .A(\vga.vs ));
 sg13g2_o21ai_1 _4071_ (.B1(_1399_),
    .Y(net24),
    .A1(net90),
    .A2(_1400_));
 sg13g2_inv_1 _4072_ (.Y(_1401_),
    .A(g0));
 sg13g2_nand2_1 _4073_ (.Y(_1402_),
    .A(net90),
    .B(b0));
 sg13g2_o21ai_1 _4074_ (.B1(_1402_),
    .Y(net26),
    .A1(net90),
    .A2(_1401_));
 sg13g2_inv_1 _4075_ (.Y(_1403_),
    .A(hs));
 sg13g2_o21ai_1 _4076_ (.B1(_1402_),
    .Y(net28),
    .A1(net90),
    .A2(_1403_));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net93),
    .D(_0006_),
    .Q_N(_2105_),
    .Q(_0026_));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net94),
    .D(_0007_),
    .Q_N(_2104_),
    .Q(_0027_));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net95),
    .D(_0085_),
    .Q_N(_2103_),
    .Q(_0030_));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net96),
    .D(_0086_),
    .Q_N(_2106_),
    .Q(_0022_));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net97),
    .D(_0002_),
    .Q_N(_2107_),
    .Q(_0021_));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net98),
    .D(_0003_),
    .Q_N(_2108_),
    .Q(_0023_));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net99),
    .D(_0010_),
    .Q_N(_2109_),
    .Q(_0032_));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net100),
    .D(_0011_),
    .Q_N(_2110_),
    .Q(_0033_));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net101),
    .D(_0000_),
    .Q_N(_2111_),
    .Q(_0018_));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net102),
    .D(_0001_),
    .Q_N(_2102_),
    .Q(_0020_));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net103),
    .D(_0087_),
    .Q_N(_2112_),
    .Q(_0017_));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net104),
    .D(_0009_),
    .Q_N(_2113_),
    .Q(_0031_));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net105),
    .D(_0012_),
    .Q_N(_2114_),
    .Q(_0034_));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net106),
    .D(_0013_),
    .Q_N(_2101_),
    .Q(_0035_));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net107),
    .D(_0088_),
    .Q_N(_2115_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net108),
    .D(_0008_),
    .Q_N(_2100_),
    .Q(_0029_));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net109),
    .D(_0089_),
    .Q_N(_2099_),
    .Q(_0028_));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net110),
    .D(_0090_),
    .Q_N(_2098_),
    .Q(_0019_));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net111),
    .D(_0091_),
    .Q_N(_2116_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net112),
    .D(_0004_),
    .Q_N(_2117_),
    .Q(_0024_));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net113),
    .D(_0005_),
    .Q_N(_2097_),
    .Q(_0025_));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net114),
    .D(_0092_),
    .Q_N(_2096_),
    .Q(_0016_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4077__93 (.L_HI(net93));
 sg13g2_buf_1 _4101_ (.A(net89),
    .X(net7));
 sg13g2_buf_1 _4102_ (.A(net89),
    .X(net8));
 sg13g2_buf_1 _4103_ (.A(net89),
    .X(net9));
 sg13g2_buf_1 _4104_ (.A(net89),
    .X(net10));
 sg13g2_buf_1 _4105_ (.A(net89),
    .X(net11));
 sg13g2_buf_1 _4106_ (.A(net89),
    .X(net12));
 sg13g2_buf_1 _4107_ (.A(net89),
    .X(net13));
 sg13g2_buf_1 _4108_ (.A(g0),
    .X(net15));
 sg13g2_buf_1 _4109_ (.A(g0),
    .X(net16));
 sg13g2_buf_1 _4110_ (.A(g0),
    .X(net17));
 sg13g2_buf_1 _4111_ (.A(g0),
    .X(net18));
 sg13g2_buf_1 _4112_ (.A(hs),
    .X(net19));
 sg13g2_buf_1 _4113_ (.A(\vga.vs ),
    .X(net20));
 sg13g2_buf_1 _4114_ (.A(net91),
    .X(uio_out[6]));
 sg13g2_buf_1 _4115_ (.A(net92),
    .X(uio_out[7]));
 sg13g2_buf_1 _4116_ (.A(g0),
    .X(net21));
 sg13g2_buf_1 _4117_ (.A(g0),
    .X(net22));
 sg13g2_buf_1 _4118_ (.A(net26),
    .X(net25));
 sg13g2_buf_1 _4119_ (.A(b0),
    .X(net27));
 sg13g2_dfrbp_1 \vga.ball_angle[0]$_SDFFE_PN1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net115),
    .D(_0093_),
    .Q_N(_0084_),
    .Q(\vga.ball_angle[0] ));
 sg13g2_dfrbp_1 \vga.ball_angle[1]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net116),
    .D(_0094_),
    .Q_N(_2095_),
    .Q(\vga.ball_angle[1] ));
 sg13g2_dfrbp_1 \vga.ball_angle[2]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net117),
    .D(_0095_),
    .Q_N(_0063_),
    .Q(\vga.ball_angle[2] ));
 sg13g2_dfrbp_1 \vga.ball_angle[3]$_SDFFE_PN1P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net118),
    .D(_0096_),
    .Q_N(_0049_),
    .Q(\vga.ball_angle[3] ));
 sg13g2_dfrbp_1 \vga.ball_motion_l$_SDFFE_PN1N_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net119),
    .D(_0097_),
    .Q_N(_0064_),
    .Q(\vga.ball_motion_l ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[0]$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net120),
    .D(_0098_),
    .Q_N(_0045_),
    .Q(\vga.ball_pos_h[0] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[1]$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net121),
    .D(_0099_),
    .Q_N(_0057_),
    .Q(\vga.ball_pos_h[1] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[2]$_SDFFE_PN1P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net122),
    .D(_0100_),
    .Q_N(_2094_),
    .Q(\vga.ball_pos_h[2] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[3]$_SDFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net123),
    .D(_0101_),
    .Q_N(_2093_),
    .Q(\vga.ball_pos_h[3] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[4]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net124),
    .D(_0102_),
    .Q_N(_2092_),
    .Q(\vga.ball_pos_h[4] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[5]$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net125),
    .D(_0103_),
    .Q_N(_0052_),
    .Q(\vga.ball_pos_h[5] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[6]$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net126),
    .D(_0104_),
    .Q_N(_2091_),
    .Q(\vga.ball_pos_h[6] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[7]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net127),
    .D(_0105_),
    .Q_N(_0046_),
    .Q(\vga.ball_pos_h[7] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[8]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net128),
    .D(_0106_),
    .Q_N(_0047_),
    .Q(\vga.ball_pos_h[8] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[9]$_SDFFE_PN1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net129),
    .D(_0107_),
    .Q_N(_0048_),
    .Q(\vga.ball_pos_h[9] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net130),
    .D(_0108_),
    .Q_N(_2090_),
    .Q(\vga.ball_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(_0109_),
    .Q_N(_2089_),
    .Q(\vga.ball_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net132),
    .D(_0110_),
    .Q_N(_2088_),
    .Q(\vga.ball_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net133),
    .D(_0111_),
    .Q_N(_0075_),
    .Q(\vga.ball_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net134),
    .D(_0112_),
    .Q_N(_2087_),
    .Q(\vga.ball_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net135),
    .D(_0113_),
    .Q_N(_0074_),
    .Q(\vga.ball_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net136),
    .D(_0114_),
    .Q_N(_0071_),
    .Q(\vga.ball_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net137),
    .D(_0115_),
    .Q_N(_0073_),
    .Q(\vga.ball_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net138),
    .D(_0116_),
    .Q_N(_0067_),
    .Q(\vga.ball_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[0]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net139),
    .D(_0117_),
    .Q_N(_2086_),
    .Q(\vga.ball_ratio[0] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[1]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net140),
    .D(_0118_),
    .Q_N(_2085_),
    .Q(\vga.ball_ratio[1] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[2]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net141),
    .D(_0119_),
    .Q_N(_2084_),
    .Q(\vga.ball_ratio[2] ));
 sg13g2_dfrbp_1 \vga.blank_h$_SDFFE_PN1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net142),
    .D(_0120_),
    .Q_N(_2083_),
    .Q(\vga.blank_h ));
 sg13g2_dfrbp_1 \vga.blank_v$_SDFFE_PN1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(_0121_),
    .Q_N(_2082_),
    .Q(\vga.blank_v ));
 sg13g2_dfrbp_1 \vga.blu$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net144),
    .D(_0122_),
    .Q_N(_2081_),
    .Q(b0));
 sg13g2_dfrbp_1 \vga.count_h[0]$_SDFF_PN1_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net145),
    .D(_0123_),
    .Q_N(_0036_),
    .Q(\vga.count_h[0] ));
 sg13g2_dfrbp_1 \vga.count_h[1]$_SDFF_PN1_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net146),
    .D(_0124_),
    .Q_N(_0051_),
    .Q(\vga.count_h[1] ));
 sg13g2_dfrbp_1 \vga.count_h[2]$_SDFF_PN1_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net147),
    .D(_0125_),
    .Q_N(_0053_),
    .Q(\vga.count_h[2] ));
 sg13g2_dfrbp_1 \vga.count_h[3]$_SDFF_PN1_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net148),
    .D(_0126_),
    .Q_N(_2080_),
    .Q(\vga.count_h[3] ));
 sg13g2_dfrbp_1 \vga.count_h[4]$_SDFF_PN1_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net149),
    .D(_0127_),
    .Q_N(_0056_),
    .Q(\vga.count_h[4] ));
 sg13g2_dfrbp_1 \vga.count_h[5]$_SDFF_PN1_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net150),
    .D(_0128_),
    .Q_N(_0058_),
    .Q(\vga.count_h[5] ));
 sg13g2_dfrbp_1 \vga.count_h[6]$_SDFF_PN1_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net151),
    .D(_0129_),
    .Q_N(_0055_),
    .Q(\vga.count_h[6] ));
 sg13g2_dfrbp_1 \vga.count_h[7]$_SDFF_PN1_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net152),
    .D(_0130_),
    .Q_N(_0050_),
    .Q(\vga.count_h[7] ));
 sg13g2_dfrbp_1 \vga.count_h[8]$_SDFF_PN1_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net153),
    .D(_0131_),
    .Q_N(_0054_),
    .Q(\vga.count_h[8] ));
 sg13g2_dfrbp_1 \vga.count_h[9]$_SDFF_PN1_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net154),
    .D(_0132_),
    .Q_N(_0066_),
    .Q(\vga.count_h[9] ));
 sg13g2_dfrbp_1 \vga.count_v[0]$_SDFFE_PN1N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net155),
    .D(_0133_),
    .Q_N(_0037_),
    .Q(\vga.count_v[0] ));
 sg13g2_dfrbp_1 \vga.count_v[1]$_SDFFE_PN1N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net156),
    .D(_0134_),
    .Q_N(_0080_),
    .Q(\vga.count_v[1] ));
 sg13g2_dfrbp_1 \vga.count_v[2]$_SDFFE_PN1N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net157),
    .D(_0135_),
    .Q_N(_0038_),
    .Q(\vga.count_v[2] ));
 sg13g2_dfrbp_1 \vga.count_v[3]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net158),
    .D(_0136_),
    .Q_N(_0039_),
    .Q(\vga.count_v[3] ));
 sg13g2_dfrbp_1 \vga.count_v[4]$_SDFFE_PN1N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net159),
    .D(_0137_),
    .Q_N(_0040_),
    .Q(\vga.count_v[4] ));
 sg13g2_dfrbp_1 \vga.count_v[5]$_SDFFE_PN1N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(_0138_),
    .Q_N(_0041_),
    .Q(\vga.count_v[5] ));
 sg13g2_dfrbp_1 \vga.count_v[6]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net161),
    .D(_0139_),
    .Q_N(_0042_),
    .Q(\vga.count_v[6] ));
 sg13g2_dfrbp_1 \vga.count_v[7]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net162),
    .D(_0140_),
    .Q_N(_0043_),
    .Q(\vga.count_v[7] ));
 sg13g2_dfrbp_1 \vga.count_v[8]$_SDFFE_PN1N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net163),
    .D(_0141_),
    .Q_N(_0044_),
    .Q(\vga.count_v[8] ));
 sg13g2_dfrbp_1 \vga.count_v[9]$_SDFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net164),
    .D(_0142_),
    .Q_N(_0065_),
    .Q(\vga.count_v[9] ));
 sg13g2_dfrbp_1 \vga.hs_out$_SDFF_PP0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net165),
    .D(_0143_),
    .Q_N(hs),
    .Q(\vga.hs_out ));
 sg13g2_dfrbp_1 \vga.interval_counter[0]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net166),
    .D(_0144_),
    .Q_N(_0083_),
    .Q(\vga.interval_counter[0] ));
 sg13g2_dfrbp_1 \vga.interval_counter[10]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net167),
    .D(_0145_),
    .Q_N(_2079_),
    .Q(\vga.interval_counter[10] ));
 sg13g2_dfrbp_1 \vga.interval_counter[11]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net168),
    .D(_0146_),
    .Q_N(_2078_),
    .Q(\vga.interval_counter[11] ));
 sg13g2_dfrbp_1 \vga.interval_counter[12]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net169),
    .D(_0147_),
    .Q_N(_2077_),
    .Q(\vga.interval_counter[12] ));
 sg13g2_dfrbp_1 \vga.interval_counter[13]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net170),
    .D(_0148_),
    .Q_N(_2076_),
    .Q(\vga.interval_counter[13] ));
 sg13g2_dfrbp_1 \vga.interval_counter[14]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net171),
    .D(_0149_),
    .Q_N(_2075_),
    .Q(\vga.interval_counter[14] ));
 sg13g2_dfrbp_1 \vga.interval_counter[15]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net172),
    .D(_0150_),
    .Q_N(_2074_),
    .Q(\vga.interval_counter[15] ));
 sg13g2_dfrbp_1 \vga.interval_counter[16]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net173),
    .D(_0151_),
    .Q_N(_2073_),
    .Q(\vga.interval_counter[16] ));
 sg13g2_dfrbp_1 \vga.interval_counter[17]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net174),
    .D(_0152_),
    .Q_N(_2072_),
    .Q(\vga.interval_counter[17] ));
 sg13g2_dfrbp_1 \vga.interval_counter[18]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net175),
    .D(_0153_),
    .Q_N(_2071_),
    .Q(\vga.interval_counter[18] ));
 sg13g2_dfrbp_1 \vga.interval_counter[19]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net176),
    .D(_0154_),
    .Q_N(_2070_),
    .Q(\vga.interval_counter[19] ));
 sg13g2_dfrbp_1 \vga.interval_counter[1]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net177),
    .D(_0155_),
    .Q_N(_2069_),
    .Q(\vga.interval_counter[1] ));
 sg13g2_dfrbp_1 \vga.interval_counter[20]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net178),
    .D(_0156_),
    .Q_N(_2068_),
    .Q(\vga.interval_counter[20] ));
 sg13g2_dfrbp_1 \vga.interval_counter[21]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net179),
    .D(_0157_),
    .Q_N(_2067_),
    .Q(\vga.interval_counter[21] ));
 sg13g2_dfrbp_1 \vga.interval_counter[22]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net180),
    .D(_0158_),
    .Q_N(_2066_),
    .Q(\vga.interval_counter[22] ));
 sg13g2_dfrbp_1 \vga.interval_counter[23]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net181),
    .D(_0159_),
    .Q_N(_2065_),
    .Q(\vga.interval_counter[23] ));
 sg13g2_dfrbp_1 \vga.interval_counter[24]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net182),
    .D(_0160_),
    .Q_N(_2064_),
    .Q(\vga.interval_counter[24] ));
 sg13g2_dfrbp_1 \vga.interval_counter[2]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net183),
    .D(_0161_),
    .Q_N(_2063_),
    .Q(\vga.interval_counter[2] ));
 sg13g2_dfrbp_1 \vga.interval_counter[3]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net184),
    .D(_0162_),
    .Q_N(_2062_),
    .Q(\vga.interval_counter[3] ));
 sg13g2_dfrbp_1 \vga.interval_counter[4]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net185),
    .D(_0163_),
    .Q_N(_2061_),
    .Q(\vga.interval_counter[4] ));
 sg13g2_dfrbp_1 \vga.interval_counter[5]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net186),
    .D(_0164_),
    .Q_N(_2060_),
    .Q(\vga.interval_counter[5] ));
 sg13g2_dfrbp_1 \vga.interval_counter[6]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net187),
    .D(_0165_),
    .Q_N(_2059_),
    .Q(\vga.interval_counter[6] ));
 sg13g2_dfrbp_1 \vga.interval_counter[7]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net188),
    .D(_0166_),
    .Q_N(_2058_),
    .Q(\vga.interval_counter[7] ));
 sg13g2_dfrbp_1 \vga.interval_counter[8]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net189),
    .D(_0167_),
    .Q_N(_2057_),
    .Q(\vga.interval_counter[8] ));
 sg13g2_dfrbp_1 \vga.interval_counter[9]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net190),
    .D(_0168_),
    .Q_N(_2056_),
    .Q(\vga.interval_counter[9] ));
 sg13g2_dfrbp_1 \vga.left_down_1d$_DFFE_PN_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net191),
    .D(_0169_),
    .Q_N(_2055_),
    .Q(\vga.left_down_1d ));
 sg13g2_dfrbp_1 \vga.left_down_pressed$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net192),
    .D(_0170_),
    .Q_N(_2054_),
    .Q(\vga.left_down_pressed ));
 sg13g2_dfrbp_1 \vga.left_up_1d$_DFFE_PN_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net193),
    .D(_0171_),
    .Q_N(_2053_),
    .Q(\vga.left_up_1d ));
 sg13g2_dfrbp_1 \vga.left_up_pressed$_SDFF_PP0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net194),
    .D(_0172_),
    .Q_N(_2052_),
    .Q(\vga.left_up_pressed ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net195),
    .D(_0173_),
    .Q_N(_0082_),
    .Q(\vga.paddle_l_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net196),
    .D(_0174_),
    .Q_N(_2051_),
    .Q(\vga.paddle_l_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net197),
    .D(_0175_),
    .Q_N(_0060_),
    .Q(\vga.paddle_l_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net198),
    .D(_0176_),
    .Q_N(_2050_),
    .Q(\vga.paddle_l_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net199),
    .D(_0177_),
    .Q_N(_0059_),
    .Q(\vga.paddle_l_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net200),
    .D(_0178_),
    .Q_N(_0077_),
    .Q(\vga.paddle_l_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net201),
    .D(_0179_),
    .Q_N(_0079_),
    .Q(\vga.paddle_l_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net202),
    .D(_0180_),
    .Q_N(_0078_),
    .Q(\vga.paddle_l_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net203),
    .D(_0181_),
    .Q_N(_0076_),
    .Q(\vga.paddle_l_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net204),
    .D(_0182_),
    .Q_N(_0081_),
    .Q(\vga.paddle_r_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net205),
    .D(_0183_),
    .Q_N(_2049_),
    .Q(\vga.paddle_r_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net206),
    .D(_0184_),
    .Q_N(_0062_),
    .Q(\vga.paddle_r_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net207),
    .D(_0185_),
    .Q_N(_2048_),
    .Q(\vga.paddle_r_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net208),
    .D(_0186_),
    .Q_N(_0061_),
    .Q(\vga.paddle_r_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net209),
    .D(_0187_),
    .Q_N(_0069_),
    .Q(\vga.paddle_r_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net210),
    .D(_0188_),
    .Q_N(_0072_),
    .Q(\vga.paddle_r_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net211),
    .D(_0189_),
    .Q_N(_0070_),
    .Q(\vga.paddle_r_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net212),
    .D(_0190_),
    .Q_N(_0068_),
    .Q(\vga.paddle_r_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.red$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net213),
    .D(_0191_),
    .Q_N(_2047_),
    .Q(g0));
 sg13g2_dfrbp_1 \vga.right_down_1d$_DFFE_PN_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net214),
    .D(_0192_),
    .Q_N(_2046_),
    .Q(\vga.right_down_1d ));
 sg13g2_dfrbp_1 \vga.right_down_pressed$_SDFF_PP0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net215),
    .D(_0193_),
    .Q_N(_2045_),
    .Q(\vga.right_down_pressed ));
 sg13g2_dfrbp_1 \vga.right_up_1d$_DFFE_PN_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net216),
    .D(_0194_),
    .Q_N(_2044_),
    .Q(\vga.right_up_1d ));
 sg13g2_dfrbp_1 \vga.right_up_pressed$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net217),
    .D(_0195_),
    .Q_N(_2043_),
    .Q(\vga.right_up_pressed ));
 sg13g2_dfrbp_1 \vga.score_l[0]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net218),
    .D(_0196_),
    .Q_N(_2042_),
    .Q(\vga.score_l[0] ));
 sg13g2_dfrbp_1 \vga.score_l[1]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net219),
    .D(_0197_),
    .Q_N(_2041_),
    .Q(\vga.score_l[1] ));
 sg13g2_dfrbp_1 \vga.score_l[2]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net220),
    .D(_0198_),
    .Q_N(_2040_),
    .Q(\vga.score_l[2] ));
 sg13g2_dfrbp_1 \vga.score_l[3]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net221),
    .D(_0199_),
    .Q_N(_2039_),
    .Q(\vga.score_l[3] ));
 sg13g2_dfrbp_1 \vga.score_l[4]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net222),
    .D(net38),
    .Q_N(_2038_),
    .Q(\vga.score_l[4] ));
 sg13g2_dfrbp_1 \vga.score_l_ten_enable$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net223),
    .D(_0201_),
    .Q_N(_2037_),
    .Q(\vga.score_l_ten_enable ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[0]$_DFFE_PP_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net224),
    .D(_0202_),
    .Q_N(_2036_),
    .Q(\vga.score_l_unit_pixels[0] ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[1]$_DFFE_PP_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net225),
    .D(_0203_),
    .Q_N(_2035_),
    .Q(\vga.score_l_unit_pixels[1] ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[2]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net226),
    .D(_0204_),
    .Q_N(_2034_),
    .Q(\vga.score_l_unit_pixels[2] ));
 sg13g2_dfrbp_1 \vga.score_r[0]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net227),
    .D(_0205_),
    .Q_N(_2033_),
    .Q(\vga.score_r[0] ));
 sg13g2_dfrbp_1 \vga.score_r[1]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net228),
    .D(_0206_),
    .Q_N(_2032_),
    .Q(\vga.score_r[1] ));
 sg13g2_dfrbp_1 \vga.score_r[2]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net229),
    .D(_0207_),
    .Q_N(_2031_),
    .Q(\vga.score_r[2] ));
 sg13g2_dfrbp_1 \vga.score_r[3]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net230),
    .D(net37),
    .Q_N(_2030_),
    .Q(\vga.score_r[3] ));
 sg13g2_dfrbp_1 \vga.score_r[4]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net231),
    .D(_0209_),
    .Q_N(_2029_),
    .Q(\vga.score_r[4] ));
 sg13g2_dfrbp_1 \vga.score_r_ten_enable$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net232),
    .D(_0210_),
    .Q_N(_2028_),
    .Q(\vga.score_r_ten_enable ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[0]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net233),
    .D(_0211_),
    .Q_N(_2027_),
    .Q(\vga.score_r_unit_pixels[0] ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[1]$_DFFE_PP_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net234),
    .D(_0212_),
    .Q_N(_2026_),
    .Q(\vga.score_r_unit_pixels[1] ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[2]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net235),
    .D(_0213_),
    .Q_N(_2025_),
    .Q(\vga.score_r_unit_pixels[2] ));
 sg13g2_dfrbp_1 \vga.speed_lsb_1d$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net236),
    .D(_0214_),
    .Q_N(_2024_),
    .Q(\vga.speed_lsb_1d ));
 sg13g2_dfrbp_1 \vga.speed_msb_1d$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net237),
    .D(_0215_),
    .Q_N(_2023_),
    .Q(\vga.speed_msb_1d ));
 sg13g2_dfrbp_1 \vga.vs_out$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net238),
    .D(_0216_),
    .Q_N(\vga.vs ),
    .Q(\vga.vs_out ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[6]));
 sg13g2_buf_1 output14 (.A(net89),
    .X(uio_oe[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[0]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[1]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[3]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[4]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[5]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[6]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout29 (.A(_1654_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1008_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0990_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0964_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1880_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1878_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0207_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0955_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0208_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0200_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1334_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1180_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0395_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0365_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1257_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1216_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1332_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1198_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1260_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1615_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1858_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1650_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1584_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0274_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0992_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0952_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0273_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1976_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1138_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0996_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0991_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0962_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1810_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1809_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1731_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1688_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1620_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1516_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1471_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1456_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1448_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1439_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0496_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0275_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1981_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1980_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1978_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1977_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1971_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1970_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1660_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1574_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1570_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1561_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1493_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1489_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1465_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1453_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1447_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1443_),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(net14),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net14),
    .X(net90));
 sg13g2_tielo _4114__91 (.L_LO(net91));
 sg13g2_tielo _4115__92 (.L_LO(net92));
 sg13g2_tiehi _4078__94 (.L_HI(net94));
 sg13g2_tiehi _4079__95 (.L_HI(net95));
 sg13g2_tiehi _4080__96 (.L_HI(net96));
 sg13g2_tiehi _4081__97 (.L_HI(net97));
 sg13g2_tiehi _4082__98 (.L_HI(net98));
 sg13g2_tiehi _4083__99 (.L_HI(net99));
 sg13g2_tiehi _4084__100 (.L_HI(net100));
 sg13g2_tiehi _4085__101 (.L_HI(net101));
 sg13g2_tiehi _4086__102 (.L_HI(net102));
 sg13g2_tiehi _4087__103 (.L_HI(net103));
 sg13g2_tiehi _4088__104 (.L_HI(net104));
 sg13g2_tiehi _4089__105 (.L_HI(net105));
 sg13g2_tiehi _4090__106 (.L_HI(net106));
 sg13g2_tiehi _4091__107 (.L_HI(net107));
 sg13g2_tiehi _4092__108 (.L_HI(net108));
 sg13g2_tiehi _4093__109 (.L_HI(net109));
 sg13g2_tiehi _4094__110 (.L_HI(net110));
 sg13g2_tiehi _4095__111 (.L_HI(net111));
 sg13g2_tiehi _4096__112 (.L_HI(net112));
 sg13g2_tiehi _4097__113 (.L_HI(net113));
 sg13g2_tiehi _4098__114 (.L_HI(net114));
 sg13g2_tiehi \vga.ball_angle[0]$_SDFFE_PN1P__115  (.L_HI(net115));
 sg13g2_tiehi \vga.ball_angle[1]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \vga.ball_angle[2]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \vga.ball_angle[3]$_SDFFE_PN1P__118  (.L_HI(net118));
 sg13g2_tiehi \vga.ball_motion_l$_SDFFE_PN1N__119  (.L_HI(net119));
 sg13g2_tiehi \vga.ball_pos_h[0]$_SDFFE_PN1P__120  (.L_HI(net120));
 sg13g2_tiehi \vga.ball_pos_h[1]$_SDFFE_PN1P__121  (.L_HI(net121));
 sg13g2_tiehi \vga.ball_pos_h[2]$_SDFFE_PN1P__122  (.L_HI(net122));
 sg13g2_tiehi \vga.ball_pos_h[3]$_SDFFE_PN1P__123  (.L_HI(net123));
 sg13g2_tiehi \vga.ball_pos_h[4]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \vga.ball_pos_h[5]$_SDFFE_PN1P__125  (.L_HI(net125));
 sg13g2_tiehi \vga.ball_pos_h[6]$_SDFFE_PN1P__126  (.L_HI(net126));
 sg13g2_tiehi \vga.ball_pos_h[7]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \vga.ball_pos_h[8]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \vga.ball_pos_h[9]$_SDFFE_PN1P__129  (.L_HI(net129));
 sg13g2_tiehi \vga.ball_pos_v[0]$_SDFFE_PN1P__130  (.L_HI(net130));
 sg13g2_tiehi \vga.ball_pos_v[1]$_SDFFE_PN1P__131  (.L_HI(net131));
 sg13g2_tiehi \vga.ball_pos_v[2]$_SDFFE_PN1P__132  (.L_HI(net132));
 sg13g2_tiehi \vga.ball_pos_v[3]$_SDFFE_PN1P__133  (.L_HI(net133));
 sg13g2_tiehi \vga.ball_pos_v[4]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \vga.ball_pos_v[5]$_SDFFE_PN1P__135  (.L_HI(net135));
 sg13g2_tiehi \vga.ball_pos_v[6]$_SDFFE_PN1P__136  (.L_HI(net136));
 sg13g2_tiehi \vga.ball_pos_v[7]$_SDFFE_PN1P__137  (.L_HI(net137));
 sg13g2_tiehi \vga.ball_pos_v[8]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \vga.ball_ratio[0]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \vga.ball_ratio[1]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \vga.ball_ratio[2]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \vga.blank_h$_SDFFE_PN1P__142  (.L_HI(net142));
 sg13g2_tiehi \vga.blank_v$_SDFFE_PN1P__143  (.L_HI(net143));
 sg13g2_tiehi \vga.blu$_SDFF_PN0__144  (.L_HI(net144));
 sg13g2_tiehi \vga.count_h[0]$_SDFF_PN1__145  (.L_HI(net145));
 sg13g2_tiehi \vga.count_h[1]$_SDFF_PN1__146  (.L_HI(net146));
 sg13g2_tiehi \vga.count_h[2]$_SDFF_PN1__147  (.L_HI(net147));
 sg13g2_tiehi \vga.count_h[3]$_SDFF_PN1__148  (.L_HI(net148));
 sg13g2_tiehi \vga.count_h[4]$_SDFF_PN1__149  (.L_HI(net149));
 sg13g2_tiehi \vga.count_h[5]$_SDFF_PN1__150  (.L_HI(net150));
 sg13g2_tiehi \vga.count_h[6]$_SDFF_PN1__151  (.L_HI(net151));
 sg13g2_tiehi \vga.count_h[7]$_SDFF_PN1__152  (.L_HI(net152));
 sg13g2_tiehi \vga.count_h[8]$_SDFF_PN1__153  (.L_HI(net153));
 sg13g2_tiehi \vga.count_h[9]$_SDFF_PN1__154  (.L_HI(net154));
 sg13g2_tiehi \vga.count_v[0]$_SDFFE_PN1N__155  (.L_HI(net155));
 sg13g2_tiehi \vga.count_v[1]$_SDFFE_PN1N__156  (.L_HI(net156));
 sg13g2_tiehi \vga.count_v[2]$_SDFFE_PN1N__157  (.L_HI(net157));
 sg13g2_tiehi \vga.count_v[3]$_SDFFE_PN1N__158  (.L_HI(net158));
 sg13g2_tiehi \vga.count_v[4]$_SDFFE_PN1N__159  (.L_HI(net159));
 sg13g2_tiehi \vga.count_v[5]$_SDFFE_PN1N__160  (.L_HI(net160));
 sg13g2_tiehi \vga.count_v[6]$_SDFFE_PN1N__161  (.L_HI(net161));
 sg13g2_tiehi \vga.count_v[7]$_SDFFE_PN1N__162  (.L_HI(net162));
 sg13g2_tiehi \vga.count_v[8]$_SDFFE_PN1N__163  (.L_HI(net163));
 sg13g2_tiehi \vga.count_v[9]$_SDFFE_PN0N__164  (.L_HI(net164));
 sg13g2_tiehi \vga.hs_out$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \vga.interval_counter[0]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \vga.interval_counter[10]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \vga.interval_counter[11]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \vga.interval_counter[12]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \vga.interval_counter[13]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \vga.interval_counter[14]$_SDFF_PP0__171  (.L_HI(net171));
 sg13g2_tiehi \vga.interval_counter[15]$_SDFF_PP0__172  (.L_HI(net172));
 sg13g2_tiehi \vga.interval_counter[16]$_SDFF_PP0__173  (.L_HI(net173));
 sg13g2_tiehi \vga.interval_counter[17]$_SDFF_PP0__174  (.L_HI(net174));
 sg13g2_tiehi \vga.interval_counter[18]$_SDFF_PP0__175  (.L_HI(net175));
 sg13g2_tiehi \vga.interval_counter[19]$_SDFF_PP0__176  (.L_HI(net176));
 sg13g2_tiehi \vga.interval_counter[1]$_SDFF_PP0__177  (.L_HI(net177));
 sg13g2_tiehi \vga.interval_counter[20]$_SDFF_PP0__178  (.L_HI(net178));
 sg13g2_tiehi \vga.interval_counter[21]$_SDFF_PP0__179  (.L_HI(net179));
 sg13g2_tiehi \vga.interval_counter[22]$_SDFF_PP0__180  (.L_HI(net180));
 sg13g2_tiehi \vga.interval_counter[23]$_SDFF_PP0__181  (.L_HI(net181));
 sg13g2_tiehi \vga.interval_counter[24]$_SDFF_PP0__182  (.L_HI(net182));
 sg13g2_tiehi \vga.interval_counter[2]$_SDFF_PP0__183  (.L_HI(net183));
 sg13g2_tiehi \vga.interval_counter[3]$_SDFF_PP0__184  (.L_HI(net184));
 sg13g2_tiehi \vga.interval_counter[4]$_SDFF_PP0__185  (.L_HI(net185));
 sg13g2_tiehi \vga.interval_counter[5]$_SDFF_PP0__186  (.L_HI(net186));
 sg13g2_tiehi \vga.interval_counter[6]$_SDFF_PP0__187  (.L_HI(net187));
 sg13g2_tiehi \vga.interval_counter[7]$_SDFF_PP0__188  (.L_HI(net188));
 sg13g2_tiehi \vga.interval_counter[8]$_SDFF_PP0__189  (.L_HI(net189));
 sg13g2_tiehi \vga.interval_counter[9]$_SDFF_PP0__190  (.L_HI(net190));
 sg13g2_tiehi \vga.left_down_1d$_DFFE_PN__191  (.L_HI(net191));
 sg13g2_tiehi \vga.left_down_pressed$_SDFF_PP0__192  (.L_HI(net192));
 sg13g2_tiehi \vga.left_up_1d$_DFFE_PN__193  (.L_HI(net193));
 sg13g2_tiehi \vga.left_up_pressed$_SDFF_PP0__194  (.L_HI(net194));
 sg13g2_tiehi \vga.paddle_l_pos_v[0]$_SDFFE_PN1P__195  (.L_HI(net195));
 sg13g2_tiehi \vga.paddle_l_pos_v[1]$_SDFFE_PN1P__196  (.L_HI(net196));
 sg13g2_tiehi \vga.paddle_l_pos_v[2]$_SDFFE_PN1P__197  (.L_HI(net197));
 sg13g2_tiehi \vga.paddle_l_pos_v[3]$_SDFFE_PN1P__198  (.L_HI(net198));
 sg13g2_tiehi \vga.paddle_l_pos_v[4]$_SDFFE_PN0P__199  (.L_HI(net199));
 sg13g2_tiehi \vga.paddle_l_pos_v[5]$_SDFFE_PN1P__200  (.L_HI(net200));
 sg13g2_tiehi \vga.paddle_l_pos_v[6]$_SDFFE_PN1P__201  (.L_HI(net201));
 sg13g2_tiehi \vga.paddle_l_pos_v[7]$_SDFFE_PN1P__202  (.L_HI(net202));
 sg13g2_tiehi \vga.paddle_l_pos_v[8]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \vga.paddle_r_pos_v[0]$_SDFFE_PN1P__204  (.L_HI(net204));
 sg13g2_tiehi \vga.paddle_r_pos_v[1]$_SDFFE_PN1P__205  (.L_HI(net205));
 sg13g2_tiehi \vga.paddle_r_pos_v[2]$_SDFFE_PN1P__206  (.L_HI(net206));
 sg13g2_tiehi \vga.paddle_r_pos_v[3]$_SDFFE_PN1P__207  (.L_HI(net207));
 sg13g2_tiehi \vga.paddle_r_pos_v[4]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \vga.paddle_r_pos_v[5]$_SDFFE_PN1P__209  (.L_HI(net209));
 sg13g2_tiehi \vga.paddle_r_pos_v[6]$_SDFFE_PN1P__210  (.L_HI(net210));
 sg13g2_tiehi \vga.paddle_r_pos_v[7]$_SDFFE_PN1P__211  (.L_HI(net211));
 sg13g2_tiehi \vga.paddle_r_pos_v[8]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \vga.red$_SDFF_PP0__213  (.L_HI(net213));
 sg13g2_tiehi \vga.right_down_1d$_DFFE_PN__214  (.L_HI(net214));
 sg13g2_tiehi \vga.right_down_pressed$_SDFF_PP0__215  (.L_HI(net215));
 sg13g2_tiehi \vga.right_up_1d$_DFFE_PN__216  (.L_HI(net216));
 sg13g2_tiehi \vga.right_up_pressed$_SDFF_PP0__217  (.L_HI(net217));
 sg13g2_tiehi \vga.score_l[0]$_SDFF_PN0__218  (.L_HI(net218));
 sg13g2_tiehi \vga.score_l[1]$_SDFF_PN0__219  (.L_HI(net219));
 sg13g2_tiehi \vga.score_l[2]$_SDFF_PN0__220  (.L_HI(net220));
 sg13g2_tiehi \vga.score_l[3]$_SDFF_PN0__221  (.L_HI(net221));
 sg13g2_tiehi \vga.score_l[4]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \vga.score_l_ten_enable$_SDFF_PN0__223  (.L_HI(net223));
 sg13g2_tiehi \vga.score_l_unit_pixels[0]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \vga.score_l_unit_pixels[1]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \vga.score_l_unit_pixels[2]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \vga.score_r[0]$_SDFF_PN0__227  (.L_HI(net227));
 sg13g2_tiehi \vga.score_r[1]$_SDFF_PN0__228  (.L_HI(net228));
 sg13g2_tiehi \vga.score_r[2]$_SDFF_PN0__229  (.L_HI(net229));
 sg13g2_tiehi \vga.score_r[3]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \vga.score_r[4]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \vga.score_r_ten_enable$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \vga.score_r_unit_pixels[0]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \vga.score_r_unit_pixels[1]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \vga.score_r_unit_pixels[2]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \vga.speed_lsb_1d$_SDFF_PN0__236  (.L_HI(net236));
 sg13g2_tiehi \vga.speed_msb_1d$_SDFF_PN0__237  (.L_HI(net237));
 sg13g2_tiehi \vga.vs_out$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_4 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_61 ();
 sg13g2_decap_8 FILLER_0_66 ();
 sg13g2_fill_2 FILLER_0_73 ();
 sg13g2_decap_8 FILLER_0_88 ();
 sg13g2_decap_8 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_8 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_87 ();
 sg13g2_decap_4 FILLER_1_114 ();
 sg13g2_fill_1 FILLER_1_118 ();
 sg13g2_decap_4 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_136 ();
 sg13g2_decap_4 FILLER_1_141 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_fill_2 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_163 ();
 sg13g2_decap_8 FILLER_1_170 ();
 sg13g2_decap_8 FILLER_1_177 ();
 sg13g2_decap_8 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_198 ();
 sg13g2_fill_2 FILLER_1_205 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_4 FILLER_1_230 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_4 FILLER_1_331 ();
 sg13g2_fill_2 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_8 FILLER_1_403 ();
 sg13g2_decap_8 FILLER_1_410 ();
 sg13g2_decap_8 FILLER_1_417 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_30 ();
 sg13g2_fill_1 FILLER_2_43 ();
 sg13g2_fill_2 FILLER_2_83 ();
 sg13g2_decap_4 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_fill_1 FILLER_2_106 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_fill_2 FILLER_2_144 ();
 sg13g2_fill_1 FILLER_2_151 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_decap_4 FILLER_2_177 ();
 sg13g2_fill_2 FILLER_2_181 ();
 sg13g2_fill_2 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_fill_1 FILLER_2_292 ();
 sg13g2_fill_2 FILLER_2_298 ();
 sg13g2_decap_4 FILLER_2_353 ();
 sg13g2_fill_2 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_18 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_fill_2 FILLER_3_44 ();
 sg13g2_fill_2 FILLER_3_64 ();
 sg13g2_fill_1 FILLER_3_69 ();
 sg13g2_fill_2 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_fill_2 FILLER_3_228 ();
 sg13g2_fill_1 FILLER_3_230 ();
 sg13g2_fill_2 FILLER_3_237 ();
 sg13g2_fill_2 FILLER_3_265 ();
 sg13g2_fill_1 FILLER_3_267 ();
 sg13g2_fill_1 FILLER_3_288 ();
 sg13g2_fill_1 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_2 FILLER_4_34 ();
 sg13g2_fill_1 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_fill_2 FILLER_4_93 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_fill_1 FILLER_4_165 ();
 sg13g2_fill_2 FILLER_4_196 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_2 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_fill_2 FILLER_4_278 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_1 FILLER_4_342 ();
 sg13g2_fill_2 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_fill_2 FILLER_5_60 ();
 sg13g2_fill_2 FILLER_5_66 ();
 sg13g2_fill_1 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_1 FILLER_5_94 ();
 sg13g2_fill_2 FILLER_5_103 ();
 sg13g2_fill_2 FILLER_5_110 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_decap_4 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_283 ();
 sg13g2_fill_2 FILLER_5_295 ();
 sg13g2_fill_1 FILLER_5_307 ();
 sg13g2_fill_1 FILLER_5_313 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_347 ();
 sg13g2_fill_1 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_1 FILLER_6_75 ();
 sg13g2_fill_2 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_111 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_fill_2 FILLER_6_129 ();
 sg13g2_fill_1 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_274 ();
 sg13g2_fill_1 FILLER_6_317 ();
 sg13g2_fill_2 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_fill_2 FILLER_7_81 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_decap_4 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_278 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_359 ();
 sg13g2_fill_2 FILLER_7_398 ();
 sg13g2_fill_1 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_404 ();
 sg13g2_decap_8 FILLER_7_411 ();
 sg13g2_decap_8 FILLER_7_418 ();
 sg13g2_decap_4 FILLER_7_425 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_fill_2 FILLER_8_57 ();
 sg13g2_fill_1 FILLER_8_113 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_202 ();
 sg13g2_fill_1 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_decap_4 FILLER_9_13 ();
 sg13g2_fill_2 FILLER_9_17 ();
 sg13g2_fill_2 FILLER_9_22 ();
 sg13g2_fill_2 FILLER_9_66 ();
 sg13g2_fill_2 FILLER_9_72 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_2 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_380 ();
 sg13g2_fill_2 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_44 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_2 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_fill_1 FILLER_10_237 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_267 ();
 sg13g2_fill_1 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_fill_2 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_26 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_207 ();
 sg13g2_fill_2 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_265 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_fill_2 FILLER_11_305 ();
 sg13g2_fill_2 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_66 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_248 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_fill_2 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_401 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_4 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_25 ();
 sg13g2_fill_2 FILLER_13_31 ();
 sg13g2_fill_1 FILLER_13_33 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_fill_1 FILLER_13_202 ();
 sg13g2_decap_4 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_344 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_267 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_32 ();
 sg13g2_fill_2 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_216 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_4 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_decap_4 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_395 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_decap_4 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_38 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_81 ();
 sg13g2_fill_2 FILLER_21_93 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_151 ();
 sg13g2_decap_4 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_2 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_414 ();
 sg13g2_fill_2 FILLER_26_423 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_46 ();
 sg13g2_fill_2 FILLER_27_52 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_28_16 ();
 sg13g2_fill_1 FILLER_28_22 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_398 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_30_5 ();
 sg13g2_fill_1 FILLER_30_43 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_6 ();
 sg13g2_fill_2 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_fill_1 FILLER_32_24 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_227 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_2 FILLER_33_34 ();
 sg13g2_fill_1 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_139 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_35_66 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_fill_2 FILLER_37_415 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_403 ();
endmodule
