module tt_um_joerdsonsilva_modem (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire clknet_0_clk;
 wire net173;
 wire demod_out;
 wire \modem._0_[0] ;
 wire \modem._0_[1] ;
 wire \modem._0_[2] ;
 wire \modem._0_[3] ;
 wire \modem._0_[4] ;
 wire \modem._0_[5] ;
 wire \modem._4_ ;
 wire \modem._5_ ;
 wire \modem._6_ ;
 wire \modem.instance1._0_ ;
 wire \modem.instance1._1_ ;
 wire \modem.instance1._2_[0] ;
 wire \modem.instance1._2_[1] ;
 wire \modem.instance1._2_[2] ;
 wire \modem.instance1._2_[3] ;
 wire \modem.instance1._2_[4] ;
 wire \modem.instance1._2_[5] ;
 wire \modem.instance1.instance1._1_ ;
 wire \modem.instance1.instance1._3_[0] ;
 wire \modem.instance1.instance1._3_[1] ;
 wire \modem.instance1.instance1._3_[2] ;
 wire \modem.instance1.instance1._3_[3] ;
 wire \modem.instance1.instance1._3_[4] ;
 wire \modem.instance1.instance1._3_[5] ;
 wire \modem.instance1.instance1._3_[6] ;
 wire \modem.instance1.instance1._6_[0] ;
 wire \modem.instance1.instance1._6_[1] ;
 wire \modem.instance1.instance1._6_[2] ;
 wire \modem.instance1.instance1._6_[3] ;
 wire \modem.instance1.instance1._6_[4] ;
 wire \modem.instance1.instance1._6_[5] ;
 wire \modem.instance1.instance1._6_[6] ;
 wire \modem.instance1.instance2._00_ ;
 wire \modem.instance1.instance2._03_ ;
 wire \modem.instance1.instance2._04_ ;
 wire \modem.instance1.instance2._05_ ;
 wire \modem.instance1.instance2._09_[0] ;
 wire \modem.instance1.instance2._09_[10] ;
 wire \modem.instance1.instance2._09_[11] ;
 wire \modem.instance1.instance2._09_[12] ;
 wire \modem.instance1.instance2._09_[13] ;
 wire \modem.instance1.instance2._09_[14] ;
 wire \modem.instance1.instance2._09_[15] ;
 wire \modem.instance1.instance2._09_[16] ;
 wire \modem.instance1.instance2._09_[17] ;
 wire \modem.instance1.instance2._09_[18] ;
 wire \modem.instance1.instance2._09_[19] ;
 wire \modem.instance1.instance2._09_[1] ;
 wire \modem.instance1.instance2._09_[20] ;
 wire \modem.instance1.instance2._09_[21] ;
 wire \modem.instance1.instance2._09_[22] ;
 wire \modem.instance1.instance2._09_[23] ;
 wire \modem.instance1.instance2._09_[24] ;
 wire \modem.instance1.instance2._09_[25] ;
 wire \modem.instance1.instance2._09_[26] ;
 wire \modem.instance1.instance2._09_[27] ;
 wire \modem.instance1.instance2._09_[28] ;
 wire \modem.instance1.instance2._09_[29] ;
 wire \modem.instance1.instance2._09_[2] ;
 wire \modem.instance1.instance2._09_[30] ;
 wire \modem.instance1.instance2._09_[31] ;
 wire \modem.instance1.instance2._09_[3] ;
 wire \modem.instance1.instance2._09_[4] ;
 wire \modem.instance1.instance2._09_[5] ;
 wire \modem.instance1.instance2._09_[6] ;
 wire \modem.instance1.instance2._09_[7] ;
 wire \modem.instance1.instance2._09_[8] ;
 wire \modem.instance1.instance2._09_[9] ;
 wire \modem.instance1.instance2._10_[0] ;
 wire \modem.instance1.instance2._10_[10] ;
 wire \modem.instance1.instance2._10_[11] ;
 wire \modem.instance1.instance2._10_[12] ;
 wire \modem.instance1.instance2._10_[13] ;
 wire \modem.instance1.instance2._10_[14] ;
 wire \modem.instance1.instance2._10_[15] ;
 wire \modem.instance1.instance2._10_[16] ;
 wire \modem.instance1.instance2._10_[17] ;
 wire \modem.instance1.instance2._10_[18] ;
 wire \modem.instance1.instance2._10_[19] ;
 wire \modem.instance1.instance2._10_[1] ;
 wire \modem.instance1.instance2._10_[20] ;
 wire \modem.instance1.instance2._10_[21] ;
 wire \modem.instance1.instance2._10_[22] ;
 wire \modem.instance1.instance2._10_[23] ;
 wire \modem.instance1.instance2._10_[24] ;
 wire \modem.instance1.instance2._10_[25] ;
 wire \modem.instance1.instance2._10_[26] ;
 wire \modem.instance1.instance2._10_[27] ;
 wire \modem.instance1.instance2._10_[28] ;
 wire \modem.instance1.instance2._10_[29] ;
 wire \modem.instance1.instance2._10_[2] ;
 wire \modem.instance1.instance2._10_[30] ;
 wire \modem.instance1.instance2._10_[31] ;
 wire \modem.instance1.instance2._10_[3] ;
 wire \modem.instance1.instance2._10_[4] ;
 wire \modem.instance1.instance2._10_[5] ;
 wire \modem.instance1.instance2._10_[6] ;
 wire \modem.instance1.instance2._10_[7] ;
 wire \modem.instance1.instance2._10_[8] ;
 wire \modem.instance1.instance2._10_[9] ;
 wire \modem.instance1.instance2.ffd0._0_ ;
 wire \modem.instance1.instance2.ffd2._0_ ;
 wire \modem.instance1.instance2.ffd3._0_ ;
 wire \modem.instance1.instance2.ffd4._0_ ;
 wire \modem.instance1.instance3._0_[1] ;
 wire \modem.instance1.instance3._3_[0] ;
 wire \modem.instance1.instance3._3_[1] ;
 wire \modem.instance1.instance3._3_[2] ;
 wire \modem.instance1.instance3._3_[3] ;
 wire \modem.instance1.instance3._3_[4] ;
 wire \modem.instance1.instance3._4_[0] ;
 wire \modem.instance1.instance3._4_[2] ;
 wire \modem.instance1.instance3._4_[3] ;
 wire \modem.instance1.instance3._4_[4] ;
 wire \modem.instance1.instance4._0_[0] ;
 wire \modem.instance1.instance4._0_[1] ;
 wire \modem.instance1.instance4._0_[2] ;
 wire \modem.instance1.instance4._0_[3] ;
 wire \modem.instance1.instance4._0_[4] ;
 wire \modem.instance1.instance4._0_[5] ;
 wire \modem.instance2._0_ ;
 wire \modem.instance2._1_ ;
 wire \modem.instance2._2_[0] ;
 wire \modem.instance2._2_[1] ;
 wire \modem.instance2._2_[2] ;
 wire \modem.instance2._2_[3] ;
 wire \modem.instance2._2_[4] ;
 wire \modem.instance2._2_[5] ;
 wire \modem.instance2._3_[0] ;
 wire \modem.instance2._3_[1] ;
 wire \modem.instance2._3_[2] ;
 wire \modem.instance2._3_[3] ;
 wire \modem.instance2._3_[4] ;
 wire \modem.instance2._3_[5] ;
 wire \modem.instance2._4_ ;
 wire \modem.instance2.instance1._1_ ;
 wire \modem.instance2.instance1._3_[0] ;
 wire \modem.instance2.instance1._3_[1] ;
 wire \modem.instance2.instance1._3_[2] ;
 wire \modem.instance2.instance1._3_[3] ;
 wire \modem.instance2.instance1._3_[4] ;
 wire \modem.instance2.instance1._3_[5] ;
 wire \modem.instance2.instance1._3_[6] ;
 wire \modem.instance2.instance1._6_[0] ;
 wire \modem.instance2.instance1._6_[1] ;
 wire \modem.instance2.instance1._6_[2] ;
 wire \modem.instance2.instance1._6_[3] ;
 wire \modem.instance2.instance1._6_[4] ;
 wire \modem.instance2.instance1._6_[5] ;
 wire \modem.instance2.instance1._6_[6] ;
 wire \modem.instance2.instance2._1_ ;
 wire \modem.instance2.instance2._3_[0] ;
 wire \modem.instance2.instance2._3_[1] ;
 wire \modem.instance2.instance2._3_[2] ;
 wire \modem.instance2.instance2._3_[3] ;
 wire \modem.instance2.instance2._3_[4] ;
 wire \modem.instance2.instance2._3_[5] ;
 wire \modem.instance2.instance2._3_[6] ;
 wire \modem.instance2.instance2._6_[0] ;
 wire \modem.instance2.instance2._6_[1] ;
 wire \modem.instance2.instance2._6_[2] ;
 wire \modem.instance2.instance2._6_[3] ;
 wire \modem.instance2.instance2._6_[4] ;
 wire \modem.instance2.instance2._6_[5] ;
 wire \modem.instance2.instance2._6_[6] ;
 wire \modem.instance2.instance3._0_[1] ;
 wire \modem.instance2.instance3._3_[0] ;
 wire \modem.instance2.instance3._3_[1] ;
 wire \modem.instance2.instance3._3_[2] ;
 wire \modem.instance2.instance3._3_[3] ;
 wire \modem.instance2.instance3._3_[4] ;
 wire \modem.instance2.instance3._4_[0] ;
 wire \modem.instance2.instance3._4_[2] ;
 wire \modem.instance2.instance3._4_[3] ;
 wire \modem.instance2.instance3._4_[4] ;
 wire \modem.instance2.instance4._0_[1] ;
 wire \modem.instance2.instance4._3_[0] ;
 wire \modem.instance2.instance4._3_[1] ;
 wire \modem.instance2.instance4._3_[2] ;
 wire \modem.instance2.instance4._3_[3] ;
 wire \modem.instance2.instance4._3_[4] ;
 wire \modem.instance2.instance4._4_[0] ;
 wire \modem.instance2.instance4._4_[2] ;
 wire \modem.instance2.instance4._4_[3] ;
 wire \modem.instance2.instance4._4_[4] ;
 wire \modem.instance2.instance5._00_ ;
 wire \modem.instance2.instance5._03_ ;
 wire \modem.instance2.instance5._04_ ;
 wire \modem.instance2.instance5._05_ ;
 wire \modem.instance2.instance5._09_[0] ;
 wire \modem.instance2.instance5._09_[10] ;
 wire \modem.instance2.instance5._09_[11] ;
 wire \modem.instance2.instance5._09_[12] ;
 wire \modem.instance2.instance5._09_[13] ;
 wire \modem.instance2.instance5._09_[14] ;
 wire \modem.instance2.instance5._09_[15] ;
 wire \modem.instance2.instance5._09_[16] ;
 wire \modem.instance2.instance5._09_[17] ;
 wire \modem.instance2.instance5._09_[18] ;
 wire \modem.instance2.instance5._09_[19] ;
 wire \modem.instance2.instance5._09_[1] ;
 wire \modem.instance2.instance5._09_[20] ;
 wire \modem.instance2.instance5._09_[21] ;
 wire \modem.instance2.instance5._09_[22] ;
 wire \modem.instance2.instance5._09_[23] ;
 wire \modem.instance2.instance5._09_[24] ;
 wire \modem.instance2.instance5._09_[25] ;
 wire \modem.instance2.instance5._09_[26] ;
 wire \modem.instance2.instance5._09_[27] ;
 wire \modem.instance2.instance5._09_[28] ;
 wire \modem.instance2.instance5._09_[29] ;
 wire \modem.instance2.instance5._09_[2] ;
 wire \modem.instance2.instance5._09_[30] ;
 wire \modem.instance2.instance5._09_[31] ;
 wire \modem.instance2.instance5._09_[3] ;
 wire \modem.instance2.instance5._09_[4] ;
 wire \modem.instance2.instance5._09_[5] ;
 wire \modem.instance2.instance5._09_[6] ;
 wire \modem.instance2.instance5._09_[7] ;
 wire \modem.instance2.instance5._09_[8] ;
 wire \modem.instance2.instance5._09_[9] ;
 wire \modem.instance2.instance5._10_[0] ;
 wire \modem.instance2.instance5._10_[10] ;
 wire \modem.instance2.instance5._10_[11] ;
 wire \modem.instance2.instance5._10_[12] ;
 wire \modem.instance2.instance5._10_[13] ;
 wire \modem.instance2.instance5._10_[14] ;
 wire \modem.instance2.instance5._10_[15] ;
 wire \modem.instance2.instance5._10_[16] ;
 wire \modem.instance2.instance5._10_[17] ;
 wire \modem.instance2.instance5._10_[18] ;
 wire \modem.instance2.instance5._10_[19] ;
 wire \modem.instance2.instance5._10_[1] ;
 wire \modem.instance2.instance5._10_[20] ;
 wire \modem.instance2.instance5._10_[21] ;
 wire \modem.instance2.instance5._10_[22] ;
 wire \modem.instance2.instance5._10_[23] ;
 wire \modem.instance2.instance5._10_[24] ;
 wire \modem.instance2.instance5._10_[25] ;
 wire \modem.instance2.instance5._10_[26] ;
 wire \modem.instance2.instance5._10_[27] ;
 wire \modem.instance2.instance5._10_[28] ;
 wire \modem.instance2.instance5._10_[29] ;
 wire \modem.instance2.instance5._10_[2] ;
 wire \modem.instance2.instance5._10_[30] ;
 wire \modem.instance2.instance5._10_[31] ;
 wire \modem.instance2.instance5._10_[3] ;
 wire \modem.instance2.instance5._10_[4] ;
 wire \modem.instance2.instance5._10_[5] ;
 wire \modem.instance2.instance5._10_[6] ;
 wire \modem.instance2.instance5._10_[7] ;
 wire \modem.instance2.instance5._10_[8] ;
 wire \modem.instance2.instance5._10_[9] ;
 wire \modem.instance2.instance5.ffd0._0_ ;
 wire \modem.instance2.instance5.ffd1._0_ ;
 wire \modem.instance2.instance5.ffd3._0_ ;
 wire \modem.instance2.instance5.ffd4._0_ ;
 wire \modem.instance3._0_ ;
 wire \modem.instance3._1_ ;
 wire \modem.instance3._2_[0] ;
 wire \modem.instance3._2_[1] ;
 wire \modem.instance3._2_[2] ;
 wire \modem.instance3._2_[3] ;
 wire \modem.instance3._2_[4] ;
 wire \modem.instance3._2_[5] ;
 wire \modem.instance3._3_[0] ;
 wire \modem.instance3._3_[1] ;
 wire \modem.instance3._3_[2] ;
 wire \modem.instance3._3_[3] ;
 wire \modem.instance3._3_[4] ;
 wire \modem.instance3._3_[5] ;
 wire \modem.instance3.instance1._1_ ;
 wire \modem.instance3.instance1._3_[0] ;
 wire \modem.instance3.instance1._3_[1] ;
 wire \modem.instance3.instance1._3_[2] ;
 wire \modem.instance3.instance1._3_[3] ;
 wire \modem.instance3.instance1._3_[4] ;
 wire \modem.instance3.instance1._3_[5] ;
 wire \modem.instance3.instance1._3_[6] ;
 wire \modem.instance3.instance1._6_[0] ;
 wire \modem.instance3.instance1._6_[1] ;
 wire \modem.instance3.instance1._6_[2] ;
 wire \modem.instance3.instance1._6_[3] ;
 wire \modem.instance3.instance1._6_[4] ;
 wire \modem.instance3.instance1._6_[5] ;
 wire \modem.instance3.instance1._6_[6] ;
 wire \modem.instance3.instance2._00_ ;
 wire \modem.instance3.instance2._03_ ;
 wire \modem.instance3.instance2._04_ ;
 wire \modem.instance3.instance2._05_ ;
 wire \modem.instance3.instance2._09_[0] ;
 wire \modem.instance3.instance2._09_[10] ;
 wire \modem.instance3.instance2._09_[11] ;
 wire \modem.instance3.instance2._09_[12] ;
 wire \modem.instance3.instance2._09_[13] ;
 wire \modem.instance3.instance2._09_[14] ;
 wire \modem.instance3.instance2._09_[15] ;
 wire \modem.instance3.instance2._09_[16] ;
 wire \modem.instance3.instance2._09_[17] ;
 wire \modem.instance3.instance2._09_[18] ;
 wire \modem.instance3.instance2._09_[19] ;
 wire \modem.instance3.instance2._09_[1] ;
 wire \modem.instance3.instance2._09_[20] ;
 wire \modem.instance3.instance2._09_[21] ;
 wire \modem.instance3.instance2._09_[22] ;
 wire \modem.instance3.instance2._09_[23] ;
 wire \modem.instance3.instance2._09_[24] ;
 wire \modem.instance3.instance2._09_[25] ;
 wire \modem.instance3.instance2._09_[26] ;
 wire \modem.instance3.instance2._09_[27] ;
 wire \modem.instance3.instance2._09_[28] ;
 wire \modem.instance3.instance2._09_[29] ;
 wire \modem.instance3.instance2._09_[2] ;
 wire \modem.instance3.instance2._09_[30] ;
 wire \modem.instance3.instance2._09_[31] ;
 wire \modem.instance3.instance2._09_[3] ;
 wire \modem.instance3.instance2._09_[4] ;
 wire \modem.instance3.instance2._09_[5] ;
 wire \modem.instance3.instance2._09_[6] ;
 wire \modem.instance3.instance2._09_[7] ;
 wire \modem.instance3.instance2._09_[8] ;
 wire \modem.instance3.instance2._09_[9] ;
 wire \modem.instance3.instance2._10_[0] ;
 wire \modem.instance3.instance2._10_[10] ;
 wire \modem.instance3.instance2._10_[11] ;
 wire \modem.instance3.instance2._10_[12] ;
 wire \modem.instance3.instance2._10_[13] ;
 wire \modem.instance3.instance2._10_[14] ;
 wire \modem.instance3.instance2._10_[15] ;
 wire \modem.instance3.instance2._10_[16] ;
 wire \modem.instance3.instance2._10_[17] ;
 wire \modem.instance3.instance2._10_[18] ;
 wire \modem.instance3.instance2._10_[19] ;
 wire \modem.instance3.instance2._10_[1] ;
 wire \modem.instance3.instance2._10_[20] ;
 wire \modem.instance3.instance2._10_[21] ;
 wire \modem.instance3.instance2._10_[22] ;
 wire \modem.instance3.instance2._10_[23] ;
 wire \modem.instance3.instance2._10_[24] ;
 wire \modem.instance3.instance2._10_[25] ;
 wire \modem.instance3.instance2._10_[26] ;
 wire \modem.instance3.instance2._10_[27] ;
 wire \modem.instance3.instance2._10_[28] ;
 wire \modem.instance3.instance2._10_[29] ;
 wire \modem.instance3.instance2._10_[2] ;
 wire \modem.instance3.instance2._10_[30] ;
 wire \modem.instance3.instance2._10_[31] ;
 wire \modem.instance3.instance2._10_[3] ;
 wire \modem.instance3.instance2._10_[4] ;
 wire \modem.instance3.instance2._10_[5] ;
 wire \modem.instance3.instance2._10_[6] ;
 wire \modem.instance3.instance2._10_[7] ;
 wire \modem.instance3.instance2._10_[8] ;
 wire \modem.instance3.instance2._10_[9] ;
 wire \modem.instance3.instance2.ffd0._0_ ;
 wire \modem.instance3.instance2.ffd1._0_ ;
 wire \modem.instance3.instance2.ffd2._0_ ;
 wire \modem.instance3.instance2.ffd4._0_ ;
 wire \modem.instance3.instance3._0_[1] ;
 wire \modem.instance3.instance3._3_[0] ;
 wire \modem.instance3.instance3._3_[1] ;
 wire \modem.instance3.instance3._3_[2] ;
 wire \modem.instance3.instance3._3_[3] ;
 wire \modem.instance3.instance3._3_[4] ;
 wire \modem.instance3.instance3._4_[0] ;
 wire \modem.instance3.instance3._4_[2] ;
 wire \modem.instance3.instance3._4_[3] ;
 wire \modem.instance3.instance3._4_[4] ;
 wire \modem.instance3.instance4._0_[1] ;
 wire \modem.instance3.instance4._3_[0] ;
 wire \modem.instance3.instance4._3_[1] ;
 wire \modem.instance3.instance4._3_[2] ;
 wire \modem.instance3.instance4._3_[3] ;
 wire \modem.instance3.instance4._3_[4] ;
 wire \modem.instance3.instance4._4_[0] ;
 wire \modem.instance3.instance4._4_[2] ;
 wire \modem.instance3.instance4._4_[3] ;
 wire \modem.instance3.instance4._4_[4] ;
 wire \modem.instance4._5_[0] ;
 wire \modem.instance4._5_[1] ;
 wire \modem.instance4._5_[2] ;
 wire \modem.instance4._5_[3] ;
 wire \modem.instance4._5_[4] ;
 wire \modem.instance4._5_[5] ;
 wire \modem.instance6._1_ ;
 wire \modem.instance7._0_[0] ;
 wire \modem.instance7._0_[1] ;
 wire \modem.instance7._0_[2] ;
 wire \modem.instance7._0_[3] ;
 wire \modem.instance7._0_[4] ;
 wire \modem.instance7._0_[5] ;
 wire \modem.instance7._1_[0] ;
 wire \modem.instance7._1_[1] ;
 wire \modem.instance7._1_[2] ;
 wire \modem.instance7._1_[3] ;
 wire \modem.instance7._1_[4] ;
 wire \modem.instance7._1_[5] ;
 wire \modem.instance7._1_[6] ;
 wire \modem.instance7.instance2._0_[1] ;
 wire \modem.instance7.instance2._3_[0] ;
 wire \modem.instance7.instance2._3_[1] ;
 wire \modem.instance7.instance2._3_[2] ;
 wire \modem.instance7.instance2._3_[3] ;
 wire \modem.instance7.instance2._3_[4] ;
 wire \modem.instance7.instance2._4_[0] ;
 wire \modem.instance7.instance2._4_[2] ;
 wire \modem.instance7.instance2._4_[3] ;
 wire \modem.instance7.instance2._4_[4] ;
 wire \modem.instance7.instance3._0_[0] ;
 wire \modem.instance7.instance3._0_[1] ;
 wire \modem.instance7.instance3._0_[2] ;
 wire \modem.instance7.instance3._0_[3] ;
 wire \modem.instance7.instance3._0_[4] ;
 wire \modem.instance7.instance3._0_[5] ;
 wire \modem.instance7.instance4._7_ ;
 wire \modem.instance7.instance4._8_[0] ;
 wire \modem.instance7.instance4._8_[10] ;
 wire \modem.instance7.instance4._8_[11] ;
 wire \modem.instance7.instance4._8_[12] ;
 wire \modem.instance7.instance4._8_[13] ;
 wire \modem.instance7.instance4._8_[14] ;
 wire \modem.instance7.instance4._8_[15] ;
 wire \modem.instance7.instance4._8_[16] ;
 wire \modem.instance7.instance4._8_[17] ;
 wire \modem.instance7.instance4._8_[18] ;
 wire \modem.instance7.instance4._8_[19] ;
 wire \modem.instance7.instance4._8_[1] ;
 wire \modem.instance7.instance4._8_[20] ;
 wire \modem.instance7.instance4._8_[21] ;
 wire \modem.instance7.instance4._8_[22] ;
 wire \modem.instance7.instance4._8_[23] ;
 wire \modem.instance7.instance4._8_[24] ;
 wire \modem.instance7.instance4._8_[25] ;
 wire \modem.instance7.instance4._8_[26] ;
 wire \modem.instance7.instance4._8_[27] ;
 wire \modem.instance7.instance4._8_[28] ;
 wire \modem.instance7.instance4._8_[29] ;
 wire \modem.instance7.instance4._8_[2] ;
 wire \modem.instance7.instance4._8_[30] ;
 wire \modem.instance7.instance4._8_[31] ;
 wire \modem.instance7.instance4._8_[3] ;
 wire \modem.instance7.instance4._8_[4] ;
 wire \modem.instance7.instance4._8_[5] ;
 wire \modem.instance7.instance4._8_[6] ;
 wire \modem.instance7.instance4._8_[7] ;
 wire \modem.instance7.instance4._8_[8] ;
 wire \modem.instance7.instance4._8_[9] ;
 wire \modem.instance7.instance4._9_[0] ;
 wire \modem.instance7.instance4._9_[10] ;
 wire \modem.instance7.instance4._9_[11] ;
 wire \modem.instance7.instance4._9_[12] ;
 wire \modem.instance7.instance4._9_[13] ;
 wire \modem.instance7.instance4._9_[14] ;
 wire \modem.instance7.instance4._9_[15] ;
 wire \modem.instance7.instance4._9_[16] ;
 wire \modem.instance7.instance4._9_[17] ;
 wire \modem.instance7.instance4._9_[18] ;
 wire \modem.instance7.instance4._9_[19] ;
 wire \modem.instance7.instance4._9_[1] ;
 wire \modem.instance7.instance4._9_[20] ;
 wire \modem.instance7.instance4._9_[21] ;
 wire \modem.instance7.instance4._9_[22] ;
 wire \modem.instance7.instance4._9_[23] ;
 wire \modem.instance7.instance4._9_[24] ;
 wire \modem.instance7.instance4._9_[25] ;
 wire \modem.instance7.instance4._9_[26] ;
 wire \modem.instance7.instance4._9_[27] ;
 wire \modem.instance7.instance4._9_[28] ;
 wire \modem.instance7.instance4._9_[29] ;
 wire \modem.instance7.instance4._9_[2] ;
 wire \modem.instance7.instance4._9_[30] ;
 wire \modem.instance7.instance4._9_[31] ;
 wire \modem.instance7.instance4._9_[3] ;
 wire \modem.instance7.instance4._9_[4] ;
 wire \modem.instance7.instance4._9_[5] ;
 wire \modem.instance7.instance4._9_[6] ;
 wire \modem.instance7.instance4._9_[7] ;
 wire \modem.instance7.instance4._9_[8] ;
 wire \modem.instance7.instance4._9_[9] ;
 wire \modem.instance8._0_[0] ;
 wire \modem.instance8._0_[1] ;
 wire \modem.instance8._0_[2] ;
 wire \modem.instance8._0_[3] ;
 wire \modem.instance8._0_[4] ;
 wire \modem.instance8._0_[5] ;
 wire \modem.instance8._1_[0] ;
 wire \modem.instance8._1_[1] ;
 wire \modem.instance8._1_[2] ;
 wire \modem.instance8._1_[3] ;
 wire \modem.instance8._1_[4] ;
 wire \modem.instance8._1_[5] ;
 wire \modem.instance8.instance2._0_[1] ;
 wire \modem.instance8.instance2._3_[0] ;
 wire \modem.instance8.instance2._3_[1] ;
 wire \modem.instance8.instance2._3_[2] ;
 wire \modem.instance8.instance2._3_[3] ;
 wire \modem.instance8.instance2._3_[4] ;
 wire \modem.instance8.instance2._4_[0] ;
 wire \modem.instance8.instance2._4_[2] ;
 wire \modem.instance8.instance2._4_[3] ;
 wire \modem.instance8.instance2._4_[4] ;
 wire \modem.instance8.instance3._0_[0] ;
 wire \modem.instance8.instance3._0_[1] ;
 wire \modem.instance8.instance3._0_[2] ;
 wire \modem.instance8.instance3._0_[3] ;
 wire \modem.instance8.instance3._0_[4] ;
 wire \modem.instance8.instance3._0_[5] ;
 wire \modem.instance8.instance5._7_ ;
 wire \modem.instance8.instance5._8_[0] ;
 wire \modem.instance8.instance5._8_[10] ;
 wire \modem.instance8.instance5._8_[11] ;
 wire \modem.instance8.instance5._8_[12] ;
 wire \modem.instance8.instance5._8_[13] ;
 wire \modem.instance8.instance5._8_[14] ;
 wire \modem.instance8.instance5._8_[15] ;
 wire \modem.instance8.instance5._8_[16] ;
 wire \modem.instance8.instance5._8_[17] ;
 wire \modem.instance8.instance5._8_[18] ;
 wire \modem.instance8.instance5._8_[19] ;
 wire \modem.instance8.instance5._8_[1] ;
 wire \modem.instance8.instance5._8_[20] ;
 wire \modem.instance8.instance5._8_[21] ;
 wire \modem.instance8.instance5._8_[22] ;
 wire \modem.instance8.instance5._8_[23] ;
 wire \modem.instance8.instance5._8_[24] ;
 wire \modem.instance8.instance5._8_[25] ;
 wire \modem.instance8.instance5._8_[26] ;
 wire \modem.instance8.instance5._8_[27] ;
 wire \modem.instance8.instance5._8_[28] ;
 wire \modem.instance8.instance5._8_[29] ;
 wire \modem.instance8.instance5._8_[2] ;
 wire \modem.instance8.instance5._8_[30] ;
 wire \modem.instance8.instance5._8_[31] ;
 wire \modem.instance8.instance5._8_[3] ;
 wire \modem.instance8.instance5._8_[4] ;
 wire \modem.instance8.instance5._8_[5] ;
 wire \modem.instance8.instance5._8_[6] ;
 wire \modem.instance8.instance5._8_[7] ;
 wire \modem.instance8.instance5._8_[8] ;
 wire \modem.instance8.instance5._8_[9] ;
 wire \modem.instance8.instance5._9_[0] ;
 wire \modem.instance8.instance5._9_[10] ;
 wire \modem.instance8.instance5._9_[11] ;
 wire \modem.instance8.instance5._9_[12] ;
 wire \modem.instance8.instance5._9_[13] ;
 wire \modem.instance8.instance5._9_[14] ;
 wire \modem.instance8.instance5._9_[15] ;
 wire \modem.instance8.instance5._9_[16] ;
 wire \modem.instance8.instance5._9_[17] ;
 wire \modem.instance8.instance5._9_[18] ;
 wire \modem.instance8.instance5._9_[19] ;
 wire \modem.instance8.instance5._9_[1] ;
 wire \modem.instance8.instance5._9_[20] ;
 wire \modem.instance8.instance5._9_[21] ;
 wire \modem.instance8.instance5._9_[22] ;
 wire \modem.instance8.instance5._9_[23] ;
 wire \modem.instance8.instance5._9_[24] ;
 wire \modem.instance8.instance5._9_[25] ;
 wire \modem.instance8.instance5._9_[26] ;
 wire \modem.instance8.instance5._9_[27] ;
 wire \modem.instance8.instance5._9_[28] ;
 wire \modem.instance8.instance5._9_[29] ;
 wire \modem.instance8.instance5._9_[2] ;
 wire \modem.instance8.instance5._9_[30] ;
 wire \modem.instance8.instance5._9_[31] ;
 wire \modem.instance8.instance5._9_[3] ;
 wire \modem.instance8.instance5._9_[4] ;
 wire \modem.instance8.instance5._9_[5] ;
 wire \modem.instance8.instance5._9_[6] ;
 wire \modem.instance8.instance5._9_[7] ;
 wire \modem.instance8.instance5._9_[8] ;
 wire \modem.instance8.instance5._9_[9] ;
 wire \modem.instance9._5_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _1479_ (.A(\modem.instance2.instance4._4_[2] ),
    .X(_0831_));
 sg13g2_buf_1 _1480_ (.A(net58),
    .X(_0832_));
 sg13g2_buf_2 _1481_ (.A(\modem.instance2.instance4._4_[4] ),
    .X(_0833_));
 sg13g2_inv_2 _1482_ (.Y(_0834_),
    .A(_0833_));
 sg13g2_buf_1 _1483_ (.A(\modem.instance2.instance4._0_[1] ),
    .X(_0835_));
 sg13g2_buf_1 _1484_ (.A(_0835_),
    .X(_0836_));
 sg13g2_buf_1 _1485_ (.A(_0052_),
    .X(_0837_));
 sg13g2_buf_1 _1486_ (.A(_0837_),
    .X(_0838_));
 sg13g2_buf_1 _1487_ (.A(\modem.instance2.instance4._4_[3] ),
    .X(_0839_));
 sg13g2_buf_1 _1488_ (.A(_0839_),
    .X(_0840_));
 sg13g2_o21ai_1 _1489_ (.B1(net25),
    .Y(_0841_),
    .A1(_0836_),
    .A2(_0838_));
 sg13g2_buf_1 _1490_ (.A(_0833_),
    .X(_0842_));
 sg13g2_and3_1 _1491_ (.X(_0843_),
    .A(net24),
    .B(_0840_),
    .C(_0838_));
 sg13g2_a21oi_1 _1492_ (.A1(_0834_),
    .A2(_0841_),
    .Y(_0844_),
    .B1(_0843_));
 sg13g2_buf_1 _1493_ (.A(\modem.instance2.instance4._4_[0] ),
    .X(_0845_));
 sg13g2_buf_1 _1494_ (.A(_0845_),
    .X(_0846_));
 sg13g2_buf_1 _1495_ (.A(_0835_),
    .X(_0847_));
 sg13g2_nand2_1 _1496_ (.Y(_0848_),
    .A(_0846_),
    .B(net22));
 sg13g2_inv_1 _1497_ (.Y(_0849_),
    .A(_0839_));
 sg13g2_a21oi_1 _1498_ (.A1(net24),
    .A2(_0848_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_nand2b_1 _1499_ (.Y(_0851_),
    .B(net26),
    .A_N(_0847_));
 sg13g2_inv_1 _1500_ (.Y(\modem.instance2.instance4._3_[0] ),
    .A(_0845_));
 sg13g2_nand2_1 _1501_ (.Y(_0852_),
    .A(\modem.instance2.instance4._3_[0] ),
    .B(net22));
 sg13g2_nand2_1 _1502_ (.Y(_0853_),
    .A(net24),
    .B(_0849_));
 sg13g2_a21oi_1 _1503_ (.A1(_0851_),
    .A2(_0852_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor3_1 _1504_ (.A(_0832_),
    .B(_0850_),
    .C(_0854_),
    .Y(_0855_));
 sg13g2_a21oi_1 _1505_ (.A1(_0832_),
    .A2(_0844_),
    .Y(_0012_),
    .B1(_0855_));
 sg13g2_nand2b_1 _1506_ (.Y(_0856_),
    .B(_0840_),
    .A_N(_0835_));
 sg13g2_nand3_1 _1507_ (.B(net22),
    .C(net26),
    .A(_0833_),
    .Y(_0857_));
 sg13g2_a21oi_1 _1508_ (.A1(_0856_),
    .A2(_0857_),
    .Y(_0858_),
    .B1(\modem.instance2.instance4._3_[0] ));
 sg13g2_nand2_1 _1509_ (.Y(_0859_),
    .A(_0835_),
    .B(_0849_));
 sg13g2_nor2b_1 _1510_ (.A(net26),
    .B_N(_0835_),
    .Y(_0860_));
 sg13g2_o21ai_1 _1511_ (.B1(net21),
    .Y(_0861_),
    .A1(_0849_),
    .A2(_0860_));
 sg13g2_a21oi_1 _1512_ (.A1(_0859_),
    .A2(_0861_),
    .Y(_0862_),
    .B1(_0834_));
 sg13g2_nor2_1 _1513_ (.A(_0845_),
    .B(_0839_),
    .Y(_0863_));
 sg13g2_a21oi_1 _1514_ (.A1(_0833_),
    .A2(net22),
    .Y(_0864_),
    .B1(_0863_));
 sg13g2_nand2b_1 _1515_ (.Y(_0865_),
    .B(net21),
    .A_N(_0859_));
 sg13g2_o21ai_1 _1516_ (.B1(_0865_),
    .Y(_0866_),
    .A1(net28),
    .A2(_0864_));
 sg13g2_nor2b_1 _1517_ (.A(_0833_),
    .B_N(net58),
    .Y(_0867_));
 sg13g2_nand2_1 _1518_ (.Y(_0868_),
    .A(_0847_),
    .B(_0837_));
 sg13g2_nand3b_1 _1519_ (.B(net25),
    .C(net23),
    .Y(_0869_),
    .A_N(_0837_));
 sg13g2_o21ai_1 _1520_ (.B1(_0869_),
    .Y(_0870_),
    .A1(net23),
    .A2(_0868_));
 sg13g2_and2_1 _1521_ (.A(_0867_),
    .B(_0870_),
    .X(_0871_));
 sg13g2_nor4_1 _1522_ (.A(_0858_),
    .B(_0862_),
    .C(_0866_),
    .D(_0871_),
    .Y(_0013_));
 sg13g2_nand4_1 _1523_ (.B(net22),
    .C(net58),
    .A(net21),
    .Y(_0872_),
    .D(net26));
 sg13g2_o21ai_1 _1524_ (.B1(_0872_),
    .Y(_0873_),
    .A1(net21),
    .A2(net26));
 sg13g2_nand2_1 _1525_ (.Y(_0874_),
    .A(_0845_),
    .B(_0837_));
 sg13g2_o21ai_1 _1526_ (.B1(_0874_),
    .Y(_0875_),
    .A1(_0835_),
    .A2(net58));
 sg13g2_nor2b_1 _1527_ (.A(net58),
    .B_N(_0845_),
    .Y(_0876_));
 sg13g2_a21o_1 _1528_ (.A2(_0875_),
    .A1(_0834_),
    .B1(_0876_),
    .X(_0877_));
 sg13g2_a21oi_1 _1529_ (.A1(net24),
    .A2(_0873_),
    .Y(_0878_),
    .B1(_0877_));
 sg13g2_nand2_1 _1530_ (.Y(_0879_),
    .A(net58),
    .B(_0849_));
 sg13g2_nand2_1 _1531_ (.Y(_0880_),
    .A(_0834_),
    .B(_0876_));
 sg13g2_o21ai_1 _1532_ (.B1(_0880_),
    .Y(_0881_),
    .A1(net23),
    .A2(_0879_));
 sg13g2_o21ai_1 _1533_ (.B1(_0839_),
    .Y(_0882_),
    .A1(_0845_),
    .A2(_0837_));
 sg13g2_nor2_1 _1534_ (.A(_0831_),
    .B(_0839_),
    .Y(_0883_));
 sg13g2_a22oi_1 _1535_ (.Y(_0884_),
    .B1(_0883_),
    .B2(net21),
    .A2(_0882_),
    .A1(_0867_));
 sg13g2_nand2_1 _1536_ (.Y(_0885_),
    .A(net27),
    .B(_0884_));
 sg13g2_o21ai_1 _1537_ (.B1(_0885_),
    .Y(_0886_),
    .A1(net27),
    .A2(_0881_));
 sg13g2_o21ai_1 _1538_ (.B1(_0886_),
    .Y(_0014_),
    .A1(_0849_),
    .A2(_0878_));
 sg13g2_nand2b_1 _1539_ (.Y(_0887_),
    .B(_0834_),
    .A_N(_0865_));
 sg13g2_nand2_1 _1540_ (.Y(_0888_),
    .A(net58),
    .B(net25));
 sg13g2_nor2_1 _1541_ (.A(_0836_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_a21oi_1 _1542_ (.A1(_0856_),
    .A2(_0879_),
    .Y(_0890_),
    .B1(net24));
 sg13g2_o21ai_1 _1543_ (.B1(_0846_),
    .Y(_0891_),
    .A1(_0889_),
    .A2(_0890_));
 sg13g2_nand2_1 _1544_ (.Y(_0892_),
    .A(net21),
    .B(net25));
 sg13g2_o21ai_1 _1545_ (.B1(_0833_),
    .Y(_0893_),
    .A1(net22),
    .A2(_0863_));
 sg13g2_o21ai_1 _1546_ (.B1(_0893_),
    .Y(_0894_),
    .A1(net24),
    .A2(_0892_));
 sg13g2_nand2b_1 _1547_ (.Y(_0895_),
    .B(_0894_),
    .A_N(net28));
 sg13g2_nand3_1 _1548_ (.B(_0891_),
    .C(_0895_),
    .A(_0887_),
    .Y(_0015_));
 sg13g2_o21ai_1 _1549_ (.B1(_0892_),
    .Y(_0896_),
    .A1(_0833_),
    .A2(net26));
 sg13g2_nand3_1 _1550_ (.B(net25),
    .C(net26),
    .A(net58),
    .Y(_0897_));
 sg13g2_nand2b_1 _1551_ (.Y(_0898_),
    .B(_0897_),
    .A_N(_0883_));
 sg13g2_a22oi_1 _1552_ (.Y(_0899_),
    .B1(_0898_),
    .B2(net24),
    .A2(_0896_),
    .A1(net28));
 sg13g2_a21oi_1 _1553_ (.A1(net23),
    .A2(net22),
    .Y(_0900_),
    .B1(net25));
 sg13g2_o21ai_1 _1554_ (.B1(_0879_),
    .Y(_0901_),
    .A1(net28),
    .A2(_0900_));
 sg13g2_nand2_1 _1555_ (.Y(_0902_),
    .A(_0834_),
    .B(_0901_));
 sg13g2_o21ai_1 _1556_ (.B1(_0902_),
    .Y(_0016_),
    .A1(net27),
    .A2(_0899_));
 sg13g2_nand2b_1 _1557_ (.Y(_0903_),
    .B(_0851_),
    .A_N(_0888_));
 sg13g2_nor4_1 _1558_ (.A(_0842_),
    .B(net27),
    .C(net26),
    .D(_0888_),
    .Y(_0904_));
 sg13g2_a21oi_1 _1559_ (.A1(_0842_),
    .A2(_0903_),
    .Y(_0017_),
    .B1(_0904_));
 sg13g2_buf_1 _1560_ (.A(\modem.instance8.instance2._4_[2] ),
    .X(_0905_));
 sg13g2_buf_1 _1561_ (.A(_0905_),
    .X(_0906_));
 sg13g2_buf_2 _1562_ (.A(\modem.instance8.instance2._4_[3] ),
    .X(_0907_));
 sg13g2_buf_1 _1563_ (.A(_0907_),
    .X(_0908_));
 sg13g2_buf_2 _1564_ (.A(_0053_),
    .X(_0909_));
 sg13g2_and2_1 _1565_ (.A(_0909_),
    .B(\modem.instance8.instance2._4_[4] ),
    .X(_0910_));
 sg13g2_buf_1 _1566_ (.A(\modem.instance8.instance2._0_[1] ),
    .X(_0911_));
 sg13g2_or2_1 _1567_ (.X(_0912_),
    .B(_0909_),
    .A(net75));
 sg13g2_buf_1 _1568_ (.A(\modem.instance8.instance2._4_[4] ),
    .X(_0913_));
 sg13g2_a21oi_1 _1569_ (.A1(net56),
    .A2(_0912_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_a21oi_1 _1570_ (.A1(net56),
    .A2(_0910_),
    .Y(_0915_),
    .B1(_0914_));
 sg13g2_buf_1 _1571_ (.A(\modem.instance8.instance2._4_[0] ),
    .X(_0916_));
 sg13g2_nand2_1 _1572_ (.Y(_0917_),
    .A(_0916_),
    .B(net56));
 sg13g2_inv_1 _1573_ (.Y(\modem.instance8.instance2._3_[0] ),
    .A(_0916_));
 sg13g2_nor2b_1 _1574_ (.A(_0907_),
    .B_N(\modem.instance8.instance2._4_[4] ),
    .Y(_0918_));
 sg13g2_nand2_1 _1575_ (.Y(_0919_),
    .A(\modem.instance8.instance2._3_[0] ),
    .B(_0918_));
 sg13g2_inv_1 _1576_ (.Y(_0920_),
    .A(net75));
 sg13g2_a21oi_1 _1577_ (.A1(_0917_),
    .A2(_0919_),
    .Y(_0921_),
    .B1(_0920_));
 sg13g2_nor2b_1 _1578_ (.A(_0913_),
    .B_N(_0907_),
    .Y(_0922_));
 sg13g2_nand2_1 _1579_ (.Y(_0923_),
    .A(_0909_),
    .B(net74));
 sg13g2_nor3_1 _1580_ (.A(_0911_),
    .B(net56),
    .C(_0923_),
    .Y(_0924_));
 sg13g2_nor4_1 _1581_ (.A(_0906_),
    .B(_0921_),
    .C(_0922_),
    .D(_0924_),
    .Y(_0925_));
 sg13g2_a21oi_1 _1582_ (.A1(_0906_),
    .A2(_0915_),
    .Y(_0036_),
    .B1(_0925_));
 sg13g2_nand2b_1 _1583_ (.Y(_0926_),
    .B(_0905_),
    .A_N(\modem.instance8.instance2._4_[4] ));
 sg13g2_nor2b_1 _1584_ (.A(_0916_),
    .B_N(\modem.instance8.instance2._0_[1] ),
    .Y(_0927_));
 sg13g2_inv_2 _1585_ (.Y(_0928_),
    .A(_0907_));
 sg13g2_nor2_1 _1586_ (.A(_0928_),
    .B(_0909_),
    .Y(_0929_));
 sg13g2_buf_1 _1587_ (.A(_0916_),
    .X(_0930_));
 sg13g2_a22oi_1 _1588_ (.Y(_0931_),
    .B1(_0929_),
    .B2(net55),
    .A2(_0927_),
    .A1(_0909_));
 sg13g2_buf_1 _1589_ (.A(net75),
    .X(_0932_));
 sg13g2_inv_1 _1590_ (.Y(_0933_),
    .A(\modem.instance8.instance2._4_[4] ));
 sg13g2_or2_1 _1591_ (.X(_0934_),
    .B(_0907_),
    .A(_0916_));
 sg13g2_o21ai_1 _1592_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_0920_),
    .A2(_0933_));
 sg13g2_inv_2 _1593_ (.Y(_0936_),
    .A(_0905_));
 sg13g2_a22oi_1 _1594_ (.Y(_0937_),
    .B1(_0935_),
    .B2(_0936_),
    .A2(_0918_),
    .A1(net54));
 sg13g2_o21ai_1 _1595_ (.B1(_0937_),
    .Y(_0938_),
    .A1(_0926_),
    .A2(_0931_));
 sg13g2_nor2_1 _1596_ (.A(net75),
    .B(_0928_),
    .Y(_0939_));
 sg13g2_a21oi_1 _1597_ (.A1(net75),
    .A2(_0910_),
    .Y(_0940_),
    .B1(_0939_));
 sg13g2_o21ai_1 _1598_ (.B1(net56),
    .Y(_0941_),
    .A1(_0909_),
    .A2(_0933_));
 sg13g2_a221oi_1 _1599_ (.B2(net75),
    .C1(net55),
    .B1(_0941_),
    .A1(_0928_),
    .Y(_0942_),
    .A2(net74));
 sg13g2_a21oi_1 _1600_ (.A1(net55),
    .A2(_0940_),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_nor2_1 _1601_ (.A(_0938_),
    .B(_0943_),
    .Y(_0037_));
 sg13g2_nor2_1 _1602_ (.A(net75),
    .B(net74),
    .Y(_0944_));
 sg13g2_o21ai_1 _1603_ (.B1(_0936_),
    .Y(_0945_),
    .A1(net55),
    .A2(_0944_));
 sg13g2_xor2_1 _1604_ (.B(net74),
    .A(_0909_),
    .X(_0946_));
 sg13g2_and2_1 _1605_ (.A(_0910_),
    .B(_0927_),
    .X(_0947_));
 sg13g2_a22oi_1 _1606_ (.Y(_0948_),
    .B1(_0947_),
    .B2(net57),
    .A2(_0946_),
    .A1(_0930_));
 sg13g2_a21o_1 _1607_ (.A2(_0948_),
    .A1(_0945_),
    .B1(_0928_),
    .X(_0949_));
 sg13g2_nand3_1 _1608_ (.B(net57),
    .C(_0928_),
    .A(\modem.instance8.instance2._3_[0] ),
    .Y(_0950_));
 sg13g2_nand3_1 _1609_ (.B(_0936_),
    .C(_0933_),
    .A(_0930_),
    .Y(_0951_));
 sg13g2_a21o_1 _1610_ (.A2(_0951_),
    .A1(_0950_),
    .B1(net54),
    .X(_0952_));
 sg13g2_nor2_1 _1611_ (.A(_0907_),
    .B(_0926_),
    .Y(_0953_));
 sg13g2_nor2_1 _1612_ (.A(_0909_),
    .B(net74),
    .Y(_0954_));
 sg13g2_nor2_1 _1613_ (.A(_0905_),
    .B(_0907_),
    .Y(_0955_));
 sg13g2_a21oi_1 _1614_ (.A1(net57),
    .A2(_0954_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_nor2_1 _1615_ (.A(net55),
    .B(_0956_),
    .Y(_0957_));
 sg13g2_o21ai_1 _1616_ (.B1(net54),
    .Y(_0958_),
    .A1(_0953_),
    .A2(_0957_));
 sg13g2_nand3_1 _1617_ (.B(_0952_),
    .C(_0958_),
    .A(_0949_),
    .Y(_0038_));
 sg13g2_nand2_1 _1618_ (.Y(_0959_),
    .A(_0936_),
    .B(net74));
 sg13g2_a21o_1 _1619_ (.A2(_0959_),
    .A1(_0939_),
    .B1(_0953_),
    .X(_0960_));
 sg13g2_o21ai_1 _1620_ (.B1(_0959_),
    .Y(_0961_),
    .A1(net74),
    .A2(_0934_));
 sg13g2_nor2_1 _1621_ (.A(_0918_),
    .B(_0922_),
    .Y(_0962_));
 sg13g2_nor3_1 _1622_ (.A(net55),
    .B(net57),
    .C(_0962_),
    .Y(_0963_));
 sg13g2_a221oi_1 _1623_ (.B2(net54),
    .C1(_0963_),
    .B1(_0961_),
    .A1(net55),
    .Y(_0964_),
    .A2(_0960_));
 sg13g2_inv_1 _1624_ (.Y(_0039_),
    .A(_0964_));
 sg13g2_nand2_1 _1625_ (.Y(_0965_),
    .A(net55),
    .B(_0923_));
 sg13g2_nand3_1 _1626_ (.B(_0939_),
    .C(_0965_),
    .A(net57),
    .Y(_0966_));
 sg13g2_nand2_1 _1627_ (.Y(_0967_),
    .A(_0916_),
    .B(_0911_));
 sg13g2_a22oi_1 _1628_ (.Y(_0968_),
    .B1(_0955_),
    .B2(_0967_),
    .A2(_0912_),
    .A1(net57));
 sg13g2_o21ai_1 _1629_ (.B1(_0926_),
    .Y(_0969_),
    .A1(net75),
    .A2(_0959_));
 sg13g2_a22oi_1 _1630_ (.Y(_0970_),
    .B1(_0969_),
    .B2(_0928_),
    .A2(_0968_),
    .A1(_0933_));
 sg13g2_nand2_1 _1631_ (.Y(_0040_),
    .A(_0966_),
    .B(_0970_));
 sg13g2_nand2_1 _1632_ (.Y(_0971_),
    .A(net57),
    .B(net56));
 sg13g2_nand3_1 _1633_ (.B(net56),
    .C(_0954_),
    .A(net57),
    .Y(_0972_));
 sg13g2_a21oi_1 _1634_ (.A1(_0923_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(net54));
 sg13g2_a21oi_1 _1635_ (.A1(net74),
    .A2(_0971_),
    .Y(_0041_),
    .B1(_0973_));
 sg13g2_buf_1 _1636_ (.A(\modem.instance7.instance2._4_[2] ),
    .X(_0974_));
 sg13g2_buf_1 _1637_ (.A(_0974_),
    .X(_0975_));
 sg13g2_buf_2 _1638_ (.A(\modem.instance7.instance2._4_[3] ),
    .X(_0976_));
 sg13g2_buf_1 _1639_ (.A(_0976_),
    .X(_0977_));
 sg13g2_buf_2 _1640_ (.A(_0054_),
    .X(_0978_));
 sg13g2_and2_1 _1641_ (.A(_0978_),
    .B(\modem.instance7.instance2._4_[4] ),
    .X(_0979_));
 sg13g2_buf_1 _1642_ (.A(\modem.instance7.instance2._0_[1] ),
    .X(_0980_));
 sg13g2_or2_1 _1643_ (.X(_0981_),
    .B(_0978_),
    .A(net73));
 sg13g2_buf_1 _1644_ (.A(\modem.instance7.instance2._4_[4] ),
    .X(_0982_));
 sg13g2_a21oi_1 _1645_ (.A1(net52),
    .A2(_0981_),
    .Y(_0983_),
    .B1(net72));
 sg13g2_a21oi_1 _1646_ (.A1(net52),
    .A2(_0979_),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_buf_1 _1647_ (.A(\modem.instance7.instance2._4_[0] ),
    .X(_0985_));
 sg13g2_nand2_1 _1648_ (.Y(_0986_),
    .A(_0985_),
    .B(_0977_));
 sg13g2_inv_1 _1649_ (.Y(\modem.instance7.instance2._3_[0] ),
    .A(_0985_));
 sg13g2_nor2b_1 _1650_ (.A(_0976_),
    .B_N(\modem.instance7.instance2._4_[4] ),
    .Y(_0987_));
 sg13g2_nand2_1 _1651_ (.Y(_0988_),
    .A(\modem.instance7.instance2._3_[0] ),
    .B(_0987_));
 sg13g2_inv_1 _1652_ (.Y(_0989_),
    .A(net73));
 sg13g2_a21oi_1 _1653_ (.A1(_0986_),
    .A2(_0988_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_nor2b_1 _1654_ (.A(net72),
    .B_N(_0976_),
    .Y(_0991_));
 sg13g2_nand2_1 _1655_ (.Y(_0992_),
    .A(_0978_),
    .B(net72));
 sg13g2_nor3_1 _1656_ (.A(net73),
    .B(net52),
    .C(_0992_),
    .Y(_0993_));
 sg13g2_nor4_1 _1657_ (.A(net53),
    .B(_0990_),
    .C(_0991_),
    .D(_0993_),
    .Y(_0994_));
 sg13g2_a21oi_1 _1658_ (.A1(net53),
    .A2(_0984_),
    .Y(_0030_),
    .B1(_0994_));
 sg13g2_nand2b_1 _1659_ (.Y(_0995_),
    .B(_0974_),
    .A_N(\modem.instance7.instance2._4_[4] ));
 sg13g2_nor2b_1 _1660_ (.A(_0985_),
    .B_N(\modem.instance7.instance2._0_[1] ),
    .Y(_0996_));
 sg13g2_inv_2 _1661_ (.Y(_0997_),
    .A(_0976_));
 sg13g2_nor2_1 _1662_ (.A(_0997_),
    .B(_0978_),
    .Y(_0998_));
 sg13g2_buf_1 _1663_ (.A(_0985_),
    .X(_0999_));
 sg13g2_a22oi_1 _1664_ (.Y(_1000_),
    .B1(_0998_),
    .B2(net51),
    .A2(_0996_),
    .A1(_0978_));
 sg13g2_buf_1 _1665_ (.A(net73),
    .X(_1001_));
 sg13g2_inv_1 _1666_ (.Y(_1002_),
    .A(\modem.instance7.instance2._4_[4] ));
 sg13g2_or2_1 _1667_ (.X(_1003_),
    .B(_0976_),
    .A(_0985_));
 sg13g2_o21ai_1 _1668_ (.B1(_1003_),
    .Y(_1004_),
    .A1(_0989_),
    .A2(_1002_));
 sg13g2_inv_1 _1669_ (.Y(_1005_),
    .A(_0974_));
 sg13g2_a22oi_1 _1670_ (.Y(_1006_),
    .B1(_1004_),
    .B2(_1005_),
    .A2(_0987_),
    .A1(net50));
 sg13g2_o21ai_1 _1671_ (.B1(_1006_),
    .Y(_1007_),
    .A1(_0995_),
    .A2(_1000_));
 sg13g2_nor2_1 _1672_ (.A(net73),
    .B(_0997_),
    .Y(_1008_));
 sg13g2_a21oi_1 _1673_ (.A1(_0980_),
    .A2(_0979_),
    .Y(_1009_),
    .B1(_1008_));
 sg13g2_o21ai_1 _1674_ (.B1(_0977_),
    .Y(_1010_),
    .A1(_0978_),
    .A2(_1002_));
 sg13g2_a221oi_1 _1675_ (.B2(_0980_),
    .C1(net51),
    .B1(_1010_),
    .A1(_0997_),
    .Y(_1011_),
    .A2(_0982_));
 sg13g2_a21oi_1 _1676_ (.A1(net51),
    .A2(_1009_),
    .Y(_1012_),
    .B1(_1011_));
 sg13g2_nor2_1 _1677_ (.A(_1007_),
    .B(_1012_),
    .Y(_0031_));
 sg13g2_nor2_1 _1678_ (.A(net73),
    .B(_0982_),
    .Y(_1013_));
 sg13g2_o21ai_1 _1679_ (.B1(_1005_),
    .Y(_1014_),
    .A1(_0999_),
    .A2(_1013_));
 sg13g2_xor2_1 _1680_ (.B(net72),
    .A(_0978_),
    .X(_1015_));
 sg13g2_and2_1 _1681_ (.A(_0979_),
    .B(_0996_),
    .X(_1016_));
 sg13g2_a22oi_1 _1682_ (.Y(_1017_),
    .B1(_1016_),
    .B2(net53),
    .A2(_1015_),
    .A1(net51));
 sg13g2_a21o_1 _1683_ (.A2(_1017_),
    .A1(_1014_),
    .B1(_0997_),
    .X(_1018_));
 sg13g2_nand3_1 _1684_ (.B(_0975_),
    .C(_0997_),
    .A(\modem.instance7.instance2._3_[0] ),
    .Y(_1019_));
 sg13g2_nand3_1 _1685_ (.B(_1005_),
    .C(_1002_),
    .A(net51),
    .Y(_1020_));
 sg13g2_a21o_1 _1686_ (.A2(_1020_),
    .A1(_1019_),
    .B1(net50),
    .X(_1021_));
 sg13g2_nor2_1 _1687_ (.A(_0976_),
    .B(_0995_),
    .Y(_1022_));
 sg13g2_nor2_1 _1688_ (.A(_0978_),
    .B(net72),
    .Y(_1023_));
 sg13g2_nor2_1 _1689_ (.A(_0974_),
    .B(_0976_),
    .Y(_1024_));
 sg13g2_a21oi_1 _1690_ (.A1(net53),
    .A2(_1023_),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_nor2_1 _1691_ (.A(_0999_),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_o21ai_1 _1692_ (.B1(_1001_),
    .Y(_1027_),
    .A1(_1022_),
    .A2(_1026_));
 sg13g2_nand3_1 _1693_ (.B(_1021_),
    .C(_1027_),
    .A(_1018_),
    .Y(_0032_));
 sg13g2_nand2_1 _1694_ (.Y(_1028_),
    .A(_1005_),
    .B(net72));
 sg13g2_a21o_1 _1695_ (.A2(_1028_),
    .A1(_1008_),
    .B1(_1022_),
    .X(_1029_));
 sg13g2_o21ai_1 _1696_ (.B1(_1028_),
    .Y(_1030_),
    .A1(net72),
    .A2(_1003_));
 sg13g2_nor2_1 _1697_ (.A(_0987_),
    .B(_0991_),
    .Y(_1031_));
 sg13g2_nor3_1 _1698_ (.A(net51),
    .B(_0975_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_a221oi_1 _1699_ (.B2(_1001_),
    .C1(_1032_),
    .B1(_1030_),
    .A1(net51),
    .Y(_1033_),
    .A2(_1029_));
 sg13g2_inv_1 _1700_ (.Y(_0033_),
    .A(_1033_));
 sg13g2_nand2_1 _1701_ (.Y(_1034_),
    .A(net51),
    .B(_0992_));
 sg13g2_nand3_1 _1702_ (.B(_1008_),
    .C(_1034_),
    .A(net53),
    .Y(_1035_));
 sg13g2_nand2_1 _1703_ (.Y(_1036_),
    .A(_0985_),
    .B(net73));
 sg13g2_a22oi_1 _1704_ (.Y(_1037_),
    .B1(_1024_),
    .B2(_1036_),
    .A2(_0981_),
    .A1(net53));
 sg13g2_o21ai_1 _1705_ (.B1(_0995_),
    .Y(_1038_),
    .A1(net73),
    .A2(_1028_));
 sg13g2_a22oi_1 _1706_ (.Y(_1039_),
    .B1(_1038_),
    .B2(_0997_),
    .A2(_1037_),
    .A1(_1002_));
 sg13g2_nand2_1 _1707_ (.Y(_0034_),
    .A(_1035_),
    .B(_1039_));
 sg13g2_nand2_1 _1708_ (.Y(_1040_),
    .A(net53),
    .B(net52));
 sg13g2_nand3_1 _1709_ (.B(net52),
    .C(_1023_),
    .A(net53),
    .Y(_1041_));
 sg13g2_a21oi_1 _1710_ (.A1(_0992_),
    .A2(_1041_),
    .Y(_1042_),
    .B1(net50));
 sg13g2_a21oi_1 _1711_ (.A1(net72),
    .A2(_1040_),
    .Y(_0035_),
    .B1(_1042_));
 sg13g2_buf_1 _1712_ (.A(\modem.instance3.instance4._4_[2] ),
    .X(_1043_));
 sg13g2_buf_1 _1713_ (.A(_1043_),
    .X(_1044_));
 sg13g2_buf_1 _1714_ (.A(_0055_),
    .X(_1045_));
 sg13g2_inv_1 _1715_ (.Y(_1046_),
    .A(net70));
 sg13g2_buf_1 _1716_ (.A(\modem.instance3.instance4._4_[4] ),
    .X(_1047_));
 sg13g2_buf_1 _1717_ (.A(net69),
    .X(_1048_));
 sg13g2_buf_1 _1718_ (.A(\modem.instance3.instance4._4_[3] ),
    .X(_1049_));
 sg13g2_buf_1 _1719_ (.A(_1049_),
    .X(_1050_));
 sg13g2_nor2b_1 _1720_ (.A(net70),
    .B_N(net69),
    .Y(_1051_));
 sg13g2_nand2_1 _1721_ (.Y(_1052_),
    .A(_1050_),
    .B(_1051_));
 sg13g2_o21ai_1 _1722_ (.B1(_1052_),
    .Y(_1053_),
    .A1(_1046_),
    .A2(_1048_));
 sg13g2_buf_2 _1723_ (.A(\modem.instance3.instance4._4_[0] ),
    .X(_1054_));
 sg13g2_buf_1 _1724_ (.A(\modem.instance3.instance4._0_[1] ),
    .X(_1055_));
 sg13g2_nor2b_1 _1725_ (.A(_1054_),
    .B_N(net68),
    .Y(_1056_));
 sg13g2_buf_1 _1726_ (.A(net47),
    .X(_1057_));
 sg13g2_nor2_1 _1727_ (.A(net70),
    .B(net69),
    .Y(_1058_));
 sg13g2_and3_1 _1728_ (.X(_1059_),
    .A(_1049_),
    .B(net70),
    .C(net69));
 sg13g2_nand2b_1 _1729_ (.Y(_1060_),
    .B(net68),
    .A_N(_1054_));
 sg13g2_o21ai_1 _1730_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_1058_),
    .A2(_1059_));
 sg13g2_o21ai_1 _1731_ (.B1(_1061_),
    .Y(_1062_),
    .A1(_1057_),
    .A2(net48));
 sg13g2_a21o_1 _1732_ (.A2(_1056_),
    .A1(_1053_),
    .B1(_1062_),
    .X(_1063_));
 sg13g2_inv_2 _1733_ (.Y(_1064_),
    .A(net69));
 sg13g2_a21oi_1 _1734_ (.A1(net68),
    .A2(_1054_),
    .Y(_1065_),
    .B1(_1064_));
 sg13g2_and2_1 _1735_ (.A(_1057_),
    .B(_1065_),
    .X(_1066_));
 sg13g2_nor2_1 _1736_ (.A(_1054_),
    .B(_1064_),
    .Y(_1067_));
 sg13g2_buf_1 _1737_ (.A(_1054_),
    .X(_1068_));
 sg13g2_a21oi_1 _1738_ (.A1(net46),
    .A2(_1064_),
    .Y(_1069_),
    .B1(net68));
 sg13g2_nor3_1 _1739_ (.A(net20),
    .B(_1067_),
    .C(_1069_),
    .Y(_1070_));
 sg13g2_nor3_1 _1740_ (.A(net49),
    .B(_1066_),
    .C(_1070_),
    .Y(_1071_));
 sg13g2_a21oi_1 _1741_ (.A1(net49),
    .A2(_1063_),
    .Y(_0024_),
    .B1(_1071_));
 sg13g2_nand2_1 _1742_ (.Y(_1072_),
    .A(net71),
    .B(_1049_));
 sg13g2_nor2_1 _1743_ (.A(net70),
    .B(_1072_),
    .Y(_1073_));
 sg13g2_xnor2_1 _1744_ (.Y(_1074_),
    .A(_1064_),
    .B(_1073_));
 sg13g2_buf_1 _1745_ (.A(net68),
    .X(_1075_));
 sg13g2_buf_1 _1746_ (.A(_0056_),
    .X(_1076_));
 sg13g2_nand2b_1 _1747_ (.Y(_1077_),
    .B(_1076_),
    .A_N(net47));
 sg13g2_nor2_1 _1748_ (.A(net45),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_inv_1 _1749_ (.Y(_1079_),
    .A(net71));
 sg13g2_nor2_1 _1750_ (.A(_1079_),
    .B(net47),
    .Y(_1080_));
 sg13g2_o21ai_1 _1751_ (.B1(net45),
    .Y(_1081_),
    .A1(_0057_),
    .A2(_1080_));
 sg13g2_nand2b_1 _1752_ (.Y(_1082_),
    .B(_1081_),
    .A_N(_1078_));
 sg13g2_inv_1 _1753_ (.Y(_1083_),
    .A(_1055_));
 sg13g2_nand2_1 _1754_ (.Y(_1084_),
    .A(_1054_),
    .B(_1049_));
 sg13g2_nand2_1 _1755_ (.Y(_1085_),
    .A(_1049_),
    .B(net69));
 sg13g2_nor2_1 _1756_ (.A(_1043_),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_nor3_1 _1757_ (.A(net46),
    .B(net47),
    .C(net48),
    .Y(_1087_));
 sg13g2_nor3_1 _1758_ (.A(net44),
    .B(_1086_),
    .C(_1087_),
    .Y(_1088_));
 sg13g2_a21oi_1 _1759_ (.A1(net44),
    .A2(_1084_),
    .Y(_1089_),
    .B1(_1088_));
 sg13g2_a21o_1 _1760_ (.A2(_1082_),
    .A1(_1074_),
    .B1(_1089_),
    .X(_0025_));
 sg13g2_nor2_1 _1761_ (.A(net71),
    .B(net20),
    .Y(_1090_));
 sg13g2_o21ai_1 _1762_ (.B1(_1060_),
    .Y(_1091_),
    .A1(net68),
    .A2(net70));
 sg13g2_nor2_1 _1763_ (.A(_1054_),
    .B(_1049_),
    .Y(_1092_));
 sg13g2_nand2b_1 _1764_ (.Y(_1093_),
    .B(_1049_),
    .A_N(_0055_));
 sg13g2_nor2_1 _1765_ (.A(net44),
    .B(_1093_),
    .Y(_1094_));
 sg13g2_a21o_1 _1766_ (.A2(_1092_),
    .A1(net44),
    .B1(_1094_),
    .X(_1095_));
 sg13g2_a21oi_1 _1767_ (.A1(net71),
    .A2(_1045_),
    .Y(_1096_),
    .B1(_1084_));
 sg13g2_a221oi_1 _1768_ (.B2(net49),
    .C1(_1096_),
    .B1(_1095_),
    .A1(_1090_),
    .Y(_1097_),
    .A2(_1091_));
 sg13g2_nand2_1 _1769_ (.Y(_1098_),
    .A(net71),
    .B(net68));
 sg13g2_nand3_1 _1770_ (.B(net47),
    .C(net70),
    .A(_1054_),
    .Y(_1099_));
 sg13g2_nand3_1 _1771_ (.B(_1098_),
    .C(_1099_),
    .A(_1077_),
    .Y(_1100_));
 sg13g2_a21oi_1 _1772_ (.A1(net45),
    .A2(_1084_),
    .Y(_1101_),
    .B1(net49));
 sg13g2_nor3_1 _1773_ (.A(_1048_),
    .B(_1100_),
    .C(_1101_),
    .Y(_1102_));
 sg13g2_a21o_1 _1774_ (.A2(_1097_),
    .A1(net48),
    .B1(_1102_),
    .X(_0026_));
 sg13g2_nand2b_1 _1775_ (.Y(_1103_),
    .B(net69),
    .A_N(_1050_));
 sg13g2_nand3b_1 _1776_ (.B(net47),
    .C(_1058_),
    .Y(_1104_),
    .A_N(net46));
 sg13g2_o21ai_1 _1777_ (.B1(_1104_),
    .Y(_1105_),
    .A1(_1046_),
    .A2(_1103_));
 sg13g2_a21o_1 _1778_ (.A2(net70),
    .A1(net47),
    .B1(_1047_),
    .X(_1106_));
 sg13g2_a22oi_1 _1779_ (.Y(_1107_),
    .B1(_1106_),
    .B2(net46),
    .A2(_1093_),
    .A1(net48));
 sg13g2_nor2_1 _1780_ (.A(net44),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _1781_ (.B1(_1044_),
    .Y(_1109_),
    .A1(_1105_),
    .A2(_1108_));
 sg13g2_nand2b_1 _1782_ (.Y(_1110_),
    .B(net71),
    .A_N(net46));
 sg13g2_o21ai_1 _1783_ (.B1(_1110_),
    .Y(_1111_),
    .A1(net49),
    .A2(_1085_));
 sg13g2_nand2_1 _1784_ (.Y(_1112_),
    .A(net45),
    .B(_1064_));
 sg13g2_o21ai_1 _1785_ (.B1(_1112_),
    .Y(_1113_),
    .A1(net20),
    .A2(_1051_));
 sg13g2_nor2b_1 _1786_ (.A(net49),
    .B_N(net46),
    .Y(_1114_));
 sg13g2_a22oi_1 _1787_ (.Y(_1115_),
    .B1(_1113_),
    .B2(_1114_),
    .A2(_1111_),
    .A1(_1083_));
 sg13g2_nand2_1 _1788_ (.Y(_0027_),
    .A(_1109_),
    .B(_1115_));
 sg13g2_nor3_1 _1789_ (.A(_1079_),
    .B(net69),
    .C(_1084_),
    .Y(_1116_));
 sg13g2_a21o_1 _1790_ (.A2(_1067_),
    .A1(_1075_),
    .B1(_1116_),
    .X(_1117_));
 sg13g2_nor4_1 _1791_ (.A(net71),
    .B(net68),
    .C(net47),
    .D(net48),
    .Y(_1118_));
 sg13g2_a21o_1 _1792_ (.A2(_1051_),
    .A1(net49),
    .B1(_1118_),
    .X(_1119_));
 sg13g2_a22oi_1 _1793_ (.Y(_1120_),
    .B1(_1119_),
    .B2(_1068_),
    .A2(_1117_),
    .A1(_1045_));
 sg13g2_o21ai_1 _1794_ (.B1(_1075_),
    .Y(_1121_),
    .A1(net48),
    .A2(_1092_));
 sg13g2_nand2_1 _1795_ (.Y(_1122_),
    .A(_1085_),
    .B(_1121_));
 sg13g2_nand3_1 _1796_ (.B(_1056_),
    .C(_1058_),
    .A(net20),
    .Y(_1123_));
 sg13g2_nand3_1 _1797_ (.B(_1103_),
    .C(_1123_),
    .A(net49),
    .Y(_1124_));
 sg13g2_o21ai_1 _1798_ (.B1(_1124_),
    .Y(_1125_),
    .A1(_1044_),
    .A2(_1122_));
 sg13g2_nand2_1 _1799_ (.Y(_0028_),
    .A(_1120_),
    .B(_1125_));
 sg13g2_nand4_1 _1800_ (.B(net45),
    .C(net20),
    .A(net71),
    .Y(_1126_),
    .D(_1076_));
 sg13g2_nor2b_1 _1801_ (.A(_1074_),
    .B_N(_1126_),
    .Y(_1127_));
 sg13g2_and3_1 _1802_ (.X(_1128_),
    .A(net20),
    .B(_1056_),
    .C(_1074_));
 sg13g2_o21ai_1 _1803_ (.B1(_1079_),
    .Y(_1129_),
    .A1(net48),
    .A2(_1078_));
 sg13g2_o21ai_1 _1804_ (.B1(_1129_),
    .Y(_0029_),
    .A1(_1127_),
    .A2(_1128_));
 sg13g2_buf_1 _1805_ (.A(\modem.instance3.instance3._4_[2] ),
    .X(_1130_));
 sg13g2_buf_1 _1806_ (.A(_1130_),
    .X(_1131_));
 sg13g2_buf_1 _1807_ (.A(\modem.instance3.instance3._4_[3] ),
    .X(_1132_));
 sg13g2_buf_1 _1808_ (.A(net67),
    .X(_1133_));
 sg13g2_buf_2 _1809_ (.A(_0058_),
    .X(_1134_));
 sg13g2_buf_1 _1810_ (.A(\modem.instance3.instance3._4_[4] ),
    .X(_1135_));
 sg13g2_and2_1 _1811_ (.A(_1134_),
    .B(_1135_),
    .X(_1136_));
 sg13g2_buf_1 _1812_ (.A(\modem.instance3.instance3._0_[1] ),
    .X(_1137_));
 sg13g2_or2_1 _1813_ (.X(_1138_),
    .B(_1134_),
    .A(_1137_));
 sg13g2_buf_1 _1814_ (.A(_1135_),
    .X(_1139_));
 sg13g2_a21oi_1 _1815_ (.A1(net42),
    .A2(_1138_),
    .Y(_1140_),
    .B1(net41));
 sg13g2_a21oi_1 _1816_ (.A1(net42),
    .A2(_1136_),
    .Y(_1141_),
    .B1(_1140_));
 sg13g2_buf_1 _1817_ (.A(\modem.instance3.instance3._4_[0] ),
    .X(_1142_));
 sg13g2_nand2_1 _1818_ (.Y(_1143_),
    .A(_1142_),
    .B(net67));
 sg13g2_inv_1 _1819_ (.Y(\modem.instance3.instance3._3_[0] ),
    .A(_1142_));
 sg13g2_nor2b_1 _1820_ (.A(net67),
    .B_N(_1135_),
    .Y(_1144_));
 sg13g2_nand2_1 _1821_ (.Y(_1145_),
    .A(\modem.instance3.instance3._3_[0] ),
    .B(_1144_));
 sg13g2_inv_1 _1822_ (.Y(_1146_),
    .A(net66));
 sg13g2_a21oi_1 _1823_ (.A1(_1143_),
    .A2(_1145_),
    .Y(_1147_),
    .B1(_1146_));
 sg13g2_nor2b_1 _1824_ (.A(net41),
    .B_N(net67),
    .Y(_1148_));
 sg13g2_nand2_1 _1825_ (.Y(_1149_),
    .A(_1134_),
    .B(net41));
 sg13g2_nor3_1 _1826_ (.A(_1137_),
    .B(net42),
    .C(_1149_),
    .Y(_1150_));
 sg13g2_nor4_1 _1827_ (.A(net43),
    .B(_1147_),
    .C(_1148_),
    .D(_1150_),
    .Y(_1151_));
 sg13g2_a21oi_1 _1828_ (.A1(_1131_),
    .A2(_1141_),
    .Y(_0018_),
    .B1(_1151_));
 sg13g2_nand2b_1 _1829_ (.Y(_1152_),
    .B(_1130_),
    .A_N(_1135_));
 sg13g2_nor2b_1 _1830_ (.A(_1142_),
    .B_N(net66),
    .Y(_1153_));
 sg13g2_inv_1 _1831_ (.Y(_1154_),
    .A(net67));
 sg13g2_nor2_1 _1832_ (.A(_1154_),
    .B(_1134_),
    .Y(_1155_));
 sg13g2_buf_1 _1833_ (.A(_1142_),
    .X(_1156_));
 sg13g2_a22oi_1 _1834_ (.Y(_1157_),
    .B1(_1155_),
    .B2(_1156_),
    .A2(_1153_),
    .A1(_1134_));
 sg13g2_buf_1 _1835_ (.A(net66),
    .X(_1158_));
 sg13g2_inv_1 _1836_ (.Y(_1159_),
    .A(_1135_));
 sg13g2_or2_1 _1837_ (.X(_1160_),
    .B(net67),
    .A(_1142_));
 sg13g2_o21ai_1 _1838_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_1146_),
    .A2(_1159_));
 sg13g2_inv_1 _1839_ (.Y(_1162_),
    .A(_1130_));
 sg13g2_a22oi_1 _1840_ (.Y(_1163_),
    .B1(_1161_),
    .B2(_1162_),
    .A2(_1144_),
    .A1(net39));
 sg13g2_o21ai_1 _1841_ (.B1(_1163_),
    .Y(_1164_),
    .A1(_1152_),
    .A2(_1157_));
 sg13g2_nor2_1 _1842_ (.A(net66),
    .B(_1154_),
    .Y(_1165_));
 sg13g2_a21oi_1 _1843_ (.A1(_1158_),
    .A2(_1136_),
    .Y(_1166_),
    .B1(_1165_));
 sg13g2_o21ai_1 _1844_ (.B1(_1132_),
    .Y(_1167_),
    .A1(_1134_),
    .A2(_1159_));
 sg13g2_a221oi_1 _1845_ (.B2(net66),
    .C1(_1156_),
    .B1(_1167_),
    .A1(_1154_),
    .Y(_1168_),
    .A2(_1139_));
 sg13g2_a21oi_1 _1846_ (.A1(net40),
    .A2(_1166_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_nor2_1 _1847_ (.A(_1164_),
    .B(_1169_),
    .Y(_0019_));
 sg13g2_nor2_1 _1848_ (.A(net66),
    .B(net41),
    .Y(_1170_));
 sg13g2_o21ai_1 _1849_ (.B1(_1162_),
    .Y(_1171_),
    .A1(_1142_),
    .A2(_1170_));
 sg13g2_xor2_1 _1850_ (.B(_1139_),
    .A(_1134_),
    .X(_1172_));
 sg13g2_and2_1 _1851_ (.A(_1136_),
    .B(_1153_),
    .X(_1173_));
 sg13g2_a22oi_1 _1852_ (.Y(_0070_),
    .B1(_1173_),
    .B2(net43),
    .A2(_1172_),
    .A1(net40));
 sg13g2_a21o_1 _1853_ (.A2(_0070_),
    .A1(_1171_),
    .B1(_1154_),
    .X(_0071_));
 sg13g2_nand3_1 _1854_ (.B(_1130_),
    .C(_1154_),
    .A(\modem.instance3.instance3._3_[0] ),
    .Y(_0072_));
 sg13g2_nand3_1 _1855_ (.B(_1162_),
    .C(_1159_),
    .A(net40),
    .Y(_0073_));
 sg13g2_a21o_1 _1856_ (.A2(_0073_),
    .A1(_0072_),
    .B1(net39),
    .X(_0074_));
 sg13g2_nor2_1 _1857_ (.A(net67),
    .B(_1152_),
    .Y(_0075_));
 sg13g2_nor2_1 _1858_ (.A(_1134_),
    .B(_1135_),
    .Y(_0076_));
 sg13g2_nor2_1 _1859_ (.A(_1130_),
    .B(net67),
    .Y(_0077_));
 sg13g2_a21oi_1 _1860_ (.A1(_1130_),
    .A2(_0076_),
    .Y(_0078_),
    .B1(_0077_));
 sg13g2_nor2_1 _1861_ (.A(net40),
    .B(_0078_),
    .Y(_0079_));
 sg13g2_o21ai_1 _1862_ (.B1(net39),
    .Y(_0080_),
    .A1(_0075_),
    .A2(_0079_));
 sg13g2_nand3_1 _1863_ (.B(_0074_),
    .C(_0080_),
    .A(_0071_),
    .Y(_0020_));
 sg13g2_nand2_1 _1864_ (.Y(_0081_),
    .A(_1162_),
    .B(_1135_));
 sg13g2_a21o_1 _1865_ (.A2(_0081_),
    .A1(_1165_),
    .B1(_0075_),
    .X(_0082_));
 sg13g2_o21ai_1 _1866_ (.B1(_0081_),
    .Y(_0083_),
    .A1(net41),
    .A2(_1160_));
 sg13g2_nor2_1 _1867_ (.A(_1144_),
    .B(_1148_),
    .Y(_0084_));
 sg13g2_nor3_1 _1868_ (.A(net40),
    .B(net43),
    .C(_0084_),
    .Y(_0085_));
 sg13g2_a221oi_1 _1869_ (.B2(net39),
    .C1(_0085_),
    .B1(_0083_),
    .A1(net40),
    .Y(_0086_),
    .A2(_0082_));
 sg13g2_inv_1 _1870_ (.Y(_0021_),
    .A(_0086_));
 sg13g2_nand2_1 _1871_ (.Y(_0087_),
    .A(net40),
    .B(_1149_));
 sg13g2_nand3_1 _1872_ (.B(_1165_),
    .C(_0087_),
    .A(_1131_),
    .Y(_0088_));
 sg13g2_nand2_1 _1873_ (.Y(_0089_),
    .A(_1142_),
    .B(net66));
 sg13g2_a22oi_1 _1874_ (.Y(_0090_),
    .B1(_0077_),
    .B2(_0089_),
    .A2(_1138_),
    .A1(net43));
 sg13g2_o21ai_1 _1875_ (.B1(_1152_),
    .Y(_0091_),
    .A1(net66),
    .A2(_0081_));
 sg13g2_a22oi_1 _1876_ (.Y(_0092_),
    .B1(_0091_),
    .B2(_1154_),
    .A2(_0090_),
    .A1(_1159_));
 sg13g2_nand2_1 _1877_ (.Y(_0022_),
    .A(_0088_),
    .B(_0092_));
 sg13g2_nand3_1 _1878_ (.B(_1133_),
    .C(_0076_),
    .A(net43),
    .Y(_0093_));
 sg13g2_a21oi_1 _1879_ (.A1(_1149_),
    .A2(_0093_),
    .Y(_0094_),
    .B1(_1158_));
 sg13g2_a21oi_1 _1880_ (.A1(net43),
    .A2(_1133_),
    .Y(_0095_),
    .B1(_1159_));
 sg13g2_nor2_1 _1881_ (.A(_0094_),
    .B(_0095_),
    .Y(_0023_));
 sg13g2_buf_1 _1882_ (.A(\modem.instance1.instance3._4_[2] ),
    .X(_0096_));
 sg13g2_buf_1 _1883_ (.A(_0096_),
    .X(_0097_));
 sg13g2_buf_1 _1884_ (.A(\modem.instance1.instance3._4_[3] ),
    .X(_0098_));
 sg13g2_inv_2 _1885_ (.Y(_0099_),
    .A(_0098_));
 sg13g2_buf_1 _1886_ (.A(\modem.instance1.instance3._0_[1] ),
    .X(_0100_));
 sg13g2_inv_1 _1887_ (.Y(_0101_),
    .A(_0100_));
 sg13g2_buf_1 _1888_ (.A(_0059_),
    .X(_0102_));
 sg13g2_nand2_1 _1889_ (.Y(_0103_),
    .A(_0101_),
    .B(net65));
 sg13g2_inv_1 _1890_ (.Y(_0104_),
    .A(\modem.instance1.instance3._4_[0] ));
 sg13g2_buf_1 _1891_ (.A(_0100_),
    .X(_0105_));
 sg13g2_nand2_1 _1892_ (.Y(_0106_),
    .A(_0104_),
    .B(_0105_));
 sg13g2_buf_1 _1893_ (.A(\modem.instance1.instance3._4_[4] ),
    .X(_0107_));
 sg13g2_inv_2 _1894_ (.Y(_0108_),
    .A(net64));
 sg13g2_a21oi_1 _1895_ (.A1(_0103_),
    .A2(_0106_),
    .Y(_0109_),
    .B1(_0108_));
 sg13g2_buf_1 _1896_ (.A(net64),
    .X(_0110_));
 sg13g2_buf_1 _1897_ (.A(\modem.instance1.instance3._4_[0] ),
    .X(_0111_));
 sg13g2_nand2_2 _1898_ (.Y(_0112_),
    .A(net63),
    .B(_0100_));
 sg13g2_a21oi_1 _1899_ (.A1(net36),
    .A2(_0112_),
    .Y(_0113_),
    .B1(_0099_));
 sg13g2_a21oi_1 _1900_ (.A1(_0099_),
    .A2(_0109_),
    .Y(_0114_),
    .B1(_0113_));
 sg13g2_buf_1 _1901_ (.A(_0098_),
    .X(_0115_));
 sg13g2_nor3_1 _1902_ (.A(net64),
    .B(net37),
    .C(_0102_),
    .Y(_0116_));
 sg13g2_nand3_1 _1903_ (.B(net35),
    .C(net65),
    .A(net64),
    .Y(_0117_));
 sg13g2_o21ai_1 _1904_ (.B1(_0117_),
    .Y(_0118_),
    .A1(net36),
    .A2(_0115_));
 sg13g2_a22oi_1 _1905_ (.Y(_0119_),
    .B1(_0118_),
    .B2(_0097_),
    .A2(_0116_),
    .A1(net35));
 sg13g2_o21ai_1 _1906_ (.B1(_0119_),
    .Y(_0000_),
    .A1(net38),
    .A2(_0114_));
 sg13g2_buf_1 _1907_ (.A(_0104_),
    .X(\modem.instance1.instance3._3_[0] ));
 sg13g2_inv_1 _1908_ (.Y(_0120_),
    .A(_0059_));
 sg13g2_nand2_1 _1909_ (.Y(_0121_),
    .A(net34),
    .B(_0120_));
 sg13g2_o21ai_1 _1910_ (.B1(_0121_),
    .Y(_0122_),
    .A1(net38),
    .A2(_0101_));
 sg13g2_inv_1 _1911_ (.Y(_0123_),
    .A(_0096_));
 sg13g2_nor2_1 _1912_ (.A(_0108_),
    .B(_0123_),
    .Y(_0124_));
 sg13g2_nand2_1 _1913_ (.Y(_0125_),
    .A(net34),
    .B(net65));
 sg13g2_o21ai_1 _1914_ (.B1(_0125_),
    .Y(_0126_),
    .A1(net65),
    .A2(_0112_));
 sg13g2_nor2_1 _1915_ (.A(net63),
    .B(_0100_),
    .Y(_0127_));
 sg13g2_a221oi_1 _1916_ (.B2(_0126_),
    .C1(_0127_),
    .B1(_0124_),
    .A1(_0108_),
    .Y(_0128_),
    .A2(_0122_));
 sg13g2_a21oi_1 _1917_ (.A1(_0096_),
    .A2(_0101_),
    .Y(_0129_),
    .B1(_0111_));
 sg13g2_nand2b_1 _1918_ (.Y(_0130_),
    .B(\modem.instance1.instance3._4_[0] ),
    .A_N(_0100_));
 sg13g2_o21ai_1 _1919_ (.B1(_0130_),
    .Y(_0131_),
    .A1(net64),
    .A2(_0129_));
 sg13g2_nor3_1 _1920_ (.A(net36),
    .B(_0120_),
    .C(_0112_),
    .Y(_0132_));
 sg13g2_a21oi_1 _1921_ (.A1(_0099_),
    .A2(_0131_),
    .Y(_0133_),
    .B1(_0132_));
 sg13g2_o21ai_1 _1922_ (.B1(_0133_),
    .Y(_0001_),
    .A1(_0099_),
    .A2(_0128_));
 sg13g2_nand4_1 _1923_ (.B(_0096_),
    .C(net37),
    .A(net34),
    .Y(_0134_),
    .D(net65));
 sg13g2_o21ai_1 _1924_ (.B1(_0134_),
    .Y(_0135_),
    .A1(net34),
    .A2(net65));
 sg13g2_a22oi_1 _1925_ (.Y(_0136_),
    .B1(net65),
    .B2(net63),
    .A2(_0101_),
    .A1(_0123_));
 sg13g2_nand2_1 _1926_ (.Y(_0137_),
    .A(net63),
    .B(_0123_));
 sg13g2_o21ai_1 _1927_ (.B1(_0137_),
    .Y(_0138_),
    .A1(net64),
    .A2(_0136_));
 sg13g2_a21oi_1 _1928_ (.A1(net36),
    .A2(_0135_),
    .Y(_0139_),
    .B1(_0138_));
 sg13g2_nand2b_1 _1929_ (.Y(_0140_),
    .B(_0108_),
    .A_N(_0130_));
 sg13g2_o21ai_1 _1930_ (.B1(_0140_),
    .Y(_0141_),
    .A1(_0115_),
    .A2(_0106_));
 sg13g2_nor2b_1 _1931_ (.A(net64),
    .B_N(_0100_),
    .Y(_0142_));
 sg13g2_o21ai_1 _1932_ (.B1(_0098_),
    .Y(_0143_),
    .A1(net63),
    .A2(_0059_));
 sg13g2_a22oi_1 _1933_ (.Y(_0144_),
    .B1(_0142_),
    .B2(_0143_),
    .A2(_0127_),
    .A1(_0099_));
 sg13g2_nand2_1 _1934_ (.Y(_0145_),
    .A(net38),
    .B(_0144_));
 sg13g2_o21ai_1 _1935_ (.B1(_0145_),
    .Y(_0146_),
    .A1(net38),
    .A2(_0141_));
 sg13g2_o21ai_1 _1936_ (.B1(_0146_),
    .Y(_0002_),
    .A1(_0099_),
    .A2(_0139_));
 sg13g2_nor2_1 _1937_ (.A(net35),
    .B(_0111_),
    .Y(_0147_));
 sg13g2_o21ai_1 _1938_ (.B1(net64),
    .Y(_0148_),
    .A1(net37),
    .A2(_0147_));
 sg13g2_nand3_1 _1939_ (.B(net35),
    .C(net34),
    .A(_0108_),
    .Y(_0149_));
 sg13g2_a21oi_1 _1940_ (.A1(_0148_),
    .A2(_0149_),
    .Y(_0150_),
    .B1(_0097_));
 sg13g2_nor2_1 _1941_ (.A(_0098_),
    .B(_0096_),
    .Y(_0151_));
 sg13g2_a21oi_1 _1942_ (.A1(_0098_),
    .A2(_0105_),
    .Y(_0152_),
    .B1(_0151_));
 sg13g2_and2_1 _1943_ (.A(_0098_),
    .B(_0096_),
    .X(_0153_));
 sg13g2_buf_2 _1944_ (.A(_0153_),
    .X(_0154_));
 sg13g2_a22oi_1 _1945_ (.Y(_0155_),
    .B1(_0154_),
    .B2(_0101_),
    .A2(_0152_),
    .A1(_0108_));
 sg13g2_nand4_1 _1946_ (.B(_0099_),
    .C(net34),
    .A(_0108_),
    .Y(_0156_),
    .D(net37));
 sg13g2_o21ai_1 _1947_ (.B1(_0156_),
    .Y(_0157_),
    .A1(\modem.instance1.instance3._3_[0] ),
    .A2(_0155_));
 sg13g2_or2_1 _1948_ (.X(_0003_),
    .B(_0157_),
    .A(_0150_));
 sg13g2_nand2_1 _1949_ (.Y(_0158_),
    .A(\modem.instance1.instance3._3_[0] ),
    .B(_0096_));
 sg13g2_o21ai_1 _1950_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_0107_),
    .A2(_0102_));
 sg13g2_a21o_1 _1951_ (.A2(_0154_),
    .A1(net65),
    .B1(_0151_),
    .X(_0160_));
 sg13g2_a22oi_1 _1952_ (.Y(_0161_),
    .B1(_0160_),
    .B2(_0110_),
    .A2(_0159_),
    .A1(net35));
 sg13g2_a21oi_1 _1953_ (.A1(_0112_),
    .A2(_0151_),
    .Y(_0162_),
    .B1(_0154_));
 sg13g2_nand2_1 _1954_ (.Y(_0163_),
    .A(_0108_),
    .B(_0162_));
 sg13g2_o21ai_1 _1955_ (.B1(_0163_),
    .Y(_0004_),
    .A1(net37),
    .A2(_0161_));
 sg13g2_nand2_1 _1956_ (.Y(_0164_),
    .A(_0103_),
    .B(_0154_));
 sg13g2_a22oi_1 _1957_ (.Y(_0005_),
    .B1(_0164_),
    .B2(_0110_),
    .A2(_0154_),
    .A1(_0116_));
 sg13g2_buf_1 _1958_ (.A(\modem.instance2.instance3._4_[2] ),
    .X(_0165_));
 sg13g2_buf_1 _1959_ (.A(_0165_),
    .X(_0166_));
 sg13g2_buf_2 _1960_ (.A(\modem.instance2.instance3._4_[3] ),
    .X(_0167_));
 sg13g2_buf_1 _1961_ (.A(_0167_),
    .X(_0168_));
 sg13g2_buf_2 _1962_ (.A(_0047_),
    .X(_0169_));
 sg13g2_and2_1 _1963_ (.A(_0169_),
    .B(\modem.instance2.instance3._4_[4] ),
    .X(_0170_));
 sg13g2_buf_1 _1964_ (.A(\modem.instance2.instance3._0_[1] ),
    .X(_0171_));
 sg13g2_or2_1 _1965_ (.X(_0172_),
    .B(_0169_),
    .A(net62));
 sg13g2_buf_1 _1966_ (.A(\modem.instance2.instance3._4_[4] ),
    .X(_0173_));
 sg13g2_a21oi_1 _1967_ (.A1(net32),
    .A2(_0172_),
    .Y(_0174_),
    .B1(net61));
 sg13g2_a21oi_1 _1968_ (.A1(net32),
    .A2(_0170_),
    .Y(_0175_),
    .B1(_0174_));
 sg13g2_buf_1 _1969_ (.A(\modem.instance2.instance3._4_[0] ),
    .X(_0176_));
 sg13g2_nand2_1 _1970_ (.Y(_0177_),
    .A(_0176_),
    .B(net32));
 sg13g2_inv_1 _1971_ (.Y(\modem.instance2.instance3._3_[0] ),
    .A(_0176_));
 sg13g2_nor2b_1 _1972_ (.A(_0167_),
    .B_N(\modem.instance2.instance3._4_[4] ),
    .Y(_0178_));
 sg13g2_nand2_1 _1973_ (.Y(_0179_),
    .A(\modem.instance2.instance3._3_[0] ),
    .B(_0178_));
 sg13g2_inv_1 _1974_ (.Y(_0180_),
    .A(net62));
 sg13g2_a21oi_1 _1975_ (.A1(_0177_),
    .A2(_0179_),
    .Y(_0181_),
    .B1(_0180_));
 sg13g2_nor2b_1 _1976_ (.A(net61),
    .B_N(_0167_),
    .Y(_0182_));
 sg13g2_nand2_1 _1977_ (.Y(_0183_),
    .A(_0169_),
    .B(net61));
 sg13g2_nor3_1 _1978_ (.A(net62),
    .B(net32),
    .C(_0183_),
    .Y(_0184_));
 sg13g2_nor4_1 _1979_ (.A(net33),
    .B(_0181_),
    .C(_0182_),
    .D(_0184_),
    .Y(_0185_));
 sg13g2_a21oi_1 _1980_ (.A1(net33),
    .A2(_0175_),
    .Y(_0006_),
    .B1(_0185_));
 sg13g2_nand2b_1 _1981_ (.Y(_0186_),
    .B(_0165_),
    .A_N(\modem.instance2.instance3._4_[4] ));
 sg13g2_nor2b_1 _1982_ (.A(_0176_),
    .B_N(\modem.instance2.instance3._0_[1] ),
    .Y(_0187_));
 sg13g2_inv_2 _1983_ (.Y(_0188_),
    .A(_0167_));
 sg13g2_nor2_1 _1984_ (.A(_0188_),
    .B(_0169_),
    .Y(_0189_));
 sg13g2_buf_1 _1985_ (.A(_0176_),
    .X(_0190_));
 sg13g2_a22oi_1 _1986_ (.Y(_0191_),
    .B1(_0189_),
    .B2(net31),
    .A2(_0187_),
    .A1(_0169_));
 sg13g2_buf_1 _1987_ (.A(net62),
    .X(_0192_));
 sg13g2_inv_1 _1988_ (.Y(_0193_),
    .A(\modem.instance2.instance3._4_[4] ));
 sg13g2_or2_1 _1989_ (.X(_0194_),
    .B(_0167_),
    .A(_0176_));
 sg13g2_o21ai_1 _1990_ (.B1(_0194_),
    .Y(_0195_),
    .A1(_0180_),
    .A2(_0193_));
 sg13g2_inv_2 _1991_ (.Y(_0196_),
    .A(_0165_));
 sg13g2_a22oi_1 _1992_ (.Y(_0197_),
    .B1(_0195_),
    .B2(_0196_),
    .A2(_0178_),
    .A1(net30));
 sg13g2_o21ai_1 _1993_ (.B1(_0197_),
    .Y(_0198_),
    .A1(_0186_),
    .A2(_0191_));
 sg13g2_nor2_1 _1994_ (.A(net62),
    .B(_0188_),
    .Y(_0199_));
 sg13g2_a21oi_1 _1995_ (.A1(net62),
    .A2(_0170_),
    .Y(_0200_),
    .B1(_0199_));
 sg13g2_o21ai_1 _1996_ (.B1(_0168_),
    .Y(_0201_),
    .A1(_0169_),
    .A2(_0193_));
 sg13g2_a221oi_1 _1997_ (.B2(_0171_),
    .C1(net31),
    .B1(_0201_),
    .A1(_0188_),
    .Y(_0202_),
    .A2(net61));
 sg13g2_a21oi_1 _1998_ (.A1(net31),
    .A2(_0200_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nor2_1 _1999_ (.A(_0198_),
    .B(_0203_),
    .Y(_0007_));
 sg13g2_nor2_1 _2000_ (.A(_0171_),
    .B(_0173_),
    .Y(_0204_));
 sg13g2_o21ai_1 _2001_ (.B1(_0196_),
    .Y(_0205_),
    .A1(net31),
    .A2(_0204_));
 sg13g2_xor2_1 _2002_ (.B(_0173_),
    .A(_0169_),
    .X(_0206_));
 sg13g2_and2_1 _2003_ (.A(_0170_),
    .B(_0187_),
    .X(_0207_));
 sg13g2_a22oi_1 _2004_ (.Y(_0208_),
    .B1(_0207_),
    .B2(net33),
    .A2(_0206_),
    .A1(_0190_));
 sg13g2_a21o_1 _2005_ (.A2(_0208_),
    .A1(_0205_),
    .B1(_0188_),
    .X(_0209_));
 sg13g2_nand3_1 _2006_ (.B(_0166_),
    .C(_0188_),
    .A(\modem.instance2.instance3._3_[0] ),
    .Y(_0210_));
 sg13g2_nand3_1 _2007_ (.B(_0196_),
    .C(_0193_),
    .A(_0190_),
    .Y(_0211_));
 sg13g2_a21o_1 _2008_ (.A2(_0211_),
    .A1(_0210_),
    .B1(_0192_),
    .X(_0212_));
 sg13g2_nor2_1 _2009_ (.A(_0167_),
    .B(_0186_),
    .Y(_0213_));
 sg13g2_nor2_1 _2010_ (.A(_0169_),
    .B(net61),
    .Y(_0214_));
 sg13g2_nor2_1 _2011_ (.A(_0165_),
    .B(_0167_),
    .Y(_0215_));
 sg13g2_a21oi_1 _2012_ (.A1(net33),
    .A2(_0214_),
    .Y(_0216_),
    .B1(_0215_));
 sg13g2_nor2_1 _2013_ (.A(net31),
    .B(_0216_),
    .Y(_0217_));
 sg13g2_o21ai_1 _2014_ (.B1(net30),
    .Y(_0218_),
    .A1(_0213_),
    .A2(_0217_));
 sg13g2_nand3_1 _2015_ (.B(_0212_),
    .C(_0218_),
    .A(_0209_),
    .Y(_0008_));
 sg13g2_nand2_1 _2016_ (.Y(_0219_),
    .A(_0196_),
    .B(net61));
 sg13g2_a21o_1 _2017_ (.A2(_0219_),
    .A1(_0199_),
    .B1(_0213_),
    .X(_0220_));
 sg13g2_o21ai_1 _2018_ (.B1(_0219_),
    .Y(_0221_),
    .A1(net61),
    .A2(_0194_));
 sg13g2_nor2_1 _2019_ (.A(_0178_),
    .B(_0182_),
    .Y(_0222_));
 sg13g2_nor3_1 _2020_ (.A(net31),
    .B(net33),
    .C(_0222_),
    .Y(_0223_));
 sg13g2_a221oi_1 _2021_ (.B2(net30),
    .C1(_0223_),
    .B1(_0221_),
    .A1(net31),
    .Y(_0224_),
    .A2(_0220_));
 sg13g2_inv_1 _2022_ (.Y(_0009_),
    .A(_0224_));
 sg13g2_nand2_1 _2023_ (.Y(_0225_),
    .A(net31),
    .B(_0183_));
 sg13g2_nand3_1 _2024_ (.B(_0199_),
    .C(_0225_),
    .A(net33),
    .Y(_0226_));
 sg13g2_nand2_1 _2025_ (.Y(_0227_),
    .A(_0176_),
    .B(net62));
 sg13g2_a22oi_1 _2026_ (.Y(_0228_),
    .B1(_0215_),
    .B2(_0227_),
    .A2(_0172_),
    .A1(net33));
 sg13g2_o21ai_1 _2027_ (.B1(_0186_),
    .Y(_0229_),
    .A1(net62),
    .A2(_0219_));
 sg13g2_a22oi_1 _2028_ (.Y(_0230_),
    .B1(_0229_),
    .B2(_0188_),
    .A2(_0228_),
    .A1(_0193_));
 sg13g2_nand2_1 _2029_ (.Y(_0010_),
    .A(_0226_),
    .B(_0230_));
 sg13g2_nand2_1 _2030_ (.Y(_0231_),
    .A(_0166_),
    .B(_0168_));
 sg13g2_nand3_1 _2031_ (.B(net32),
    .C(_0214_),
    .A(net33),
    .Y(_0232_));
 sg13g2_a21oi_1 _2032_ (.A1(_0183_),
    .A2(_0232_),
    .Y(_0233_),
    .B1(net30));
 sg13g2_a21oi_1 _2033_ (.A1(net61),
    .A2(_0231_),
    .Y(_0011_),
    .B1(_0233_));
 sg13g2_or2_1 _2034_ (.X(_0234_),
    .B(\modem.instance1.instance1._6_[2] ),
    .A(\modem.instance1.instance1._6_[1] ));
 sg13g2_buf_2 _2035_ (.A(\modem.instance1.instance1._6_[3] ),
    .X(_0235_));
 sg13g2_nand2_1 _2036_ (.Y(_0236_),
    .A(_0235_),
    .B(\modem.instance1.instance1._6_[4] ));
 sg13g2_nor4_2 _2037_ (.A(\modem.instance1.instance1._6_[5] ),
    .B(\modem.instance1.instance1._6_[6] ),
    .C(_0234_),
    .Y(_0237_),
    .D(_0236_));
 sg13g2_nand2_1 _2038_ (.Y(_0238_),
    .A(\modem.instance1.instance1._6_[0] ),
    .B(_0237_));
 sg13g2_mux2_1 _2039_ (.A0(net97),
    .A1(\modem.instance1._0_ ),
    .S(_0238_),
    .X(_0063_));
 sg13g2_buf_2 _2040_ (.A(\modem.instance1._1_ ),
    .X(_0239_));
 sg13g2_buf_1 _2041_ (.A(\modem.instance1.instance2._10_[23] ),
    .X(_0240_));
 sg13g2_nor4_1 _2042_ (.A(\modem.instance1.instance2._10_[16] ),
    .B(\modem.instance1.instance2._10_[21] ),
    .C(\modem.instance1.instance2._10_[22] ),
    .D(_0240_),
    .Y(_0241_));
 sg13g2_nor4_1 _2043_ (.A(\modem.instance1.instance2._10_[17] ),
    .B(\modem.instance1.instance2._10_[18] ),
    .C(\modem.instance1.instance2._10_[19] ),
    .D(\modem.instance1.instance2._10_[20] ),
    .Y(_0242_));
 sg13g2_nor4_1 _2044_ (.A(\modem.instance1.instance2._10_[24] ),
    .B(\modem.instance1.instance2._10_[29] ),
    .C(\modem.instance1.instance2._10_[30] ),
    .D(\modem.instance1.instance2._10_[31] ),
    .Y(_0243_));
 sg13g2_nor4_1 _2045_ (.A(\modem.instance1.instance2._10_[25] ),
    .B(\modem.instance1.instance2._10_[26] ),
    .C(\modem.instance1.instance2._10_[27] ),
    .D(\modem.instance1.instance2._10_[28] ),
    .Y(_0244_));
 sg13g2_nand4_1 _2046_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0245_),
    .D(_0244_));
 sg13g2_nor4_1 _2047_ (.A(\modem.instance1.instance2._10_[7] ),
    .B(\modem.instance1.instance2._10_[12] ),
    .C(\modem.instance1.instance2._10_[13] ),
    .D(\modem.instance1.instance2._10_[14] ),
    .Y(_0246_));
 sg13g2_nor4_1 _2048_ (.A(\modem.instance1.instance2._10_[8] ),
    .B(\modem.instance1.instance2._10_[9] ),
    .C(\modem.instance1.instance2._10_[10] ),
    .D(\modem.instance1.instance2._10_[11] ),
    .Y(_0247_));
 sg13g2_buf_1 _2049_ (.A(\modem.instance1.instance2._10_[6] ),
    .X(_0248_));
 sg13g2_nor4_1 _2050_ (.A(\modem.instance1.instance2._10_[4] ),
    .B(\modem.instance1.instance2._10_[5] ),
    .C(_0248_),
    .D(\modem.instance1.instance2._10_[15] ),
    .Y(_0249_));
 sg13g2_inv_1 _2051_ (.Y(\modem.instance1.instance2._09_[0] ),
    .A(\modem.instance1.instance2._10_[0] ));
 sg13g2_nor4_1 _2052_ (.A(\modem.instance1.instance2._10_[1] ),
    .B(\modem.instance1.instance2._09_[0] ),
    .C(\modem.instance1.instance2._10_[2] ),
    .D(\modem.instance1.instance2._10_[3] ),
    .Y(_0250_));
 sg13g2_nand4_1 _2053_ (.B(_0247_),
    .C(_0249_),
    .A(_0246_),
    .Y(_0251_),
    .D(_0250_));
 sg13g2_nor2_1 _2054_ (.A(_0245_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_mux2_1 _2055_ (.A0(_0239_),
    .A1(\modem.instance1.instance2._05_ ),
    .S(_0252_),
    .X(_0064_));
 sg13g2_buf_1 _2056_ (.A(\modem.instance2.instance1._6_[1] ),
    .X(_0253_));
 sg13g2_buf_1 _2057_ (.A(\modem.instance2.instance1._6_[0] ),
    .X(_0254_));
 sg13g2_nand3_1 _2058_ (.B(\modem.instance2.instance1._6_[3] ),
    .C(\modem.instance2.instance1._6_[4] ),
    .A(_0254_),
    .Y(_0255_));
 sg13g2_or4_1 _2059_ (.A(\modem.instance2.instance1._6_[2] ),
    .B(\modem.instance2.instance1._6_[5] ),
    .C(\modem.instance2.instance1._6_[6] ),
    .D(_0255_),
    .X(_0256_));
 sg13g2_buf_1 _2060_ (.A(_0256_),
    .X(_0257_));
 sg13g2_nor2_1 _2061_ (.A(net60),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_mux2_1 _2062_ (.A0(\modem.instance2._0_ ),
    .A1(net89),
    .S(_0258_),
    .X(_0065_));
 sg13g2_inv_1 _2063_ (.Y(_0259_),
    .A(\modem.instance2.instance2._6_[3] ));
 sg13g2_nor4_1 _2064_ (.A(\modem.instance2.instance2._6_[2] ),
    .B(\modem.instance2.instance2._6_[5] ),
    .C(\modem.instance2.instance2._6_[4] ),
    .D(\modem.instance2.instance2._6_[6] ),
    .Y(_0260_));
 sg13g2_and2_1 _2065_ (.A(_0259_),
    .B(_0260_),
    .X(_0261_));
 sg13g2_nand3b_1 _2066_ (.B(\modem.instance2.instance2._6_[0] ),
    .C(_0261_),
    .Y(_0262_),
    .A_N(\modem.instance2.instance2._6_[1] ));
 sg13g2_mux2_1 _2067_ (.A0(\modem.instance2.instance2._1_ ),
    .A1(net83),
    .S(_0262_),
    .X(_0066_));
 sg13g2_buf_1 _2068_ (.A(\modem.instance2._4_ ),
    .X(_0263_));
 sg13g2_buf_1 _2069_ (.A(\modem.instance2.instance5._10_[23] ),
    .X(_0264_));
 sg13g2_nor4_1 _2070_ (.A(\modem.instance2.instance5._10_[16] ),
    .B(\modem.instance2.instance5._10_[21] ),
    .C(\modem.instance2.instance5._10_[22] ),
    .D(_0264_),
    .Y(_0265_));
 sg13g2_buf_1 _2071_ (.A(\modem.instance2.instance5._10_[18] ),
    .X(_0266_));
 sg13g2_nor4_1 _2072_ (.A(\modem.instance2.instance5._10_[17] ),
    .B(_0266_),
    .C(\modem.instance2.instance5._10_[19] ),
    .D(\modem.instance2.instance5._10_[20] ),
    .Y(_0267_));
 sg13g2_nor4_1 _2073_ (.A(\modem.instance2.instance5._10_[24] ),
    .B(\modem.instance2.instance5._10_[29] ),
    .C(\modem.instance2.instance5._10_[30] ),
    .D(\modem.instance2.instance5._10_[31] ),
    .Y(_0268_));
 sg13g2_buf_1 _2074_ (.A(\modem.instance2.instance5._10_[27] ),
    .X(_0269_));
 sg13g2_nor4_1 _2075_ (.A(\modem.instance2.instance5._10_[25] ),
    .B(\modem.instance2.instance5._10_[26] ),
    .C(_0269_),
    .D(\modem.instance2.instance5._10_[28] ),
    .Y(_0270_));
 sg13g2_nand4_1 _2076_ (.B(_0267_),
    .C(_0268_),
    .A(_0265_),
    .Y(_0271_),
    .D(_0270_));
 sg13g2_buf_1 _2077_ (.A(\modem.instance2.instance5._10_[14] ),
    .X(_0272_));
 sg13g2_nor4_1 _2078_ (.A(\modem.instance2.instance5._10_[7] ),
    .B(\modem.instance2.instance5._10_[12] ),
    .C(\modem.instance2.instance5._10_[13] ),
    .D(_0272_),
    .Y(_0273_));
 sg13g2_nor4_1 _2079_ (.A(\modem.instance2.instance5._10_[8] ),
    .B(\modem.instance2.instance5._10_[9] ),
    .C(\modem.instance2.instance5._10_[10] ),
    .D(\modem.instance2.instance5._10_[11] ),
    .Y(_0274_));
 sg13g2_buf_1 _2080_ (.A(\modem.instance2.instance5._10_[4] ),
    .X(_0275_));
 sg13g2_nor4_1 _2081_ (.A(_0275_),
    .B(\modem.instance2.instance5._10_[5] ),
    .C(\modem.instance2.instance5._10_[6] ),
    .D(\modem.instance2.instance5._10_[15] ),
    .Y(_0276_));
 sg13g2_inv_1 _2082_ (.Y(\modem.instance2.instance5._09_[0] ),
    .A(\modem.instance2.instance5._10_[0] ));
 sg13g2_nor4_1 _2083_ (.A(\modem.instance2.instance5._09_[0] ),
    .B(\modem.instance2.instance5._10_[1] ),
    .C(\modem.instance2.instance5._10_[2] ),
    .D(\modem.instance2.instance5._10_[3] ),
    .Y(_0277_));
 sg13g2_nand4_1 _2084_ (.B(_0274_),
    .C(_0276_),
    .A(_0273_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nor2_1 _2085_ (.A(_0271_),
    .B(_0278_),
    .Y(_0279_));
 sg13g2_mux2_1 _2086_ (.A0(_0263_),
    .A1(\modem.instance2.instance5._05_ ),
    .S(_0279_),
    .X(_0067_));
 sg13g2_buf_1 _2087_ (.A(\modem.instance3.instance1._6_[1] ),
    .X(_0280_));
 sg13g2_inv_1 _2088_ (.Y(\modem.instance3.instance1._3_[0] ),
    .A(\modem.instance3.instance1._6_[0] ));
 sg13g2_nor4_1 _2089_ (.A(\modem.instance3.instance1._3_[0] ),
    .B(\modem.instance3.instance1._6_[2] ),
    .C(\modem.instance3.instance1._6_[5] ),
    .D(\modem.instance3.instance1._6_[6] ),
    .Y(_0281_));
 sg13g2_nand3_1 _2090_ (.B(\modem.instance3.instance1._6_[4] ),
    .C(_0281_),
    .A(\modem.instance3.instance1._6_[3] ),
    .Y(_0282_));
 sg13g2_nor2_1 _2091_ (.A(net59),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_mux2_1 _2092_ (.A0(\modem.instance3._0_ ),
    .A1(net82),
    .S(_0283_),
    .X(_0068_));
 sg13g2_buf_2 _2093_ (.A(\modem.instance3._1_ ),
    .X(_0284_));
 sg13g2_nor4_1 _2094_ (.A(\modem.instance3.instance2._10_[17] ),
    .B(\modem.instance3.instance2._10_[20] ),
    .C(\modem.instance3.instance2._10_[23] ),
    .D(\modem.instance3.instance2._10_[22] ),
    .Y(_0285_));
 sg13g2_buf_1 _2095_ (.A(\modem.instance3.instance2._10_[16] ),
    .X(_0286_));
 sg13g2_nor4_1 _2096_ (.A(_0286_),
    .B(\modem.instance3.instance2._10_[19] ),
    .C(\modem.instance3.instance2._10_[18] ),
    .D(\modem.instance3.instance2._10_[21] ),
    .Y(_0287_));
 sg13g2_nor4_1 _2097_ (.A(\modem.instance3.instance2._10_[25] ),
    .B(\modem.instance3.instance2._10_[28] ),
    .C(\modem.instance3.instance2._10_[31] ),
    .D(\modem.instance3.instance2._10_[30] ),
    .Y(_0288_));
 sg13g2_nor4_1 _2098_ (.A(\modem.instance3.instance2._10_[24] ),
    .B(\modem.instance3.instance2._10_[27] ),
    .C(\modem.instance3.instance2._10_[26] ),
    .D(\modem.instance3.instance2._10_[29] ),
    .Y(_0289_));
 sg13g2_nand4_1 _2099_ (.B(_0287_),
    .C(_0288_),
    .A(_0285_),
    .Y(_0290_),
    .D(_0289_));
 sg13g2_nor4_1 _2100_ (.A(\modem.instance3.instance2._10_[6] ),
    .B(\modem.instance3.instance2._10_[13] ),
    .C(\modem.instance3.instance2._10_[12] ),
    .D(\modem.instance3.instance2._10_[15] ),
    .Y(_0291_));
 sg13g2_buf_1 _2101_ (.A(\modem.instance3.instance2._10_[8] ),
    .X(_0292_));
 sg13g2_nor4_1 _2102_ (.A(\modem.instance3.instance2._10_[9] ),
    .B(_0292_),
    .C(\modem.instance3.instance2._10_[11] ),
    .D(\modem.instance3.instance2._10_[10] ),
    .Y(_0293_));
 sg13g2_buf_2 _2103_ (.A(\modem.instance3.instance2._10_[4] ),
    .X(_0294_));
 sg13g2_nor4_1 _2104_ (.A(\modem.instance3.instance2._10_[5] ),
    .B(_0294_),
    .C(\modem.instance3.instance2._10_[7] ),
    .D(\modem.instance3.instance2._10_[14] ),
    .Y(_0295_));
 sg13g2_buf_8 _2105_ (.A(\modem.instance3.instance2._10_[1] ),
    .X(_0296_));
 sg13g2_buf_8 _2106_ (.A(\modem.instance3.instance2._10_[0] ),
    .X(_0297_));
 sg13g2_inv_1 _2107_ (.Y(\modem.instance3.instance2._09_[0] ),
    .A(_0297_));
 sg13g2_nor4_1 _2108_ (.A(_0296_),
    .B(\modem.instance3.instance2._09_[0] ),
    .C(\modem.instance3.instance2._10_[3] ),
    .D(\modem.instance3.instance2._10_[2] ),
    .Y(_0298_));
 sg13g2_nand4_1 _2109_ (.B(_0293_),
    .C(_0295_),
    .A(_0291_),
    .Y(_0299_),
    .D(_0298_));
 sg13g2_nor2_1 _2110_ (.A(_0290_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_mux2_1 _2111_ (.A0(_0284_),
    .A1(\modem.instance3.instance2._05_ ),
    .S(_0300_),
    .X(_0069_));
 sg13g2_xnor2_1 _2112_ (.Y(_0060_),
    .A(\modem.instance1.instance2._05_ ),
    .B(\modem.instance1.instance2._04_ ));
 sg13g2_xnor2_1 _2113_ (.Y(_0061_),
    .A(\modem.instance2.instance5._05_ ),
    .B(\modem.instance2.instance5._04_ ));
 sg13g2_xnor2_1 _2114_ (.Y(_0062_),
    .A(\modem.instance3.instance2._05_ ),
    .B(\modem.instance3.instance2._04_ ));
 sg13g2_inv_1 _2115_ (.Y(\modem.instance1.instance1._3_[0] ),
    .A(\modem.instance1.instance1._6_[0] ));
 sg13g2_nor3_1 _2116_ (.A(\modem.instance1.instance1._3_[0] ),
    .B(\modem.instance1.instance1._6_[1] ),
    .C(_0237_),
    .Y(_0301_));
 sg13g2_a21o_1 _2117_ (.A2(\modem.instance1.instance1._6_[1] ),
    .A1(\modem.instance1.instance1._3_[0] ),
    .B1(_0301_),
    .X(\modem.instance1.instance1._3_[1] ));
 sg13g2_nand2_1 _2118_ (.Y(_0302_),
    .A(\modem.instance1.instance1._6_[0] ),
    .B(\modem.instance1.instance1._6_[1] ));
 sg13g2_xnor2_1 _2119_ (.Y(\modem.instance1.instance1._3_[2] ),
    .A(\modem.instance1.instance1._6_[2] ),
    .B(_0302_));
 sg13g2_nand2_1 _2120_ (.Y(_0303_),
    .A(\modem.instance1.instance1._6_[1] ),
    .B(\modem.instance1.instance1._6_[2] ));
 sg13g2_nor3_1 _2121_ (.A(\modem.instance1.instance1._3_[0] ),
    .B(_0235_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_a21oi_1 _2122_ (.A1(_0235_),
    .A2(_0303_),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_nand2_1 _2123_ (.Y(_0306_),
    .A(\modem.instance1.instance1._3_[0] ),
    .B(_0235_));
 sg13g2_o21ai_1 _2124_ (.B1(_0306_),
    .Y(\modem.instance1.instance1._3_[3] ),
    .A1(_0237_),
    .A2(_0305_));
 sg13g2_and2_1 _2125_ (.A(\modem.instance1.instance1._6_[1] ),
    .B(\modem.instance1.instance1._6_[2] ),
    .X(_0307_));
 sg13g2_nand3_1 _2126_ (.B(_0235_),
    .C(_0307_),
    .A(\modem.instance1.instance1._6_[0] ),
    .Y(_0308_));
 sg13g2_a21oi_1 _2127_ (.A1(_0235_),
    .A2(_0307_),
    .Y(_0309_),
    .B1(_0237_));
 sg13g2_o21ai_1 _2128_ (.B1(\modem.instance1.instance1._6_[4] ),
    .Y(_0310_),
    .A1(\modem.instance1.instance1._3_[0] ),
    .A2(_0309_));
 sg13g2_o21ai_1 _2129_ (.B1(_0310_),
    .Y(\modem.instance1.instance1._3_[4] ),
    .A1(\modem.instance1.instance1._6_[4] ),
    .A2(_0308_));
 sg13g2_nand4_1 _2130_ (.B(_0235_),
    .C(\modem.instance1.instance1._6_[4] ),
    .A(\modem.instance1.instance1._6_[0] ),
    .Y(_0311_),
    .D(_0307_));
 sg13g2_xnor2_1 _2131_ (.Y(\modem.instance1.instance1._3_[5] ),
    .A(\modem.instance1.instance1._6_[5] ),
    .B(_0311_));
 sg13g2_inv_1 _2132_ (.Y(_0312_),
    .A(\modem.instance1.instance1._6_[5] ));
 sg13g2_nor2_1 _2133_ (.A(_0312_),
    .B(_0311_),
    .Y(_0313_));
 sg13g2_xor2_1 _2134_ (.B(_0313_),
    .A(\modem.instance1.instance1._6_[6] ),
    .X(\modem.instance1.instance1._3_[6] ));
 sg13g2_and4_1 _2135_ (.A(\modem.instance1.instance2._10_[1] ),
    .B(\modem.instance1.instance2._10_[0] ),
    .C(\modem.instance1.instance2._10_[2] ),
    .D(\modem.instance1.instance2._10_[3] ),
    .X(_0314_));
 sg13g2_buf_1 _2136_ (.A(_0314_),
    .X(_0315_));
 sg13g2_and4_1 _2137_ (.A(\modem.instance1.instance2._10_[5] ),
    .B(_0248_),
    .C(\modem.instance1.instance2._10_[7] ),
    .D(\modem.instance1.instance2._10_[8] ),
    .X(_0316_));
 sg13g2_nand4_1 _2138_ (.B(\modem.instance1.instance2._10_[9] ),
    .C(_0315_),
    .A(\modem.instance1.instance2._10_[4] ),
    .Y(_0317_),
    .D(_0316_));
 sg13g2_buf_2 _2139_ (.A(_0317_),
    .X(_0318_));
 sg13g2_xnor2_1 _2140_ (.Y(\modem.instance1.instance2._09_[10] ),
    .A(\modem.instance1.instance2._10_[10] ),
    .B(_0318_));
 sg13g2_inv_1 _2141_ (.Y(_0319_),
    .A(_0318_));
 sg13g2_nand2_1 _2142_ (.Y(_0320_),
    .A(\modem.instance1.instance2._10_[10] ),
    .B(_0319_));
 sg13g2_xnor2_1 _2143_ (.Y(\modem.instance1.instance2._09_[11] ),
    .A(\modem.instance1.instance2._10_[11] ),
    .B(_0320_));
 sg13g2_and3_1 _2144_ (.X(_0321_),
    .A(\modem.instance1.instance2._10_[10] ),
    .B(\modem.instance1.instance2._10_[11] ),
    .C(_0319_));
 sg13g2_xor2_1 _2145_ (.B(_0321_),
    .A(\modem.instance1.instance2._10_[12] ),
    .X(\modem.instance1.instance2._09_[12] ));
 sg13g2_nand3_1 _2146_ (.B(\modem.instance1.instance2._10_[11] ),
    .C(\modem.instance1.instance2._10_[12] ),
    .A(\modem.instance1.instance2._10_[10] ),
    .Y(_0322_));
 sg13g2_nor2_2 _2147_ (.A(_0318_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_xor2_1 _2148_ (.B(_0323_),
    .A(\modem.instance1.instance2._10_[13] ),
    .X(\modem.instance1.instance2._09_[13] ));
 sg13g2_nand2_1 _2149_ (.Y(_0324_),
    .A(\modem.instance1.instance2._10_[13] ),
    .B(_0323_));
 sg13g2_xnor2_1 _2150_ (.Y(\modem.instance1.instance2._09_[14] ),
    .A(\modem.instance1.instance2._10_[14] ),
    .B(_0324_));
 sg13g2_and3_1 _2151_ (.X(_0325_),
    .A(\modem.instance1.instance2._10_[13] ),
    .B(\modem.instance1.instance2._10_[14] ),
    .C(_0323_));
 sg13g2_xor2_1 _2152_ (.B(_0325_),
    .A(\modem.instance1.instance2._10_[15] ),
    .X(\modem.instance1.instance2._09_[15] ));
 sg13g2_and3_1 _2153_ (.X(_0326_),
    .A(\modem.instance1.instance2._10_[13] ),
    .B(\modem.instance1.instance2._10_[14] ),
    .C(\modem.instance1.instance2._10_[15] ));
 sg13g2_buf_1 _2154_ (.A(_0326_),
    .X(_0327_));
 sg13g2_nand2_1 _2155_ (.Y(_0328_),
    .A(_0323_),
    .B(_0327_));
 sg13g2_xnor2_1 _2156_ (.Y(\modem.instance1.instance2._09_[16] ),
    .A(\modem.instance1.instance2._10_[16] ),
    .B(_0328_));
 sg13g2_nand3_1 _2157_ (.B(_0323_),
    .C(_0327_),
    .A(\modem.instance1.instance2._10_[16] ),
    .Y(_0329_));
 sg13g2_xnor2_1 _2158_ (.Y(\modem.instance1.instance2._09_[17] ),
    .A(\modem.instance1.instance2._10_[17] ),
    .B(_0329_));
 sg13g2_and4_1 _2159_ (.A(\modem.instance1.instance2._10_[16] ),
    .B(\modem.instance1.instance2._10_[17] ),
    .C(_0323_),
    .D(_0327_),
    .X(_0330_));
 sg13g2_xor2_1 _2160_ (.B(_0330_),
    .A(\modem.instance1.instance2._10_[18] ),
    .X(\modem.instance1.instance2._09_[18] ));
 sg13g2_inv_1 _2161_ (.Y(_0331_),
    .A(\modem.instance1.instance2._10_[19] ));
 sg13g2_nand4_1 _2162_ (.B(\modem.instance1.instance2._10_[17] ),
    .C(\modem.instance1.instance2._10_[18] ),
    .A(\modem.instance1.instance2._10_[16] ),
    .Y(_0332_),
    .D(_0327_));
 sg13g2_nor3_1 _2163_ (.A(_0318_),
    .B(_0322_),
    .C(_0332_),
    .Y(_0333_));
 sg13g2_xnor2_1 _2164_ (.Y(\modem.instance1.instance2._09_[19] ),
    .A(_0331_),
    .B(_0333_));
 sg13g2_xnor2_1 _2165_ (.Y(_0334_),
    .A(\modem.instance1.instance2._10_[1] ),
    .B(\modem.instance1.instance2._10_[0] ));
 sg13g2_nor2_1 _2166_ (.A(_0252_),
    .B(_0334_),
    .Y(\modem.instance1.instance2._09_[1] ));
 sg13g2_nor4_2 _2167_ (.A(_0331_),
    .B(_0318_),
    .C(_0322_),
    .Y(_0335_),
    .D(_0332_));
 sg13g2_xor2_1 _2168_ (.B(_0335_),
    .A(\modem.instance1.instance2._10_[20] ),
    .X(\modem.instance1.instance2._09_[20] ));
 sg13g2_nand2_1 _2169_ (.Y(_0336_),
    .A(\modem.instance1.instance2._10_[20] ),
    .B(_0335_));
 sg13g2_xnor2_1 _2170_ (.Y(\modem.instance1.instance2._09_[21] ),
    .A(\modem.instance1.instance2._10_[21] ),
    .B(_0336_));
 sg13g2_nand3_1 _2171_ (.B(\modem.instance1.instance2._10_[21] ),
    .C(_0335_),
    .A(\modem.instance1.instance2._10_[20] ),
    .Y(_0337_));
 sg13g2_xnor2_1 _2172_ (.Y(\modem.instance1.instance2._09_[22] ),
    .A(\modem.instance1.instance2._10_[22] ),
    .B(_0337_));
 sg13g2_nand4_1 _2173_ (.B(\modem.instance1.instance2._10_[20] ),
    .C(\modem.instance1.instance2._10_[21] ),
    .A(\modem.instance1.instance2._10_[19] ),
    .Y(_0338_),
    .D(\modem.instance1.instance2._10_[22] ));
 sg13g2_nor4_1 _2174_ (.A(_0318_),
    .B(_0322_),
    .C(_0332_),
    .D(_0338_),
    .Y(_0339_));
 sg13g2_buf_1 _2175_ (.A(_0339_),
    .X(_0340_));
 sg13g2_xor2_1 _2176_ (.B(net10),
    .A(_0240_),
    .X(\modem.instance1.instance2._09_[23] ));
 sg13g2_nand2_1 _2177_ (.Y(_0341_),
    .A(_0240_),
    .B(net10));
 sg13g2_xnor2_1 _2178_ (.Y(\modem.instance1.instance2._09_[24] ),
    .A(\modem.instance1.instance2._10_[24] ),
    .B(_0341_));
 sg13g2_nand3_1 _2179_ (.B(\modem.instance1.instance2._10_[24] ),
    .C(net10),
    .A(_0240_),
    .Y(_0342_));
 sg13g2_xnor2_1 _2180_ (.Y(\modem.instance1.instance2._09_[25] ),
    .A(\modem.instance1.instance2._10_[25] ),
    .B(_0342_));
 sg13g2_nand4_1 _2181_ (.B(\modem.instance1.instance2._10_[24] ),
    .C(\modem.instance1.instance2._10_[25] ),
    .A(_0240_),
    .Y(_0343_),
    .D(_0340_));
 sg13g2_xnor2_1 _2182_ (.Y(\modem.instance1.instance2._09_[26] ),
    .A(\modem.instance1.instance2._10_[26] ),
    .B(_0343_));
 sg13g2_and4_1 _2183_ (.A(_0240_),
    .B(\modem.instance1.instance2._10_[24] ),
    .C(\modem.instance1.instance2._10_[25] ),
    .D(\modem.instance1.instance2._10_[26] ),
    .X(_0344_));
 sg13g2_nand2_1 _2184_ (.Y(_0345_),
    .A(net10),
    .B(_0344_));
 sg13g2_xnor2_1 _2185_ (.Y(\modem.instance1.instance2._09_[27] ),
    .A(\modem.instance1.instance2._10_[27] ),
    .B(_0345_));
 sg13g2_nand3_1 _2186_ (.B(net10),
    .C(_0344_),
    .A(\modem.instance1.instance2._10_[27] ),
    .Y(_0346_));
 sg13g2_xnor2_1 _2187_ (.Y(\modem.instance1.instance2._09_[28] ),
    .A(\modem.instance1.instance2._10_[28] ),
    .B(_0346_));
 sg13g2_and3_1 _2188_ (.X(_0347_),
    .A(\modem.instance1.instance2._10_[27] ),
    .B(\modem.instance1.instance2._10_[28] ),
    .C(_0344_));
 sg13g2_and2_1 _2189_ (.A(net10),
    .B(_0347_),
    .X(_0348_));
 sg13g2_xor2_1 _2190_ (.B(_0348_),
    .A(\modem.instance1.instance2._10_[29] ),
    .X(\modem.instance1.instance2._09_[29] ));
 sg13g2_nand2_1 _2191_ (.Y(_0349_),
    .A(\modem.instance1.instance2._10_[1] ),
    .B(\modem.instance1.instance2._10_[0] ));
 sg13g2_xnor2_1 _2192_ (.Y(\modem.instance1.instance2._09_[2] ),
    .A(\modem.instance1.instance2._10_[2] ),
    .B(_0349_));
 sg13g2_nand3_1 _2193_ (.B(net10),
    .C(_0347_),
    .A(\modem.instance1.instance2._10_[29] ),
    .Y(_0350_));
 sg13g2_xnor2_1 _2194_ (.Y(\modem.instance1.instance2._09_[30] ),
    .A(\modem.instance1.instance2._10_[30] ),
    .B(_0350_));
 sg13g2_nand4_1 _2195_ (.B(\modem.instance1.instance2._10_[30] ),
    .C(net10),
    .A(\modem.instance1.instance2._10_[29] ),
    .Y(_0351_),
    .D(_0347_));
 sg13g2_xnor2_1 _2196_ (.Y(\modem.instance1.instance2._09_[31] ),
    .A(\modem.instance1.instance2._10_[31] ),
    .B(_0351_));
 sg13g2_nand3_1 _2197_ (.B(\modem.instance1.instance2._10_[0] ),
    .C(\modem.instance1.instance2._10_[2] ),
    .A(\modem.instance1.instance2._10_[1] ),
    .Y(_0352_));
 sg13g2_xnor2_1 _2198_ (.Y(\modem.instance1.instance2._09_[3] ),
    .A(\modem.instance1.instance2._10_[3] ),
    .B(_0352_));
 sg13g2_xor2_1 _2199_ (.B(_0315_),
    .A(\modem.instance1.instance2._10_[4] ),
    .X(\modem.instance1.instance2._09_[4] ));
 sg13g2_nand2_1 _2200_ (.Y(_0353_),
    .A(\modem.instance1.instance2._10_[4] ),
    .B(_0315_));
 sg13g2_xnor2_1 _2201_ (.Y(\modem.instance1.instance2._09_[5] ),
    .A(\modem.instance1.instance2._10_[5] ),
    .B(_0353_));
 sg13g2_and3_1 _2202_ (.X(_0354_),
    .A(\modem.instance1.instance2._10_[4] ),
    .B(\modem.instance1.instance2._10_[5] ),
    .C(_0315_));
 sg13g2_buf_1 _2203_ (.A(_0354_),
    .X(_0355_));
 sg13g2_xor2_1 _2204_ (.B(_0355_),
    .A(_0248_),
    .X(\modem.instance1.instance2._09_[6] ));
 sg13g2_nand2_1 _2205_ (.Y(_0356_),
    .A(_0248_),
    .B(_0355_));
 sg13g2_xnor2_1 _2206_ (.Y(\modem.instance1.instance2._09_[7] ),
    .A(\modem.instance1.instance2._10_[7] ),
    .B(_0356_));
 sg13g2_nand3_1 _2207_ (.B(\modem.instance1.instance2._10_[7] ),
    .C(_0355_),
    .A(_0248_),
    .Y(_0357_));
 sg13g2_xnor2_1 _2208_ (.Y(\modem.instance1.instance2._09_[8] ),
    .A(\modem.instance1.instance2._10_[8] ),
    .B(_0357_));
 sg13g2_nand4_1 _2209_ (.B(\modem.instance1.instance2._10_[7] ),
    .C(\modem.instance1.instance2._10_[8] ),
    .A(_0248_),
    .Y(_0358_),
    .D(_0355_));
 sg13g2_xnor2_1 _2210_ (.Y(\modem.instance1.instance2._09_[9] ),
    .A(\modem.instance1.instance2._10_[9] ),
    .B(_0358_));
 sg13g2_a21o_1 _2211_ (.A2(_0154_),
    .A1(net36),
    .B1(_0130_),
    .X(_0359_));
 sg13g2_nand2_1 _2212_ (.Y(\modem.instance1.instance3._3_[1] ),
    .A(_0106_),
    .B(_0359_));
 sg13g2_a21oi_1 _2213_ (.A1(net36),
    .A2(net35),
    .Y(_0360_),
    .B1(net37));
 sg13g2_o21ai_1 _2214_ (.B1(net38),
    .Y(_0361_),
    .A1(net34),
    .A2(_0360_));
 sg13g2_o21ai_1 _2215_ (.B1(_0361_),
    .Y(\modem.instance1.instance3._3_[2] ),
    .A1(net38),
    .A2(_0112_));
 sg13g2_nand3_1 _2216_ (.B(net38),
    .C(net37),
    .A(net63),
    .Y(_0362_));
 sg13g2_nor2_1 _2217_ (.A(net36),
    .B(net37),
    .Y(_0363_));
 sg13g2_nand2_1 _2218_ (.Y(_0364_),
    .A(net63),
    .B(net38));
 sg13g2_o21ai_1 _2219_ (.B1(net35),
    .Y(_0365_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_o21ai_1 _2220_ (.B1(_0365_),
    .Y(\modem.instance1.instance3._3_[3] ),
    .A1(net35),
    .A2(_0362_));
 sg13g2_nand2_1 _2221_ (.Y(_0366_),
    .A(net63),
    .B(_0154_));
 sg13g2_mux2_1 _2222_ (.A0(_0142_),
    .A1(net36),
    .S(_0366_),
    .X(\modem.instance1.instance3._3_[4] ));
 sg13g2_and2_1 _2223_ (.A(_0239_),
    .B(\modem.instance1._2_[0] ),
    .X(\modem.instance1.instance4._0_[0] ));
 sg13g2_nand2b_1 _2224_ (.Y(\modem.instance1.instance4._0_[1] ),
    .B(_0239_),
    .A_N(\modem.instance1._2_[1] ));
 sg13g2_nand2b_1 _2225_ (.Y(\modem.instance1.instance4._0_[2] ),
    .B(_0239_),
    .A_N(\modem.instance1._2_[2] ));
 sg13g2_nand2b_1 _2226_ (.Y(\modem.instance1.instance4._0_[3] ),
    .B(_0239_),
    .A_N(\modem.instance1._2_[3] ));
 sg13g2_nand2b_1 _2227_ (.Y(\modem.instance1.instance4._0_[4] ),
    .B(_0239_),
    .A_N(\modem.instance1._2_[4] ));
 sg13g2_and2_1 _2228_ (.A(_0239_),
    .B(\modem.instance1._2_[5] ),
    .X(\modem.instance1.instance4._0_[5] ));
 sg13g2_inv_1 _2229_ (.Y(\modem.instance2.instance1._3_[0] ),
    .A(_0254_));
 sg13g2_nand2_1 _2230_ (.Y(_0367_),
    .A(_0254_),
    .B(_0257_));
 sg13g2_nand2_1 _2231_ (.Y(_0368_),
    .A(net60),
    .B(\modem.instance2.instance1._3_[0] ));
 sg13g2_o21ai_1 _2232_ (.B1(_0368_),
    .Y(\modem.instance2.instance1._3_[1] ),
    .A1(net60),
    .A2(_0367_));
 sg13g2_nand2_1 _2233_ (.Y(_0369_),
    .A(net60),
    .B(_0254_));
 sg13g2_xnor2_1 _2234_ (.Y(\modem.instance2.instance1._3_[2] ),
    .A(\modem.instance2.instance1._6_[2] ),
    .B(_0369_));
 sg13g2_nand2_1 _2235_ (.Y(_0370_),
    .A(\modem.instance2.instance1._6_[3] ),
    .B(_0257_));
 sg13g2_nand2_1 _2236_ (.Y(_0371_),
    .A(_0254_),
    .B(\modem.instance2.instance1._6_[2] ));
 sg13g2_xnor2_1 _2237_ (.Y(_0372_),
    .A(\modem.instance2.instance1._6_[3] ),
    .B(_0371_));
 sg13g2_nand2_1 _2238_ (.Y(_0373_),
    .A(net60),
    .B(_0372_));
 sg13g2_o21ai_1 _2239_ (.B1(_0373_),
    .Y(\modem.instance2.instance1._3_[3] ),
    .A1(net60),
    .A2(_0370_));
 sg13g2_nand2_1 _2240_ (.Y(_0374_),
    .A(\modem.instance2.instance1._6_[4] ),
    .B(_0257_));
 sg13g2_nand3_1 _2241_ (.B(\modem.instance2.instance1._6_[2] ),
    .C(\modem.instance2.instance1._6_[3] ),
    .A(_0254_),
    .Y(_0375_));
 sg13g2_xnor2_1 _2242_ (.Y(_0376_),
    .A(\modem.instance2.instance1._6_[4] ),
    .B(_0375_));
 sg13g2_nand2_1 _2243_ (.Y(_0377_),
    .A(net60),
    .B(_0376_));
 sg13g2_o21ai_1 _2244_ (.B1(_0377_),
    .Y(\modem.instance2.instance1._3_[4] ),
    .A1(net60),
    .A2(_0374_));
 sg13g2_nand2_1 _2245_ (.Y(_0378_),
    .A(_0253_),
    .B(\modem.instance2.instance1._6_[2] ));
 sg13g2_nor2_1 _2246_ (.A(_0255_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_xor2_1 _2247_ (.B(_0379_),
    .A(\modem.instance2.instance1._6_[5] ),
    .X(\modem.instance2.instance1._3_[5] ));
 sg13g2_nand2_1 _2248_ (.Y(_0380_),
    .A(\modem.instance2.instance1._6_[5] ),
    .B(_0379_));
 sg13g2_xnor2_1 _2249_ (.Y(\modem.instance2.instance1._3_[6] ),
    .A(\modem.instance2.instance1._6_[6] ),
    .B(_0380_));
 sg13g2_inv_1 _2250_ (.Y(\modem.instance2.instance2._3_[0] ),
    .A(\modem.instance2.instance2._6_[0] ));
 sg13g2_nor3_1 _2251_ (.A(\modem.instance2.instance2._6_[1] ),
    .B(\modem.instance2.instance2._3_[0] ),
    .C(_0261_),
    .Y(_0381_));
 sg13g2_a21o_1 _2252_ (.A2(\modem.instance2.instance2._3_[0] ),
    .A1(\modem.instance2.instance2._6_[1] ),
    .B1(_0381_),
    .X(\modem.instance2.instance2._3_[1] ));
 sg13g2_nand2_1 _2253_ (.Y(_0382_),
    .A(\modem.instance2.instance2._6_[1] ),
    .B(\modem.instance2.instance2._6_[0] ));
 sg13g2_xnor2_1 _2254_ (.Y(\modem.instance2.instance2._3_[2] ),
    .A(\modem.instance2.instance2._6_[2] ),
    .B(_0382_));
 sg13g2_nand3_1 _2255_ (.B(\modem.instance2.instance2._6_[0] ),
    .C(\modem.instance2.instance2._6_[2] ),
    .A(\modem.instance2.instance2._6_[1] ),
    .Y(_0383_));
 sg13g2_xnor2_1 _2256_ (.Y(\modem.instance2.instance2._3_[3] ),
    .A(\modem.instance2.instance2._6_[3] ),
    .B(_0383_));
 sg13g2_nor2_1 _2257_ (.A(_0259_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_xor2_1 _2258_ (.B(_0384_),
    .A(\modem.instance2.instance2._6_[4] ),
    .X(\modem.instance2.instance2._3_[4] ));
 sg13g2_nand2_1 _2259_ (.Y(_0385_),
    .A(\modem.instance2.instance2._6_[4] ),
    .B(_0384_));
 sg13g2_xnor2_1 _2260_ (.Y(\modem.instance2.instance2._3_[5] ),
    .A(\modem.instance2.instance2._6_[5] ),
    .B(_0385_));
 sg13g2_nand3_1 _2261_ (.B(\modem.instance2.instance2._6_[4] ),
    .C(_0384_),
    .A(\modem.instance2.instance2._6_[5] ),
    .Y(_0386_));
 sg13g2_xnor2_1 _2262_ (.Y(\modem.instance2.instance2._3_[6] ),
    .A(\modem.instance2.instance2._6_[6] ),
    .B(_0386_));
 sg13g2_nor2_1 _2263_ (.A(\modem.instance2.instance3._3_[0] ),
    .B(_0192_),
    .Y(_0387_));
 sg13g2_o21ai_1 _2264_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0050_),
    .A2(_0231_));
 sg13g2_nand2b_1 _2265_ (.Y(\modem.instance2.instance3._3_[1] ),
    .B(_0388_),
    .A_N(_0187_));
 sg13g2_inv_1 _2266_ (.Y(_0389_),
    .A(_0050_));
 sg13g2_a21o_1 _2267_ (.A2(_0389_),
    .A1(net32),
    .B1(net30),
    .X(_0390_));
 sg13g2_nor2_1 _2268_ (.A(\modem.instance2.instance3._3_[0] ),
    .B(_0196_),
    .Y(_0391_));
 sg13g2_a22oi_1 _2269_ (.Y(\modem.instance2.instance3._3_[2] ),
    .B1(_0390_),
    .B2(_0391_),
    .A2(_0227_),
    .A1(_0196_));
 sg13g2_nand2_1 _2270_ (.Y(_0392_),
    .A(net30),
    .B(_0391_));
 sg13g2_nand2_1 _2271_ (.Y(_0393_),
    .A(_0176_),
    .B(_0165_));
 sg13g2_nor2_1 _2272_ (.A(net30),
    .B(_0389_),
    .Y(_0394_));
 sg13g2_o21ai_1 _2273_ (.B1(net32),
    .Y(_0395_),
    .A1(_0393_),
    .A2(_0394_));
 sg13g2_o21ai_1 _2274_ (.B1(_0395_),
    .Y(\modem.instance2.instance3._3_[3] ),
    .A1(net32),
    .A2(_0392_));
 sg13g2_nor2_1 _2275_ (.A(_0188_),
    .B(_0393_),
    .Y(_0396_));
 sg13g2_nand3_1 _2276_ (.B(_0050_),
    .C(_0396_),
    .A(net30),
    .Y(_0397_));
 sg13g2_o21ai_1 _2277_ (.B1(_0397_),
    .Y(\modem.instance2.instance3._3_[4] ),
    .A1(_0050_),
    .A2(_0396_));
 sg13g2_nor2_1 _2278_ (.A(net21),
    .B(net27),
    .Y(_0398_));
 sg13g2_o21ai_1 _2279_ (.B1(_0398_),
    .Y(_0399_),
    .A1(_0834_),
    .A2(_0888_));
 sg13g2_nand2_1 _2280_ (.Y(\modem.instance2.instance4._3_[1] ),
    .A(_0852_),
    .B(_0399_));
 sg13g2_a21oi_1 _2281_ (.A1(_0833_),
    .A2(net25),
    .Y(_0400_),
    .B1(net22));
 sg13g2_nand2b_1 _2282_ (.Y(_0401_),
    .B(net23),
    .A_N(_0400_));
 sg13g2_a22oi_1 _2283_ (.Y(_0402_),
    .B1(_0401_),
    .B2(net28),
    .A2(_0876_),
    .A1(net27));
 sg13g2_inv_1 _2284_ (.Y(\modem.instance2.instance4._3_[2] ),
    .A(_0402_));
 sg13g2_nand3_1 _2285_ (.B(net27),
    .C(net28),
    .A(net23),
    .Y(_0403_));
 sg13g2_nand2_1 _2286_ (.Y(_0404_),
    .A(net23),
    .B(net28));
 sg13g2_nor3_1 _2287_ (.A(_0051_),
    .B(_0400_),
    .C(_0404_),
    .Y(_0405_));
 sg13g2_a21oi_1 _2288_ (.A1(_0051_),
    .A2(_0403_),
    .Y(\modem.instance2.instance4._3_[3] ),
    .B1(_0405_));
 sg13g2_nand3_1 _2289_ (.B(net28),
    .C(net25),
    .A(net23),
    .Y(_0406_));
 sg13g2_nand2_1 _2290_ (.Y(_0407_),
    .A(_0834_),
    .B(net27));
 sg13g2_nand2_1 _2291_ (.Y(_0408_),
    .A(net24),
    .B(_0406_));
 sg13g2_o21ai_1 _2292_ (.B1(_0408_),
    .Y(\modem.instance2.instance4._3_[4] ),
    .A1(_0406_),
    .A2(_0407_));
 sg13g2_inv_1 _2293_ (.Y(_0409_),
    .A(\modem.instance2.instance5._10_[10] ));
 sg13g2_inv_1 _2294_ (.Y(_0410_),
    .A(\modem.instance2.instance5._10_[9] ));
 sg13g2_and4_1 _2295_ (.A(\modem.instance2.instance5._10_[0] ),
    .B(\modem.instance2.instance5._10_[1] ),
    .C(\modem.instance2.instance5._10_[2] ),
    .D(\modem.instance2.instance5._10_[3] ),
    .X(_0411_));
 sg13g2_buf_1 _2296_ (.A(_0411_),
    .X(_0412_));
 sg13g2_and4_1 _2297_ (.A(_0275_),
    .B(\modem.instance2.instance5._10_[5] ),
    .C(\modem.instance2.instance5._10_[6] ),
    .D(\modem.instance2.instance5._10_[7] ),
    .X(_0413_));
 sg13g2_nand3_1 _2298_ (.B(_0412_),
    .C(_0413_),
    .A(\modem.instance2.instance5._10_[8] ),
    .Y(_0414_));
 sg13g2_buf_2 _2299_ (.A(_0414_),
    .X(_0415_));
 sg13g2_nor2_1 _2300_ (.A(_0410_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_xnor2_1 _2301_ (.Y(\modem.instance2.instance5._09_[10] ),
    .A(_0409_),
    .B(_0416_));
 sg13g2_nor3_1 _2302_ (.A(_0410_),
    .B(_0409_),
    .C(_0415_),
    .Y(_0417_));
 sg13g2_xor2_1 _2303_ (.B(_0417_),
    .A(\modem.instance2.instance5._10_[11] ),
    .X(\modem.instance2.instance5._09_[11] ));
 sg13g2_and2_1 _2304_ (.A(\modem.instance2.instance5._10_[11] ),
    .B(_0417_),
    .X(_0418_));
 sg13g2_xor2_1 _2305_ (.B(_0418_),
    .A(\modem.instance2.instance5._10_[12] ),
    .X(\modem.instance2.instance5._09_[12] ));
 sg13g2_and4_1 _2306_ (.A(\modem.instance2.instance5._10_[9] ),
    .B(\modem.instance2.instance5._10_[10] ),
    .C(\modem.instance2.instance5._10_[11] ),
    .D(\modem.instance2.instance5._10_[12] ),
    .X(_0419_));
 sg13g2_nor2b_1 _2307_ (.A(_0415_),
    .B_N(_0419_),
    .Y(_0420_));
 sg13g2_xor2_1 _2308_ (.B(_0420_),
    .A(\modem.instance2.instance5._10_[13] ),
    .X(\modem.instance2.instance5._09_[13] ));
 sg13g2_nand2_1 _2309_ (.Y(_0421_),
    .A(\modem.instance2.instance5._10_[13] ),
    .B(_0419_));
 sg13g2_nor2_2 _2310_ (.A(_0415_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_xor2_1 _2311_ (.B(_0422_),
    .A(_0272_),
    .X(\modem.instance2.instance5._09_[14] ));
 sg13g2_nand2_1 _2312_ (.Y(_0423_),
    .A(_0272_),
    .B(_0422_));
 sg13g2_xnor2_1 _2313_ (.Y(\modem.instance2.instance5._09_[15] ),
    .A(\modem.instance2.instance5._10_[15] ),
    .B(_0423_));
 sg13g2_nand3_1 _2314_ (.B(\modem.instance2.instance5._10_[15] ),
    .C(_0422_),
    .A(_0272_),
    .Y(_0424_));
 sg13g2_xnor2_1 _2315_ (.Y(\modem.instance2.instance5._09_[16] ),
    .A(\modem.instance2.instance5._10_[16] ),
    .B(_0424_));
 sg13g2_nand4_1 _2316_ (.B(\modem.instance2.instance5._10_[15] ),
    .C(\modem.instance2.instance5._10_[16] ),
    .A(_0272_),
    .Y(_0425_),
    .D(_0422_));
 sg13g2_xnor2_1 _2317_ (.Y(\modem.instance2.instance5._09_[17] ),
    .A(\modem.instance2.instance5._10_[17] ),
    .B(_0425_));
 sg13g2_and4_1 _2318_ (.A(_0272_),
    .B(\modem.instance2.instance5._10_[15] ),
    .C(\modem.instance2.instance5._10_[16] ),
    .D(\modem.instance2.instance5._10_[17] ),
    .X(_0426_));
 sg13g2_nand3_1 _2319_ (.B(_0419_),
    .C(_0426_),
    .A(\modem.instance2.instance5._10_[13] ),
    .Y(_0427_));
 sg13g2_nor2_2 _2320_ (.A(_0415_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_xor2_1 _2321_ (.B(_0428_),
    .A(_0266_),
    .X(\modem.instance2.instance5._09_[18] ));
 sg13g2_nand2_1 _2322_ (.Y(_0429_),
    .A(_0266_),
    .B(_0428_));
 sg13g2_xnor2_1 _2323_ (.Y(\modem.instance2.instance5._09_[19] ),
    .A(\modem.instance2.instance5._10_[19] ),
    .B(_0429_));
 sg13g2_xnor2_1 _2324_ (.Y(_0430_),
    .A(\modem.instance2.instance5._10_[0] ),
    .B(\modem.instance2.instance5._10_[1] ));
 sg13g2_nor2_1 _2325_ (.A(_0279_),
    .B(_0430_),
    .Y(\modem.instance2.instance5._09_[1] ));
 sg13g2_nand3_1 _2326_ (.B(\modem.instance2.instance5._10_[19] ),
    .C(_0428_),
    .A(_0266_),
    .Y(_0431_));
 sg13g2_xnor2_1 _2327_ (.Y(\modem.instance2.instance5._09_[20] ),
    .A(\modem.instance2.instance5._10_[20] ),
    .B(_0431_));
 sg13g2_nand4_1 _2328_ (.B(\modem.instance2.instance5._10_[19] ),
    .C(\modem.instance2.instance5._10_[20] ),
    .A(_0266_),
    .Y(_0432_),
    .D(_0428_));
 sg13g2_xnor2_1 _2329_ (.Y(\modem.instance2.instance5._09_[21] ),
    .A(\modem.instance2.instance5._10_[21] ),
    .B(_0432_));
 sg13g2_and4_1 _2330_ (.A(_0266_),
    .B(\modem.instance2.instance5._10_[19] ),
    .C(\modem.instance2.instance5._10_[20] ),
    .D(\modem.instance2.instance5._10_[21] ),
    .X(_0433_));
 sg13g2_nand2_1 _2331_ (.Y(_0434_),
    .A(_0428_),
    .B(_0433_));
 sg13g2_xnor2_1 _2332_ (.Y(\modem.instance2.instance5._09_[22] ),
    .A(\modem.instance2.instance5._10_[22] ),
    .B(_0434_));
 sg13g2_nand2_1 _2333_ (.Y(_0435_),
    .A(\modem.instance2.instance5._10_[22] ),
    .B(_0433_));
 sg13g2_nor3_1 _2334_ (.A(_0415_),
    .B(_0427_),
    .C(_0435_),
    .Y(_0436_));
 sg13g2_buf_1 _2335_ (.A(_0436_),
    .X(_0437_));
 sg13g2_xor2_1 _2336_ (.B(net9),
    .A(_0264_),
    .X(\modem.instance2.instance5._09_[23] ));
 sg13g2_nand2_1 _2337_ (.Y(_0438_),
    .A(_0264_),
    .B(net9));
 sg13g2_xnor2_1 _2338_ (.Y(\modem.instance2.instance5._09_[24] ),
    .A(\modem.instance2.instance5._10_[24] ),
    .B(_0438_));
 sg13g2_nand3_1 _2339_ (.B(\modem.instance2.instance5._10_[24] ),
    .C(net9),
    .A(_0264_),
    .Y(_0439_));
 sg13g2_xnor2_1 _2340_ (.Y(\modem.instance2.instance5._09_[25] ),
    .A(\modem.instance2.instance5._10_[25] ),
    .B(_0439_));
 sg13g2_nand4_1 _2341_ (.B(\modem.instance2.instance5._10_[24] ),
    .C(\modem.instance2.instance5._10_[25] ),
    .A(_0264_),
    .Y(_0440_),
    .D(net9));
 sg13g2_xnor2_1 _2342_ (.Y(\modem.instance2.instance5._09_[26] ),
    .A(\modem.instance2.instance5._10_[26] ),
    .B(_0440_));
 sg13g2_and4_1 _2343_ (.A(_0264_),
    .B(\modem.instance2.instance5._10_[24] ),
    .C(\modem.instance2.instance5._10_[25] ),
    .D(\modem.instance2.instance5._10_[26] ),
    .X(_0441_));
 sg13g2_buf_1 _2344_ (.A(_0441_),
    .X(_0442_));
 sg13g2_nand2_1 _2345_ (.Y(_0443_),
    .A(_0437_),
    .B(_0442_));
 sg13g2_xnor2_1 _2346_ (.Y(\modem.instance2.instance5._09_[27] ),
    .A(_0269_),
    .B(_0443_));
 sg13g2_nand3_1 _2347_ (.B(net9),
    .C(_0442_),
    .A(_0269_),
    .Y(_0444_));
 sg13g2_xnor2_1 _2348_ (.Y(\modem.instance2.instance5._09_[28] ),
    .A(\modem.instance2.instance5._10_[28] ),
    .B(_0444_));
 sg13g2_nand4_1 _2349_ (.B(\modem.instance2.instance5._10_[28] ),
    .C(net9),
    .A(_0269_),
    .Y(_0445_),
    .D(_0442_));
 sg13g2_xnor2_1 _2350_ (.Y(\modem.instance2.instance5._09_[29] ),
    .A(\modem.instance2.instance5._10_[29] ),
    .B(_0445_));
 sg13g2_nand2_1 _2351_ (.Y(_0446_),
    .A(\modem.instance2.instance5._10_[0] ),
    .B(\modem.instance2.instance5._10_[1] ));
 sg13g2_xnor2_1 _2352_ (.Y(\modem.instance2.instance5._09_[2] ),
    .A(\modem.instance2.instance5._10_[2] ),
    .B(_0446_));
 sg13g2_and2_1 _2353_ (.A(\modem.instance2.instance5._10_[28] ),
    .B(\modem.instance2.instance5._10_[29] ),
    .X(_0447_));
 sg13g2_nand4_1 _2354_ (.B(net9),
    .C(_0442_),
    .A(_0269_),
    .Y(_0448_),
    .D(_0447_));
 sg13g2_xnor2_1 _2355_ (.Y(\modem.instance2.instance5._09_[30] ),
    .A(\modem.instance2.instance5._10_[30] ),
    .B(_0448_));
 sg13g2_and2_1 _2356_ (.A(\modem.instance2.instance5._10_[30] ),
    .B(_0447_),
    .X(_0449_));
 sg13g2_nand4_1 _2357_ (.B(net9),
    .C(_0442_),
    .A(_0269_),
    .Y(_0450_),
    .D(_0449_));
 sg13g2_xnor2_1 _2358_ (.Y(\modem.instance2.instance5._09_[31] ),
    .A(\modem.instance2.instance5._10_[31] ),
    .B(_0450_));
 sg13g2_nand3_1 _2359_ (.B(\modem.instance2.instance5._10_[1] ),
    .C(\modem.instance2.instance5._10_[2] ),
    .A(\modem.instance2.instance5._10_[0] ),
    .Y(_0451_));
 sg13g2_xnor2_1 _2360_ (.Y(\modem.instance2.instance5._09_[3] ),
    .A(\modem.instance2.instance5._10_[3] ),
    .B(_0451_));
 sg13g2_xor2_1 _2361_ (.B(_0412_),
    .A(_0275_),
    .X(\modem.instance2.instance5._09_[4] ));
 sg13g2_nand2_1 _2362_ (.Y(_0452_),
    .A(_0275_),
    .B(_0412_));
 sg13g2_xnor2_1 _2363_ (.Y(\modem.instance2.instance5._09_[5] ),
    .A(\modem.instance2.instance5._10_[5] ),
    .B(_0452_));
 sg13g2_nand3_1 _2364_ (.B(\modem.instance2.instance5._10_[5] ),
    .C(_0412_),
    .A(_0275_),
    .Y(_0453_));
 sg13g2_xnor2_1 _2365_ (.Y(\modem.instance2.instance5._09_[6] ),
    .A(\modem.instance2.instance5._10_[6] ),
    .B(_0453_));
 sg13g2_nand4_1 _2366_ (.B(\modem.instance2.instance5._10_[5] ),
    .C(\modem.instance2.instance5._10_[6] ),
    .A(_0275_),
    .Y(_0454_),
    .D(_0412_));
 sg13g2_xnor2_1 _2367_ (.Y(\modem.instance2.instance5._09_[7] ),
    .A(\modem.instance2.instance5._10_[7] ),
    .B(_0454_));
 sg13g2_nand2_1 _2368_ (.Y(_0455_),
    .A(_0412_),
    .B(_0413_));
 sg13g2_xnor2_1 _2369_ (.Y(\modem.instance2.instance5._09_[8] ),
    .A(\modem.instance2.instance5._10_[8] ),
    .B(_0455_));
 sg13g2_xnor2_1 _2370_ (.Y(\modem.instance2.instance5._09_[9] ),
    .A(\modem.instance2.instance5._10_[9] ),
    .B(_0415_));
 sg13g2_nand2_1 _2371_ (.Y(_0456_),
    .A(\modem.instance3.instance1._6_[0] ),
    .B(_0282_));
 sg13g2_nand2_1 _2372_ (.Y(_0457_),
    .A(_0280_),
    .B(\modem.instance3.instance1._3_[0] ));
 sg13g2_o21ai_1 _2373_ (.B1(_0457_),
    .Y(\modem.instance3.instance1._3_[1] ),
    .A1(net59),
    .A2(_0456_));
 sg13g2_nand2_1 _2374_ (.Y(_0458_),
    .A(net59),
    .B(\modem.instance3.instance1._6_[0] ));
 sg13g2_xnor2_1 _2375_ (.Y(\modem.instance3.instance1._3_[2] ),
    .A(\modem.instance3.instance1._6_[2] ),
    .B(_0458_));
 sg13g2_nand2_1 _2376_ (.Y(_0459_),
    .A(\modem.instance3.instance1._6_[3] ),
    .B(_0282_));
 sg13g2_and2_1 _2377_ (.A(\modem.instance3.instance1._6_[0] ),
    .B(\modem.instance3.instance1._6_[2] ),
    .X(_0460_));
 sg13g2_xor2_1 _2378_ (.B(_0460_),
    .A(\modem.instance3.instance1._6_[3] ),
    .X(_0461_));
 sg13g2_nand2_1 _2379_ (.Y(_0462_),
    .A(net59),
    .B(_0461_));
 sg13g2_o21ai_1 _2380_ (.B1(_0462_),
    .Y(\modem.instance3.instance1._3_[3] ),
    .A1(net59),
    .A2(_0459_));
 sg13g2_nand2_1 _2381_ (.Y(_0463_),
    .A(\modem.instance3.instance1._6_[4] ),
    .B(_0282_));
 sg13g2_nand2_1 _2382_ (.Y(_0464_),
    .A(\modem.instance3.instance1._6_[3] ),
    .B(_0460_));
 sg13g2_xnor2_1 _2383_ (.Y(_0465_),
    .A(\modem.instance3.instance1._6_[4] ),
    .B(_0464_));
 sg13g2_nand2_1 _2384_ (.Y(_0466_),
    .A(net59),
    .B(_0465_));
 sg13g2_o21ai_1 _2385_ (.B1(_0466_),
    .Y(\modem.instance3.instance1._3_[4] ),
    .A1(net59),
    .A2(_0463_));
 sg13g2_nand4_1 _2386_ (.B(\modem.instance3.instance1._6_[3] ),
    .C(\modem.instance3.instance1._6_[4] ),
    .A(net59),
    .Y(_0467_),
    .D(_0460_));
 sg13g2_xnor2_1 _2387_ (.Y(\modem.instance3.instance1._3_[5] ),
    .A(\modem.instance3.instance1._6_[5] ),
    .B(_0467_));
 sg13g2_inv_1 _2388_ (.Y(_0468_),
    .A(\modem.instance3.instance1._6_[5] ));
 sg13g2_or2_1 _2389_ (.X(_0469_),
    .B(_0467_),
    .A(_0468_));
 sg13g2_xnor2_1 _2390_ (.Y(\modem.instance3.instance1._3_[6] ),
    .A(\modem.instance3.instance1._6_[6] ),
    .B(_0469_));
 sg13g2_nand4_1 _2391_ (.B(_0297_),
    .C(\modem.instance3.instance2._10_[3] ),
    .A(_0296_),
    .Y(_0470_),
    .D(\modem.instance3.instance2._10_[2] ));
 sg13g2_nand4_1 _2392_ (.B(_0294_),
    .C(\modem.instance3.instance2._10_[7] ),
    .A(\modem.instance3.instance2._10_[5] ),
    .Y(_0471_),
    .D(\modem.instance3.instance2._10_[6] ));
 sg13g2_nor2_2 _2393_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nand3_1 _2394_ (.B(_0292_),
    .C(_0472_),
    .A(\modem.instance3.instance2._10_[9] ),
    .Y(_0473_));
 sg13g2_xnor2_1 _2395_ (.Y(\modem.instance3.instance2._09_[10] ),
    .A(\modem.instance3.instance2._10_[10] ),
    .B(_0473_));
 sg13g2_nand4_1 _2396_ (.B(_0292_),
    .C(\modem.instance3.instance2._10_[10] ),
    .A(\modem.instance3.instance2._10_[9] ),
    .Y(_0474_),
    .D(_0472_));
 sg13g2_xnor2_1 _2397_ (.Y(\modem.instance3.instance2._09_[11] ),
    .A(\modem.instance3.instance2._10_[11] ),
    .B(_0474_));
 sg13g2_nand2_1 _2398_ (.Y(_0475_),
    .A(\modem.instance3.instance2._10_[11] ),
    .B(\modem.instance3.instance2._10_[10] ));
 sg13g2_nor2_1 _2399_ (.A(_0473_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_xor2_1 _2400_ (.B(_0476_),
    .A(\modem.instance3.instance2._10_[12] ),
    .X(\modem.instance3.instance2._09_[12] ));
 sg13g2_inv_1 _2401_ (.Y(_0477_),
    .A(\modem.instance3.instance2._10_[9] ));
 sg13g2_nand4_1 _2402_ (.B(\modem.instance3.instance2._10_[11] ),
    .C(\modem.instance3.instance2._10_[10] ),
    .A(_0292_),
    .Y(_0478_),
    .D(\modem.instance3.instance2._10_[12] ));
 sg13g2_nor4_2 _2403_ (.A(_0477_),
    .B(_0470_),
    .C(_0471_),
    .Y(_0479_),
    .D(_0478_));
 sg13g2_xor2_1 _2404_ (.B(_0479_),
    .A(\modem.instance3.instance2._10_[13] ),
    .X(\modem.instance3.instance2._09_[13] ));
 sg13g2_nand2_1 _2405_ (.Y(_0480_),
    .A(\modem.instance3.instance2._10_[13] ),
    .B(_0479_));
 sg13g2_xnor2_1 _2406_ (.Y(\modem.instance3.instance2._09_[14] ),
    .A(\modem.instance3.instance2._10_[14] ),
    .B(_0480_));
 sg13g2_nand3_1 _2407_ (.B(\modem.instance3.instance2._10_[14] ),
    .C(_0479_),
    .A(\modem.instance3.instance2._10_[13] ),
    .Y(_0481_));
 sg13g2_xnor2_1 _2408_ (.Y(\modem.instance3.instance2._09_[15] ),
    .A(\modem.instance3.instance2._10_[15] ),
    .B(_0481_));
 sg13g2_and3_1 _2409_ (.X(_0482_),
    .A(\modem.instance3.instance2._10_[13] ),
    .B(\modem.instance3.instance2._10_[15] ),
    .C(\modem.instance3.instance2._10_[14] ));
 sg13g2_buf_1 _2410_ (.A(_0482_),
    .X(_0483_));
 sg13g2_nand2_1 _2411_ (.Y(_0484_),
    .A(_0479_),
    .B(_0483_));
 sg13g2_xnor2_1 _2412_ (.Y(\modem.instance3.instance2._09_[16] ),
    .A(_0286_),
    .B(_0484_));
 sg13g2_nand3_1 _2413_ (.B(_0479_),
    .C(_0483_),
    .A(_0286_),
    .Y(_0485_));
 sg13g2_buf_1 _2414_ (.A(_0485_),
    .X(_0486_));
 sg13g2_xnor2_1 _2415_ (.Y(\modem.instance3.instance2._09_[17] ),
    .A(\modem.instance3.instance2._10_[17] ),
    .B(_0486_));
 sg13g2_nand4_1 _2416_ (.B(_0286_),
    .C(_0479_),
    .A(\modem.instance3.instance2._10_[17] ),
    .Y(_0487_),
    .D(_0483_));
 sg13g2_xnor2_1 _2417_ (.Y(\modem.instance3.instance2._09_[18] ),
    .A(\modem.instance3.instance2._10_[18] ),
    .B(_0487_));
 sg13g2_inv_1 _2418_ (.Y(_0488_),
    .A(\modem.instance3.instance2._10_[19] ));
 sg13g2_nand2_1 _2419_ (.Y(_0489_),
    .A(\modem.instance3.instance2._10_[17] ),
    .B(\modem.instance3.instance2._10_[18] ));
 sg13g2_nor2_1 _2420_ (.A(_0486_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_xnor2_1 _2421_ (.Y(\modem.instance3.instance2._09_[19] ),
    .A(_0488_),
    .B(_0490_));
 sg13g2_xnor2_1 _2422_ (.Y(_0491_),
    .A(_0296_),
    .B(_0297_));
 sg13g2_nor2_1 _2423_ (.A(_0300_),
    .B(_0491_),
    .Y(\modem.instance3.instance2._09_[1] ));
 sg13g2_nor3_1 _2424_ (.A(_0488_),
    .B(_0486_),
    .C(_0489_),
    .Y(_0492_));
 sg13g2_xor2_1 _2425_ (.B(_0492_),
    .A(\modem.instance3.instance2._10_[20] ),
    .X(\modem.instance3.instance2._09_[20] ));
 sg13g2_inv_1 _2426_ (.Y(_0493_),
    .A(\modem.instance3.instance2._10_[21] ));
 sg13g2_nand4_1 _2427_ (.B(\modem.instance3.instance2._10_[19] ),
    .C(\modem.instance3.instance2._10_[18] ),
    .A(\modem.instance3.instance2._10_[17] ),
    .Y(_0494_),
    .D(\modem.instance3.instance2._10_[20] ));
 sg13g2_nor2_1 _2428_ (.A(_0486_),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_xnor2_1 _2429_ (.Y(\modem.instance3.instance2._09_[21] ),
    .A(_0493_),
    .B(_0495_));
 sg13g2_nor3_1 _2430_ (.A(_0493_),
    .B(_0486_),
    .C(_0494_),
    .Y(_0496_));
 sg13g2_xor2_1 _2431_ (.B(_0496_),
    .A(\modem.instance3.instance2._10_[22] ),
    .X(\modem.instance3.instance2._09_[22] ));
 sg13g2_nand2_1 _2432_ (.Y(_0497_),
    .A(\modem.instance3.instance2._10_[21] ),
    .B(\modem.instance3.instance2._10_[22] ));
 sg13g2_nor2_1 _2433_ (.A(_0494_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_and4_1 _2434_ (.A(_0286_),
    .B(_0479_),
    .C(_0483_),
    .D(_0498_),
    .X(_0499_));
 sg13g2_xor2_1 _2435_ (.B(_0499_),
    .A(\modem.instance3.instance2._10_[23] ),
    .X(\modem.instance3.instance2._09_[23] ));
 sg13g2_nand2_1 _2436_ (.Y(_0500_),
    .A(\modem.instance3.instance2._10_[23] ),
    .B(_0499_));
 sg13g2_xnor2_1 _2437_ (.Y(\modem.instance3.instance2._09_[24] ),
    .A(\modem.instance3.instance2._10_[24] ),
    .B(_0500_));
 sg13g2_nand3_1 _2438_ (.B(\modem.instance3.instance2._10_[24] ),
    .C(_0499_),
    .A(\modem.instance3.instance2._10_[23] ),
    .Y(_0501_));
 sg13g2_xnor2_1 _2439_ (.Y(\modem.instance3.instance2._09_[25] ),
    .A(\modem.instance3.instance2._10_[25] ),
    .B(_0501_));
 sg13g2_nand4_1 _2440_ (.B(\modem.instance3.instance2._10_[23] ),
    .C(\modem.instance3.instance2._10_[25] ),
    .A(_0286_),
    .Y(_0502_),
    .D(\modem.instance3.instance2._10_[24] ));
 sg13g2_nor3_1 _2441_ (.A(_0494_),
    .B(_0497_),
    .C(_0502_),
    .Y(_0503_));
 sg13g2_nand3_1 _2442_ (.B(_0483_),
    .C(_0503_),
    .A(_0479_),
    .Y(_0504_));
 sg13g2_buf_2 _2443_ (.A(_0504_),
    .X(_0505_));
 sg13g2_xnor2_1 _2444_ (.Y(\modem.instance3.instance2._09_[26] ),
    .A(\modem.instance3.instance2._10_[26] ),
    .B(_0505_));
 sg13g2_inv_1 _2445_ (.Y(_0506_),
    .A(\modem.instance3.instance2._10_[26] ));
 sg13g2_nor2_1 _2446_ (.A(_0506_),
    .B(_0505_),
    .Y(_0507_));
 sg13g2_xor2_1 _2447_ (.B(_0507_),
    .A(\modem.instance3.instance2._10_[27] ),
    .X(\modem.instance3.instance2._09_[27] ));
 sg13g2_inv_1 _2448_ (.Y(_0508_),
    .A(\modem.instance3.instance2._10_[28] ));
 sg13g2_nand2_1 _2449_ (.Y(_0509_),
    .A(\modem.instance3.instance2._10_[27] ),
    .B(\modem.instance3.instance2._10_[26] ));
 sg13g2_nor2_1 _2450_ (.A(_0505_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_xnor2_1 _2451_ (.Y(\modem.instance3.instance2._09_[28] ),
    .A(_0508_),
    .B(_0510_));
 sg13g2_nor3_1 _2452_ (.A(_0508_),
    .B(_0505_),
    .C(_0509_),
    .Y(_0511_));
 sg13g2_xor2_1 _2453_ (.B(_0511_),
    .A(\modem.instance3.instance2._10_[29] ),
    .X(\modem.instance3.instance2._09_[29] ));
 sg13g2_nand2_1 _2454_ (.Y(_0512_),
    .A(_0296_),
    .B(_0297_));
 sg13g2_xnor2_1 _2455_ (.Y(\modem.instance3.instance2._09_[2] ),
    .A(\modem.instance3.instance2._10_[2] ),
    .B(_0512_));
 sg13g2_inv_1 _2456_ (.Y(_0513_),
    .A(\modem.instance3.instance2._10_[30] ));
 sg13g2_nand4_1 _2457_ (.B(\modem.instance3.instance2._10_[26] ),
    .C(\modem.instance3.instance2._10_[29] ),
    .A(\modem.instance3.instance2._10_[27] ),
    .Y(_0514_),
    .D(\modem.instance3.instance2._10_[28] ));
 sg13g2_nor2_1 _2458_ (.A(_0505_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_xnor2_1 _2459_ (.Y(\modem.instance3.instance2._09_[30] ),
    .A(_0513_),
    .B(_0515_));
 sg13g2_nor3_1 _2460_ (.A(_0513_),
    .B(_0505_),
    .C(_0514_),
    .Y(_0516_));
 sg13g2_xor2_1 _2461_ (.B(_0516_),
    .A(\modem.instance3.instance2._10_[31] ),
    .X(\modem.instance3.instance2._09_[31] ));
 sg13g2_nand3_1 _2462_ (.B(_0297_),
    .C(\modem.instance3.instance2._10_[2] ),
    .A(_0296_),
    .Y(_0517_));
 sg13g2_xnor2_1 _2463_ (.Y(\modem.instance3.instance2._09_[3] ),
    .A(\modem.instance3.instance2._10_[3] ),
    .B(_0517_));
 sg13g2_xnor2_1 _2464_ (.Y(\modem.instance3.instance2._09_[4] ),
    .A(_0294_),
    .B(_0470_));
 sg13g2_and4_1 _2465_ (.A(_0296_),
    .B(_0297_),
    .C(\modem.instance3.instance2._10_[3] ),
    .D(\modem.instance3.instance2._10_[2] ),
    .X(_0518_));
 sg13g2_nand2_1 _2466_ (.Y(_0519_),
    .A(_0294_),
    .B(_0518_));
 sg13g2_xnor2_1 _2467_ (.Y(\modem.instance3.instance2._09_[5] ),
    .A(\modem.instance3.instance2._10_[5] ),
    .B(_0519_));
 sg13g2_nand3_1 _2468_ (.B(_0294_),
    .C(_0518_),
    .A(\modem.instance3.instance2._10_[5] ),
    .Y(_0520_));
 sg13g2_xnor2_1 _2469_ (.Y(\modem.instance3.instance2._09_[6] ),
    .A(\modem.instance3.instance2._10_[6] ),
    .B(_0520_));
 sg13g2_nand4_1 _2470_ (.B(_0294_),
    .C(\modem.instance3.instance2._10_[6] ),
    .A(\modem.instance3.instance2._10_[5] ),
    .Y(_0521_),
    .D(_0518_));
 sg13g2_xnor2_1 _2471_ (.Y(\modem.instance3.instance2._09_[7] ),
    .A(\modem.instance3.instance2._10_[7] ),
    .B(_0521_));
 sg13g2_xor2_1 _2472_ (.B(_0472_),
    .A(_0292_),
    .X(\modem.instance3.instance2._09_[8] ));
 sg13g2_nand2_1 _2473_ (.Y(_0522_),
    .A(_0292_),
    .B(_0472_));
 sg13g2_xnor2_1 _2474_ (.Y(\modem.instance3.instance2._09_[9] ),
    .A(\modem.instance3.instance2._10_[9] ),
    .B(_0522_));
 sg13g2_nor2_1 _2475_ (.A(\modem.instance3.instance3._3_[0] ),
    .B(net39),
    .Y(_0523_));
 sg13g2_nand3_1 _2476_ (.B(net42),
    .C(net41),
    .A(net43),
    .Y(_0524_));
 sg13g2_a21o_1 _2477_ (.A2(_0524_),
    .A1(_0523_),
    .B1(_1153_),
    .X(\modem.instance3.instance3._3_[1] ));
 sg13g2_a21o_1 _2478_ (.A2(net41),
    .A1(net42),
    .B1(net39),
    .X(_0525_));
 sg13g2_nor2_1 _2479_ (.A(\modem.instance3.instance3._3_[0] ),
    .B(_1162_),
    .Y(_0526_));
 sg13g2_a22oi_1 _2480_ (.Y(\modem.instance3.instance3._3_[2] ),
    .B1(_0525_),
    .B2(_0526_),
    .A2(_0089_),
    .A1(_1162_));
 sg13g2_nand2_1 _2481_ (.Y(_0527_),
    .A(net39),
    .B(_0526_));
 sg13g2_nand2_1 _2482_ (.Y(_0528_),
    .A(net40),
    .B(net43));
 sg13g2_o21ai_1 _2483_ (.B1(net42),
    .Y(_0529_),
    .A1(_1170_),
    .A2(_0528_));
 sg13g2_o21ai_1 _2484_ (.B1(_0529_),
    .Y(\modem.instance3.instance3._3_[3] ),
    .A1(net42),
    .A2(_0527_));
 sg13g2_nand2_1 _2485_ (.Y(_0530_),
    .A(net42),
    .B(_0526_));
 sg13g2_nand2_1 _2486_ (.Y(_0531_),
    .A(net39),
    .B(_1159_));
 sg13g2_nand2_1 _2487_ (.Y(_0532_),
    .A(net41),
    .B(_0530_));
 sg13g2_o21ai_1 _2488_ (.B1(_0532_),
    .Y(\modem.instance3.instance3._3_[4] ),
    .A1(_0530_),
    .A2(_0531_));
 sg13g2_nor3_1 _2489_ (.A(_1064_),
    .B(_1076_),
    .C(_1072_),
    .Y(_0533_));
 sg13g2_a21oi_1 _2490_ (.A1(net44),
    .A2(_0533_),
    .Y(\modem.instance3.instance4._3_[0] ),
    .B1(net46));
 sg13g2_nand2_1 _2491_ (.Y(_0534_),
    .A(_1083_),
    .B(_1068_));
 sg13g2_o21ai_1 _2492_ (.B1(_1060_),
    .Y(\modem.instance3.instance4._3_[1] ),
    .A1(_0533_),
    .A2(_0534_));
 sg13g2_xor2_1 _2493_ (.B(_0057_),
    .A(net46),
    .X(_0535_));
 sg13g2_or3_1 _2494_ (.A(net45),
    .B(_0057_),
    .C(_0533_),
    .X(_0536_));
 sg13g2_o21ai_1 _2495_ (.B1(_0536_),
    .Y(\modem.instance3.instance4._3_[2] ),
    .A1(net44),
    .A2(_0535_));
 sg13g2_nor2_1 _2496_ (.A(_1079_),
    .B(_1076_),
    .Y(_0537_));
 sg13g2_o21ai_1 _2497_ (.B1(_0537_),
    .Y(_0538_),
    .A1(net45),
    .A2(net48));
 sg13g2_nor3_1 _2498_ (.A(net20),
    .B(_1076_),
    .C(_1098_),
    .Y(_0539_));
 sg13g2_a21o_1 _2499_ (.A2(_0538_),
    .A1(net20),
    .B1(_0539_),
    .X(\modem.instance3.instance4._3_[3] ));
 sg13g2_a21oi_1 _2500_ (.A1(net44),
    .A2(_1076_),
    .Y(_0540_),
    .B1(_1072_));
 sg13g2_o21ai_1 _2501_ (.B1(net45),
    .Y(_0541_),
    .A1(_1067_),
    .A2(_1116_));
 sg13g2_o21ai_1 _2502_ (.B1(_0541_),
    .Y(\modem.instance3.instance4._3_[4] ),
    .A1(_1064_),
    .A2(_0540_));
 sg13g2_nor2b_1 _2503_ (.A(net29),
    .B_N(\modem.instance2._3_[0] ),
    .Y(_0542_));
 sg13g2_a21oi_1 _2504_ (.A1(\modem.instance2._2_[0] ),
    .A2(net29),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_buf_2 _2505_ (.A(ui_in[0]),
    .X(_0544_));
 sg13g2_buf_2 _2506_ (.A(ui_in[1]),
    .X(_0545_));
 sg13g2_nand2b_1 _2507_ (.Y(_0546_),
    .B(_0545_),
    .A_N(_0544_));
 sg13g2_buf_2 _2508_ (.A(_0546_),
    .X(_0547_));
 sg13g2_mux2_1 _2509_ (.A0(\modem.instance3._3_[0] ),
    .A1(\modem.instance3._2_[0] ),
    .S(_0284_),
    .X(_0548_));
 sg13g2_mux2_1 _2510_ (.A0(\modem._0_[0] ),
    .A1(_0548_),
    .S(_0545_),
    .X(_0549_));
 sg13g2_nand2_1 _2511_ (.Y(_0550_),
    .A(_0544_),
    .B(_0549_));
 sg13g2_o21ai_1 _2512_ (.B1(_0550_),
    .Y(\modem.instance4._5_[0] ),
    .A1(_0543_),
    .A2(_0547_));
 sg13g2_nor2b_1 _2513_ (.A(net29),
    .B_N(\modem.instance2._3_[1] ),
    .Y(_0551_));
 sg13g2_a21oi_1 _2514_ (.A1(net29),
    .A2(\modem.instance2._2_[1] ),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_mux2_1 _2515_ (.A0(\modem.instance3._3_[1] ),
    .A1(\modem.instance3._2_[1] ),
    .S(_0284_),
    .X(_0553_));
 sg13g2_mux2_1 _2516_ (.A0(\modem._0_[1] ),
    .A1(_0553_),
    .S(_0545_),
    .X(_0554_));
 sg13g2_nand2_1 _2517_ (.Y(_0555_),
    .A(_0544_),
    .B(_0554_));
 sg13g2_o21ai_1 _2518_ (.B1(_0555_),
    .Y(\modem.instance4._5_[1] ),
    .A1(_0547_),
    .A2(_0552_));
 sg13g2_nor2b_1 _2519_ (.A(net29),
    .B_N(\modem.instance2._3_[2] ),
    .Y(_0556_));
 sg13g2_a21oi_1 _2520_ (.A1(_0263_),
    .A2(\modem.instance2._2_[2] ),
    .Y(_0557_),
    .B1(_0556_));
 sg13g2_mux2_1 _2521_ (.A0(\modem.instance3._3_[2] ),
    .A1(\modem.instance3._2_[2] ),
    .S(_0284_),
    .X(_0558_));
 sg13g2_mux2_1 _2522_ (.A0(\modem._0_[2] ),
    .A1(_0558_),
    .S(_0545_),
    .X(_0559_));
 sg13g2_nand2_1 _2523_ (.Y(_0560_),
    .A(_0544_),
    .B(_0559_));
 sg13g2_o21ai_1 _2524_ (.B1(_0560_),
    .Y(\modem.instance4._5_[2] ),
    .A1(_0547_),
    .A2(_0557_));
 sg13g2_nor2b_1 _2525_ (.A(\modem.instance2._4_ ),
    .B_N(\modem.instance2._3_[3] ),
    .Y(_0561_));
 sg13g2_a21oi_1 _2526_ (.A1(net29),
    .A2(\modem.instance2._2_[3] ),
    .Y(_0562_),
    .B1(_0561_));
 sg13g2_mux2_1 _2527_ (.A0(\modem.instance3._3_[3] ),
    .A1(\modem.instance3._2_[3] ),
    .S(_0284_),
    .X(_0563_));
 sg13g2_mux2_1 _2528_ (.A0(\modem._0_[3] ),
    .A1(_0563_),
    .S(_0545_),
    .X(_0564_));
 sg13g2_nand2_1 _2529_ (.Y(_0565_),
    .A(_0544_),
    .B(_0564_));
 sg13g2_o21ai_1 _2530_ (.B1(_0565_),
    .Y(\modem.instance4._5_[3] ),
    .A1(_0547_),
    .A2(_0562_));
 sg13g2_nor2b_1 _2531_ (.A(\modem.instance2._4_ ),
    .B_N(\modem.instance2._3_[4] ),
    .Y(_0566_));
 sg13g2_a21oi_1 _2532_ (.A1(net29),
    .A2(\modem.instance2._2_[4] ),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_mux2_1 _2533_ (.A0(\modem.instance3._3_[4] ),
    .A1(\modem.instance3._2_[4] ),
    .S(_0284_),
    .X(_0568_));
 sg13g2_mux2_1 _2534_ (.A0(\modem._0_[4] ),
    .A1(_0568_),
    .S(_0545_),
    .X(_0569_));
 sg13g2_nand2_1 _2535_ (.Y(_0570_),
    .A(_0544_),
    .B(_0569_));
 sg13g2_o21ai_1 _2536_ (.B1(_0570_),
    .Y(\modem.instance4._5_[4] ),
    .A1(_0547_),
    .A2(_0567_));
 sg13g2_nor2b_1 _2537_ (.A(\modem.instance2._4_ ),
    .B_N(\modem.instance2._3_[5] ),
    .Y(_0571_));
 sg13g2_a21oi_1 _2538_ (.A1(net29),
    .A2(\modem.instance2._2_[5] ),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_mux2_1 _2539_ (.A0(\modem.instance3._3_[5] ),
    .A1(\modem.instance3._2_[5] ),
    .S(_0284_),
    .X(_0573_));
 sg13g2_mux2_1 _2540_ (.A0(\modem._0_[5] ),
    .A1(_0573_),
    .S(_0545_),
    .X(_0574_));
 sg13g2_nand2_1 _2541_ (.Y(_0575_),
    .A(_0544_),
    .B(_0574_));
 sg13g2_o21ai_1 _2542_ (.B1(_0575_),
    .Y(\modem.instance4._5_[5] ),
    .A1(_0547_),
    .A2(_0572_));
 sg13g2_nor2b_1 _2543_ (.A(\modem._0_[0] ),
    .B_N(\modem._0_[1] ),
    .Y(_0576_));
 sg13g2_nor2b_1 _2544_ (.A(\modem._0_[5] ),
    .B_N(\modem._0_[4] ),
    .Y(_0577_));
 sg13g2_nand4_1 _2545_ (.B(\modem._0_[2] ),
    .C(_0576_),
    .A(\modem._0_[3] ),
    .Y(\modem.instance6._1_ ),
    .D(_0577_));
 sg13g2_nor2_1 _2546_ (.A(\modem.instance7.instance2._3_[0] ),
    .B(net50),
    .Y(_0578_));
 sg13g2_o21ai_1 _2547_ (.B1(_0578_),
    .Y(_0579_),
    .A1(_0046_),
    .A2(_1040_));
 sg13g2_nand2b_1 _2548_ (.Y(\modem.instance7.instance2._3_[1] ),
    .B(_0579_),
    .A_N(_0996_));
 sg13g2_inv_1 _2549_ (.Y(_0580_),
    .A(_0046_));
 sg13g2_a21o_1 _2550_ (.A2(_0580_),
    .A1(net52),
    .B1(net50),
    .X(_0581_));
 sg13g2_nor2_1 _2551_ (.A(\modem.instance7.instance2._3_[0] ),
    .B(_1005_),
    .Y(_0582_));
 sg13g2_a22oi_1 _2552_ (.Y(\modem.instance7.instance2._3_[2] ),
    .B1(_0581_),
    .B2(_0582_),
    .A2(_1036_),
    .A1(_1005_));
 sg13g2_nand2_1 _2553_ (.Y(_0583_),
    .A(net50),
    .B(_0582_));
 sg13g2_nand2_1 _2554_ (.Y(_0584_),
    .A(_0985_),
    .B(_0974_));
 sg13g2_nor2_1 _2555_ (.A(net50),
    .B(_0580_),
    .Y(_0585_));
 sg13g2_o21ai_1 _2556_ (.B1(net52),
    .Y(_0586_),
    .A1(_0584_),
    .A2(_0585_));
 sg13g2_o21ai_1 _2557_ (.B1(_0586_),
    .Y(\modem.instance7.instance2._3_[3] ),
    .A1(net52),
    .A2(_0583_));
 sg13g2_nor2_1 _2558_ (.A(_0997_),
    .B(_0584_),
    .Y(_0587_));
 sg13g2_nand3_1 _2559_ (.B(_0046_),
    .C(_0587_),
    .A(net50),
    .Y(_0588_));
 sg13g2_o21ai_1 _2560_ (.B1(_0588_),
    .Y(\modem.instance7.instance2._3_[4] ),
    .A1(_0046_),
    .A2(_0587_));
 sg13g2_xor2_1 _2561_ (.B(_0543_),
    .A(\modem.instance7._0_[0] ),
    .X(\modem.instance7.instance3._0_[0] ));
 sg13g2_xor2_1 _2562_ (.B(_0552_),
    .A(\modem.instance7._0_[1] ),
    .X(\modem.instance7.instance3._0_[1] ));
 sg13g2_xor2_1 _2563_ (.B(_0557_),
    .A(\modem.instance7._0_[2] ),
    .X(\modem.instance7.instance3._0_[2] ));
 sg13g2_xor2_1 _2564_ (.B(_0562_),
    .A(\modem.instance7._0_[3] ),
    .X(\modem.instance7.instance3._0_[3] ));
 sg13g2_xor2_1 _2565_ (.B(_0567_),
    .A(\modem.instance7._0_[4] ),
    .X(\modem.instance7.instance3._0_[4] ));
 sg13g2_xor2_1 _2566_ (.B(_0572_),
    .A(\modem.instance7._0_[5] ),
    .X(\modem.instance7.instance3._0_[5] ));
 sg13g2_buf_1 _2567_ (.A(\modem.instance7.instance4._9_[23] ),
    .X(_0589_));
 sg13g2_nor4_1 _2568_ (.A(\modem.instance7.instance4._9_[16] ),
    .B(_0589_),
    .C(\modem.instance7.instance4._9_[22] ),
    .D(\modem.instance7.instance4._9_[24] ),
    .Y(_0590_));
 sg13g2_nor4_1 _2569_ (.A(\modem.instance7.instance4._9_[19] ),
    .B(\modem.instance7.instance4._9_[18] ),
    .C(\modem.instance7.instance4._9_[21] ),
    .D(\modem.instance7.instance4._9_[20] ),
    .Y(_0591_));
 sg13g2_nor4_1 _2570_ (.A(\modem.instance7.instance4._9_[3] ),
    .B(\modem.instance7.instance4._9_[25] ),
    .C(\modem.instance7.instance4._9_[31] ),
    .D(\modem.instance7.instance4._9_[30] ),
    .Y(_0592_));
 sg13g2_nor4_1 _2571_ (.A(\modem.instance7.instance4._9_[27] ),
    .B(\modem.instance7.instance4._9_[26] ),
    .C(\modem.instance7.instance4._9_[29] ),
    .D(\modem.instance7.instance4._9_[28] ),
    .Y(_0593_));
 sg13g2_nand4_1 _2572_ (.B(_0591_),
    .C(_0592_),
    .A(_0590_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_buf_1 _2573_ (.A(\modem.instance7.instance4._9_[15] ),
    .X(_0595_));
 sg13g2_nor2_1 _2574_ (.A(_0595_),
    .B(\modem.instance7.instance4._9_[14] ),
    .Y(_0596_));
 sg13g2_nor4_1 _2575_ (.A(\modem.instance7.instance4._9_[8] ),
    .B(\modem.instance7.instance4._9_[10] ),
    .C(\modem.instance7.instance4._9_[13] ),
    .D(\modem.instance7.instance4._9_[12] ),
    .Y(_0597_));
 sg13g2_nor4_1 _2576_ (.A(\modem.instance7.instance4._9_[6] ),
    .B(\modem.instance7.instance4._9_[9] ),
    .C(\modem.instance7.instance4._9_[11] ),
    .D(\modem.instance7.instance4._9_[17] ),
    .Y(_0598_));
 sg13g2_buf_2 _2577_ (.A(\modem.instance7.instance4._9_[2] ),
    .X(_0599_));
 sg13g2_nor4_1 _2578_ (.A(_0599_),
    .B(\modem.instance7.instance4._9_[5] ),
    .C(\modem.instance7.instance4._9_[4] ),
    .D(\modem.instance7.instance4._9_[7] ),
    .Y(_0600_));
 sg13g2_nand4_1 _2579_ (.B(_0597_),
    .C(_0598_),
    .A(_0596_),
    .Y(_0601_),
    .D(_0600_));
 sg13g2_nor2_1 _2580_ (.A(_0594_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_buf_1 _2581_ (.A(\modem.instance7.instance4._9_[0] ),
    .X(_0603_));
 sg13g2_buf_2 _2582_ (.A(\modem.instance7.instance4._9_[1] ),
    .X(_0604_));
 sg13g2_nand2_1 _2583_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_a21oi_1 _2584_ (.A1(_0602_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(_0049_));
 sg13g2_nor2b_1 _2585_ (.A(_0604_),
    .B_N(_0049_),
    .Y(_0607_));
 sg13g2_inv_1 _2586_ (.Y(_0608_),
    .A(_0043_));
 sg13g2_and4_1 _2587_ (.A(\modem.instance7._1_[2] ),
    .B(\modem.instance7._1_[3] ),
    .C(\modem.instance7._1_[4] ),
    .D(\modem.instance7._1_[5] ),
    .X(_0609_));
 sg13g2_nand4_1 _2588_ (.B(\modem.instance7._1_[0] ),
    .C(\modem.instance7._1_[1] ),
    .A(_0608_),
    .Y(_0610_),
    .D(_0609_));
 sg13g2_buf_1 _2589_ (.A(_0610_),
    .X(_0611_));
 sg13g2_a21oi_1 _2590_ (.A1(_0602_),
    .A2(_0607_),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_nor2b_1 _2591_ (.A(_0606_),
    .B_N(_0612_),
    .Y(\modem.instance7.instance4._7_ ));
 sg13g2_buf_1 _2592_ (.A(_0611_),
    .X(_0613_));
 sg13g2_nor2_1 _2593_ (.A(_0603_),
    .B(_0613_),
    .Y(\modem.instance7.instance4._8_[0] ));
 sg13g2_nand2_2 _2594_ (.Y(_0614_),
    .A(\modem.instance7.instance4._9_[5] ),
    .B(\modem.instance7.instance4._9_[4] ));
 sg13g2_nand4_1 _2595_ (.B(_0604_),
    .C(\modem.instance7.instance4._9_[3] ),
    .A(_0603_),
    .Y(_0615_),
    .D(_0599_));
 sg13g2_buf_2 _2596_ (.A(_0615_),
    .X(_0616_));
 sg13g2_nand3_1 _2597_ (.B(\modem.instance7.instance4._9_[6] ),
    .C(\modem.instance7.instance4._9_[8] ),
    .A(\modem.instance7.instance4._9_[7] ),
    .Y(_0617_));
 sg13g2_nor3_2 _2598_ (.A(_0614_),
    .B(_0616_),
    .C(_0617_),
    .Y(_0618_));
 sg13g2_nand2_1 _2599_ (.Y(_0619_),
    .A(\modem.instance7.instance4._9_[9] ),
    .B(_0618_));
 sg13g2_xor2_1 _2600_ (.B(_0619_),
    .A(\modem.instance7.instance4._9_[10] ),
    .X(_0620_));
 sg13g2_nor2_1 _2601_ (.A(net18),
    .B(_0620_),
    .Y(\modem.instance7.instance4._8_[10] ));
 sg13g2_nand2_1 _2602_ (.Y(_0621_),
    .A(\modem.instance7.instance4._9_[9] ),
    .B(\modem.instance7.instance4._9_[10] ));
 sg13g2_nor4_2 _2603_ (.A(_0614_),
    .B(_0616_),
    .C(_0617_),
    .Y(_0622_),
    .D(_0621_));
 sg13g2_xnor2_1 _2604_ (.Y(_0623_),
    .A(\modem.instance7.instance4._9_[11] ),
    .B(_0622_));
 sg13g2_nor2_1 _2605_ (.A(net18),
    .B(_0623_),
    .Y(\modem.instance7.instance4._8_[11] ));
 sg13g2_nand2_1 _2606_ (.Y(_0624_),
    .A(\modem.instance7.instance4._9_[11] ),
    .B(_0622_));
 sg13g2_xor2_1 _2607_ (.B(_0624_),
    .A(\modem.instance7.instance4._9_[12] ),
    .X(_0625_));
 sg13g2_nor2_1 _2608_ (.A(net18),
    .B(_0625_),
    .Y(\modem.instance7.instance4._8_[12] ));
 sg13g2_nand3_1 _2609_ (.B(\modem.instance7.instance4._9_[12] ),
    .C(_0622_),
    .A(\modem.instance7.instance4._9_[11] ),
    .Y(_0626_));
 sg13g2_xor2_1 _2610_ (.B(_0626_),
    .A(\modem.instance7.instance4._9_[13] ),
    .X(_0627_));
 sg13g2_nor2_1 _2611_ (.A(net18),
    .B(_0627_),
    .Y(\modem.instance7.instance4._8_[13] ));
 sg13g2_nand3_1 _2612_ (.B(\modem.instance7.instance4._9_[13] ),
    .C(\modem.instance7.instance4._9_[12] ),
    .A(\modem.instance7.instance4._9_[11] ),
    .Y(_0628_));
 sg13g2_nor2_1 _2613_ (.A(_0621_),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_nand2_1 _2614_ (.Y(_0630_),
    .A(_0618_),
    .B(_0629_));
 sg13g2_xor2_1 _2615_ (.B(_0630_),
    .A(\modem.instance7.instance4._9_[14] ),
    .X(_0631_));
 sg13g2_nor2_1 _2616_ (.A(net18),
    .B(_0631_),
    .Y(\modem.instance7.instance4._8_[14] ));
 sg13g2_and4_1 _2617_ (.A(_0603_),
    .B(_0604_),
    .C(\modem.instance7.instance4._9_[3] ),
    .D(_0599_),
    .X(_0632_));
 sg13g2_buf_1 _2618_ (.A(_0632_),
    .X(_0633_));
 sg13g2_buf_1 _2619_ (.A(_0633_),
    .X(_0634_));
 sg13g2_nand3_1 _2620_ (.B(\modem.instance7.instance4._9_[4] ),
    .C(\modem.instance7.instance4._9_[14] ),
    .A(\modem.instance7.instance4._9_[5] ),
    .Y(_0635_));
 sg13g2_nor4_2 _2621_ (.A(_0617_),
    .B(_0621_),
    .C(_0628_),
    .Y(_0636_),
    .D(_0635_));
 sg13g2_buf_1 _2622_ (.A(_0636_),
    .X(_0637_));
 sg13g2_nand2_1 _2623_ (.Y(_0638_),
    .A(net17),
    .B(net19));
 sg13g2_xor2_1 _2624_ (.B(_0638_),
    .A(_0595_),
    .X(_0639_));
 sg13g2_nor2_1 _2625_ (.A(net18),
    .B(_0639_),
    .Y(\modem.instance7.instance4._8_[15] ));
 sg13g2_nand3_1 _2626_ (.B(net17),
    .C(net19),
    .A(_0595_),
    .Y(_0640_));
 sg13g2_xor2_1 _2627_ (.B(_0640_),
    .A(\modem.instance7.instance4._9_[16] ),
    .X(_0641_));
 sg13g2_nor2_1 _2628_ (.A(net18),
    .B(_0641_),
    .Y(\modem.instance7.instance4._8_[16] ));
 sg13g2_inv_1 _2629_ (.Y(_0642_),
    .A(_0048_));
 sg13g2_and4_1 _2630_ (.A(_0604_),
    .B(_0595_),
    .C(\modem.instance7.instance4._9_[16] ),
    .D(_0642_),
    .X(_0643_));
 sg13g2_nand4_1 _2631_ (.B(_0599_),
    .C(_0636_),
    .A(\modem.instance7.instance4._9_[3] ),
    .Y(_0644_),
    .D(_0643_));
 sg13g2_xor2_1 _2632_ (.B(_0644_),
    .A(\modem.instance7.instance4._9_[17] ),
    .X(_0645_));
 sg13g2_nor2_1 _2633_ (.A(_0613_),
    .B(_0645_),
    .Y(\modem.instance7.instance4._8_[17] ));
 sg13g2_and3_1 _2634_ (.X(_0646_),
    .A(_0595_),
    .B(\modem.instance7.instance4._9_[17] ),
    .C(\modem.instance7.instance4._9_[16] ));
 sg13g2_nand3_1 _2635_ (.B(net19),
    .C(_0646_),
    .A(net17),
    .Y(_0647_));
 sg13g2_xor2_1 _2636_ (.B(_0647_),
    .A(\modem.instance7.instance4._9_[18] ),
    .X(_0648_));
 sg13g2_nor2_1 _2637_ (.A(net18),
    .B(_0648_),
    .Y(\modem.instance7.instance4._8_[18] ));
 sg13g2_buf_1 _2638_ (.A(_0611_),
    .X(_0649_));
 sg13g2_nand4_1 _2639_ (.B(net17),
    .C(_0636_),
    .A(\modem.instance7.instance4._9_[18] ),
    .Y(_0650_),
    .D(_0646_));
 sg13g2_xor2_1 _2640_ (.B(_0650_),
    .A(\modem.instance7.instance4._9_[19] ),
    .X(_0651_));
 sg13g2_nor2_1 _2641_ (.A(net16),
    .B(_0651_),
    .Y(\modem.instance7.instance4._8_[19] ));
 sg13g2_xnor2_1 _2642_ (.Y(_0652_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_nor2_1 _2643_ (.A(net16),
    .B(_0652_),
    .Y(\modem.instance7.instance4._8_[1] ));
 sg13g2_and3_1 _2644_ (.X(_0653_),
    .A(\modem.instance7.instance4._9_[19] ),
    .B(\modem.instance7.instance4._9_[18] ),
    .C(_0646_));
 sg13g2_nand3_1 _2645_ (.B(_0636_),
    .C(_0653_),
    .A(_0633_),
    .Y(_0654_));
 sg13g2_xor2_1 _2646_ (.B(_0654_),
    .A(\modem.instance7.instance4._9_[20] ),
    .X(_0655_));
 sg13g2_nor2_1 _2647_ (.A(net16),
    .B(_0655_),
    .Y(\modem.instance7.instance4._8_[20] ));
 sg13g2_nand4_1 _2648_ (.B(_0633_),
    .C(_0636_),
    .A(\modem.instance7.instance4._9_[20] ),
    .Y(_0656_),
    .D(_0653_));
 sg13g2_xor2_1 _2649_ (.B(_0656_),
    .A(\modem.instance7.instance4._9_[21] ),
    .X(_0657_));
 sg13g2_nor2_1 _2650_ (.A(net16),
    .B(_0657_),
    .Y(\modem.instance7.instance4._8_[21] ));
 sg13g2_nand2_1 _2651_ (.Y(_0658_),
    .A(\modem.instance7.instance4._9_[21] ),
    .B(\modem.instance7.instance4._9_[20] ));
 sg13g2_o21ai_1 _2652_ (.B1(\modem.instance7.instance4._9_[22] ),
    .Y(_0659_),
    .A1(_0654_),
    .A2(_0658_));
 sg13g2_or3_1 _2653_ (.A(\modem.instance7.instance4._9_[22] ),
    .B(_0654_),
    .C(_0658_),
    .X(_0660_));
 sg13g2_a21oi_1 _2654_ (.A1(_0659_),
    .A2(_0660_),
    .Y(\modem.instance7.instance4._8_[22] ),
    .B1(_0611_));
 sg13g2_nand4_1 _2655_ (.B(\modem.instance7.instance4._9_[17] ),
    .C(\modem.instance7.instance4._9_[16] ),
    .A(_0595_),
    .Y(_0661_),
    .D(\modem.instance7.instance4._9_[22] ));
 sg13g2_nand4_1 _2656_ (.B(\modem.instance7.instance4._9_[18] ),
    .C(\modem.instance7.instance4._9_[21] ),
    .A(\modem.instance7.instance4._9_[19] ),
    .Y(_0662_),
    .D(\modem.instance7.instance4._9_[20] ));
 sg13g2_nor2_1 _2657_ (.A(_0661_),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_nand3_1 _2658_ (.B(net19),
    .C(_0663_),
    .A(_0634_),
    .Y(_0664_));
 sg13g2_xor2_1 _2659_ (.B(_0664_),
    .A(_0589_),
    .X(_0665_));
 sg13g2_nor2_1 _2660_ (.A(_0649_),
    .B(_0665_),
    .Y(\modem.instance7.instance4._8_[23] ));
 sg13g2_nand4_1 _2661_ (.B(_0633_),
    .C(_0636_),
    .A(_0589_),
    .Y(_0666_),
    .D(_0663_));
 sg13g2_xor2_1 _2662_ (.B(_0666_),
    .A(\modem.instance7.instance4._9_[24] ),
    .X(_0667_));
 sg13g2_nor2_1 _2663_ (.A(net16),
    .B(_0667_),
    .Y(\modem.instance7.instance4._8_[24] ));
 sg13g2_and2_1 _2664_ (.A(_0589_),
    .B(\modem.instance7.instance4._9_[24] ),
    .X(_0668_));
 sg13g2_nand4_1 _2665_ (.B(_0637_),
    .C(_0663_),
    .A(_0634_),
    .Y(_0669_),
    .D(_0668_));
 sg13g2_xor2_1 _2666_ (.B(_0669_),
    .A(\modem.instance7.instance4._9_[25] ),
    .X(_0670_));
 sg13g2_nor2_1 _2667_ (.A(_0649_),
    .B(_0670_),
    .Y(\modem.instance7.instance4._8_[25] ));
 sg13g2_nand3_1 _2668_ (.B(\modem.instance7.instance4._9_[25] ),
    .C(\modem.instance7.instance4._9_[24] ),
    .A(_0589_),
    .Y(_0671_));
 sg13g2_nor2_1 _2669_ (.A(_0616_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_nand3_1 _2670_ (.B(_0663_),
    .C(_0672_),
    .A(net19),
    .Y(_0673_));
 sg13g2_xor2_1 _2671_ (.B(_0673_),
    .A(\modem.instance7.instance4._9_[26] ),
    .X(_0674_));
 sg13g2_nor2_1 _2672_ (.A(net16),
    .B(_0674_),
    .Y(\modem.instance7.instance4._8_[26] ));
 sg13g2_nand4_1 _2673_ (.B(\modem.instance7.instance4._9_[25] ),
    .C(\modem.instance7.instance4._9_[24] ),
    .A(_0589_),
    .Y(_0675_),
    .D(\modem.instance7.instance4._9_[26] ));
 sg13g2_nor4_2 _2674_ (.A(_0616_),
    .B(_0661_),
    .C(_0662_),
    .Y(_0676_),
    .D(_0675_));
 sg13g2_nand2_1 _2675_ (.Y(_0677_),
    .A(_0637_),
    .B(_0676_));
 sg13g2_xor2_1 _2676_ (.B(_0677_),
    .A(\modem.instance7.instance4._9_[27] ),
    .X(_0678_));
 sg13g2_nor2_1 _2677_ (.A(net16),
    .B(_0678_),
    .Y(\modem.instance7.instance4._8_[27] ));
 sg13g2_nand3_1 _2678_ (.B(net19),
    .C(_0676_),
    .A(\modem.instance7.instance4._9_[27] ),
    .Y(_0679_));
 sg13g2_xor2_1 _2679_ (.B(_0679_),
    .A(\modem.instance7.instance4._9_[28] ),
    .X(_0680_));
 sg13g2_nor2_1 _2680_ (.A(net16),
    .B(_0680_),
    .Y(\modem.instance7.instance4._8_[28] ));
 sg13g2_buf_1 _2681_ (.A(_0611_),
    .X(_0681_));
 sg13g2_nand4_1 _2682_ (.B(\modem.instance7.instance4._9_[28] ),
    .C(_0636_),
    .A(\modem.instance7.instance4._9_[27] ),
    .Y(_0682_),
    .D(_0676_));
 sg13g2_xor2_1 _2683_ (.B(_0682_),
    .A(\modem.instance7.instance4._9_[29] ),
    .X(_0683_));
 sg13g2_nor2_1 _2684_ (.A(net15),
    .B(_0683_),
    .Y(\modem.instance7.instance4._8_[29] ));
 sg13g2_xor2_1 _2685_ (.B(_0605_),
    .A(_0599_),
    .X(_0684_));
 sg13g2_nor2_1 _2686_ (.A(net15),
    .B(_0684_),
    .Y(\modem.instance7.instance4._8_[2] ));
 sg13g2_nand4_1 _2687_ (.B(\modem.instance7.instance4._9_[26] ),
    .C(\modem.instance7.instance4._9_[29] ),
    .A(\modem.instance7.instance4._9_[27] ),
    .Y(_0685_),
    .D(\modem.instance7.instance4._9_[28] ));
 sg13g2_nor4_1 _2688_ (.A(_0661_),
    .B(_0662_),
    .C(_0671_),
    .D(_0685_),
    .Y(_0686_));
 sg13g2_nand3_1 _2689_ (.B(net19),
    .C(_0686_),
    .A(net17),
    .Y(_0687_));
 sg13g2_xor2_1 _2690_ (.B(_0687_),
    .A(\modem.instance7.instance4._9_[30] ),
    .X(_0688_));
 sg13g2_nor2_1 _2691_ (.A(net15),
    .B(_0688_),
    .Y(\modem.instance7.instance4._8_[30] ));
 sg13g2_nand4_1 _2692_ (.B(net17),
    .C(net19),
    .A(\modem.instance7.instance4._9_[30] ),
    .Y(_0689_),
    .D(_0686_));
 sg13g2_xnor2_1 _2693_ (.Y(_0690_),
    .A(_0049_),
    .B(_0689_));
 sg13g2_nor2_1 _2694_ (.A(_0681_),
    .B(_0690_),
    .Y(\modem.instance7.instance4._8_[31] ));
 sg13g2_nand3_1 _2695_ (.B(_0604_),
    .C(_0599_),
    .A(_0603_),
    .Y(_0691_));
 sg13g2_xor2_1 _2696_ (.B(_0691_),
    .A(\modem.instance7.instance4._9_[3] ),
    .X(_0692_));
 sg13g2_nor2_1 _2697_ (.A(_0681_),
    .B(_0692_),
    .Y(\modem.instance7.instance4._8_[3] ));
 sg13g2_xnor2_1 _2698_ (.Y(_0693_),
    .A(\modem.instance7.instance4._9_[4] ),
    .B(net17));
 sg13g2_nor2_1 _2699_ (.A(net15),
    .B(_0693_),
    .Y(\modem.instance7.instance4._8_[4] ));
 sg13g2_nand2_1 _2700_ (.Y(_0694_),
    .A(\modem.instance7.instance4._9_[4] ),
    .B(net17));
 sg13g2_xor2_1 _2701_ (.B(_0694_),
    .A(\modem.instance7.instance4._9_[5] ),
    .X(_0695_));
 sg13g2_nor2_1 _2702_ (.A(net15),
    .B(_0695_),
    .Y(\modem.instance7.instance4._8_[5] ));
 sg13g2_nor2_1 _2703_ (.A(_0614_),
    .B(_0616_),
    .Y(_0696_));
 sg13g2_xnor2_1 _2704_ (.Y(_0697_),
    .A(\modem.instance7.instance4._9_[6] ),
    .B(_0696_));
 sg13g2_nor2_1 _2705_ (.A(net15),
    .B(_0697_),
    .Y(\modem.instance7.instance4._8_[6] ));
 sg13g2_nand2_1 _2706_ (.Y(_0698_),
    .A(\modem.instance7.instance4._9_[6] ),
    .B(_0696_));
 sg13g2_xor2_1 _2707_ (.B(_0698_),
    .A(\modem.instance7.instance4._9_[7] ),
    .X(_0699_));
 sg13g2_nor2_1 _2708_ (.A(net15),
    .B(_0699_),
    .Y(\modem.instance7.instance4._8_[7] ));
 sg13g2_nand3_1 _2709_ (.B(\modem.instance7.instance4._9_[6] ),
    .C(_0696_),
    .A(\modem.instance7.instance4._9_[7] ),
    .Y(_0700_));
 sg13g2_xor2_1 _2710_ (.B(_0700_),
    .A(\modem.instance7.instance4._9_[8] ),
    .X(_0701_));
 sg13g2_nor2_1 _2711_ (.A(net15),
    .B(_0701_),
    .Y(\modem.instance7.instance4._8_[8] ));
 sg13g2_xnor2_1 _2712_ (.Y(_0702_),
    .A(\modem.instance7.instance4._9_[9] ),
    .B(_0618_));
 sg13g2_nor2_1 _2713_ (.A(_0611_),
    .B(_0702_),
    .Y(\modem.instance7.instance4._8_[9] ));
 sg13g2_nor2_1 _2714_ (.A(\modem.instance8.instance2._3_[0] ),
    .B(_0932_),
    .Y(_0703_));
 sg13g2_o21ai_1 _2715_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0042_),
    .A2(_0971_));
 sg13g2_nand2b_1 _2716_ (.Y(\modem.instance8.instance2._3_[1] ),
    .B(_0704_),
    .A_N(_0927_));
 sg13g2_inv_1 _2717_ (.Y(_0705_),
    .A(_0042_));
 sg13g2_a21o_1 _2718_ (.A2(_0705_),
    .A1(_0908_),
    .B1(net54),
    .X(_0706_));
 sg13g2_nor2_1 _2719_ (.A(\modem.instance8.instance2._3_[0] ),
    .B(_0936_),
    .Y(_0707_));
 sg13g2_a22oi_1 _2720_ (.Y(\modem.instance8.instance2._3_[2] ),
    .B1(_0706_),
    .B2(_0707_),
    .A2(_0967_),
    .A1(_0936_));
 sg13g2_nand2_1 _2721_ (.Y(_0708_),
    .A(net54),
    .B(_0707_));
 sg13g2_nand2_1 _2722_ (.Y(_0709_),
    .A(_0916_),
    .B(_0905_));
 sg13g2_nor2_1 _2723_ (.A(net54),
    .B(_0705_),
    .Y(_0710_));
 sg13g2_o21ai_1 _2724_ (.B1(_0908_),
    .Y(_0711_),
    .A1(_0709_),
    .A2(_0710_));
 sg13g2_o21ai_1 _2725_ (.B1(_0711_),
    .Y(\modem.instance8.instance2._3_[3] ),
    .A1(net56),
    .A2(_0708_));
 sg13g2_nor2_1 _2726_ (.A(_0928_),
    .B(_0709_),
    .Y(_0712_));
 sg13g2_nand3_1 _2727_ (.B(_0042_),
    .C(_0712_),
    .A(_0932_),
    .Y(_0713_));
 sg13g2_o21ai_1 _2728_ (.B1(_0713_),
    .Y(\modem.instance8.instance2._3_[4] ),
    .A1(_0042_),
    .A2(_0712_));
 sg13g2_xnor2_1 _2729_ (.Y(\modem.instance8.instance3._0_[0] ),
    .A(\modem.instance8._0_[0] ),
    .B(_0548_));
 sg13g2_xnor2_1 _2730_ (.Y(\modem.instance8.instance3._0_[1] ),
    .A(\modem.instance8._0_[1] ),
    .B(_0553_));
 sg13g2_xnor2_1 _2731_ (.Y(\modem.instance8.instance3._0_[2] ),
    .A(\modem.instance8._0_[2] ),
    .B(_0558_));
 sg13g2_xnor2_1 _2732_ (.Y(\modem.instance8.instance3._0_[3] ),
    .A(\modem.instance8._0_[3] ),
    .B(_0563_));
 sg13g2_xnor2_1 _2733_ (.Y(\modem.instance8.instance3._0_[4] ),
    .A(\modem.instance8._0_[4] ),
    .B(_0568_));
 sg13g2_xnor2_1 _2734_ (.Y(\modem.instance8.instance3._0_[5] ),
    .A(\modem.instance8._0_[5] ),
    .B(_0573_));
 sg13g2_and4_1 _2735_ (.A(\modem.instance8._1_[3] ),
    .B(\modem.instance8._1_[4] ),
    .C(\modem.instance8._1_[5] ),
    .D(_0608_),
    .X(_0714_));
 sg13g2_nand4_1 _2736_ (.B(\modem.instance8._1_[1] ),
    .C(\modem.instance8._1_[2] ),
    .A(\modem.instance8._1_[0] ),
    .Y(_0715_),
    .D(_0714_));
 sg13g2_buf_1 _2737_ (.A(_0715_),
    .X(_0716_));
 sg13g2_buf_2 _2738_ (.A(\modem.instance8.instance5._9_[1] ),
    .X(_0717_));
 sg13g2_inv_1 _2739_ (.Y(_0718_),
    .A(_0045_));
 sg13g2_buf_2 _2740_ (.A(\modem.instance8.instance5._9_[16] ),
    .X(_0719_));
 sg13g2_nor4_1 _2741_ (.A(_0719_),
    .B(\modem.instance8.instance5._9_[23] ),
    .C(\modem.instance8.instance5._9_[22] ),
    .D(\modem.instance8.instance5._9_[24] ),
    .Y(_0720_));
 sg13g2_nor4_1 _2742_ (.A(\modem.instance8.instance5._9_[19] ),
    .B(\modem.instance8.instance5._9_[18] ),
    .C(\modem.instance8.instance5._9_[21] ),
    .D(\modem.instance8.instance5._9_[20] ),
    .Y(_0721_));
 sg13g2_buf_2 _2743_ (.A(\modem.instance8.instance5._9_[25] ),
    .X(_0722_));
 sg13g2_nor4_1 _2744_ (.A(\modem.instance8.instance5._9_[3] ),
    .B(_0722_),
    .C(\modem.instance8.instance5._9_[31] ),
    .D(\modem.instance8.instance5._9_[30] ),
    .Y(_0723_));
 sg13g2_nor4_1 _2745_ (.A(\modem.instance8.instance5._9_[27] ),
    .B(\modem.instance8.instance5._9_[26] ),
    .C(\modem.instance8.instance5._9_[29] ),
    .D(\modem.instance8.instance5._9_[28] ),
    .Y(_0724_));
 sg13g2_nand4_1 _2746_ (.B(_0721_),
    .C(_0723_),
    .A(_0720_),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_buf_2 _2747_ (.A(\modem.instance8.instance5._9_[15] ),
    .X(_0726_));
 sg13g2_nor2_1 _2748_ (.A(_0726_),
    .B(\modem.instance8.instance5._9_[14] ),
    .Y(_0727_));
 sg13g2_nor4_1 _2749_ (.A(\modem.instance8.instance5._9_[8] ),
    .B(\modem.instance8.instance5._9_[10] ),
    .C(\modem.instance8.instance5._9_[13] ),
    .D(\modem.instance8.instance5._9_[12] ),
    .Y(_0728_));
 sg13g2_buf_1 _2750_ (.A(\modem.instance8.instance5._9_[11] ),
    .X(_0729_));
 sg13g2_nor4_1 _2751_ (.A(\modem.instance8.instance5._9_[6] ),
    .B(\modem.instance8.instance5._9_[9] ),
    .C(_0729_),
    .D(\modem.instance8.instance5._9_[17] ),
    .Y(_0730_));
 sg13g2_nor4_1 _2752_ (.A(\modem.instance8.instance5._9_[2] ),
    .B(\modem.instance8.instance5._9_[5] ),
    .C(\modem.instance8.instance5._9_[4] ),
    .D(\modem.instance8.instance5._9_[7] ),
    .Y(_0731_));
 sg13g2_nand4_1 _2753_ (.B(_0728_),
    .C(_0730_),
    .A(_0727_),
    .Y(_0732_),
    .D(_0731_));
 sg13g2_nor4_1 _2754_ (.A(_0717_),
    .B(_0718_),
    .C(_0725_),
    .D(_0732_),
    .Y(_0733_));
 sg13g2_nor2_1 _2755_ (.A(_0725_),
    .B(_0732_),
    .Y(_0734_));
 sg13g2_buf_1 _2756_ (.A(\modem.instance8.instance5._9_[0] ),
    .X(_0735_));
 sg13g2_nand2_2 _2757_ (.Y(_0736_),
    .A(_0735_),
    .B(_0717_));
 sg13g2_a21oi_1 _2758_ (.A1(_0734_),
    .A2(_0736_),
    .Y(_0737_),
    .B1(_0045_));
 sg13g2_nor3_1 _2759_ (.A(_0716_),
    .B(_0733_),
    .C(_0737_),
    .Y(\modem.instance8.instance5._7_ ));
 sg13g2_buf_1 _2760_ (.A(_0716_),
    .X(_0738_));
 sg13g2_nor2_1 _2761_ (.A(_0735_),
    .B(_0738_),
    .Y(\modem.instance8.instance5._8_[0] ));
 sg13g2_nand4_1 _2762_ (.B(\modem.instance8.instance5._9_[2] ),
    .C(\modem.instance8.instance5._9_[5] ),
    .A(\modem.instance8.instance5._9_[3] ),
    .Y(_0739_),
    .D(\modem.instance8.instance5._9_[4] ));
 sg13g2_buf_1 _2763_ (.A(_0739_),
    .X(_0740_));
 sg13g2_nand3_1 _2764_ (.B(\modem.instance8.instance5._9_[6] ),
    .C(\modem.instance8.instance5._9_[8] ),
    .A(\modem.instance8.instance5._9_[7] ),
    .Y(_0741_));
 sg13g2_nor3_2 _2765_ (.A(_0736_),
    .B(_0740_),
    .C(_0741_),
    .Y(_0742_));
 sg13g2_buf_1 _2766_ (.A(_0742_),
    .X(_0743_));
 sg13g2_nand2_1 _2767_ (.Y(_0744_),
    .A(\modem.instance8.instance5._9_[9] ),
    .B(_0743_));
 sg13g2_xor2_1 _2768_ (.B(_0744_),
    .A(\modem.instance8.instance5._9_[10] ),
    .X(_0745_));
 sg13g2_nor2_1 _2769_ (.A(net13),
    .B(_0745_),
    .Y(\modem.instance8.instance5._8_[10] ));
 sg13g2_and2_1 _2770_ (.A(\modem.instance8.instance5._9_[9] ),
    .B(\modem.instance8.instance5._9_[10] ),
    .X(_0746_));
 sg13g2_buf_1 _2771_ (.A(_0746_),
    .X(_0747_));
 sg13g2_nand2_1 _2772_ (.Y(_0748_),
    .A(net14),
    .B(_0747_));
 sg13g2_xor2_1 _2773_ (.B(_0748_),
    .A(_0729_),
    .X(_0749_));
 sg13g2_nor2_1 _2774_ (.A(net13),
    .B(_0749_),
    .Y(\modem.instance8.instance5._8_[11] ));
 sg13g2_nand3_1 _2775_ (.B(net14),
    .C(_0747_),
    .A(_0729_),
    .Y(_0750_));
 sg13g2_xor2_1 _2776_ (.B(_0750_),
    .A(\modem.instance8.instance5._9_[12] ),
    .X(_0751_));
 sg13g2_nor2_1 _2777_ (.A(net13),
    .B(_0751_),
    .Y(\modem.instance8.instance5._8_[12] ));
 sg13g2_nand4_1 _2778_ (.B(\modem.instance8.instance5._9_[12] ),
    .C(_0742_),
    .A(_0729_),
    .Y(_0752_),
    .D(_0747_));
 sg13g2_xor2_1 _2779_ (.B(_0752_),
    .A(\modem.instance8.instance5._9_[13] ),
    .X(_0753_));
 sg13g2_nor2_1 _2780_ (.A(net13),
    .B(_0753_),
    .Y(\modem.instance8.instance5._8_[13] ));
 sg13g2_and3_1 _2781_ (.X(_0754_),
    .A(_0729_),
    .B(\modem.instance8.instance5._9_[13] ),
    .C(\modem.instance8.instance5._9_[12] ));
 sg13g2_nand3_1 _2782_ (.B(_0747_),
    .C(_0754_),
    .A(net14),
    .Y(_0755_));
 sg13g2_xor2_1 _2783_ (.B(_0755_),
    .A(\modem.instance8.instance5._9_[14] ),
    .X(_0756_));
 sg13g2_nor2_1 _2784_ (.A(net13),
    .B(_0756_),
    .Y(\modem.instance8.instance5._8_[14] ));
 sg13g2_and3_1 _2785_ (.X(_0757_),
    .A(\modem.instance8.instance5._9_[14] ),
    .B(_0747_),
    .C(_0754_));
 sg13g2_buf_2 _2786_ (.A(_0757_),
    .X(_0758_));
 sg13g2_nand2_1 _2787_ (.Y(_0759_),
    .A(net14),
    .B(_0758_));
 sg13g2_xor2_1 _2788_ (.B(_0759_),
    .A(_0726_),
    .X(_0760_));
 sg13g2_nor2_1 _2789_ (.A(net13),
    .B(_0760_),
    .Y(\modem.instance8.instance5._8_[15] ));
 sg13g2_nand3_1 _2790_ (.B(net14),
    .C(_0758_),
    .A(_0726_),
    .Y(_0761_));
 sg13g2_xor2_1 _2791_ (.B(_0761_),
    .A(_0719_),
    .X(_0762_));
 sg13g2_nor2_1 _2792_ (.A(net13),
    .B(_0762_),
    .Y(\modem.instance8.instance5._8_[16] ));
 sg13g2_nand2b_1 _2793_ (.Y(_0763_),
    .B(_0719_),
    .A_N(_0044_));
 sg13g2_nand2_1 _2794_ (.Y(_0764_),
    .A(_0717_),
    .B(_0726_));
 sg13g2_nor4_1 _2795_ (.A(_0740_),
    .B(_0741_),
    .C(_0763_),
    .D(_0764_),
    .Y(_0765_));
 sg13g2_nand2_1 _2796_ (.Y(_0766_),
    .A(_0758_),
    .B(_0765_));
 sg13g2_xor2_1 _2797_ (.B(_0766_),
    .A(\modem.instance8.instance5._9_[17] ),
    .X(_0767_));
 sg13g2_nor2_1 _2798_ (.A(_0738_),
    .B(_0767_),
    .Y(\modem.instance8.instance5._8_[17] ));
 sg13g2_and2_1 _2799_ (.A(_0726_),
    .B(\modem.instance8.instance5._9_[17] ),
    .X(_0768_));
 sg13g2_nand4_1 _2800_ (.B(_0742_),
    .C(_0758_),
    .A(_0719_),
    .Y(_0769_),
    .D(_0768_));
 sg13g2_xor2_1 _2801_ (.B(_0769_),
    .A(\modem.instance8.instance5._9_[18] ),
    .X(_0770_));
 sg13g2_nor2_1 _2802_ (.A(net13),
    .B(_0770_),
    .Y(\modem.instance8.instance5._8_[18] ));
 sg13g2_buf_1 _2803_ (.A(_0716_),
    .X(_0771_));
 sg13g2_and3_1 _2804_ (.X(_0772_),
    .A(_0719_),
    .B(\modem.instance8.instance5._9_[18] ),
    .C(_0768_));
 sg13g2_nand3_1 _2805_ (.B(_0758_),
    .C(_0772_),
    .A(net14),
    .Y(_0773_));
 sg13g2_xor2_1 _2806_ (.B(_0773_),
    .A(\modem.instance8.instance5._9_[19] ),
    .X(_0774_));
 sg13g2_nor2_1 _2807_ (.A(net12),
    .B(_0774_),
    .Y(\modem.instance8.instance5._8_[19] ));
 sg13g2_xnor2_1 _2808_ (.Y(_0775_),
    .A(_0735_),
    .B(_0717_));
 sg13g2_nor2_1 _2809_ (.A(net12),
    .B(_0775_),
    .Y(\modem.instance8.instance5._8_[1] ));
 sg13g2_nand4_1 _2810_ (.B(_0742_),
    .C(_0758_),
    .A(\modem.instance8.instance5._9_[19] ),
    .Y(_0776_),
    .D(_0772_));
 sg13g2_xor2_1 _2811_ (.B(_0776_),
    .A(\modem.instance8.instance5._9_[20] ),
    .X(_0777_));
 sg13g2_nor2_1 _2812_ (.A(net12),
    .B(_0777_),
    .Y(\modem.instance8.instance5._8_[20] ));
 sg13g2_nand4_1 _2813_ (.B(\modem.instance8.instance5._9_[17] ),
    .C(_0719_),
    .A(_0726_),
    .Y(_0778_),
    .D(\modem.instance8.instance5._9_[18] ));
 sg13g2_nand2_1 _2814_ (.Y(_0779_),
    .A(\modem.instance8.instance5._9_[19] ),
    .B(\modem.instance8.instance5._9_[20] ));
 sg13g2_nor2_1 _2815_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_nand3_1 _2816_ (.B(_0758_),
    .C(_0780_),
    .A(net14),
    .Y(_0781_));
 sg13g2_xor2_1 _2817_ (.B(_0781_),
    .A(\modem.instance8.instance5._9_[21] ),
    .X(_0782_));
 sg13g2_nor2_1 _2818_ (.A(net12),
    .B(_0782_),
    .Y(\modem.instance8.instance5._8_[21] ));
 sg13g2_nand4_1 _2819_ (.B(_0742_),
    .C(_0758_),
    .A(\modem.instance8.instance5._9_[21] ),
    .Y(_0783_),
    .D(_0780_));
 sg13g2_xor2_1 _2820_ (.B(_0783_),
    .A(\modem.instance8.instance5._9_[22] ),
    .X(_0784_));
 sg13g2_nor2_1 _2821_ (.A(net12),
    .B(_0784_),
    .Y(\modem.instance8.instance5._8_[22] ));
 sg13g2_nand4_1 _2822_ (.B(_0729_),
    .C(\modem.instance8.instance5._9_[10] ),
    .A(\modem.instance8.instance5._9_[9] ),
    .Y(_0785_),
    .D(\modem.instance8.instance5._9_[12] ));
 sg13g2_nand4_1 _2823_ (.B(\modem.instance8.instance5._9_[14] ),
    .C(\modem.instance8.instance5._9_[21] ),
    .A(\modem.instance8.instance5._9_[13] ),
    .Y(_0786_),
    .D(\modem.instance8.instance5._9_[22] ));
 sg13g2_nor4_2 _2824_ (.A(_0778_),
    .B(_0779_),
    .C(_0785_),
    .Y(_0787_),
    .D(_0786_));
 sg13g2_nand2_1 _2825_ (.Y(_0788_),
    .A(net14),
    .B(_0787_));
 sg13g2_xor2_1 _2826_ (.B(_0788_),
    .A(\modem.instance8.instance5._9_[23] ),
    .X(_0789_));
 sg13g2_nor2_1 _2827_ (.A(net12),
    .B(_0789_),
    .Y(\modem.instance8.instance5._8_[23] ));
 sg13g2_nand3_1 _2828_ (.B(_0742_),
    .C(_0787_),
    .A(\modem.instance8.instance5._9_[23] ),
    .Y(_0790_));
 sg13g2_xor2_1 _2829_ (.B(_0790_),
    .A(\modem.instance8.instance5._9_[24] ),
    .X(_0791_));
 sg13g2_nor2_1 _2830_ (.A(net12),
    .B(_0791_),
    .Y(\modem.instance8.instance5._8_[24] ));
 sg13g2_nand2_1 _2831_ (.Y(_0792_),
    .A(\modem.instance8.instance5._9_[23] ),
    .B(\modem.instance8.instance5._9_[24] ));
 sg13g2_nor4_2 _2832_ (.A(_0736_),
    .B(_0740_),
    .C(_0741_),
    .Y(_0793_),
    .D(_0792_));
 sg13g2_and2_1 _2833_ (.A(_0787_),
    .B(_0793_),
    .X(_0794_));
 sg13g2_xnor2_1 _2834_ (.Y(_0795_),
    .A(_0722_),
    .B(_0794_));
 sg13g2_nor2_1 _2835_ (.A(_0771_),
    .B(_0795_),
    .Y(\modem.instance8.instance5._8_[25] ));
 sg13g2_nand3_1 _2836_ (.B(_0787_),
    .C(_0793_),
    .A(_0722_),
    .Y(_0796_));
 sg13g2_xor2_1 _2837_ (.B(_0796_),
    .A(\modem.instance8.instance5._9_[26] ),
    .X(_0797_));
 sg13g2_nor2_1 _2838_ (.A(net12),
    .B(_0797_),
    .Y(\modem.instance8.instance5._8_[26] ));
 sg13g2_nand4_1 _2839_ (.B(\modem.instance8.instance5._9_[26] ),
    .C(_0787_),
    .A(_0722_),
    .Y(_0798_),
    .D(_0793_));
 sg13g2_xor2_1 _2840_ (.B(_0798_),
    .A(\modem.instance8.instance5._9_[27] ),
    .X(_0799_));
 sg13g2_nor2_1 _2841_ (.A(_0771_),
    .B(_0799_),
    .Y(\modem.instance8.instance5._8_[27] ));
 sg13g2_buf_1 _2842_ (.A(_0716_),
    .X(_0800_));
 sg13g2_and2_1 _2843_ (.A(\modem.instance8.instance5._9_[27] ),
    .B(\modem.instance8.instance5._9_[26] ),
    .X(_0801_));
 sg13g2_nand4_1 _2844_ (.B(_0787_),
    .C(_0793_),
    .A(_0722_),
    .Y(_0802_),
    .D(_0801_));
 sg13g2_xor2_1 _2845_ (.B(_0802_),
    .A(\modem.instance8.instance5._9_[28] ),
    .X(_0803_));
 sg13g2_nor2_1 _2846_ (.A(_0800_),
    .B(_0803_),
    .Y(\modem.instance8.instance5._8_[28] ));
 sg13g2_and2_1 _2847_ (.A(_0722_),
    .B(\modem.instance8.instance5._9_[28] ),
    .X(_0804_));
 sg13g2_nand4_1 _2848_ (.B(_0793_),
    .C(_0801_),
    .A(_0787_),
    .Y(_0805_),
    .D(_0804_));
 sg13g2_xor2_1 _2849_ (.B(_0805_),
    .A(\modem.instance8.instance5._9_[29] ),
    .X(_0806_));
 sg13g2_nor2_1 _2850_ (.A(net11),
    .B(_0806_),
    .Y(\modem.instance8.instance5._8_[29] ));
 sg13g2_xor2_1 _2851_ (.B(_0736_),
    .A(\modem.instance8.instance5._9_[2] ),
    .X(_0807_));
 sg13g2_nor2_1 _2852_ (.A(net11),
    .B(_0807_),
    .Y(\modem.instance8.instance5._8_[2] ));
 sg13g2_inv_1 _2853_ (.Y(_0808_),
    .A(\modem.instance8.instance5._9_[30] ));
 sg13g2_and4_1 _2854_ (.A(_0722_),
    .B(\modem.instance8.instance5._9_[29] ),
    .C(\modem.instance8.instance5._9_[28] ),
    .D(_0801_),
    .X(_0809_));
 sg13g2_nand3_1 _2855_ (.B(_0793_),
    .C(_0809_),
    .A(_0787_),
    .Y(_0810_));
 sg13g2_xnor2_1 _2856_ (.Y(_0811_),
    .A(_0808_),
    .B(_0810_));
 sg13g2_nor2_1 _2857_ (.A(_0800_),
    .B(_0811_),
    .Y(\modem.instance8.instance5._8_[30] ));
 sg13g2_o21ai_1 _2858_ (.B1(_0718_),
    .Y(_0812_),
    .A1(_0808_),
    .A2(_0810_));
 sg13g2_nand4_1 _2859_ (.B(_0045_),
    .C(_0794_),
    .A(\modem.instance8.instance5._9_[30] ),
    .Y(_0813_),
    .D(_0809_));
 sg13g2_a21oi_1 _2860_ (.A1(_0812_),
    .A2(_0813_),
    .Y(\modem.instance8.instance5._8_[31] ),
    .B1(_0716_));
 sg13g2_nand3_1 _2861_ (.B(_0717_),
    .C(\modem.instance8.instance5._9_[2] ),
    .A(_0735_),
    .Y(_0814_));
 sg13g2_xor2_1 _2862_ (.B(_0814_),
    .A(\modem.instance8.instance5._9_[3] ),
    .X(_0815_));
 sg13g2_nor2_1 _2863_ (.A(net11),
    .B(_0815_),
    .Y(\modem.instance8.instance5._8_[3] ));
 sg13g2_inv_1 _2864_ (.Y(_0816_),
    .A(\modem.instance8.instance5._9_[4] ));
 sg13g2_nand4_1 _2865_ (.B(_0717_),
    .C(\modem.instance8.instance5._9_[3] ),
    .A(_0735_),
    .Y(_0817_),
    .D(\modem.instance8.instance5._9_[2] ));
 sg13g2_xnor2_1 _2866_ (.Y(_0818_),
    .A(_0816_),
    .B(_0817_));
 sg13g2_nor2_1 _2867_ (.A(net11),
    .B(_0818_),
    .Y(\modem.instance8.instance5._8_[4] ));
 sg13g2_nor2_1 _2868_ (.A(_0816_),
    .B(_0817_),
    .Y(_0819_));
 sg13g2_xnor2_1 _2869_ (.Y(_0820_),
    .A(\modem.instance8.instance5._9_[5] ),
    .B(_0819_));
 sg13g2_nor2_1 _2870_ (.A(net11),
    .B(_0820_),
    .Y(\modem.instance8.instance5._8_[5] ));
 sg13g2_nor2_1 _2871_ (.A(_0736_),
    .B(_0740_),
    .Y(_0821_));
 sg13g2_xnor2_1 _2872_ (.Y(_0822_),
    .A(\modem.instance8.instance5._9_[6] ),
    .B(_0821_));
 sg13g2_nor2_1 _2873_ (.A(net11),
    .B(_0822_),
    .Y(\modem.instance8.instance5._8_[6] ));
 sg13g2_nand2_1 _2874_ (.Y(_0823_),
    .A(\modem.instance8.instance5._9_[6] ),
    .B(_0821_));
 sg13g2_xor2_1 _2875_ (.B(_0823_),
    .A(\modem.instance8.instance5._9_[7] ),
    .X(_0824_));
 sg13g2_nor2_1 _2876_ (.A(net11),
    .B(_0824_),
    .Y(\modem.instance8.instance5._8_[7] ));
 sg13g2_nand3_1 _2877_ (.B(\modem.instance8.instance5._9_[6] ),
    .C(_0821_),
    .A(\modem.instance8.instance5._9_[7] ),
    .Y(_0825_));
 sg13g2_xor2_1 _2878_ (.B(_0825_),
    .A(\modem.instance8.instance5._9_[8] ),
    .X(_0826_));
 sg13g2_nor2_1 _2879_ (.A(net11),
    .B(_0826_),
    .Y(\modem.instance8.instance5._8_[8] ));
 sg13g2_xnor2_1 _2880_ (.Y(_0827_),
    .A(\modem.instance8.instance5._9_[9] ),
    .B(_0743_));
 sg13g2_nor2_1 _2881_ (.A(_0716_),
    .B(_0827_),
    .Y(\modem.instance8.instance5._8_[9] ));
 sg13g2_inv_1 _2882_ (.Y(_0828_),
    .A(_0547_));
 sg13g2_mux2_1 _2883_ (.A0(\modem._4_ ),
    .A1(\modem._6_ ),
    .S(_0545_),
    .X(_0829_));
 sg13g2_a22oi_1 _2884_ (.Y(_0830_),
    .B1(_0829_),
    .B2(_0544_),
    .A2(_0828_),
    .A1(\modem._5_ ));
 sg13g2_inv_1 _2885_ (.Y(\modem.instance9._5_ ),
    .A(_0830_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \modem.instance1.instance2.ffd0._1_$_DFF_N__173  (.L_HI(net173));
 sg13g2_buf_1 _2888_ (.A(net156),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2889_ (.A(net157),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2890_ (.A(net158),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2891_ (.A(net159),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2892_ (.A(net160),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2893_ (.A(net161),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2894_ (.A(net162),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2895_ (.A(net163),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2896_ (.A(net164),
    .X(uio_out[0]));
 sg13g2_buf_1 _2897_ (.A(net165),
    .X(uio_out[1]));
 sg13g2_buf_1 _2898_ (.A(net166),
    .X(uio_out[2]));
 sg13g2_buf_1 _2899_ (.A(net167),
    .X(uio_out[3]));
 sg13g2_buf_1 _2900_ (.A(net168),
    .X(uio_out[4]));
 sg13g2_buf_1 _2901_ (.A(net169),
    .X(uio_out[5]));
 sg13g2_buf_1 _2902_ (.A(net170),
    .X(uio_out[6]));
 sg13g2_buf_1 _2903_ (.A(net171),
    .X(uio_out[7]));
 sg13g2_buf_1 _2904_ (.A(net172),
    .X(uo_out[6]));
 sg13g2_buf_1 _2905_ (.A(demod_out),
    .X(net8));
 sg13g2_dfrbp_1 \modem.instance1.instance1._5_$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net110),
    .D(_0063_),
    .Q_N(\modem.instance1.instance1._1_ ),
    .Q(\modem.instance1._0_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[0]$_DFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net110),
    .D(\modem.instance1.instance1._3_[0] ),
    .Q_N(_1289_),
    .Q(\modem.instance1.instance1._6_[0] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[1]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance1.instance1._3_[1] ),
    .Q_N(_1290_),
    .Q(\modem.instance1.instance1._6_[1] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[2]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance1.instance1._3_[2] ),
    .Q_N(_1291_),
    .Q(\modem.instance1.instance1._6_[2] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[3]$_DFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net111),
    .D(\modem.instance1.instance1._3_[3] ),
    .Q_N(_1292_),
    .Q(\modem.instance1.instance1._6_[3] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[4]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance1.instance1._3_[4] ),
    .Q_N(_1293_),
    .Q(\modem.instance1.instance1._6_[4] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[5]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance1.instance1._3_[5] ),
    .Q_N(_1294_),
    .Q(\modem.instance1.instance1._6_[5] ));
 sg13g2_dfrbp_1 \modem.instance1.instance1._6_[6]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net130),
    .D(\modem.instance1.instance1._3_[6] ),
    .Q_N(_1288_),
    .Q(\modem.instance1.instance1._6_[6] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._02_$_DFFE_NN0N_  (.CLK(net96),
    .RESET_B(net131),
    .D(_0064_),
    .Q_N(_1287_),
    .Q(\modem.instance1._1_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[0]$_DFF_NN0_  (.CLK(net95),
    .RESET_B(net102),
    .D(\modem.instance1.instance2._09_[0] ),
    .Q_N(_1286_),
    .Q(\modem.instance1.instance2._10_[0] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[10]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[10] ),
    .Q_N(_1285_),
    .Q(\modem.instance1.instance2._10_[10] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[11]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[11] ),
    .Q_N(_1284_),
    .Q(\modem.instance1.instance2._10_[11] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[12]$_DFF_NN0_  (.CLK(net93),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[12] ),
    .Q_N(_1283_),
    .Q(\modem.instance1.instance2._10_[12] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[13]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[13] ),
    .Q_N(_1282_),
    .Q(\modem.instance1.instance2._10_[13] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[14]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[14] ),
    .Q_N(_1281_),
    .Q(\modem.instance1.instance2._10_[14] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[15]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[15] ),
    .Q_N(_1280_),
    .Q(\modem.instance1.instance2._10_[15] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[16]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[16] ),
    .Q_N(_1279_),
    .Q(\modem.instance1.instance2._10_[16] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[17]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[17] ),
    .Q_N(_1278_),
    .Q(\modem.instance1.instance2._10_[17] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[18]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[18] ),
    .Q_N(_1277_),
    .Q(\modem.instance1.instance2._10_[18] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[19]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[19] ),
    .Q_N(_1276_),
    .Q(\modem.instance1.instance2._10_[19] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[1]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[1] ),
    .Q_N(_1275_),
    .Q(\modem.instance1.instance2._10_[1] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[20]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[20] ),
    .Q_N(_1274_),
    .Q(\modem.instance1.instance2._10_[20] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[21]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[21] ),
    .Q_N(_1273_),
    .Q(\modem.instance1.instance2._10_[21] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[22]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net101),
    .D(\modem.instance1.instance2._09_[22] ),
    .Q_N(_1272_),
    .Q(\modem.instance1.instance2._10_[22] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[23]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[23] ),
    .Q_N(_1271_),
    .Q(\modem.instance1.instance2._10_[23] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[24]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[24] ),
    .Q_N(_1270_),
    .Q(\modem.instance1.instance2._10_[24] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[25]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[25] ),
    .Q_N(_1269_),
    .Q(\modem.instance1.instance2._10_[25] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[26]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[26] ),
    .Q_N(_1268_),
    .Q(\modem.instance1.instance2._10_[26] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[27]$_DFF_NN0_  (.CLK(net97),
    .RESET_B(net110),
    .D(\modem.instance1.instance2._09_[27] ),
    .Q_N(_1267_),
    .Q(\modem.instance1.instance2._10_[27] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[28]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net110),
    .D(\modem.instance1.instance2._09_[28] ),
    .Q_N(_1266_),
    .Q(\modem.instance1.instance2._10_[28] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[29]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[29] ),
    .Q_N(_1265_),
    .Q(\modem.instance1.instance2._10_[29] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[2]$_DFF_NN0_  (.CLK(net94),
    .RESET_B(net102),
    .D(\modem.instance1.instance2._09_[2] ),
    .Q_N(_1264_),
    .Q(\modem.instance1.instance2._10_[2] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[30]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[30] ),
    .Q_N(_1263_),
    .Q(\modem.instance1.instance2._10_[30] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[31]$_DFF_NN0_  (.CLK(net98),
    .RESET_B(net108),
    .D(\modem.instance1.instance2._09_[31] ),
    .Q_N(_1262_),
    .Q(\modem.instance1.instance2._10_[31] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[3]$_DFF_NN0_  (.CLK(net95),
    .RESET_B(net102),
    .D(\modem.instance1.instance2._09_[3] ),
    .Q_N(_1261_),
    .Q(\modem.instance1.instance2._10_[3] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[4]$_DFF_NN0_  (.CLK(net93),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[4] ),
    .Q_N(_1260_),
    .Q(\modem.instance1.instance2._10_[4] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[5]$_DFF_NN0_  (.CLK(net93),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[5] ),
    .Q_N(_1259_),
    .Q(\modem.instance1.instance2._10_[5] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[6]$_DFF_NN0_  (.CLK(net93),
    .RESET_B(net100),
    .D(\modem.instance1.instance2._09_[6] ),
    .Q_N(_1258_),
    .Q(\modem.instance1.instance2._10_[6] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[7]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net99),
    .D(\modem.instance1.instance2._09_[7] ),
    .Q_N(_1257_),
    .Q(\modem.instance1.instance2._10_[7] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[8]$_DFF_NN0_  (.CLK(net92),
    .RESET_B(net100),
    .D(\modem.instance1.instance2._09_[8] ),
    .Q_N(_1256_),
    .Q(\modem.instance1.instance2._10_[8] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2._10_[9]$_DFF_NN0_  (.CLK(net93),
    .RESET_B(net100),
    .D(\modem.instance1.instance2._09_[9] ),
    .Q_N(_1255_),
    .Q(\modem.instance1.instance2._10_[9] ));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd0._0_$_DFF_NN1_  (.CLK(net96),
    .RESET_B(net111),
    .D(_0060_),
    .Q_N(\modem.instance1.instance2.ffd0._0_ ),
    .Q(_1465_));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd0._1_$_DFF_N_  (.CLK(net96),
    .RESET_B(net173),
    .D(\modem.instance1.instance2.ffd0._0_ ),
    .Q_N(_1254_),
    .Q(\modem.instance1.instance2._00_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd2._0_$_DFF_NN1_  (.CLK(net96),
    .RESET_B(net111),
    .D(_1254_),
    .Q_N(\modem.instance1.instance2.ffd2._0_ ),
    .Q(_1466_));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd2._1_$_DFF_N_  (.CLK(net96),
    .RESET_B(net174),
    .D(\modem.instance1.instance2.ffd2._0_ ),
    .Q_N(_1253_),
    .Q(\modem.instance1.instance2._03_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd3._0_$_DFF_NN1_  (.CLK(net97),
    .RESET_B(net111),
    .D(_1253_),
    .Q_N(\modem.instance1.instance2.ffd3._0_ ),
    .Q(_1467_));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd3._1_$_DFF_N_  (.CLK(net96),
    .RESET_B(net175),
    .D(\modem.instance1.instance2.ffd3._0_ ),
    .Q_N(_1252_),
    .Q(\modem.instance1.instance2._04_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd4._0_$_DFF_NN1_  (.CLK(net96),
    .RESET_B(net130),
    .D(_1252_),
    .Q_N(\modem.instance1.instance2.ffd4._0_ ),
    .Q(_1468_));
 sg13g2_dfrbp_1 \modem.instance1.instance2.ffd4._1_$_DFF_N_  (.CLK(net96),
    .RESET_B(net176),
    .D(\modem.instance1.instance2.ffd4._0_ ),
    .Q_N(_1295_),
    .Q(\modem.instance1.instance2._05_ ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._4_[0]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(net34),
    .Q_N(_1296_),
    .Q(\modem.instance1.instance3._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._4_[1]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(\modem.instance1.instance3._3_[1] ),
    .Q_N(_0059_),
    .Q(\modem.instance1.instance3._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._4_[2]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net131),
    .D(\modem.instance1.instance3._3_[2] ),
    .Q_N(_1297_),
    .Q(\modem.instance1.instance3._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._4_[3]$_DFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net115),
    .D(\modem.instance1.instance3._3_[3] ),
    .Q_N(_1298_),
    .Q(\modem.instance1.instance3._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._4_[4]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(\modem.instance1.instance3._3_[4] ),
    .Q_N(_1299_),
    .Q(\modem.instance1.instance3._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[0]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(_0000_),
    .Q_N(_1300_),
    .Q(\modem.instance1._2_[0] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[1]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net131),
    .D(_0001_),
    .Q_N(_1301_),
    .Q(\modem.instance1._2_[1] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[2]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net132),
    .D(_0002_),
    .Q_N(_1302_),
    .Q(\modem.instance1._2_[2] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[3]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net132),
    .D(_0003_),
    .Q_N(_1303_),
    .Q(\modem.instance1._2_[3] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[4]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net132),
    .D(_0004_),
    .Q_N(_1304_),
    .Q(\modem.instance1._2_[4] ));
 sg13g2_dfrbp_1 \modem.instance1.instance3._5_[5]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net136),
    .D(_0005_),
    .Q_N(_1305_),
    .Q(\modem.instance1._2_[5] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[0]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net142),
    .D(\modem.instance1.instance4._0_[0] ),
    .Q_N(_1306_),
    .Q(\modem._0_[0] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[1]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net142),
    .D(\modem.instance1.instance4._0_[1] ),
    .Q_N(_1307_),
    .Q(\modem._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[2]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net142),
    .D(\modem.instance1.instance4._0_[2] ),
    .Q_N(_1308_),
    .Q(\modem._0_[2] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[3]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net132),
    .D(\modem.instance1.instance4._0_[3] ),
    .Q_N(_1309_),
    .Q(\modem._0_[3] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[4]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net142),
    .D(\modem.instance1.instance4._0_[4] ),
    .Q_N(_1310_),
    .Q(\modem._0_[4] ));
 sg13g2_dfrbp_1 \modem.instance1.instance4._1_[5]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net136),
    .D(\modem.instance1.instance4._0_[5] ),
    .Q_N(_1251_),
    .Q(\modem._0_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._5_$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net113),
    .D(_0065_),
    .Q_N(\modem.instance2.instance1._1_ ),
    .Q(\modem.instance2._0_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[0]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net111),
    .D(\modem.instance2.instance1._3_[0] ),
    .Q_N(_1311_),
    .Q(\modem.instance2.instance1._6_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[1]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net109),
    .D(\modem.instance2.instance1._3_[1] ),
    .Q_N(_1312_),
    .Q(\modem.instance2.instance1._6_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[2]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net111),
    .D(\modem.instance2.instance1._3_[2] ),
    .Q_N(_1313_),
    .Q(\modem.instance2.instance1._6_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[3]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net109),
    .D(\modem.instance2.instance1._3_[3] ),
    .Q_N(_1314_),
    .Q(\modem.instance2.instance1._6_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[4]$_DFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net109),
    .D(\modem.instance2.instance1._3_[4] ),
    .Q_N(_1315_),
    .Q(\modem.instance2.instance1._6_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[5]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net109),
    .D(\modem.instance2.instance1._3_[5] ),
    .Q_N(_1316_),
    .Q(\modem.instance2.instance1._6_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance1._6_[6]$_DFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net110),
    .D(\modem.instance2.instance1._3_[6] ),
    .Q_N(_1250_),
    .Q(\modem.instance2.instance1._6_[6] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._5_$_DFFE_PN0N_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net130),
    .D(_0066_),
    .Q_N(\modem.instance2.instance2._1_ ),
    .Q(\modem.instance2._1_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[0]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance2.instance2._3_[0] ),
    .Q_N(_1317_),
    .Q(\modem.instance2.instance2._6_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[1]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net130),
    .D(\modem.instance2.instance2._3_[1] ),
    .Q_N(_1318_),
    .Q(\modem.instance2.instance2._6_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[2]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance2.instance2._3_[2] ),
    .Q_N(_1319_),
    .Q(\modem.instance2.instance2._6_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[3]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net129),
    .D(\modem.instance2.instance2._3_[3] ),
    .Q_N(_1320_),
    .Q(\modem.instance2.instance2._6_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[4]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net110),
    .D(\modem.instance2.instance2._3_[4] ),
    .Q_N(_1321_),
    .Q(\modem.instance2.instance2._6_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[5]$_DFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net110),
    .D(\modem.instance2.instance2._3_[5] ),
    .Q_N(_1322_),
    .Q(\modem.instance2.instance2._6_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance2._6_[6]$_DFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net110),
    .D(\modem.instance2.instance2._3_[6] ),
    .Q_N(_1323_),
    .Q(\modem.instance2.instance2._6_[6] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._4_[0]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net134),
    .D(\modem.instance2.instance3._3_[0] ),
    .Q_N(_1324_),
    .Q(\modem.instance2.instance3._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._4_[1]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net135),
    .D(\modem.instance2.instance3._3_[1] ),
    .Q_N(_0047_),
    .Q(\modem.instance2.instance3._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._4_[2]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net134),
    .D(\modem.instance2.instance3._3_[2] ),
    .Q_N(_1325_),
    .Q(\modem.instance2.instance3._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._4_[3]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net134),
    .D(\modem.instance2.instance3._3_[3] ),
    .Q_N(_1326_),
    .Q(\modem.instance2.instance3._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._4_[4]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net135),
    .D(\modem.instance2.instance3._3_[4] ),
    .Q_N(_0050_),
    .Q(\modem.instance2.instance3._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[0]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net134),
    .D(_0006_),
    .Q_N(_1327_),
    .Q(\modem.instance2._2_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[1]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net135),
    .D(_0007_),
    .Q_N(_1328_),
    .Q(\modem.instance2._2_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[2]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net135),
    .D(_0008_),
    .Q_N(_1329_),
    .Q(\modem.instance2._2_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[3]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net136),
    .D(_0009_),
    .Q_N(_1330_),
    .Q(\modem.instance2._2_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[4]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net135),
    .D(_0010_),
    .Q_N(_1331_),
    .Q(\modem.instance2._2_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance3._5_[5]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net134),
    .D(_0011_),
    .Q_N(_1332_),
    .Q(\modem.instance2._2_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._4_[0]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net130),
    .D(net21),
    .Q_N(_1333_),
    .Q(\modem.instance2.instance4._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._4_[1]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net134),
    .D(\modem.instance2.instance4._3_[1] ),
    .Q_N(_0052_),
    .Q(\modem.instance2.instance4._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._4_[2]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net129),
    .D(\modem.instance2.instance4._3_[2] ),
    .Q_N(_1334_),
    .Q(\modem.instance2.instance4._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._4_[3]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net130),
    .D(\modem.instance2.instance4._3_[3] ),
    .Q_N(_0051_),
    .Q(\modem.instance2.instance4._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._4_[4]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net130),
    .D(\modem.instance2.instance4._3_[4] ),
    .Q_N(_1335_),
    .Q(\modem.instance2.instance4._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[0]$_DFF_PN0_  (.CLK(net84),
    .RESET_B(net134),
    .D(_0012_),
    .Q_N(_1336_),
    .Q(\modem.instance2._3_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[1]$_DFF_PN0_  (.CLK(net84),
    .RESET_B(net133),
    .D(_0013_),
    .Q_N(_1337_),
    .Q(\modem.instance2._3_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[2]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net133),
    .D(_0014_),
    .Q_N(_1338_),
    .Q(\modem.instance2._3_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[3]$_DFF_PN0_  (.CLK(net84),
    .RESET_B(net132),
    .D(_0015_),
    .Q_N(_1339_),
    .Q(\modem.instance2._3_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[4]$_DFF_PN0_  (.CLK(net83),
    .RESET_B(net133),
    .D(_0016_),
    .Q_N(_1340_),
    .Q(\modem.instance2._3_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance4._5_[5]$_DFF_PN0_  (.CLK(net84),
    .RESET_B(net134),
    .D(_0017_),
    .Q_N(_1249_),
    .Q(\modem.instance2._3_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._02_$_DFFE_NN0N_  (.CLK(net90),
    .RESET_B(net115),
    .D(_0067_),
    .Q_N(_1248_),
    .Q(\modem.instance2._4_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[0]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net113),
    .D(\modem.instance2.instance5._09_[0] ),
    .Q_N(_1247_),
    .Q(\modem.instance2.instance5._10_[0] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[10]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[10] ),
    .Q_N(_1246_),
    .Q(\modem.instance2.instance5._10_[10] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[11]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[11] ),
    .Q_N(_1245_),
    .Q(\modem.instance2.instance5._10_[11] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[12]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[12] ),
    .Q_N(_1244_),
    .Q(\modem.instance2.instance5._10_[12] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[13]$_DFF_NN0_  (.CLK(net86),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[13] ),
    .Q_N(_1243_),
    .Q(\modem.instance2.instance5._10_[13] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[14]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[14] ),
    .Q_N(_1242_),
    .Q(\modem.instance2.instance5._10_[14] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[15]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[15] ),
    .Q_N(_1241_),
    .Q(\modem.instance2.instance5._10_[15] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[16]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[16] ),
    .Q_N(_1240_),
    .Q(\modem.instance2.instance5._10_[16] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[17]$_DFF_NN0_  (.CLK(net88),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[17] ),
    .Q_N(_1239_),
    .Q(\modem.instance2.instance5._10_[17] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[18]$_DFF_NN0_  (.CLK(net86),
    .RESET_B(net105),
    .D(\modem.instance2.instance5._09_[18] ),
    .Q_N(_1238_),
    .Q(\modem.instance2.instance5._10_[18] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[19]$_DFF_NN0_  (.CLK(net86),
    .RESET_B(net105),
    .D(\modem.instance2.instance5._09_[19] ),
    .Q_N(_1237_),
    .Q(\modem.instance2.instance5._10_[19] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[1]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net113),
    .D(\modem.instance2.instance5._09_[1] ),
    .Q_N(_1236_),
    .Q(\modem.instance2.instance5._10_[1] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[20]$_DFF_NN0_  (.CLK(net86),
    .RESET_B(net105),
    .D(\modem.instance2.instance5._09_[20] ),
    .Q_N(_1235_),
    .Q(\modem.instance2.instance5._10_[20] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[21]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net105),
    .D(\modem.instance2.instance5._09_[21] ),
    .Q_N(_1234_),
    .Q(\modem.instance2.instance5._10_[21] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[22]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[22] ),
    .Q_N(_1233_),
    .Q(\modem.instance2.instance5._10_[22] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[23]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[23] ),
    .Q_N(_1232_),
    .Q(\modem.instance2.instance5._10_[23] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[24]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[24] ),
    .Q_N(_1231_),
    .Q(\modem.instance2.instance5._10_[24] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[25]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net107),
    .D(\modem.instance2.instance5._09_[25] ),
    .Q_N(_1230_),
    .Q(\modem.instance2.instance5._10_[25] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[26]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net107),
    .D(\modem.instance2.instance5._09_[26] ),
    .Q_N(_1229_),
    .Q(\modem.instance2.instance5._10_[26] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[27]$_DFF_NN0_  (.CLK(net90),
    .RESET_B(net114),
    .D(\modem.instance2.instance5._09_[27] ),
    .Q_N(_1228_),
    .Q(\modem.instance2.instance5._10_[27] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[28]$_DFF_NN0_  (.CLK(net90),
    .RESET_B(net114),
    .D(\modem.instance2.instance5._09_[28] ),
    .Q_N(_1227_),
    .Q(\modem.instance2.instance5._10_[28] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[29]$_DFF_NN0_  (.CLK(net91),
    .RESET_B(net113),
    .D(\modem.instance2.instance5._09_[29] ),
    .Q_N(_1226_),
    .Q(\modem.instance2.instance5._10_[29] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[2]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net102),
    .D(\modem.instance2.instance5._09_[2] ),
    .Q_N(_1225_),
    .Q(\modem.instance2.instance5._10_[2] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[30]$_DFF_NN0_  (.CLK(net91),
    .RESET_B(net113),
    .D(\modem.instance2.instance5._09_[30] ),
    .Q_N(_1224_),
    .Q(\modem.instance2.instance5._10_[30] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[31]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net113),
    .D(\modem.instance2.instance5._09_[31] ),
    .Q_N(_1223_),
    .Q(\modem.instance2.instance5._10_[31] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[3]$_DFF_NN0_  (.CLK(net89),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[3] ),
    .Q_N(_1222_),
    .Q(\modem.instance2.instance5._10_[3] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[4]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net106),
    .D(\modem.instance2.instance5._09_[4] ),
    .Q_N(_1221_),
    .Q(\modem.instance2.instance5._10_[4] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[5]$_DFF_NN0_  (.CLK(net87),
    .RESET_B(net102),
    .D(\modem.instance2.instance5._09_[5] ),
    .Q_N(_1220_),
    .Q(\modem.instance2.instance5._10_[5] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[6]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[6] ),
    .Q_N(_1219_),
    .Q(\modem.instance2.instance5._10_[6] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[7]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[7] ),
    .Q_N(_1218_),
    .Q(\modem.instance2.instance5._10_[7] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[8]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net100),
    .D(\modem.instance2.instance5._09_[8] ),
    .Q_N(_1217_),
    .Q(\modem.instance2.instance5._10_[8] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5._10_[9]$_DFF_NN0_  (.CLK(net85),
    .RESET_B(net104),
    .D(\modem.instance2.instance5._09_[9] ),
    .Q_N(_1216_),
    .Q(\modem.instance2.instance5._10_[9] ));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd0._0_$_DFF_NN1_  (.CLK(net90),
    .RESET_B(net113),
    .D(_1214_),
    .Q_N(\modem.instance2.instance5.ffd0._0_ ),
    .Q(_1469_));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd0._1_$_DFF_N_  (.CLK(net91),
    .RESET_B(net177),
    .D(\modem.instance2.instance5.ffd0._0_ ),
    .Q_N(_1215_),
    .Q(\modem.instance2.instance5._03_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd1._0_$_DFF_NN1_  (.CLK(net90),
    .RESET_B(net113),
    .D(_0061_),
    .Q_N(\modem.instance2.instance5.ffd1._0_ ),
    .Q(_1470_));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd1._1_$_DFF_N_  (.CLK(net90),
    .RESET_B(net178),
    .D(\modem.instance2.instance5.ffd1._0_ ),
    .Q_N(_1214_),
    .Q(\modem.instance2.instance5._00_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd3._0_$_DFF_NN1_  (.CLK(net91),
    .RESET_B(net115),
    .D(_1215_),
    .Q_N(\modem.instance2.instance5.ffd3._0_ ),
    .Q(_1471_));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd3._1_$_DFF_N_  (.CLK(net90),
    .RESET_B(net179),
    .D(\modem.instance2.instance5.ffd3._0_ ),
    .Q_N(_1213_),
    .Q(\modem.instance2.instance5._04_ ));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd4._0_$_DFF_NN1_  (.CLK(net90),
    .RESET_B(net115),
    .D(_1213_),
    .Q_N(\modem.instance2.instance5.ffd4._0_ ),
    .Q(_1472_));
 sg13g2_dfrbp_1 \modem.instance2.instance5.ffd4._1_$_DFF_N_  (.CLK(net91),
    .RESET_B(net180),
    .D(\modem.instance2.instance5.ffd4._0_ ),
    .Q_N(_1212_),
    .Q(\modem.instance2.instance5._05_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._5_$_DFFE_PN0N_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net121),
    .D(_0068_),
    .Q_N(\modem.instance3.instance1._1_ ),
    .Q(\modem.instance3._0_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[0]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net121),
    .D(\modem.instance3.instance1._3_[0] ),
    .Q_N(_1341_),
    .Q(\modem.instance3.instance1._6_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[1]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net121),
    .D(\modem.instance3.instance1._3_[1] ),
    .Q_N(_1342_),
    .Q(\modem.instance3.instance1._6_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[2]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net122),
    .D(\modem.instance3.instance1._3_[2] ),
    .Q_N(_1343_),
    .Q(\modem.instance3.instance1._6_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[3]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net122),
    .D(\modem.instance3.instance1._3_[3] ),
    .Q_N(_1344_),
    .Q(\modem.instance3.instance1._6_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[4]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net122),
    .D(\modem.instance3.instance1._3_[4] ),
    .Q_N(_1345_),
    .Q(\modem.instance3.instance1._6_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[5]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net123),
    .D(\modem.instance3.instance1._3_[5] ),
    .Q_N(_1346_),
    .Q(\modem.instance3.instance1._6_[5] ));
 sg13g2_dfrbp_1 \modem.instance3.instance1._6_[6]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net123),
    .D(\modem.instance3.instance1._3_[6] ),
    .Q_N(_1211_),
    .Q(\modem.instance3.instance1._6_[6] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._02_$_DFFE_NN0N_  (.CLK(net80),
    .RESET_B(net124),
    .D(_0069_),
    .Q_N(_1210_),
    .Q(\modem.instance3._1_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[0]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net107),
    .D(\modem.instance3.instance2._09_[0] ),
    .Q_N(_1209_),
    .Q(\modem.instance3.instance2._10_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[10]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[10] ),
    .Q_N(_1208_),
    .Q(\modem.instance3.instance2._10_[10] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[11]$_DFF_NN0_  (.CLK(net77),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[11] ),
    .Q_N(_1207_),
    .Q(\modem.instance3.instance2._10_[11] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[12]$_DFF_NN0_  (.CLK(net77),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[12] ),
    .Q_N(_1206_),
    .Q(\modem.instance3.instance2._10_[12] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[13]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[13] ),
    .Q_N(_1205_),
    .Q(\modem.instance3.instance2._10_[13] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[14]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[14] ),
    .Q_N(_1204_),
    .Q(\modem.instance3.instance2._10_[14] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[15]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[15] ),
    .Q_N(_1203_),
    .Q(\modem.instance3.instance2._10_[15] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[16]$_DFF_NN0_  (.CLK(net77),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[16] ),
    .Q_N(_1202_),
    .Q(\modem.instance3.instance2._10_[16] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[17]$_DFF_NN0_  (.CLK(net82),
    .RESET_B(net121),
    .D(\modem.instance3.instance2._09_[17] ),
    .Q_N(_1201_),
    .Q(\modem.instance3.instance2._10_[17] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[18]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[18] ),
    .Q_N(_1200_),
    .Q(\modem.instance3.instance2._10_[18] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[19]$_DFF_NN0_  (.CLK(net82),
    .RESET_B(net120),
    .D(\modem.instance3.instance2._09_[19] ),
    .Q_N(_1199_),
    .Q(\modem.instance3.instance2._10_[19] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[1]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[1] ),
    .Q_N(_1198_),
    .Q(\modem.instance3.instance2._10_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[20]$_DFF_NN0_  (.CLK(net82),
    .RESET_B(net120),
    .D(\modem.instance3.instance2._09_[20] ),
    .Q_N(_1197_),
    .Q(\modem.instance3.instance2._10_[20] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[21]$_DFF_NN0_  (.CLK(net82),
    .RESET_B(net121),
    .D(\modem.instance3.instance2._09_[21] ),
    .Q_N(_1196_),
    .Q(\modem.instance3.instance2._10_[21] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[22]$_DFF_NN0_  (.CLK(net82),
    .RESET_B(net121),
    .D(\modem.instance3.instance2._09_[22] ),
    .Q_N(_1195_),
    .Q(\modem.instance3.instance2._10_[22] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[23]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net118),
    .D(\modem.instance3.instance2._09_[23] ),
    .Q_N(_1194_),
    .Q(\modem.instance3.instance2._10_[23] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[24]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net118),
    .D(\modem.instance3.instance2._09_[24] ),
    .Q_N(_1193_),
    .Q(\modem.instance3.instance2._10_[24] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[25]$_DFF_NN0_  (.CLK(net79),
    .RESET_B(net118),
    .D(\modem.instance3.instance2._09_[25] ),
    .Q_N(_1192_),
    .Q(\modem.instance3.instance2._10_[25] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[26]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net118),
    .D(\modem.instance3.instance2._09_[26] ),
    .Q_N(_1191_),
    .Q(\modem.instance3.instance2._10_[26] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[27]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net122),
    .D(\modem.instance3.instance2._09_[27] ),
    .Q_N(_1190_),
    .Q(\modem.instance3.instance2._10_[27] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[28]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net122),
    .D(\modem.instance3.instance2._09_[28] ),
    .Q_N(_1189_),
    .Q(\modem.instance3.instance2._10_[28] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[29]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net122),
    .D(\modem.instance3.instance2._09_[29] ),
    .Q_N(_1188_),
    .Q(\modem.instance3.instance2._10_[29] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[2]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net105),
    .D(\modem.instance3.instance2._09_[2] ),
    .Q_N(_1187_),
    .Q(\modem.instance3.instance2._10_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[30]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net122),
    .D(\modem.instance3.instance2._09_[30] ),
    .Q_N(_1186_),
    .Q(\modem.instance3.instance2._10_[30] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[31]$_DFF_NN0_  (.CLK(net78),
    .RESET_B(net122),
    .D(\modem.instance3.instance2._09_[31] ),
    .Q_N(_1185_),
    .Q(\modem.instance3.instance2._10_[31] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[3]$_DFF_NN0_  (.CLK(net77),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[3] ),
    .Q_N(_1184_),
    .Q(\modem.instance3.instance2._10_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[4]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[4] ),
    .Q_N(_1183_),
    .Q(\modem.instance3.instance2._10_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[5]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[5] ),
    .Q_N(_1182_),
    .Q(\modem.instance3.instance2._10_[5] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[6]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[6] ),
    .Q_N(_1181_),
    .Q(\modem.instance3.instance2._10_[6] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[7]$_DFF_NN0_  (.CLK(net76),
    .RESET_B(net117),
    .D(\modem.instance3.instance2._09_[7] ),
    .Q_N(_1180_),
    .Q(\modem.instance3.instance2._10_[7] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[8]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[8] ),
    .Q_N(_1179_),
    .Q(\modem.instance3.instance2._10_[8] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2._10_[9]$_DFF_NN0_  (.CLK(net81),
    .RESET_B(net119),
    .D(\modem.instance3.instance2._09_[9] ),
    .Q_N(_1178_),
    .Q(\modem.instance3.instance2._10_[9] ));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd0._0_$_DFF_NN1_  (.CLK(net80),
    .RESET_B(net124),
    .D(_1175_),
    .Q_N(\modem.instance3.instance2.ffd0._0_ ),
    .Q(_1473_));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd0._1_$_DFF_N_  (.CLK(net80),
    .RESET_B(net181),
    .D(\modem.instance3.instance2.ffd0._0_ ),
    .Q_N(_1177_),
    .Q(\modem.instance3.instance2._04_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd1._0_$_DFF_NN1_  (.CLK(net80),
    .RESET_B(net114),
    .D(_0062_),
    .Q_N(\modem.instance3.instance2.ffd1._0_ ),
    .Q(_1474_));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd1._1_$_DFF_N_  (.CLK(net80),
    .RESET_B(net182),
    .D(\modem.instance3.instance2.ffd1._0_ ),
    .Q_N(_1176_),
    .Q(\modem.instance3.instance2._00_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd2._0_$_DFF_NN1_  (.CLK(net80),
    .RESET_B(net114),
    .D(_1176_),
    .Q_N(\modem.instance3.instance2.ffd2._0_ ),
    .Q(_1475_));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd2._1_$_DFF_N_  (.CLK(net80),
    .RESET_B(net183),
    .D(\modem.instance3.instance2.ffd2._0_ ),
    .Q_N(_1175_),
    .Q(\modem.instance3.instance2._03_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd4._0_$_DFF_NN1_  (.CLK(net81),
    .RESET_B(net124),
    .D(_1177_),
    .Q_N(\modem.instance3.instance2.ffd4._0_ ),
    .Q(_1476_));
 sg13g2_dfrbp_1 \modem.instance3.instance2.ffd4._1_$_DFF_N_  (.CLK(net80),
    .RESET_B(net184),
    .D(\modem.instance3.instance2.ffd4._0_ ),
    .Q_N(_1347_),
    .Q(\modem.instance3.instance2._05_ ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._4_[0]$_DFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net124),
    .D(\modem.instance3.instance3._3_[0] ),
    .Q_N(_1348_),
    .Q(\modem.instance3.instance3._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._4_[1]$_DFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net124),
    .D(\modem.instance3.instance3._3_[1] ),
    .Q_N(_0058_),
    .Q(\modem.instance3.instance3._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._4_[2]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net124),
    .D(\modem.instance3.instance3._3_[2] ),
    .Q_N(_1349_),
    .Q(\modem.instance3.instance3._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._4_[3]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net124),
    .D(\modem.instance3.instance3._3_[3] ),
    .Q_N(_1350_),
    .Q(\modem.instance3.instance3._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._4_[4]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net124),
    .D(\modem.instance3.instance3._3_[4] ),
    .Q_N(_1351_),
    .Q(\modem.instance3.instance3._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[0]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0018_),
    .Q_N(_1352_),
    .Q(\modem.instance3._2_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[1]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0019_),
    .Q_N(_1353_),
    .Q(\modem.instance3._2_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[2]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net140),
    .D(_0020_),
    .Q_N(_1354_),
    .Q(\modem.instance3._2_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[3]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net141),
    .D(_0021_),
    .Q_N(_1355_),
    .Q(\modem.instance3._2_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[4]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net141),
    .D(_0022_),
    .Q_N(_1356_),
    .Q(\modem.instance3._2_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance3._5_[5]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net127),
    .D(_0023_),
    .Q_N(_1357_),
    .Q(\modem.instance3._2_[5] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._4_[0]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net115),
    .D(\modem.instance3.instance4._3_[0] ),
    .Q_N(_0056_),
    .Q(\modem.instance3.instance4._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._4_[1]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net131),
    .D(\modem.instance3.instance4._3_[1] ),
    .Q_N(_0055_),
    .Q(\modem.instance3.instance4._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._4_[2]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net115),
    .D(\modem.instance3.instance4._3_[2] ),
    .Q_N(_0057_),
    .Q(\modem.instance3.instance4._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._4_[3]$_DFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net114),
    .D(\modem.instance3.instance4._3_[3] ),
    .Q_N(_1358_),
    .Q(\modem.instance3.instance4._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._4_[4]$_DFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net127),
    .D(\modem.instance3.instance4._3_[4] ),
    .Q_N(_1359_),
    .Q(\modem.instance3.instance4._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[0]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0024_),
    .Q_N(_1360_),
    .Q(\modem.instance3._3_[0] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[1]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net140),
    .D(_0025_),
    .Q_N(_1361_),
    .Q(\modem.instance3._3_[1] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[2]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0026_),
    .Q_N(_1362_),
    .Q(\modem.instance3._3_[2] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[3]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0027_),
    .Q_N(_1363_),
    .Q(\modem.instance3._3_[3] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[4]$_DFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net140),
    .D(_0028_),
    .Q_N(_1364_),
    .Q(\modem.instance3._3_[4] ));
 sg13g2_dfrbp_1 \modem.instance3.instance4._5_[5]$_DFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net127),
    .D(_0029_),
    .Q_N(_1365_),
    .Q(\modem.instance3._3_[5] ));
 sg13g2_dfrbp_1 \modem.instance4._6_[0]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[0] ),
    .Q_N(_1366_),
    .Q(net2));
 sg13g2_dfrbp_1 \modem.instance4._6_[1]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[1] ),
    .Q_N(_1367_),
    .Q(net3));
 sg13g2_dfrbp_1 \modem.instance4._6_[2]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[2] ),
    .Q_N(_1368_),
    .Q(net4));
 sg13g2_dfrbp_1 \modem.instance4._6_[3]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[3] ),
    .Q_N(_1369_),
    .Q(net5));
 sg13g2_dfrbp_1 \modem.instance4._6_[4]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[4] ),
    .Q_N(_1370_),
    .Q(net6));
 sg13g2_dfrbp_1 \modem.instance4._6_[5]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance4._5_[5] ),
    .Q_N(_1371_),
    .Q(net7));
 sg13g2_dfrbp_1 \modem.instance6._2_$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net150),
    .D(\modem.instance6._1_ ),
    .Q_N(_1372_),
    .Q(\modem._4_ ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._4_[0]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net137),
    .D(\modem.instance7.instance2._3_[0] ),
    .Q_N(_1373_),
    .Q(\modem.instance7.instance2._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._4_[1]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net136),
    .D(\modem.instance7.instance2._3_[1] ),
    .Q_N(_0054_),
    .Q(\modem.instance7.instance2._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._4_[2]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(\modem.instance7.instance2._3_[2] ),
    .Q_N(_1374_),
    .Q(\modem.instance7.instance2._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._4_[3]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net137),
    .D(\modem.instance7.instance2._3_[3] ),
    .Q_N(_1375_),
    .Q(\modem.instance7.instance2._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._4_[4]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(\modem.instance7.instance2._3_[4] ),
    .Q_N(_0046_),
    .Q(\modem.instance7.instance2._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[0]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(_0030_),
    .Q_N(_1376_),
    .Q(\modem.instance7._0_[0] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[1]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(_0031_),
    .Q_N(_1377_),
    .Q(\modem.instance7._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[2]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(_0032_),
    .Q_N(_1378_),
    .Q(\modem.instance7._0_[2] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[3]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net136),
    .D(_0033_),
    .Q_N(_1379_),
    .Q(\modem.instance7._0_[3] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[4]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(_0034_),
    .Q_N(_1380_),
    .Q(\modem.instance7._0_[4] ));
 sg13g2_dfrbp_1 \modem.instance7.instance2._5_[5]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(_0035_),
    .Q_N(_1381_),
    .Q(\modem.instance7._0_[5] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[0]$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net150),
    .D(\modem.instance7.instance3._0_[0] ),
    .Q_N(_1382_),
    .Q(\modem.instance7._1_[0] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[1]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance7.instance3._0_[1] ),
    .Q_N(_1383_),
    .Q(\modem.instance7._1_[1] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[2]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(\modem.instance7.instance3._0_[2] ),
    .Q_N(_1384_),
    .Q(\modem.instance7._1_[2] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[3]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net138),
    .D(\modem.instance7.instance3._0_[3] ),
    .Q_N(_1385_),
    .Q(\modem.instance7._1_[3] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[4]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net137),
    .D(\modem.instance7.instance3._0_[4] ),
    .Q_N(_1386_),
    .Q(\modem.instance7._1_[4] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[5]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net138),
    .D(\modem.instance7.instance3._0_[5] ),
    .Q_N(_1387_),
    .Q(\modem.instance7._1_[5] ));
 sg13g2_dfrbp_1 \modem.instance7.instance3._1_[6]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net142),
    .D(net185),
    .Q_N(_0043_),
    .Q(\modem.instance7._1_[6] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._1_$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net149),
    .D(\modem.instance7.instance4._7_ ),
    .Q_N(_1388_),
    .Q(\modem._5_ ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[0]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[0] ),
    .Q_N(_0048_),
    .Q(\modem.instance7.instance4._9_[0] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[10]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net150),
    .D(\modem.instance7.instance4._8_[10] ),
    .Q_N(_1389_),
    .Q(\modem.instance7.instance4._9_[10] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[11]$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[11] ),
    .Q_N(_1390_),
    .Q(\modem.instance7.instance4._9_[11] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[12]$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[12] ),
    .Q_N(_1391_),
    .Q(\modem.instance7.instance4._9_[12] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[13]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[13] ),
    .Q_N(_1392_),
    .Q(\modem.instance7.instance4._9_[13] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[14]$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net150),
    .D(\modem.instance7.instance4._8_[14] ),
    .Q_N(_1393_),
    .Q(\modem.instance7.instance4._9_[14] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[15]$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[15] ),
    .Q_N(_1394_),
    .Q(\modem.instance7.instance4._9_[15] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[16]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[16] ),
    .Q_N(_1395_),
    .Q(\modem.instance7.instance4._9_[16] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[17]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[17] ),
    .Q_N(_1396_),
    .Q(\modem.instance7.instance4._9_[17] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[18]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance7.instance4._8_[18] ),
    .Q_N(_1397_),
    .Q(\modem.instance7.instance4._9_[18] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[19]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net147),
    .D(\modem.instance7.instance4._8_[19] ),
    .Q_N(_1398_),
    .Q(\modem.instance7.instance4._9_[19] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[1]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[1] ),
    .Q_N(_1399_),
    .Q(\modem.instance7.instance4._9_[1] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[20]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[20] ),
    .Q_N(_1400_),
    .Q(\modem.instance7.instance4._9_[20] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[21]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[21] ),
    .Q_N(_1401_),
    .Q(\modem.instance7.instance4._9_[21] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[22]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[22] ),
    .Q_N(_1402_),
    .Q(\modem.instance7.instance4._9_[22] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[23]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[23] ),
    .Q_N(_1403_),
    .Q(\modem.instance7.instance4._9_[23] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[24]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net153),
    .D(\modem.instance7.instance4._8_[24] ),
    .Q_N(_1404_),
    .Q(\modem.instance7.instance4._9_[24] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[25]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[25] ),
    .Q_N(_1405_),
    .Q(\modem.instance7.instance4._9_[25] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[26]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[26] ),
    .Q_N(_1406_),
    .Q(\modem.instance7.instance4._9_[26] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[27]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[27] ),
    .Q_N(_1407_),
    .Q(\modem.instance7.instance4._9_[27] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[28]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[28] ),
    .Q_N(_1408_),
    .Q(\modem.instance7.instance4._9_[28] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[29]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[29] ),
    .Q_N(_1409_),
    .Q(\modem.instance7.instance4._9_[29] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[2]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[2] ),
    .Q_N(_1410_),
    .Q(\modem.instance7.instance4._9_[2] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[30]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(\modem.instance7.instance4._8_[30] ),
    .Q_N(_1411_),
    .Q(\modem.instance7.instance4._9_[30] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[31]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[31] ),
    .Q_N(_0049_),
    .Q(\modem.instance7.instance4._9_[31] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[3]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[3] ),
    .Q_N(_1412_),
    .Q(\modem.instance7.instance4._9_[3] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[4]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[4] ),
    .Q_N(_1413_),
    .Q(\modem.instance7.instance4._9_[4] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[5]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[5] ),
    .Q_N(_1414_),
    .Q(\modem.instance7.instance4._9_[5] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[6]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[6] ),
    .Q_N(_1415_),
    .Q(\modem.instance7.instance4._9_[6] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[7]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[7] ),
    .Q_N(_1416_),
    .Q(\modem.instance7.instance4._9_[7] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[8]$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net151),
    .D(\modem.instance7.instance4._8_[8] ),
    .Q_N(_1417_),
    .Q(\modem.instance7.instance4._9_[8] ));
 sg13g2_dfrbp_1 \modem.instance7.instance4._9_[9]$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net150),
    .D(\modem.instance7.instance4._8_[9] ),
    .Q_N(_1418_),
    .Q(\modem.instance7.instance4._9_[9] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._4_[0]$_DFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net149),
    .D(\modem.instance8.instance2._3_[0] ),
    .Q_N(_1419_),
    .Q(\modem.instance8.instance2._4_[0] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._4_[1]$_DFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(\modem.instance8.instance2._3_[1] ),
    .Q_N(_0053_),
    .Q(\modem.instance8.instance2._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._4_[2]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net149),
    .D(\modem.instance8.instance2._3_[2] ),
    .Q_N(_1420_),
    .Q(\modem.instance8.instance2._4_[2] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._4_[3]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net149),
    .D(\modem.instance8.instance2._3_[3] ),
    .Q_N(_1421_),
    .Q(\modem.instance8.instance2._4_[3] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._4_[4]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net149),
    .D(\modem.instance8.instance2._3_[4] ),
    .Q_N(_0042_),
    .Q(\modem.instance8.instance2._4_[4] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[0]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(_0036_),
    .Q_N(_1422_),
    .Q(\modem.instance8._0_[0] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[1]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net141),
    .D(_0037_),
    .Q_N(_1423_),
    .Q(\modem.instance8._0_[1] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[2]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net143),
    .D(_0038_),
    .Q_N(_1424_),
    .Q(\modem.instance8._0_[2] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[3]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net142),
    .D(_0039_),
    .Q_N(_1425_),
    .Q(\modem.instance8._0_[3] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[4]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net142),
    .D(_0040_),
    .Q_N(_1426_),
    .Q(\modem.instance8._0_[4] ));
 sg13g2_dfrbp_1 \modem.instance8.instance2._5_[5]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net142),
    .D(_0041_),
    .Q_N(_1427_),
    .Q(\modem.instance8._0_[5] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[0]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[0] ),
    .Q_N(_1428_),
    .Q(\modem.instance8._1_[0] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[1]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[1] ),
    .Q_N(_1429_),
    .Q(\modem.instance8._1_[1] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[2]$_DFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[2] ),
    .Q_N(_1430_),
    .Q(\modem.instance8._1_[2] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[3]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[3] ),
    .Q_N(_1431_),
    .Q(\modem.instance8._1_[3] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[4]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[4] ),
    .Q_N(_1432_),
    .Q(\modem.instance8._1_[4] ));
 sg13g2_dfrbp_1 \modem.instance8.instance3._1_[5]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net143),
    .D(\modem.instance8.instance3._0_[5] ),
    .Q_N(_1433_),
    .Q(\modem.instance8._1_[5] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._1_$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net141),
    .D(\modem.instance8.instance5._7_ ),
    .Q_N(_1434_),
    .Q(\modem._6_ ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[0]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[0] ),
    .Q_N(_0044_),
    .Q(\modem.instance8.instance5._9_[0] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[10]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[10] ),
    .Q_N(_1435_),
    .Q(\modem.instance8.instance5._9_[10] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[11]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net121),
    .D(\modem.instance8.instance5._8_[11] ),
    .Q_N(_1436_),
    .Q(\modem.instance8.instance5._9_[11] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[12]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[12] ),
    .Q_N(_1437_),
    .Q(\modem.instance8.instance5._9_[12] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[13]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[13] ),
    .Q_N(_1438_),
    .Q(\modem.instance8.instance5._9_[13] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[14]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net121),
    .D(\modem.instance8.instance5._8_[14] ),
    .Q_N(_1439_),
    .Q(\modem.instance8.instance5._9_[14] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[15]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net123),
    .D(\modem.instance8.instance5._8_[15] ),
    .Q_N(_1440_),
    .Q(\modem.instance8.instance5._9_[15] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[16]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[16] ),
    .Q_N(_1441_),
    .Q(\modem.instance8.instance5._9_[16] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[17]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[17] ),
    .Q_N(_1442_),
    .Q(\modem.instance8.instance5._9_[17] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[18]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[18] ),
    .Q_N(_1443_),
    .Q(\modem.instance8.instance5._9_[18] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[19]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[19] ),
    .Q_N(_1444_),
    .Q(\modem.instance8.instance5._9_[19] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[1]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[1] ),
    .Q_N(_1445_),
    .Q(\modem.instance8.instance5._9_[1] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[20]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net126),
    .D(\modem.instance8.instance5._8_[20] ),
    .Q_N(_1446_),
    .Q(\modem.instance8.instance5._9_[20] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[21]$_DFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[21] ),
    .Q_N(_1447_),
    .Q(\modem.instance8.instance5._9_[21] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[22]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[22] ),
    .Q_N(_1448_),
    .Q(\modem.instance8.instance5._9_[22] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[23]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[23] ),
    .Q_N(_1449_),
    .Q(\modem.instance8.instance5._9_[23] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[24]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net127),
    .D(\modem.instance8.instance5._8_[24] ),
    .Q_N(_1450_),
    .Q(\modem.instance8.instance5._9_[24] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[25]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net147),
    .D(\modem.instance8.instance5._8_[25] ),
    .Q_N(_1451_),
    .Q(\modem.instance8.instance5._9_[25] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[26]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[26] ),
    .Q_N(_1452_),
    .Q(\modem.instance8.instance5._9_[26] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[27]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[27] ),
    .Q_N(_1453_),
    .Q(\modem.instance8.instance5._9_[27] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[28]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net147),
    .D(\modem.instance8.instance5._8_[28] ),
    .Q_N(_1454_),
    .Q(\modem.instance8.instance5._9_[28] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[29]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net147),
    .D(\modem.instance8.instance5._8_[29] ),
    .Q_N(_1455_),
    .Q(\modem.instance8.instance5._9_[29] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[2]$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[2] ),
    .Q_N(_1456_),
    .Q(\modem.instance8.instance5._9_[2] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[30]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance8.instance5._8_[30] ),
    .Q_N(_1457_),
    .Q(\modem.instance8.instance5._9_[30] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[31]$_DFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[31] ),
    .Q_N(_0045_),
    .Q(\modem.instance8.instance5._9_[31] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[3]$_DFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net146),
    .D(\modem.instance8.instance5._8_[3] ),
    .Q_N(_1458_),
    .Q(\modem.instance8.instance5._9_[3] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[4]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[4] ),
    .Q_N(_1459_),
    .Q(\modem.instance8.instance5._9_[4] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[5]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[5] ),
    .Q_N(_1460_),
    .Q(\modem.instance8.instance5._9_[5] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[6]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[6] ),
    .Q_N(_1461_),
    .Q(\modem.instance8.instance5._9_[6] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[7]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(\modem.instance8.instance5._8_[7] ),
    .Q_N(_1462_),
    .Q(\modem.instance8.instance5._9_[7] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[8]$_DFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[8] ),
    .Q_N(_1463_),
    .Q(\modem.instance8.instance5._9_[8] ));
 sg13g2_dfrbp_1 \modem.instance8.instance5._9_[9]$_DFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net125),
    .D(\modem.instance8.instance5._8_[9] ),
    .Q_N(_1464_),
    .Q(\modem.instance8.instance5._9_[9] ));
 sg13g2_dfrbp_1 \modem.instance9._6_$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net138),
    .D(\modem.instance9._5_ ),
    .Q_N(_1174_),
    .Q(demod_out));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout9 (.A(_0437_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_0340_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0800_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0771_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0738_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0743_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0681_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0649_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0634_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0613_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0637_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1057_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(\modem.instance2.instance4._3_[0] ),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0847_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0846_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0842_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0840_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0838_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0836_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0832_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0263_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0192_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0190_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0168_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0166_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(\modem.instance1.instance3._3_[0] ),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0115_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0110_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0105_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0097_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1158_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1156_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1139_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1133_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1131_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1083_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1075_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1068_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1050_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1048_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1044_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1001_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0999_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0977_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0975_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0932_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0930_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0908_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0906_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0831_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0280_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0253_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0173_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0171_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0111_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0107_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0102_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1137_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1132_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1055_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1047_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1045_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1043_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0982_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0980_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0913_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0911_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net79),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net79),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net79),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(\modem.instance3.instance1._1_ ),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net82),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(\modem.instance3.instance1._1_ ),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(\modem.instance2._1_ ),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(\modem.instance2._1_ ),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(net88),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net88),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(\modem.instance2.instance1._1_ ),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net91),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(\modem.instance2.instance1._1_ ),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net95),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(\modem.instance1.instance1._1_ ),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(\modem.instance1.instance1._1_ ),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(\modem.instance1.instance1._1_ ),
    .X(net98));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net103));
 sg13g2_buf_2 fanout100 (.A(net103),
    .X(net100));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net103));
 sg13g2_buf_2 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(net116),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net107));
 sg13g2_buf_2 fanout105 (.A(net107),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net107));
 sg13g2_buf_2 fanout107 (.A(net116),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net112));
 sg13g2_buf_2 fanout109 (.A(net112),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net112));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(net116),
    .X(net112));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(net115));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net116));
 sg13g2_buf_1 fanout116 (.A(net155),
    .X(net116));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net120));
 sg13g2_buf_2 fanout118 (.A(net120),
    .X(net118));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(net120));
 sg13g2_buf_2 fanout120 (.A(net128),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net123));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net128));
 sg13g2_buf_2 fanout123 (.A(net128),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net127));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(net126));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(net127));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net155),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net130));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net133));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net133));
 sg13g2_buf_2 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net139),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net139));
 sg13g2_buf_2 fanout135 (.A(net139),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net138));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net138));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net155),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net144));
 sg13g2_buf_2 fanout141 (.A(net144),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net144));
 sg13g2_buf_1 fanout144 (.A(net154),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net147));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net147));
 sg13g2_buf_2 fanout147 (.A(net154),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net150));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net154));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net154));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(net153));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net154));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net1),
    .X(net155));
 sg13g2_tielo _2888__156 (.L_LO(net156));
 sg13g2_tielo _2889__157 (.L_LO(net157));
 sg13g2_tielo _2890__158 (.L_LO(net158));
 sg13g2_tielo _2891__159 (.L_LO(net159));
 sg13g2_tielo _2892__160 (.L_LO(net160));
 sg13g2_tielo _2893__161 (.L_LO(net161));
 sg13g2_tielo _2894__162 (.L_LO(net162));
 sg13g2_tielo _2895__163 (.L_LO(net163));
 sg13g2_tielo _2896__164 (.L_LO(net164));
 sg13g2_tielo _2897__165 (.L_LO(net165));
 sg13g2_tielo _2898__166 (.L_LO(net166));
 sg13g2_tielo _2899__167 (.L_LO(net167));
 sg13g2_tielo _2900__168 (.L_LO(net168));
 sg13g2_tielo _2901__169 (.L_LO(net169));
 sg13g2_tielo _2902__170 (.L_LO(net170));
 sg13g2_tielo _2903__171 (.L_LO(net171));
 sg13g2_tielo _2904__172 (.L_LO(net172));
 sg13g2_tiehi \modem.instance1.instance2.ffd2._1_$_DFF_N__174  (.L_HI(net174));
 sg13g2_tiehi \modem.instance1.instance2.ffd3._1_$_DFF_N__175  (.L_HI(net175));
 sg13g2_tiehi \modem.instance1.instance2.ffd4._1_$_DFF_N__176  (.L_HI(net176));
 sg13g2_tiehi \modem.instance2.instance5.ffd0._1_$_DFF_N__177  (.L_HI(net177));
 sg13g2_tiehi \modem.instance2.instance5.ffd1._1_$_DFF_N__178  (.L_HI(net178));
 sg13g2_tiehi \modem.instance2.instance5.ffd3._1_$_DFF_N__179  (.L_HI(net179));
 sg13g2_tiehi \modem.instance2.instance5.ffd4._1_$_DFF_N__180  (.L_HI(net180));
 sg13g2_tiehi \modem.instance3.instance2.ffd0._1_$_DFF_N__181  (.L_HI(net181));
 sg13g2_tiehi \modem.instance3.instance2.ffd1._1_$_DFF_N__182  (.L_HI(net182));
 sg13g2_tiehi \modem.instance3.instance2.ffd2._1_$_DFF_N__183  (.L_HI(net183));
 sg13g2_tiehi \modem.instance3.instance2.ffd4._1_$_DFF_N__184  (.L_HI(net184));
 sg13g2_tiehi \modem.instance7.instance3._1_[6]$_DFF_PN0__185  (.L_HI(net185));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_4 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_decap_4 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_decap_8 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_decap_8 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_265 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_12_419 ();
 sg13g2_decap_4 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_4 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_decap_8 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_13_414 ();
 sg13g2_decap_8 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_4 FILLER_14_285 ();
 sg13g2_fill_1 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_4 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_decap_4 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_411 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_33 ();
 sg13g2_decap_8 FILLER_16_66 ();
 sg13g2_decap_8 FILLER_16_73 ();
 sg13g2_decap_4 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_148 ();
 sg13g2_decap_8 FILLER_16_155 ();
 sg13g2_decap_4 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_2 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_17 ();
 sg13g2_decap_4 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_decap_8 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_decap_4 FILLER_17_163 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_4 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_8 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_decap_8 FILLER_18_36 ();
 sg13g2_decap_8 FILLER_18_43 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_decap_4 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_106 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_4 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_16 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_106 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_decap_4 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_decap_4 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_78 ();
 sg13g2_decap_8 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_decap_4 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_57 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_122 ();
 sg13g2_decap_4 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_4 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_285 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_85 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_decap_8 FILLER_22_124 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_8 FILLER_22_153 ();
 sg13g2_decap_4 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_217 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_4 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_decap_8 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_31 ();
 sg13g2_decap_4 FILLER_23_38 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_56 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_decap_4 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_8 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_decap_8 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_4 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_decap_8 FILLER_24_106 ();
 sg13g2_decap_4 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_decap_4 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_24_414 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_51 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_4 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_4 FILLER_26_32 ();
 sg13g2_fill_1 FILLER_26_41 ();
 sg13g2_decap_4 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_2 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_206 ();
 sg13g2_fill_2 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_decap_4 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_decap_4 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_33 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_decap_8 FILLER_27_80 ();
 sg13g2_decap_8 FILLER_27_87 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_decap_4 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_127 ();
 sg13g2_decap_4 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_97 ();
 sg13g2_decap_8 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_4 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_decap_4 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_134 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_decap_8 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_decap_4 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_4 FILLER_29_283 ();
 sg13g2_fill_2 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_318 ();
 sg13g2_decap_4 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_4 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_8 ();
 sg13g2_decap_8 FILLER_30_15 ();
 sg13g2_decap_8 FILLER_30_22 ();
 sg13g2_decap_8 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_decap_8 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_decap_8 FILLER_30_239 ();
 sg13g2_decap_8 FILLER_30_246 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_324 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_decap_8 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_30_414 ();
 sg13g2_decap_8 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_4 FILLER_31_30 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_93 ();
 sg13g2_decap_8 FILLER_31_100 ();
 sg13g2_decap_4 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_decap_8 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_143 ();
 sg13g2_decap_4 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_178 ();
 sg13g2_decap_8 FILLER_32_185 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_32_412 ();
 sg13g2_decap_8 FILLER_32_419 ();
 sg13g2_decap_4 FILLER_32_426 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_decap_8 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_decap_4 FILLER_33_72 ();
 sg13g2_fill_2 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_decap_4 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_decap_8 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_33_414 ();
 sg13g2_decap_8 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_15 ();
 sg13g2_fill_2 FILLER_34_22 ();
 sg13g2_decap_8 FILLER_34_30 ();
 sg13g2_decap_4 FILLER_34_45 ();
 sg13g2_decap_4 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_decap_4 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_34_404 ();
 sg13g2_decap_8 FILLER_34_411 ();
 sg13g2_decap_8 FILLER_34_418 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_decap_8 FILLER_35_64 ();
 sg13g2_decap_4 FILLER_35_71 ();
 sg13g2_fill_2 FILLER_35_75 ();
 sg13g2_decap_8 FILLER_35_139 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_423 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_37 ();
 sg13g2_decap_8 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_53 ();
 sg13g2_decap_4 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_128 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_4 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_404 ();
 sg13g2_decap_8 FILLER_36_411 ();
 sg13g2_decap_8 FILLER_36_418 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_9 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_4 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_4 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_4 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_decap_4 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_1 FILLER_38_149 ();
 sg13g2_decap_4 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_decap_4 FILLER_38_213 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_4 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_352 ();
 sg13g2_fill_2 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_2 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_4 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_33 ();
 sg13g2_decap_8 FILLER_39_40 ();
 sg13g2_fill_1 FILLER_39_47 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_decap_8 FILLER_39_67 ();
 sg13g2_decap_4 FILLER_39_74 ();
 sg13g2_decap_8 FILLER_39_150 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_195 ();
 sg13g2_decap_4 FILLER_39_202 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_decap_4 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_229 ();
 sg13g2_fill_2 FILLER_39_236 ();
 sg13g2_decap_8 FILLER_39_242 ();
 sg13g2_decap_8 FILLER_39_249 ();
 sg13g2_fill_2 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_282 ();
 sg13g2_decap_4 FILLER_39_287 ();
 sg13g2_fill_2 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_54 ();
 sg13g2_fill_2 FILLER_40_61 ();
 sg13g2_decap_8 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_104 ();
 sg13g2_decap_4 FILLER_40_111 ();
 sg13g2_decap_4 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_123 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_decap_8 FILLER_40_177 ();
 sg13g2_decap_4 FILLER_40_184 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_decap_8 FILLER_40_234 ();
 sg13g2_decap_8 FILLER_40_241 ();
 sg13g2_decap_8 FILLER_40_248 ();
 sg13g2_decap_8 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_262 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_decap_4 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_313 ();
 sg13g2_decap_8 FILLER_40_320 ();
 sg13g2_decap_4 FILLER_40_327 ();
 sg13g2_fill_1 FILLER_40_331 ();
 sg13g2_fill_2 FILLER_40_336 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_365 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_422 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_fill_1 FILLER_41_30 ();
 sg13g2_fill_2 FILLER_41_57 ();
 sg13g2_fill_1 FILLER_41_59 ();
 sg13g2_decap_8 FILLER_41_64 ();
 sg13g2_decap_8 FILLER_41_71 ();
 sg13g2_decap_8 FILLER_41_78 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_decap_8 FILLER_41_99 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_decap_8 FILLER_41_120 ();
 sg13g2_decap_8 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_decap_4 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_209 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_233 ();
 sg13g2_decap_8 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_decap_4 FILLER_41_261 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_2 FILLER_41_293 ();
 sg13g2_decap_8 FILLER_41_310 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_decap_4 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_342 ();
 sg13g2_decap_8 FILLER_41_354 ();
 sg13g2_decap_8 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_368 ();
 sg13g2_fill_2 FILLER_41_375 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_8 FILLER_41_404 ();
 sg13g2_decap_8 FILLER_41_411 ();
 sg13g2_decap_8 FILLER_41_418 ();
 sg13g2_decap_4 FILLER_41_425 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_128 ();
 sg13g2_fill_1 FILLER_42_139 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_fill_2 FILLER_42_150 ();
 sg13g2_decap_4 FILLER_42_160 ();
 sg13g2_fill_2 FILLER_42_164 ();
 sg13g2_fill_2 FILLER_42_228 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_decap_4 FILLER_42_264 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_300 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_decap_8 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_fill_2 FILLER_42_374 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_decap_8 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_decap_4 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_37 ();
 sg13g2_decap_4 FILLER_43_44 ();
 sg13g2_fill_1 FILLER_43_48 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_4 FILLER_43_175 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_196 ();
 sg13g2_fill_1 FILLER_43_202 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_2 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_268 ();
 sg13g2_fill_1 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_306 ();
 sg13g2_decap_4 FILLER_43_315 ();
 sg13g2_fill_2 FILLER_43_319 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_fill_2 FILLER_43_340 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_369 ();
 sg13g2_fill_2 FILLER_43_396 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_decap_8 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_410 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_decap_4 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_4 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_decap_8 FILLER_44_25 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_65 ();
 sg13g2_fill_1 FILLER_44_72 ();
 sg13g2_fill_2 FILLER_44_118 ();
 sg13g2_decap_4 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_132 ();
 sg13g2_decap_8 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_1 FILLER_44_162 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_4 FILLER_44_245 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_decap_4 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_264 ();
 sg13g2_fill_2 FILLER_44_300 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_fill_2 FILLER_44_315 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_decap_4 FILLER_44_376 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_decap_4 FILLER_45_45 ();
 sg13g2_decap_4 FILLER_45_66 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_decap_8 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_128 ();
 sg13g2_decap_8 FILLER_45_135 ();
 sg13g2_fill_2 FILLER_45_142 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_fill_2 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_198 ();
 sg13g2_decap_8 FILLER_45_229 ();
 sg13g2_decap_8 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_decap_8 FILLER_45_302 ();
 sg13g2_decap_8 FILLER_45_309 ();
 sg13g2_decap_8 FILLER_45_316 ();
 sg13g2_fill_1 FILLER_45_323 ();
 sg13g2_decap_4 FILLER_45_336 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_decap_4 FILLER_45_360 ();
 sg13g2_fill_2 FILLER_45_364 ();
 sg13g2_fill_2 FILLER_45_371 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_399 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_36 ();
 sg13g2_decap_8 FILLER_46_43 ();
 sg13g2_fill_2 FILLER_46_50 ();
 sg13g2_decap_8 FILLER_46_65 ();
 sg13g2_decap_8 FILLER_46_72 ();
 sg13g2_decap_4 FILLER_46_79 ();
 sg13g2_fill_2 FILLER_46_83 ();
 sg13g2_decap_4 FILLER_46_111 ();
 sg13g2_fill_2 FILLER_46_115 ();
 sg13g2_decap_8 FILLER_46_148 ();
 sg13g2_decap_8 FILLER_46_155 ();
 sg13g2_decap_8 FILLER_46_162 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_decap_8 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_2 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_201 ();
 sg13g2_fill_2 FILLER_46_208 ();
 sg13g2_decap_4 FILLER_46_234 ();
 sg13g2_fill_1 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_265 ();
 sg13g2_decap_4 FILLER_46_272 ();
 sg13g2_fill_1 FILLER_46_276 ();
 sg13g2_decap_8 FILLER_46_303 ();
 sg13g2_decap_8 FILLER_46_310 ();
 sg13g2_decap_4 FILLER_46_317 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_4 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_355 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_387 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_8 FILLER_46_403 ();
 sg13g2_decap_8 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_decap_8 FILLER_47_19 ();
 sg13g2_decap_8 FILLER_47_26 ();
 sg13g2_decap_8 FILLER_47_33 ();
 sg13g2_fill_2 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_fill_2 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_2 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_fill_1 FILLER_47_215 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_281 ();
 sg13g2_decap_8 FILLER_47_288 ();
 sg13g2_decap_8 FILLER_47_295 ();
 sg13g2_decap_8 FILLER_47_302 ();
 sg13g2_decap_8 FILLER_47_309 ();
 sg13g2_fill_2 FILLER_47_316 ();
 sg13g2_decap_4 FILLER_47_344 ();
 sg13g2_fill_1 FILLER_47_348 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_fill_2 FILLER_47_364 ();
 sg13g2_fill_2 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_9 ();
 sg13g2_fill_2 FILLER_48_27 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_4 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_109 ();
 sg13g2_decap_8 FILLER_48_114 ();
 sg13g2_decap_8 FILLER_48_121 ();
 sg13g2_decap_8 FILLER_48_128 ();
 sg13g2_decap_4 FILLER_48_135 ();
 sg13g2_fill_1 FILLER_48_149 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_4 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_fill_1 FILLER_48_177 ();
 sg13g2_decap_4 FILLER_48_182 ();
 sg13g2_fill_1 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_237 ();
 sg13g2_fill_2 FILLER_48_265 ();
 sg13g2_decap_8 FILLER_48_303 ();
 sg13g2_decap_8 FILLER_48_310 ();
 sg13g2_decap_4 FILLER_48_317 ();
 sg13g2_fill_1 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_337 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_decap_8 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_48_414 ();
 sg13g2_decap_8 FILLER_48_421 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_fill_2 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_31 ();
 sg13g2_fill_1 FILLER_49_33 ();
 sg13g2_fill_2 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_78 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_110 ();
 sg13g2_decap_8 FILLER_49_117 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_decap_4 FILLER_49_131 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_decap_4 FILLER_49_164 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_fill_1 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_308 ();
 sg13g2_fill_2 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_377 ();
 sg13g2_decap_8 FILLER_49_384 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_decap_4 FILLER_49_424 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_decap_4 FILLER_50_29 ();
 sg13g2_fill_2 FILLER_50_33 ();
 sg13g2_decap_4 FILLER_50_61 ();
 sg13g2_fill_2 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_75 ();
 sg13g2_decap_8 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_90 ();
 sg13g2_decap_8 FILLER_50_97 ();
 sg13g2_decap_8 FILLER_50_104 ();
 sg13g2_decap_8 FILLER_50_111 ();
 sg13g2_decap_8 FILLER_50_118 ();
 sg13g2_decap_8 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_146 ();
 sg13g2_decap_8 FILLER_50_164 ();
 sg13g2_fill_1 FILLER_50_171 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_fill_2 FILLER_50_204 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_240 ();
 sg13g2_decap_8 FILLER_50_247 ();
 sg13g2_decap_8 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_272 ();
 sg13g2_decap_4 FILLER_50_279 ();
 sg13g2_fill_1 FILLER_50_283 ();
 sg13g2_decap_8 FILLER_50_292 ();
 sg13g2_decap_8 FILLER_50_299 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_decap_8 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_320 ();
 sg13g2_decap_4 FILLER_50_337 ();
 sg13g2_fill_2 FILLER_50_341 ();
 sg13g2_decap_4 FILLER_50_348 ();
 sg13g2_fill_1 FILLER_50_352 ();
 sg13g2_decap_8 FILLER_50_363 ();
 sg13g2_fill_1 FILLER_50_370 ();
 sg13g2_fill_2 FILLER_50_385 ();
 sg13g2_fill_1 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_50_409 ();
 sg13g2_decap_8 FILLER_50_416 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_4 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_60 ();
 sg13g2_decap_8 FILLER_51_88 ();
 sg13g2_decap_8 FILLER_51_95 ();
 sg13g2_decap_4 FILLER_51_102 ();
 sg13g2_fill_2 FILLER_51_106 ();
 sg13g2_fill_2 FILLER_51_134 ();
 sg13g2_fill_1 FILLER_51_136 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_157 ();
 sg13g2_fill_2 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_fill_2 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_fill_2 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_308 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_354 ();
 sg13g2_decap_4 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_372 ();
 sg13g2_decap_4 FILLER_51_387 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_decap_8 FILLER_51_416 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_79 ();
 sg13g2_decap_8 FILLER_52_86 ();
 sg13g2_decap_8 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_100 ();
 sg13g2_decap_8 FILLER_52_109 ();
 sg13g2_decap_8 FILLER_52_116 ();
 sg13g2_decap_4 FILLER_52_123 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_138 ();
 sg13g2_fill_1 FILLER_52_143 ();
 sg13g2_fill_2 FILLER_52_151 ();
 sg13g2_fill_1 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_180 ();
 sg13g2_decap_8 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_decap_8 FILLER_52_295 ();
 sg13g2_decap_8 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_52_389 ();
 sg13g2_fill_2 FILLER_52_395 ();
 sg13g2_fill_1 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_424 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_decap_8 FILLER_53_61 ();
 sg13g2_decap_8 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_155 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_decap_8 FILLER_53_184 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_fill_1 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_fill_1 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_230 ();
 sg13g2_decap_8 FILLER_53_236 ();
 sg13g2_decap_8 FILLER_53_243 ();
 sg13g2_decap_8 FILLER_53_250 ();
 sg13g2_decap_8 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_274 ();
 sg13g2_fill_2 FILLER_53_285 ();
 sg13g2_decap_8 FILLER_53_318 ();
 sg13g2_decap_8 FILLER_53_325 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_decap_8 FILLER_53_339 ();
 sg13g2_fill_1 FILLER_53_346 ();
 sg13g2_fill_2 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_53_412 ();
 sg13g2_decap_8 FILLER_53_419 ();
 sg13g2_decap_4 FILLER_53_426 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_2 FILLER_54_39 ();
 sg13g2_fill_2 FILLER_54_71 ();
 sg13g2_fill_2 FILLER_54_105 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_decap_8 FILLER_54_113 ();
 sg13g2_decap_8 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_139 ();
 sg13g2_fill_2 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_202 ();
 sg13g2_decap_8 FILLER_54_209 ();
 sg13g2_decap_4 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_225 ();
 sg13g2_decap_8 FILLER_54_232 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_8 FILLER_54_246 ();
 sg13g2_decap_8 FILLER_54_253 ();
 sg13g2_fill_2 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_262 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_4 FILLER_54_315 ();
 sg13g2_fill_2 FILLER_54_319 ();
 sg13g2_decap_8 FILLER_54_325 ();
 sg13g2_decap_8 FILLER_54_332 ();
 sg13g2_fill_2 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_404 ();
 sg13g2_decap_8 FILLER_54_411 ();
 sg13g2_decap_8 FILLER_54_418 ();
 sg13g2_decap_4 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_decap_4 FILLER_55_11 ();
 sg13g2_decap_8 FILLER_55_22 ();
 sg13g2_decap_8 FILLER_55_29 ();
 sg13g2_decap_4 FILLER_55_36 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_1 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_fill_2 FILLER_55_96 ();
 sg13g2_decap_8 FILLER_55_124 ();
 sg13g2_decap_4 FILLER_55_131 ();
 sg13g2_fill_1 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_2 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_158 ();
 sg13g2_decap_8 FILLER_55_164 ();
 sg13g2_decap_8 FILLER_55_171 ();
 sg13g2_decap_8 FILLER_55_178 ();
 sg13g2_decap_8 FILLER_55_185 ();
 sg13g2_decap_8 FILLER_55_192 ();
 sg13g2_decap_8 FILLER_55_199 ();
 sg13g2_decap_8 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_213 ();
 sg13g2_decap_8 FILLER_55_220 ();
 sg13g2_decap_8 FILLER_55_227 ();
 sg13g2_decap_8 FILLER_55_234 ();
 sg13g2_decap_8 FILLER_55_241 ();
 sg13g2_decap_8 FILLER_55_248 ();
 sg13g2_decap_8 FILLER_55_255 ();
 sg13g2_decap_8 FILLER_55_262 ();
 sg13g2_decap_8 FILLER_55_269 ();
 sg13g2_decap_8 FILLER_55_276 ();
 sg13g2_decap_8 FILLER_55_283 ();
 sg13g2_decap_4 FILLER_55_290 ();
 sg13g2_decap_8 FILLER_55_320 ();
 sg13g2_decap_4 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_365 ();
 sg13g2_decap_4 FILLER_55_371 ();
 sg13g2_fill_2 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_396 ();
 sg13g2_decap_8 FILLER_55_403 ();
 sg13g2_decap_8 FILLER_55_410 ();
 sg13g2_decap_8 FILLER_55_417 ();
 sg13g2_decap_4 FILLER_55_424 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_23 ();
 sg13g2_fill_1 FILLER_56_50 ();
 sg13g2_decap_4 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_81 ();
 sg13g2_decap_8 FILLER_56_87 ();
 sg13g2_decap_8 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_101 ();
 sg13g2_decap_4 FILLER_56_108 ();
 sg13g2_decap_8 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_decap_8 FILLER_56_157 ();
 sg13g2_decap_4 FILLER_56_164 ();
 sg13g2_fill_2 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_205 ();
 sg13g2_decap_8 FILLER_56_212 ();
 sg13g2_decap_8 FILLER_56_219 ();
 sg13g2_decap_4 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_decap_4 FILLER_56_295 ();
 sg13g2_decap_8 FILLER_56_325 ();
 sg13g2_decap_8 FILLER_56_332 ();
 sg13g2_decap_8 FILLER_56_339 ();
 sg13g2_decap_4 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_376 ();
 sg13g2_decap_8 FILLER_56_403 ();
 sg13g2_decap_8 FILLER_56_410 ();
 sg13g2_decap_8 FILLER_56_417 ();
 sg13g2_decap_4 FILLER_56_424 ();
 sg13g2_fill_2 FILLER_56_428 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_18 ();
 sg13g2_decap_8 FILLER_57_29 ();
 sg13g2_decap_4 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_54 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_fill_1 FILLER_57_67 ();
 sg13g2_fill_2 FILLER_57_75 ();
 sg13g2_fill_1 FILLER_57_77 ();
 sg13g2_decap_4 FILLER_57_93 ();
 sg13g2_decap_8 FILLER_57_123 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_fill_1 FILLER_57_132 ();
 sg13g2_fill_2 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_fill_2 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_159 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_decap_8 FILLER_57_178 ();
 sg13g2_decap_8 FILLER_57_185 ();
 sg13g2_fill_2 FILLER_57_192 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_1 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_232 ();
 sg13g2_decap_8 FILLER_57_239 ();
 sg13g2_decap_4 FILLER_57_246 ();
 sg13g2_decap_8 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_309 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_decap_8 FILLER_57_324 ();
 sg13g2_decap_8 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_57_338 ();
 sg13g2_decap_8 FILLER_57_345 ();
 sg13g2_decap_8 FILLER_57_352 ();
 sg13g2_decap_8 FILLER_57_359 ();
 sg13g2_decap_8 FILLER_57_366 ();
 sg13g2_decap_8 FILLER_57_373 ();
 sg13g2_decap_8 FILLER_57_380 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_decap_8 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_422 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_decap_8 FILLER_58_36 ();
 sg13g2_decap_8 FILLER_58_43 ();
 sg13g2_fill_2 FILLER_58_50 ();
 sg13g2_fill_2 FILLER_58_66 ();
 sg13g2_fill_2 FILLER_58_71 ();
 sg13g2_fill_1 FILLER_58_77 ();
 sg13g2_fill_1 FILLER_58_88 ();
 sg13g2_decap_8 FILLER_58_94 ();
 sg13g2_decap_8 FILLER_58_101 ();
 sg13g2_decap_8 FILLER_58_108 ();
 sg13g2_decap_8 FILLER_58_115 ();
 sg13g2_decap_8 FILLER_58_122 ();
 sg13g2_fill_2 FILLER_58_129 ();
 sg13g2_fill_2 FILLER_58_171 ();
 sg13g2_fill_1 FILLER_58_204 ();
 sg13g2_fill_2 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_fill_1 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_decap_8 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_58_415 ();
 sg13g2_decap_8 FILLER_58_422 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_47 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_71 ();
 sg13g2_decap_4 FILLER_59_100 ();
 sg13g2_decap_8 FILLER_59_108 ();
 sg13g2_decap_4 FILLER_59_115 ();
 sg13g2_fill_1 FILLER_59_119 ();
 sg13g2_decap_4 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_decap_8 FILLER_59_180 ();
 sg13g2_decap_8 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_fill_2 FILLER_59_201 ();
 sg13g2_decap_8 FILLER_59_229 ();
 sg13g2_decap_8 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_243 ();
 sg13g2_decap_8 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_257 ();
 sg13g2_fill_2 FILLER_59_292 ();
 sg13g2_decap_8 FILLER_59_302 ();
 sg13g2_decap_8 FILLER_59_309 ();
 sg13g2_decap_4 FILLER_59_316 ();
 sg13g2_decap_8 FILLER_59_377 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_8 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_59_412 ();
 sg13g2_decap_8 FILLER_59_419 ();
 sg13g2_decap_4 FILLER_59_426 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_51 ();
 sg13g2_fill_2 FILLER_60_58 ();
 sg13g2_fill_1 FILLER_60_65 ();
 sg13g2_fill_2 FILLER_60_70 ();
 sg13g2_fill_1 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_fill_2 FILLER_60_171 ();
 sg13g2_decap_8 FILLER_60_204 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_decap_8 FILLER_60_218 ();
 sg13g2_decap_8 FILLER_60_225 ();
 sg13g2_decap_4 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_236 ();
 sg13g2_decap_4 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_303 ();
 sg13g2_decap_8 FILLER_60_310 ();
 sg13g2_decap_4 FILLER_60_317 ();
 sg13g2_decap_4 FILLER_60_325 ();
 sg13g2_decap_4 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_341 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_decap_4 FILLER_60_365 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_fill_2 FILLER_60_374 ();
 sg13g2_decap_4 FILLER_60_384 ();
 sg13g2_fill_1 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_427 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_4 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_46 ();
 sg13g2_fill_1 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_decap_4 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_decap_8 FILLER_61_130 ();
 sg13g2_decap_8 FILLER_61_137 ();
 sg13g2_fill_2 FILLER_61_144 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_decap_4 FILLER_61_152 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_decap_4 FILLER_61_204 ();
 sg13g2_fill_1 FILLER_61_208 ();
 sg13g2_decap_8 FILLER_61_235 ();
 sg13g2_decap_4 FILLER_61_271 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_fill_1 FILLER_61_311 ();
 sg13g2_fill_1 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_347 ();
 sg13g2_fill_2 FILLER_61_375 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_decap_8 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_61_414 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_fill_2 FILLER_62_64 ();
 sg13g2_fill_1 FILLER_62_76 ();
 sg13g2_decap_8 FILLER_62_92 ();
 sg13g2_decap_8 FILLER_62_99 ();
 sg13g2_decap_8 FILLER_62_106 ();
 sg13g2_decap_8 FILLER_62_113 ();
 sg13g2_fill_2 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_122 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_fill_2 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_186 ();
 sg13g2_decap_8 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_decap_8 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_242 ();
 sg13g2_decap_8 FILLER_62_249 ();
 sg13g2_decap_8 FILLER_62_264 ();
 sg13g2_decap_8 FILLER_62_271 ();
 sg13g2_decap_8 FILLER_62_278 ();
 sg13g2_decap_8 FILLER_62_285 ();
 sg13g2_fill_2 FILLER_62_292 ();
 sg13g2_decap_8 FILLER_62_298 ();
 sg13g2_fill_2 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_348 ();
 sg13g2_fill_1 FILLER_62_353 ();
 sg13g2_fill_1 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_371 ();
 sg13g2_decap_4 FILLER_62_379 ();
 sg13g2_fill_1 FILLER_62_383 ();
 sg13g2_fill_2 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_30 ();
 sg13g2_decap_8 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_decap_8 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_144 ();
 sg13g2_decap_4 FILLER_63_212 ();
 sg13g2_fill_1 FILLER_63_216 ();
 sg13g2_decap_8 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_261 ();
 sg13g2_fill_2 FILLER_63_265 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_2 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_313 ();
 sg13g2_decap_8 FILLER_63_320 ();
 sg13g2_fill_2 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_338 ();
 sg13g2_decap_8 FILLER_63_345 ();
 sg13g2_decap_8 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_decap_8 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_401 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_4 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_46 ();
 sg13g2_fill_2 FILLER_64_83 ();
 sg13g2_decap_8 FILLER_64_96 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_decap_8 FILLER_64_110 ();
 sg13g2_decap_8 FILLER_64_117 ();
 sg13g2_decap_8 FILLER_64_124 ();
 sg13g2_decap_4 FILLER_64_131 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_fill_1 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_188 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_decap_8 FILLER_64_209 ();
 sg13g2_fill_1 FILLER_64_216 ();
 sg13g2_fill_2 FILLER_64_275 ();
 sg13g2_fill_1 FILLER_64_277 ();
 sg13g2_fill_2 FILLER_64_287 ();
 sg13g2_decap_4 FILLER_64_296 ();
 sg13g2_decap_8 FILLER_64_326 ();
 sg13g2_decap_8 FILLER_64_333 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_2 FILLER_64_375 ();
 sg13g2_fill_1 FILLER_64_377 ();
 sg13g2_decap_4 FILLER_64_395 ();
 sg13g2_fill_1 FILLER_64_399 ();
 sg13g2_decap_8 FILLER_64_404 ();
 sg13g2_decap_8 FILLER_64_411 ();
 sg13g2_decap_8 FILLER_64_418 ();
 sg13g2_decap_4 FILLER_64_425 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_84 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_151 ();
 sg13g2_decap_4 FILLER_65_157 ();
 sg13g2_decap_8 FILLER_65_164 ();
 sg13g2_decap_8 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_decap_4 FILLER_65_185 ();
 sg13g2_decap_8 FILLER_65_197 ();
 sg13g2_decap_8 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_223 ();
 sg13g2_decap_4 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_decap_4 FILLER_65_245 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_281 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_decap_4 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_307 ();
 sg13g2_fill_2 FILLER_65_313 ();
 sg13g2_decap_4 FILLER_65_334 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_fill_2 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_356 ();
 sg13g2_fill_2 FILLER_65_369 ();
 sg13g2_fill_1 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_8 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_4 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_58 ();
 sg13g2_decap_8 FILLER_66_65 ();
 sg13g2_decap_8 FILLER_66_72 ();
 sg13g2_decap_8 FILLER_66_79 ();
 sg13g2_decap_8 FILLER_66_86 ();
 sg13g2_decap_8 FILLER_66_93 ();
 sg13g2_decap_8 FILLER_66_100 ();
 sg13g2_decap_8 FILLER_66_107 ();
 sg13g2_decap_4 FILLER_66_114 ();
 sg13g2_decap_8 FILLER_66_123 ();
 sg13g2_decap_4 FILLER_66_130 ();
 sg13g2_fill_2 FILLER_66_191 ();
 sg13g2_fill_1 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_220 ();
 sg13g2_decap_8 FILLER_66_227 ();
 sg13g2_decap_8 FILLER_66_234 ();
 sg13g2_decap_8 FILLER_66_241 ();
 sg13g2_decap_4 FILLER_66_248 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_298 ();
 sg13g2_decap_4 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_309 ();
 sg13g2_fill_2 FILLER_66_346 ();
 sg13g2_decap_4 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_356 ();
 sg13g2_decap_4 FILLER_66_368 ();
 sg13g2_fill_2 FILLER_66_372 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_fill_2 FILLER_66_394 ();
 sg13g2_decap_4 FILLER_66_426 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_32 ();
 sg13g2_decap_8 FILLER_67_64 ();
 sg13g2_decap_8 FILLER_67_71 ();
 sg13g2_decap_8 FILLER_67_78 ();
 sg13g2_decap_8 FILLER_67_85 ();
 sg13g2_fill_2 FILLER_67_92 ();
 sg13g2_fill_1 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_142 ();
 sg13g2_fill_1 FILLER_67_144 ();
 sg13g2_fill_2 FILLER_67_150 ();
 sg13g2_fill_1 FILLER_67_152 ();
 sg13g2_fill_1 FILLER_67_171 ();
 sg13g2_fill_2 FILLER_67_176 ();
 sg13g2_decap_8 FILLER_67_220 ();
 sg13g2_decap_8 FILLER_67_227 ();
 sg13g2_decap_8 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_241 ();
 sg13g2_decap_8 FILLER_67_248 ();
 sg13g2_decap_4 FILLER_67_283 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_344 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_fill_2 FILLER_67_378 ();
 sg13g2_fill_1 FILLER_67_380 ();
 sg13g2_fill_2 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_decap_8 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_422 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_4 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_53 ();
 sg13g2_fill_2 FILLER_68_68 ();
 sg13g2_fill_1 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_90 ();
 sg13g2_decap_8 FILLER_68_97 ();
 sg13g2_decap_8 FILLER_68_104 ();
 sg13g2_decap_8 FILLER_68_111 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_fill_2 FILLER_68_145 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_decap_8 FILLER_68_253 ();
 sg13g2_decap_4 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_287 ();
 sg13g2_decap_4 FILLER_68_297 ();
 sg13g2_fill_2 FILLER_68_301 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_fill_1 FILLER_68_309 ();
 sg13g2_fill_1 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_323 ();
 sg13g2_fill_1 FILLER_68_334 ();
 sg13g2_fill_2 FILLER_68_347 ();
 sg13g2_fill_2 FILLER_68_353 ();
 sg13g2_fill_1 FILLER_68_355 ();
 sg13g2_fill_2 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_398 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_49 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_2 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_decap_4 FILLER_69_134 ();
 sg13g2_fill_2 FILLER_69_143 ();
 sg13g2_fill_1 FILLER_69_145 ();
 sg13g2_fill_1 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_178 ();
 sg13g2_decap_8 FILLER_69_185 ();
 sg13g2_decap_8 FILLER_69_192 ();
 sg13g2_decap_8 FILLER_69_199 ();
 sg13g2_decap_8 FILLER_69_206 ();
 sg13g2_decap_8 FILLER_69_213 ();
 sg13g2_fill_2 FILLER_69_220 ();
 sg13g2_decap_4 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_decap_8 FILLER_69_249 ();
 sg13g2_decap_4 FILLER_69_256 ();
 sg13g2_decap_4 FILLER_69_264 ();
 sg13g2_fill_2 FILLER_69_273 ();
 sg13g2_fill_1 FILLER_69_275 ();
 sg13g2_decap_4 FILLER_69_291 ();
 sg13g2_fill_2 FILLER_69_326 ();
 sg13g2_fill_2 FILLER_69_333 ();
 sg13g2_fill_1 FILLER_69_335 ();
 sg13g2_decap_8 FILLER_69_347 ();
 sg13g2_decap_4 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_fill_2 FILLER_69_384 ();
 sg13g2_fill_1 FILLER_69_386 ();
 sg13g2_fill_2 FILLER_69_391 ();
 sg13g2_decap_4 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_decap_8 FILLER_69_415 ();
 sg13g2_decap_8 FILLER_69_422 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_41 ();
 sg13g2_fill_2 FILLER_70_57 ();
 sg13g2_fill_1 FILLER_70_89 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_decap_8 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_decap_8 FILLER_70_115 ();
 sg13g2_decap_8 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_129 ();
 sg13g2_fill_1 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_181 ();
 sg13g2_decap_8 FILLER_70_188 ();
 sg13g2_decap_8 FILLER_70_195 ();
 sg13g2_decap_8 FILLER_70_202 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_decap_8 FILLER_70_225 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_fill_1 FILLER_70_234 ();
 sg13g2_decap_8 FILLER_70_240 ();
 sg13g2_decap_8 FILLER_70_247 ();
 sg13g2_fill_2 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_256 ();
 sg13g2_fill_1 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_278 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_decap_8 FILLER_70_298 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_4 FILLER_70_319 ();
 sg13g2_fill_1 FILLER_70_323 ();
 sg13g2_fill_2 FILLER_70_333 ();
 sg13g2_decap_4 FILLER_70_341 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_decap_4 FILLER_70_350 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_decap_8 FILLER_70_361 ();
 sg13g2_decap_8 FILLER_70_368 ();
 sg13g2_decap_4 FILLER_70_375 ();
 sg13g2_decap_8 FILLER_70_411 ();
 sg13g2_decap_8 FILLER_70_418 ();
 sg13g2_decap_4 FILLER_70_425 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_4 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_39 ();
 sg13g2_fill_1 FILLER_71_53 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_decap_4 FILLER_71_85 ();
 sg13g2_fill_1 FILLER_71_89 ();
 sg13g2_fill_2 FILLER_71_94 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_2 FILLER_71_123 ();
 sg13g2_fill_1 FILLER_71_125 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_147 ();
 sg13g2_fill_1 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_163 ();
 sg13g2_decap_4 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_270 ();
 sg13g2_fill_1 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_334 ();
 sg13g2_decap_4 FILLER_71_351 ();
 sg13g2_decap_4 FILLER_71_359 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_49 ();
 sg13g2_fill_1 FILLER_72_51 ();
 sg13g2_fill_2 FILLER_72_60 ();
 sg13g2_fill_2 FILLER_72_65 ();
 sg13g2_fill_2 FILLER_72_99 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_fill_2 FILLER_72_119 ();
 sg13g2_fill_1 FILLER_72_121 ();
 sg13g2_fill_1 FILLER_72_127 ();
 sg13g2_fill_1 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_140 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_fill_2 FILLER_72_176 ();
 sg13g2_fill_1 FILLER_72_178 ();
 sg13g2_fill_2 FILLER_72_213 ();
 sg13g2_decap_4 FILLER_72_220 ();
 sg13g2_fill_2 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_4 FILLER_72_238 ();
 sg13g2_fill_2 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_decap_4 FILLER_72_254 ();
 sg13g2_fill_1 FILLER_72_258 ();
 sg13g2_decap_4 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_decap_4 FILLER_72_341 ();
 sg13g2_fill_2 FILLER_72_350 ();
 sg13g2_fill_1 FILLER_72_352 ();
 sg13g2_fill_2 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_72_412 ();
 sg13g2_decap_8 FILLER_72_419 ();
 sg13g2_decap_4 FILLER_72_426 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_4 FILLER_73_35 ();
 sg13g2_fill_2 FILLER_73_39 ();
 sg13g2_decap_4 FILLER_73_51 ();
 sg13g2_fill_1 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_94 ();
 sg13g2_fill_2 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_163 ();
 sg13g2_fill_1 FILLER_73_170 ();
 sg13g2_fill_2 FILLER_73_214 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_2 FILLER_73_353 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_fill_2 FILLER_73_380 ();
 sg13g2_fill_1 FILLER_73_382 ();
 sg13g2_decap_4 FILLER_73_394 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_fill_2 FILLER_74_59 ();
 sg13g2_fill_2 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_139 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_181 ();
 sg13g2_decap_8 FILLER_74_188 ();
 sg13g2_decap_8 FILLER_74_195 ();
 sg13g2_decap_8 FILLER_74_202 ();
 sg13g2_decap_8 FILLER_74_209 ();
 sg13g2_decap_8 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_4 FILLER_74_252 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_fill_2 FILLER_74_272 ();
 sg13g2_fill_1 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_313 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_331 ();
 sg13g2_decap_4 FILLER_74_342 ();
 sg13g2_fill_1 FILLER_74_355 ();
 sg13g2_fill_2 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_74_376 ();
 sg13g2_fill_1 FILLER_74_378 ();
 sg13g2_decap_4 FILLER_74_384 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_decap_8 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_74_414 ();
 sg13g2_decap_8 FILLER_74_421 ();
 sg13g2_fill_2 FILLER_74_428 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_fill_2 FILLER_75_51 ();
 sg13g2_fill_1 FILLER_75_53 ();
 sg13g2_fill_2 FILLER_75_58 ();
 sg13g2_fill_1 FILLER_75_60 ();
 sg13g2_fill_1 FILLER_75_64 ();
 sg13g2_fill_2 FILLER_75_69 ();
 sg13g2_fill_1 FILLER_75_81 ();
 sg13g2_fill_1 FILLER_75_86 ();
 sg13g2_decap_8 FILLER_75_92 ();
 sg13g2_decap_8 FILLER_75_99 ();
 sg13g2_decap_8 FILLER_75_106 ();
 sg13g2_decap_8 FILLER_75_113 ();
 sg13g2_decap_8 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_140 ();
 sg13g2_fill_1 FILLER_75_142 ();
 sg13g2_fill_1 FILLER_75_157 ();
 sg13g2_fill_1 FILLER_75_163 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_179 ();
 sg13g2_fill_1 FILLER_75_181 ();
 sg13g2_decap_4 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_fill_1 FILLER_75_288 ();
 sg13g2_decap_8 FILLER_75_293 ();
 sg13g2_decap_8 FILLER_75_300 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_decap_8 FILLER_75_314 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_decap_4 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_4 FILLER_75_350 ();
 sg13g2_fill_1 FILLER_75_354 ();
 sg13g2_decap_4 FILLER_75_381 ();
 sg13g2_fill_1 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_4 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_51 ();
 sg13g2_fill_2 FILLER_76_65 ();
 sg13g2_fill_1 FILLER_76_72 ();
 sg13g2_fill_2 FILLER_76_78 ();
 sg13g2_decap_8 FILLER_76_85 ();
 sg13g2_decap_8 FILLER_76_92 ();
 sg13g2_decap_8 FILLER_76_99 ();
 sg13g2_decap_8 FILLER_76_106 ();
 sg13g2_decap_8 FILLER_76_113 ();
 sg13g2_decap_8 FILLER_76_120 ();
 sg13g2_decap_8 FILLER_76_127 ();
 sg13g2_fill_2 FILLER_76_134 ();
 sg13g2_fill_1 FILLER_76_136 ();
 sg13g2_fill_1 FILLER_76_144 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_decap_8 FILLER_76_180 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_decap_8 FILLER_76_194 ();
 sg13g2_decap_4 FILLER_76_201 ();
 sg13g2_fill_2 FILLER_76_205 ();
 sg13g2_decap_4 FILLER_76_210 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_4 FILLER_76_256 ();
 sg13g2_fill_1 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_296 ();
 sg13g2_decap_8 FILLER_76_303 ();
 sg13g2_fill_2 FILLER_76_310 ();
 sg13g2_fill_1 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_317 ();
 sg13g2_fill_1 FILLER_76_324 ();
 sg13g2_decap_4 FILLER_76_329 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_decap_4 FILLER_76_343 ();
 sg13g2_fill_2 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_fill_2 FILLER_76_373 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_decap_4 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_fill_1 FILLER_76_394 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_4 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_32 ();
 sg13g2_fill_1 FILLER_77_59 ();
 sg13g2_fill_1 FILLER_77_64 ();
 sg13g2_fill_1 FILLER_77_81 ();
 sg13g2_fill_1 FILLER_77_88 ();
 sg13g2_decap_8 FILLER_77_115 ();
 sg13g2_fill_1 FILLER_77_122 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_fill_2 FILLER_77_177 ();
 sg13g2_decap_4 FILLER_77_205 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_decap_8 FILLER_77_236 ();
 sg13g2_decap_8 FILLER_77_243 ();
 sg13g2_fill_2 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_252 ();
 sg13g2_fill_1 FILLER_77_339 ();
 sg13g2_decap_8 FILLER_77_344 ();
 sg13g2_fill_2 FILLER_77_351 ();
 sg13g2_decap_4 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_366 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_378 ();
 sg13g2_fill_1 FILLER_77_383 ();
 sg13g2_fill_2 FILLER_77_392 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_fill_2 FILLER_78_85 ();
 sg13g2_fill_1 FILLER_78_87 ();
 sg13g2_decap_8 FILLER_78_96 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_decap_8 FILLER_78_110 ();
 sg13g2_fill_1 FILLER_78_117 ();
 sg13g2_fill_2 FILLER_78_149 ();
 sg13g2_fill_2 FILLER_78_155 ();
 sg13g2_fill_2 FILLER_78_164 ();
 sg13g2_decap_8 FILLER_78_171 ();
 sg13g2_fill_2 FILLER_78_178 ();
 sg13g2_fill_1 FILLER_78_180 ();
 sg13g2_fill_2 FILLER_78_186 ();
 sg13g2_fill_1 FILLER_78_188 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_203 ();
 sg13g2_decap_4 FILLER_78_208 ();
 sg13g2_fill_1 FILLER_78_310 ();
 sg13g2_fill_1 FILLER_78_315 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_4 FILLER_78_424 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_57 ();
 sg13g2_fill_2 FILLER_79_61 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_fill_1 FILLER_79_73 ();
 sg13g2_fill_1 FILLER_79_79 ();
 sg13g2_decap_8 FILLER_79_93 ();
 sg13g2_fill_2 FILLER_79_100 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_decap_8 FILLER_79_111 ();
 sg13g2_decap_8 FILLER_79_118 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_127 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_8 FILLER_79_139 ();
 sg13g2_decap_4 FILLER_79_146 ();
 sg13g2_fill_2 FILLER_79_150 ();
 sg13g2_decap_4 FILLER_79_156 ();
 sg13g2_fill_2 FILLER_79_160 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_218 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_2 FILLER_79_266 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_fill_2 FILLER_79_274 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_288 ();
 sg13g2_fill_1 FILLER_79_290 ();
 sg13g2_decap_4 FILLER_79_304 ();
 sg13g2_decap_4 FILLER_79_334 ();
 sg13g2_fill_1 FILLER_79_338 ();
 sg13g2_fill_2 FILLER_79_373 ();
 sg13g2_fill_1 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_410 ();
 sg13g2_decap_8 FILLER_79_417 ();
 sg13g2_decap_4 FILLER_79_424 ();
 sg13g2_fill_2 FILLER_79_428 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_72 ();
 sg13g2_decap_4 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_89 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_fill_1 FILLER_80_103 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_fill_1 FILLER_80_110 ();
 sg13g2_fill_2 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_125 ();
 sg13g2_fill_2 FILLER_80_130 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_149 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_168 ();
 sg13g2_fill_2 FILLER_80_175 ();
 sg13g2_fill_1 FILLER_80_177 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_fill_2 FILLER_80_193 ();
 sg13g2_fill_1 FILLER_80_195 ();
 sg13g2_fill_2 FILLER_80_204 ();
 sg13g2_decap_8 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_225 ();
 sg13g2_fill_2 FILLER_80_232 ();
 sg13g2_fill_1 FILLER_80_234 ();
 sg13g2_fill_1 FILLER_80_239 ();
 sg13g2_decap_4 FILLER_80_244 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_fill_1 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_decap_4 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_369 ();
 sg13g2_fill_2 FILLER_80_376 ();
 sg13g2_fill_1 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
