module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_inv ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _14753_ (.A(\cpu.dec.r_op[5] ),
    .X(_08051_));
 sg13g2_buf_1 _14754_ (.A(_08051_),
    .X(_08052_));
 sg13g2_buf_8 _14755_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08053_));
 sg13g2_buf_1 _14756_ (.A(net1096),
    .X(_08054_));
 sg13g2_buf_8 _14757_ (.A(\cpu.ex.pc[12] ),
    .X(_08055_));
 sg13g2_buf_4 _14758_ (.X(_08056_),
    .A(_08055_));
 sg13g2_buf_2 _14759_ (.A(_08056_),
    .X(_08057_));
 sg13g2_buf_8 _14760_ (.A(\cpu.ex.pc[13] ),
    .X(_08058_));
 sg13g2_buf_1 _14761_ (.A(net1095),
    .X(_08059_));
 sg13g2_buf_1 _14762_ (.A(net1041),
    .X(_08060_));
 sg13g2_mux4_1 _14763_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net913),
    .X(_08061_));
 sg13g2_mux4_1 _14764_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net913),
    .X(_08062_));
 sg13g2_buf_2 _14765_ (.A(_08056_),
    .X(_08063_));
 sg13g2_buf_1 _14766_ (.A(net1041),
    .X(_08064_));
 sg13g2_mux4_1 _14767_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(net911),
    .X(_08065_));
 sg13g2_buf_2 _14768_ (.A(_08056_),
    .X(_08066_));
 sg13g2_buf_1 _14769_ (.A(net1041),
    .X(_08067_));
 sg13g2_mux4_1 _14770_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net909),
    .X(_08068_));
 sg13g2_buf_1 _14771_ (.A(\cpu.ex.pc[15] ),
    .X(_08069_));
 sg13g2_inv_2 _14772_ (.Y(_08070_),
    .A(net1094));
 sg13g2_buf_2 _14773_ (.A(_08070_),
    .X(_08071_));
 sg13g2_buf_8 _14774_ (.A(\cpu.ex.pc[14] ),
    .X(_08072_));
 sg13g2_buf_8 _14775_ (.A(_08072_),
    .X(_08073_));
 sg13g2_buf_1 _14776_ (.A(net1040),
    .X(_08074_));
 sg13g2_mux4_1 _14777_ (.S0(net908),
    .A0(_08061_),
    .A1(_08062_),
    .A2(_08065_),
    .A3(_08068_),
    .S1(net907),
    .X(_08075_));
 sg13g2_mux4_1 _14778_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net909),
    .X(_08076_));
 sg13g2_mux4_1 _14779_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net913),
    .X(_08077_));
 sg13g2_mux4_1 _14780_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net911),
    .X(_08078_));
 sg13g2_mux4_1 _14781_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net911),
    .X(_08079_));
 sg13g2_mux4_1 _14782_ (.S0(net908),
    .A0(_08076_),
    .A1(_08077_),
    .A2(_08078_),
    .A3(_08079_),
    .S1(net907),
    .X(_08080_));
 sg13g2_buf_8 _14783_ (.A(\cpu.dec.supmode ),
    .X(_08081_));
 sg13g2_buf_1 _14784_ (.A(_08081_),
    .X(_08082_));
 sg13g2_mux2_1 _14785_ (.A0(_08075_),
    .A1(_08080_),
    .S(_08082_),
    .X(_08083_));
 sg13g2_inv_1 _14786_ (.Y(_08084_),
    .A(net1095));
 sg13g2_nor2_1 _14787_ (.A(_08084_),
    .B(net1042),
    .Y(_08085_));
 sg13g2_a21oi_1 _14788_ (.A1(net1042),
    .A2(_08083_),
    .Y(_08086_),
    .B1(_08085_));
 sg13g2_buf_1 _14789_ (.A(_08086_),
    .X(_08087_));
 sg13g2_buf_1 _14790_ (.A(_00190_),
    .X(_08088_));
 sg13g2_buf_1 _14791_ (.A(\cpu.ex.pc[3] ),
    .X(_08089_));
 sg13g2_inv_2 _14792_ (.Y(_08090_),
    .A(net1092));
 sg13g2_buf_1 _14793_ (.A(\cpu.ex.pc[4] ),
    .X(_08091_));
 sg13g2_buf_1 _14794_ (.A(_08091_),
    .X(_08092_));
 sg13g2_inv_2 _14795_ (.Y(_08093_),
    .A(_08091_));
 sg13g2_buf_2 _14796_ (.A(\cpu.ex.pc[2] ),
    .X(_08094_));
 sg13g2_a21oi_1 _14797_ (.A1(net1092),
    .A2(_08093_),
    .Y(_08095_),
    .B1(_08094_));
 sg13g2_a21o_1 _14798_ (.A2(_08092_),
    .A1(_08090_),
    .B1(_08095_),
    .X(_08096_));
 sg13g2_nand2_1 _14799_ (.Y(_08097_),
    .A(net1093),
    .B(_08096_));
 sg13g2_buf_2 _14800_ (.A(_08097_),
    .X(_08098_));
 sg13g2_buf_1 _14801_ (.A(_08098_),
    .X(_08099_));
 sg13g2_buf_1 _14802_ (.A(_08099_),
    .X(_08100_));
 sg13g2_buf_1 _14803_ (.A(net477),
    .X(_08101_));
 sg13g2_buf_1 _14804_ (.A(_08098_),
    .X(_08102_));
 sg13g2_buf_1 _14805_ (.A(net547),
    .X(_08103_));
 sg13g2_buf_1 _14806_ (.A(_08103_),
    .X(_08104_));
 sg13g2_inv_2 _14807_ (.Y(_08105_),
    .A(net1093));
 sg13g2_buf_1 _14808_ (.A(_08105_),
    .X(_08106_));
 sg13g2_buf_1 _14809_ (.A(net906),
    .X(_08107_));
 sg13g2_buf_1 _14810_ (.A(_08094_),
    .X(_08108_));
 sg13g2_buf_2 _14811_ (.A(_08108_),
    .X(_08109_));
 sg13g2_buf_1 _14812_ (.A(net1092),
    .X(_08110_));
 sg13g2_buf_2 _14813_ (.A(net1036),
    .X(_08111_));
 sg13g2_buf_1 _14814_ (.A(net904),
    .X(_08112_));
 sg13g2_buf_1 _14815_ (.A(_08112_),
    .X(_08113_));
 sg13g2_mux4_1 _14816_ (.S0(net905),
    .A0(\cpu.icache.r_tag[4][13] ),
    .A1(\cpu.icache.r_tag[5][13] ),
    .A2(\cpu.icache.r_tag[6][13] ),
    .A3(\cpu.icache.r_tag[7][13] ),
    .S1(net703),
    .X(_08114_));
 sg13g2_nand2_1 _14817_ (.Y(_08115_),
    .A(net777),
    .B(_08114_));
 sg13g2_nor2_1 _14818_ (.A(_08094_),
    .B(_08090_),
    .Y(_08116_));
 sg13g2_buf_2 _14819_ (.A(_08116_),
    .X(_08117_));
 sg13g2_and2_1 _14820_ (.A(_08093_),
    .B(_08117_),
    .X(_08118_));
 sg13g2_buf_2 _14821_ (.A(_08118_),
    .X(_08119_));
 sg13g2_buf_1 _14822_ (.A(_08119_),
    .X(_08120_));
 sg13g2_buf_1 _14823_ (.A(net546),
    .X(_08121_));
 sg13g2_nand2_1 _14824_ (.Y(_08122_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(net475));
 sg13g2_inv_1 _14825_ (.Y(_08123_),
    .A(_08094_));
 sg13g2_nor3_1 _14826_ (.A(_08123_),
    .B(net1092),
    .C(_08092_),
    .Y(_08124_));
 sg13g2_buf_2 _14827_ (.A(_08124_),
    .X(_08125_));
 sg13g2_buf_1 _14828_ (.A(_08125_),
    .X(_08126_));
 sg13g2_buf_1 _14829_ (.A(net702),
    .X(_08127_));
 sg13g2_nand2_1 _14830_ (.Y(_08128_),
    .A(_08094_),
    .B(net1092));
 sg13g2_buf_1 _14831_ (.A(_08128_),
    .X(_08129_));
 sg13g2_nor2_1 _14832_ (.A(_08105_),
    .B(_08129_),
    .Y(_08130_));
 sg13g2_buf_1 _14833_ (.A(_08130_),
    .X(_08131_));
 sg13g2_buf_1 _14834_ (.A(_08131_),
    .X(_08132_));
 sg13g2_buf_1 _14835_ (.A(net598),
    .X(_08133_));
 sg13g2_a22oi_1 _14836_ (.Y(_08134_),
    .B1(net545),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(net599),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_nand4_1 _14837_ (.B(_08115_),
    .C(_08122_),
    .A(net410),
    .Y(_08135_),
    .D(_08134_));
 sg13g2_o21ai_1 _14838_ (.B1(_08135_),
    .Y(_08136_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net411));
 sg13g2_xnor2_1 _14839_ (.Y(_08137_),
    .A(net478),
    .B(_08136_));
 sg13g2_mux4_1 _14840_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net909),
    .X(_08138_));
 sg13g2_mux4_1 _14841_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net913),
    .X(_08139_));
 sg13g2_mux4_1 _14842_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(net911),
    .X(_08140_));
 sg13g2_mux4_1 _14843_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(net911),
    .X(_08141_));
 sg13g2_mux4_1 _14844_ (.S0(net908),
    .A0(_08138_),
    .A1(_08139_),
    .A2(_08140_),
    .A3(_08141_),
    .S1(net907),
    .X(_08142_));
 sg13g2_mux4_1 _14845_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net909),
    .X(_08143_));
 sg13g2_mux4_1 _14846_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net909),
    .X(_08144_));
 sg13g2_mux4_1 _14847_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net911),
    .X(_08145_));
 sg13g2_mux4_1 _14848_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net911),
    .X(_08146_));
 sg13g2_mux4_1 _14849_ (.S0(net908),
    .A0(_08143_),
    .A1(_08144_),
    .A2(_08145_),
    .A3(_08146_),
    .S1(net907),
    .X(_08147_));
 sg13g2_mux2_1 _14850_ (.A0(_08142_),
    .A1(_08147_),
    .S(net1039),
    .X(_08148_));
 sg13g2_inv_2 _14851_ (.Y(_08149_),
    .A(_08055_));
 sg13g2_nor2_1 _14852_ (.A(_08149_),
    .B(net1042),
    .Y(_08150_));
 sg13g2_a21oi_1 _14853_ (.A1(net1042),
    .A2(_08148_),
    .Y(_08151_),
    .B1(_08150_));
 sg13g2_buf_1 _14854_ (.A(_08151_),
    .X(_08152_));
 sg13g2_and2_1 _14855_ (.A(_08105_),
    .B(_08117_),
    .X(_08153_));
 sg13g2_buf_1 _14856_ (.A(_08153_),
    .X(_08154_));
 sg13g2_buf_1 _14857_ (.A(_08154_),
    .X(_08155_));
 sg13g2_a22oi_1 _14858_ (.Y(_08156_),
    .B1(_08155_),
    .B2(\cpu.icache.r_tag[6][12] ),
    .A2(net475),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_buf_1 _14859_ (.A(_08133_),
    .X(_08157_));
 sg13g2_a22oi_1 _14860_ (.Y(_08158_),
    .B1(net473),
    .B2(\cpu.icache.r_tag[3][12] ),
    .A2(_08127_),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_buf_1 _14861_ (.A(_08088_),
    .X(_08159_));
 sg13g2_buf_1 _14862_ (.A(net1035),
    .X(_08160_));
 sg13g2_buf_1 _14863_ (.A(net903),
    .X(_08161_));
 sg13g2_buf_1 _14864_ (.A(net775),
    .X(_08162_));
 sg13g2_buf_1 _14865_ (.A(net1036),
    .X(_08163_));
 sg13g2_mux2_1 _14866_ (.A0(\cpu.icache.r_tag[5][12] ),
    .A1(\cpu.icache.r_tag[7][12] ),
    .S(net902),
    .X(_08164_));
 sg13g2_nor2_1 _14867_ (.A(net905),
    .B(net776),
    .Y(_08165_));
 sg13g2_a22oi_1 _14868_ (.Y(_08166_),
    .B1(_08165_),
    .B2(\cpu.icache.r_tag[4][12] ),
    .A2(_08164_),
    .A1(net905));
 sg13g2_or2_1 _14869_ (.X(_08167_),
    .B(_08166_),
    .A(net701));
 sg13g2_nand4_1 _14870_ (.B(_08156_),
    .C(_08158_),
    .A(net410),
    .Y(_08168_),
    .D(_08167_));
 sg13g2_o21ai_1 _14871_ (.B1(_08168_),
    .Y(_08169_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net411));
 sg13g2_xnor2_1 _14872_ (.Y(_08170_),
    .A(net474),
    .B(_08169_));
 sg13g2_nand2_1 _14873_ (.Y(_08171_),
    .A(_08137_),
    .B(_08170_));
 sg13g2_buf_4 _14874_ (.X(_08172_),
    .A(_00192_));
 sg13g2_buf_2 _14875_ (.A(_08172_),
    .X(_08173_));
 sg13g2_buf_2 _14876_ (.A(_08055_),
    .X(_08174_));
 sg13g2_buf_2 _14877_ (.A(_08174_),
    .X(_08175_));
 sg13g2_buf_1 _14878_ (.A(net1095),
    .X(_08176_));
 sg13g2_buf_1 _14879_ (.A(_08176_),
    .X(_08177_));
 sg13g2_buf_1 _14880_ (.A(_08177_),
    .X(_08178_));
 sg13g2_mux4_1 _14881_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net774),
    .X(_08179_));
 sg13g2_mux4_1 _14882_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net774),
    .X(_08180_));
 sg13g2_mux4_1 _14883_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net774),
    .X(_08181_));
 sg13g2_mux4_1 _14884_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net774),
    .X(_08182_));
 sg13g2_buf_2 _14885_ (.A(net908),
    .X(_08183_));
 sg13g2_buf_1 _14886_ (.A(net1040),
    .X(_08184_));
 sg13g2_mux4_1 _14887_ (.S0(net773),
    .A0(_08179_),
    .A1(_08180_),
    .A2(_08181_),
    .A3(_08182_),
    .S1(net899),
    .X(_08185_));
 sg13g2_mux4_1 _14888_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net774),
    .X(_08186_));
 sg13g2_mux4_1 _14889_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net774),
    .X(_08187_));
 sg13g2_buf_2 _14890_ (.A(_08056_),
    .X(_08188_));
 sg13g2_buf_1 _14891_ (.A(_08059_),
    .X(_08189_));
 sg13g2_mux4_1 _14892_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net897),
    .X(_08190_));
 sg13g2_mux4_1 _14893_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net897),
    .X(_08191_));
 sg13g2_mux4_1 _14894_ (.S0(net773),
    .A0(_08186_),
    .A1(_08187_),
    .A2(_08190_),
    .A3(_08191_),
    .S1(net899),
    .X(_08192_));
 sg13g2_buf_1 _14895_ (.A(net1039),
    .X(_08193_));
 sg13g2_mux2_1 _14896_ (.A0(_08185_),
    .A1(_08192_),
    .S(net896),
    .X(_08194_));
 sg13g2_nand2b_1 _14897_ (.Y(_08195_),
    .B(_08194_),
    .A_N(net1034));
 sg13g2_buf_1 _14898_ (.A(_08195_),
    .X(_08196_));
 sg13g2_nor2_1 _14899_ (.A(net1092),
    .B(net1093),
    .Y(_08197_));
 sg13g2_and2_1 _14900_ (.A(_08094_),
    .B(_08197_),
    .X(_08198_));
 sg13g2_buf_2 _14901_ (.A(_08198_),
    .X(_08199_));
 sg13g2_buf_1 _14902_ (.A(_08199_),
    .X(_08200_));
 sg13g2_a22oi_1 _14903_ (.Y(_08201_),
    .B1(net700),
    .B2(\cpu.icache.r_tag[5][18] ),
    .A2(net475),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_nor3_2 _14904_ (.A(_08094_),
    .B(net1092),
    .C(net1093),
    .Y(_08202_));
 sg13g2_buf_1 _14905_ (.A(_08202_),
    .X(_08203_));
 sg13g2_buf_1 _14906_ (.A(net895),
    .X(_08204_));
 sg13g2_buf_1 _14907_ (.A(_08204_),
    .X(_08205_));
 sg13g2_a22oi_1 _14908_ (.Y(_08206_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][18] ),
    .A2(net544),
    .A1(\cpu.icache.r_tag[6][18] ));
 sg13g2_buf_1 _14909_ (.A(_08125_),
    .X(_08207_));
 sg13g2_buf_1 _14910_ (.A(net698),
    .X(_08208_));
 sg13g2_nor2_1 _14911_ (.A(net1093),
    .B(_08129_),
    .Y(_08209_));
 sg13g2_buf_1 _14912_ (.A(_08209_),
    .X(_08210_));
 sg13g2_and2_1 _14913_ (.A(\cpu.icache.r_tag[7][18] ),
    .B(net697),
    .X(_08211_));
 sg13g2_a221oi_1 _14914_ (.B2(\cpu.icache.r_tag[3][18] ),
    .C1(_08211_),
    .B1(net545),
    .A1(\cpu.icache.r_tag[1][18] ),
    .Y(_08212_),
    .A2(net596));
 sg13g2_nand4_1 _14915_ (.B(_08201_),
    .C(_08206_),
    .A(net410),
    .Y(_08213_),
    .D(_08212_));
 sg13g2_o21ai_1 _14916_ (.B1(_08213_),
    .Y(_08214_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net411));
 sg13g2_xnor2_1 _14917_ (.Y(_08215_),
    .A(net409),
    .B(_08214_));
 sg13g2_mux4_1 _14918_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net774),
    .X(_08216_));
 sg13g2_mux4_1 _14919_ (.S0(net901),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net774),
    .X(_08217_));
 sg13g2_mux4_1 _14920_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net897),
    .X(_08218_));
 sg13g2_mux4_1 _14921_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(net897),
    .X(_08219_));
 sg13g2_mux4_1 _14922_ (.S0(net773),
    .A0(_08216_),
    .A1(_08217_),
    .A2(_08218_),
    .A3(_08219_),
    .S1(net899),
    .X(_08220_));
 sg13g2_mux4_1 _14923_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net897),
    .X(_08221_));
 sg13g2_mux4_1 _14924_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net897),
    .X(_08222_));
 sg13g2_mux4_1 _14925_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net913),
    .X(_08223_));
 sg13g2_mux4_1 _14926_ (.S0(_08057_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(_08060_),
    .X(_08224_));
 sg13g2_mux4_1 _14927_ (.S0(net773),
    .A0(_08221_),
    .A1(_08222_),
    .A2(_08223_),
    .A3(_08224_),
    .S1(net899),
    .X(_08225_));
 sg13g2_mux2_1 _14928_ (.A0(_08220_),
    .A1(_08225_),
    .S(net896),
    .X(_08226_));
 sg13g2_nand2b_1 _14929_ (.Y(_08227_),
    .B(_08226_),
    .A_N(net1034));
 sg13g2_buf_1 _14930_ (.A(_08227_),
    .X(_08228_));
 sg13g2_buf_1 _14931_ (.A(_08119_),
    .X(_08229_));
 sg13g2_buf_1 _14932_ (.A(net543),
    .X(_08230_));
 sg13g2_a22oi_1 _14933_ (.Y(_08231_),
    .B1(net599),
    .B2(\cpu.icache.r_tag[1][21] ),
    .A2(net472),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_a22oi_1 _14934_ (.Y(_08232_),
    .B1(net700),
    .B2(\cpu.icache.r_tag[5][21] ),
    .A2(net544),
    .A1(\cpu.icache.r_tag[6][21] ));
 sg13g2_mux2_1 _14935_ (.A0(\cpu.icache.r_tag[7][21] ),
    .A1(\cpu.icache.r_tag[3][21] ),
    .S(net775),
    .X(_08233_));
 sg13g2_nor2_1 _14936_ (.A(_08123_),
    .B(_08090_),
    .Y(_08234_));
 sg13g2_buf_2 _14937_ (.A(_08234_),
    .X(_08235_));
 sg13g2_buf_1 _14938_ (.A(_08235_),
    .X(_08236_));
 sg13g2_a22oi_1 _14939_ (.Y(_08237_),
    .B1(_08233_),
    .B2(net696),
    .A2(net772),
    .A1(\cpu.icache.r_tag[4][21] ));
 sg13g2_nand4_1 _14940_ (.B(_08231_),
    .C(_08232_),
    .A(net477),
    .Y(_08238_),
    .D(_08237_));
 sg13g2_o21ai_1 _14941_ (.B1(_08238_),
    .Y(_08239_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net411));
 sg13g2_xnor2_1 _14942_ (.Y(_08240_),
    .A(net408),
    .B(_08239_));
 sg13g2_mux4_1 _14943_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(net897),
    .X(_08241_));
 sg13g2_mux4_1 _14944_ (.S0(net898),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net897),
    .X(_08242_));
 sg13g2_mux4_1 _14945_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(net909),
    .X(_08243_));
 sg13g2_mux4_1 _14946_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net913),
    .X(_08244_));
 sg13g2_mux4_1 _14947_ (.S0(net773),
    .A0(_08241_),
    .A1(_08242_),
    .A2(_08243_),
    .A3(_08244_),
    .S1(net899),
    .X(_08245_));
 sg13g2_mux4_1 _14948_ (.S0(_08188_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(_08189_),
    .X(_08246_));
 sg13g2_mux4_1 _14949_ (.S0(_08188_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(_08189_),
    .X(_08247_));
 sg13g2_mux4_1 _14950_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net909),
    .X(_08248_));
 sg13g2_mux4_1 _14951_ (.S0(_08066_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(_08067_),
    .X(_08249_));
 sg13g2_mux4_1 _14952_ (.S0(_08183_),
    .A0(_08246_),
    .A1(_08247_),
    .A2(_08248_),
    .A3(_08249_),
    .S1(net899),
    .X(_08250_));
 sg13g2_mux2_1 _14953_ (.A0(_08245_),
    .A1(_08250_),
    .S(net896),
    .X(_08251_));
 sg13g2_nand2b_1 _14954_ (.Y(_08252_),
    .B(_08251_),
    .A_N(net1034));
 sg13g2_buf_1 _14955_ (.A(_08252_),
    .X(_08253_));
 sg13g2_a22oi_1 _14956_ (.Y(_08254_),
    .B1(net700),
    .B2(\cpu.icache.r_tag[5][22] ),
    .A2(net472),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_a22oi_1 _14957_ (.Y(_08255_),
    .B1(net545),
    .B2(\cpu.icache.r_tag[3][22] ),
    .A2(net596),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_mux2_1 _14958_ (.A0(\cpu.icache.r_tag[4][22] ),
    .A1(\cpu.icache.r_tag[6][22] ),
    .S(net902),
    .X(_08256_));
 sg13g2_buf_2 _14959_ (.A(_08123_),
    .X(_08257_));
 sg13g2_buf_1 _14960_ (.A(_08257_),
    .X(_08258_));
 sg13g2_a22oi_1 _14961_ (.Y(_08259_),
    .B1(_08256_),
    .B2(net771),
    .A2(net696),
    .A1(\cpu.icache.r_tag[7][22] ));
 sg13g2_or2_1 _14962_ (.X(_08260_),
    .B(_08259_),
    .A(net701));
 sg13g2_nand4_1 _14963_ (.B(_08254_),
    .C(_08255_),
    .A(net477),
    .Y(_08261_),
    .D(_08260_));
 sg13g2_o21ai_1 _14964_ (.B1(_08261_),
    .Y(_08262_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(net411));
 sg13g2_xnor2_1 _14965_ (.Y(_08263_),
    .A(net471),
    .B(_08262_));
 sg13g2_mux4_1 _14966_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net913),
    .X(_08264_));
 sg13g2_mux4_1 _14967_ (.S0(net914),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net913),
    .X(_08265_));
 sg13g2_mux4_1 _14968_ (.S0(net912),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net911),
    .X(_08266_));
 sg13g2_mux4_1 _14969_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(net909),
    .X(_08267_));
 sg13g2_mux4_1 _14970_ (.S0(net773),
    .A0(_08264_),
    .A1(_08265_),
    .A2(_08266_),
    .A3(_08267_),
    .S1(net907),
    .X(_08268_));
 sg13g2_mux4_1 _14971_ (.S0(_08066_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(_08067_),
    .X(_08269_));
 sg13g2_mux4_1 _14972_ (.S0(_08057_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(_08060_),
    .X(_08270_));
 sg13g2_mux4_1 _14973_ (.S0(_08063_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(_08064_),
    .X(_08271_));
 sg13g2_mux4_1 _14974_ (.S0(_08063_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(_08064_),
    .X(_08272_));
 sg13g2_mux4_1 _14975_ (.S0(net908),
    .A0(_08269_),
    .A1(_08270_),
    .A2(_08271_),
    .A3(_08272_),
    .S1(net907),
    .X(_08273_));
 sg13g2_mux2_1 _14976_ (.A0(_08268_),
    .A1(_08273_),
    .S(_08193_),
    .X(_08274_));
 sg13g2_nand2b_1 _14977_ (.Y(_08275_),
    .B(_08274_),
    .A_N(net1034));
 sg13g2_buf_1 _14978_ (.A(_08275_),
    .X(_08276_));
 sg13g2_a22oi_1 _14979_ (.Y(_08277_),
    .B1(net544),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(net596),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_a22oi_1 _14980_ (.Y(_08278_),
    .B1(net772),
    .B2(\cpu.icache.r_tag[4][16] ),
    .A2(net472),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_buf_1 _14981_ (.A(_08197_),
    .X(_08279_));
 sg13g2_mux2_1 _14982_ (.A0(\cpu.icache.r_tag[7][16] ),
    .A1(\cpu.icache.r_tag[3][16] ),
    .S(net903),
    .X(_08280_));
 sg13g2_a22oi_1 _14983_ (.Y(_08281_),
    .B1(_08280_),
    .B2(net703),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_buf_1 _14984_ (.A(net905),
    .X(_08282_));
 sg13g2_nand2b_1 _14985_ (.Y(_08283_),
    .B(net770),
    .A_N(_08281_));
 sg13g2_nand4_1 _14986_ (.B(_08277_),
    .C(_08278_),
    .A(net477),
    .Y(_08284_),
    .D(_08283_));
 sg13g2_o21ai_1 _14987_ (.B1(_08284_),
    .Y(_08285_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net411));
 sg13g2_xnor2_1 _14988_ (.Y(_08286_),
    .A(_08276_),
    .B(_08285_));
 sg13g2_nand4_1 _14989_ (.B(_08240_),
    .C(_08263_),
    .A(_08215_),
    .Y(_08287_),
    .D(_08286_));
 sg13g2_buf_2 _14990_ (.A(_08055_),
    .X(_08288_));
 sg13g2_buf_2 _14991_ (.A(net1031),
    .X(_08289_));
 sg13g2_buf_2 _14992_ (.A(_08289_),
    .X(_08290_));
 sg13g2_buf_2 _14993_ (.A(net1032),
    .X(_08291_));
 sg13g2_buf_1 _14994_ (.A(_08291_),
    .X(_08292_));
 sg13g2_mux4_1 _14995_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net768),
    .X(_08293_));
 sg13g2_mux4_1 _14996_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net768),
    .X(_08294_));
 sg13g2_mux4_1 _14997_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(net768),
    .X(_08295_));
 sg13g2_mux4_1 _14998_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net768),
    .X(_08296_));
 sg13g2_mux4_1 _14999_ (.S0(_08183_),
    .A0(_08293_),
    .A1(_08294_),
    .A2(_08295_),
    .A3(_08296_),
    .S1(net899),
    .X(_08297_));
 sg13g2_mux4_1 _15000_ (.S0(_08290_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(_08292_),
    .X(_08298_));
 sg13g2_mux4_1 _15001_ (.S0(_08290_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(_08292_),
    .X(_08299_));
 sg13g2_mux4_1 _15002_ (.S0(_08175_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(_08178_),
    .X(_08300_));
 sg13g2_mux4_1 _15003_ (.S0(_08175_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(_08178_),
    .X(_08301_));
 sg13g2_mux4_1 _15004_ (.S0(net773),
    .A0(_08298_),
    .A1(_08299_),
    .A2(_08300_),
    .A3(_08301_),
    .S1(net899),
    .X(_08302_));
 sg13g2_mux2_1 _15005_ (.A0(_08297_),
    .A1(_08302_),
    .S(_08193_),
    .X(_08303_));
 sg13g2_nand2b_1 _15006_ (.Y(_08304_),
    .B(_08303_),
    .A_N(net1034));
 sg13g2_buf_1 _15007_ (.A(_08304_),
    .X(_08305_));
 sg13g2_buf_1 _15008_ (.A(net903),
    .X(_08306_));
 sg13g2_mux2_1 _15009_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(net767),
    .X(_08307_));
 sg13g2_a22oi_1 _15010_ (.Y(_08308_),
    .B1(_08307_),
    .B2(net696),
    .A2(net772),
    .A1(\cpu.icache.r_tag[4][20] ));
 sg13g2_buf_1 _15011_ (.A(_08200_),
    .X(_08309_));
 sg13g2_a22oi_1 _15012_ (.Y(_08310_),
    .B1(net595),
    .B2(\cpu.icache.r_tag[5][20] ),
    .A2(net475),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_a22oi_1 _15013_ (.Y(_08311_),
    .B1(net544),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(net599),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_nand4_1 _15014_ (.B(_08308_),
    .C(_08310_),
    .A(net410),
    .Y(_08312_),
    .D(_08311_));
 sg13g2_o21ai_1 _15015_ (.B1(_08312_),
    .Y(_08313_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net411));
 sg13g2_xnor2_1 _15016_ (.Y(_08314_),
    .A(net407),
    .B(_08313_));
 sg13g2_mux4_1 _15017_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1032),
    .X(_08315_));
 sg13g2_mux4_1 _15018_ (.S0(_08288_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net1041),
    .X(_08316_));
 sg13g2_mux4_1 _15019_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1032),
    .X(_08317_));
 sg13g2_mux4_1 _15020_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(net1032),
    .X(_08318_));
 sg13g2_mux4_1 _15021_ (.S0(_08070_),
    .A0(_08315_),
    .A1(_08316_),
    .A2(_08317_),
    .A3(_08318_),
    .S1(net1040),
    .X(_08319_));
 sg13g2_mux4_1 _15022_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1032),
    .X(_08320_));
 sg13g2_mux4_1 _15023_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net1032),
    .X(_08321_));
 sg13g2_mux4_1 _15024_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(_08176_),
    .X(_08322_));
 sg13g2_mux4_1 _15025_ (.S0(net1031),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net1032),
    .X(_08323_));
 sg13g2_mux4_1 _15026_ (.S0(_08070_),
    .A0(_08320_),
    .A1(_08321_),
    .A2(_08322_),
    .A3(_08323_),
    .S1(net1040),
    .X(_08324_));
 sg13g2_mux2_1 _15027_ (.A0(_08319_),
    .A1(_08324_),
    .S(net1039),
    .X(_08325_));
 sg13g2_nand2b_2 _15028_ (.Y(_08326_),
    .B(_08325_),
    .A_N(net1034));
 sg13g2_buf_1 _15029_ (.A(_08326_),
    .X(_08327_));
 sg13g2_a22oi_1 _15030_ (.Y(_08328_),
    .B1(net772),
    .B2(\cpu.icache.r_tag[4][23] ),
    .A2(net544),
    .A1(\cpu.icache.r_tag[6][23] ));
 sg13g2_a22oi_1 _15031_ (.Y(_08329_),
    .B1(net596),
    .B2(\cpu.icache.r_tag[1][23] ),
    .A2(net472),
    .A1(\cpu.icache.r_tag[2][23] ));
 sg13g2_mux2_1 _15032_ (.A0(\cpu.icache.r_tag[7][23] ),
    .A1(\cpu.icache.r_tag[3][23] ),
    .S(net1035),
    .X(_08330_));
 sg13g2_a22oi_1 _15033_ (.Y(_08331_),
    .B1(_08330_),
    .B2(net776),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][23] ));
 sg13g2_nand2b_1 _15034_ (.Y(_08332_),
    .B(net770),
    .A_N(_08331_));
 sg13g2_nand4_1 _15035_ (.B(_08328_),
    .C(_08329_),
    .A(net476),
    .Y(_08333_),
    .D(_08332_));
 sg13g2_o21ai_1 _15036_ (.B1(_08333_),
    .Y(_08334_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net477));
 sg13g2_xor2_1 _15037_ (.B(_08334_),
    .A(net542),
    .X(_08335_));
 sg13g2_buf_2 _15038_ (.A(_08288_),
    .X(_08336_));
 sg13g2_buf_1 _15039_ (.A(net1032),
    .X(_08337_));
 sg13g2_mux4_1 _15040_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net889),
    .X(_08338_));
 sg13g2_mux4_1 _15041_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net889),
    .X(_08339_));
 sg13g2_mux4_1 _15042_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net891),
    .X(_08340_));
 sg13g2_mux4_1 _15043_ (.S0(_08289_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(_08291_),
    .X(_08341_));
 sg13g2_mux4_1 _15044_ (.S0(net1094),
    .A0(_08338_),
    .A1(_08339_),
    .A2(_08340_),
    .A3(_08341_),
    .S1(_08082_),
    .X(_08342_));
 sg13g2_a21oi_1 _15045_ (.A1(net1042),
    .A2(_08342_),
    .Y(_08343_),
    .B1(_08184_));
 sg13g2_inv_2 _15046_ (.Y(_08344_),
    .A(_08073_));
 sg13g2_inv_2 _15047_ (.Y(_08345_),
    .A(net1096));
 sg13g2_mux4_1 _15048_ (.S0(_08336_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(_08337_),
    .X(_08346_));
 sg13g2_mux4_1 _15049_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net889),
    .X(_08347_));
 sg13g2_mux4_1 _15050_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net889),
    .X(_08348_));
 sg13g2_mux4_1 _15051_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net889),
    .X(_08349_));
 sg13g2_mux4_1 _15052_ (.S0(net1094),
    .A0(_08346_),
    .A1(_08347_),
    .A2(_08348_),
    .A3(_08349_),
    .S1(net1039),
    .X(_08350_));
 sg13g2_nor3_1 _15053_ (.A(_08344_),
    .B(_08345_),
    .C(_08350_),
    .Y(_08351_));
 sg13g2_or2_1 _15054_ (.X(_08352_),
    .B(_08351_),
    .A(_08343_));
 sg13g2_buf_1 _15055_ (.A(_08352_),
    .X(_08353_));
 sg13g2_a22oi_1 _15056_ (.Y(_08354_),
    .B1(\cpu.icache.r_tag[1][14] ),
    .B2(_08093_),
    .A2(\cpu.icache.r_tag[5][14] ),
    .A1(net777));
 sg13g2_nor2_2 _15057_ (.A(_08090_),
    .B(_08105_),
    .Y(_08355_));
 sg13g2_nand2_1 _15058_ (.Y(_08356_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(_08355_));
 sg13g2_o21ai_1 _15059_ (.B1(_08356_),
    .Y(_08357_),
    .A1(net703),
    .A2(_08354_));
 sg13g2_mux2_1 _15060_ (.A0(\cpu.icache.r_tag[4][14] ),
    .A1(\cpu.icache.r_tag[6][14] ),
    .S(net902),
    .X(_08358_));
 sg13g2_a22oi_1 _15061_ (.Y(_08359_),
    .B1(_08358_),
    .B2(net771),
    .A2(net696),
    .A1(\cpu.icache.r_tag[7][14] ));
 sg13g2_and2_1 _15062_ (.A(net1035),
    .B(_08096_),
    .X(_08360_));
 sg13g2_buf_1 _15063_ (.A(_08360_),
    .X(_08361_));
 sg13g2_buf_1 _15064_ (.A(_08361_),
    .X(_08362_));
 sg13g2_nand2_1 _15065_ (.Y(_08363_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net541));
 sg13g2_o21ai_1 _15066_ (.B1(_08363_),
    .Y(_08364_),
    .A1(net701),
    .A2(_08359_));
 sg13g2_a221oi_1 _15067_ (.B2(net770),
    .C1(_08364_),
    .B1(_08357_),
    .A1(\cpu.icache.r_tag[2][14] ),
    .Y(_08365_),
    .A2(net475));
 sg13g2_xor2_1 _15068_ (.B(_08365_),
    .A(net469),
    .X(_08366_));
 sg13g2_nor2_1 _15069_ (.A(_08335_),
    .B(_08366_),
    .Y(_08367_));
 sg13g2_mux4_1 _15070_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(net891),
    .X(_08368_));
 sg13g2_mux4_1 _15071_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net891),
    .X(_08369_));
 sg13g2_mux4_1 _15072_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net900),
    .X(_08370_));
 sg13g2_mux4_1 _15073_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net900),
    .X(_08371_));
 sg13g2_mux4_1 _15074_ (.S0(net908),
    .A0(_08368_),
    .A1(_08369_),
    .A2(_08370_),
    .A3(_08371_),
    .S1(net907),
    .X(_08372_));
 sg13g2_mux4_1 _15075_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net900),
    .X(_08373_));
 sg13g2_mux4_1 _15076_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net900),
    .X(_08374_));
 sg13g2_mux4_1 _15077_ (.S0(_08056_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net1041),
    .X(_08375_));
 sg13g2_mux4_1 _15078_ (.S0(_08056_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net1041),
    .X(_08376_));
 sg13g2_mux4_1 _15079_ (.S0(_08071_),
    .A0(_08373_),
    .A1(_08374_),
    .A2(_08375_),
    .A3(_08376_),
    .S1(_08074_),
    .X(_08377_));
 sg13g2_mux2_1 _15080_ (.A0(_08372_),
    .A1(_08377_),
    .S(net1039),
    .X(_08378_));
 sg13g2_nand2b_1 _15081_ (.Y(_08379_),
    .B(_08378_),
    .A_N(net1034));
 sg13g2_buf_1 _15082_ (.A(_08379_),
    .X(_08380_));
 sg13g2_a22oi_1 _15083_ (.Y(_08381_),
    .B1(net697),
    .B2(\cpu.icache.r_tag[7][19] ),
    .A2(net546),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_a22oi_1 _15084_ (.Y(_08382_),
    .B1(net545),
    .B2(\cpu.icache.r_tag[3][19] ),
    .A2(net702),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_nor2_2 _15085_ (.A(net894),
    .B(net1036),
    .Y(_08383_));
 sg13g2_mux2_1 _15086_ (.A0(\cpu.icache.r_tag[4][19] ),
    .A1(\cpu.icache.r_tag[6][19] ),
    .S(net904),
    .X(_08384_));
 sg13g2_buf_1 _15087_ (.A(net894),
    .X(_08385_));
 sg13g2_a22oi_1 _15088_ (.Y(_08386_),
    .B1(_08384_),
    .B2(net766),
    .A2(_08383_),
    .A1(\cpu.icache.r_tag[5][19] ));
 sg13g2_or2_1 _15089_ (.X(_08387_),
    .B(_08386_),
    .A(net775));
 sg13g2_nand4_1 _15090_ (.B(_08381_),
    .C(_08382_),
    .A(net476),
    .Y(_08388_),
    .D(_08387_));
 sg13g2_o21ai_1 _15091_ (.B1(_08388_),
    .Y(_08389_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(net477));
 sg13g2_xor2_1 _15092_ (.B(_08389_),
    .A(net468),
    .X(_08390_));
 sg13g2_mux4_1 _15093_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net900),
    .X(_08391_));
 sg13g2_mux4_1 _15094_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net891),
    .X(_08392_));
 sg13g2_mux4_1 _15095_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net900),
    .X(_08393_));
 sg13g2_mux4_1 _15096_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net900),
    .X(_08394_));
 sg13g2_mux4_1 _15097_ (.S0(net908),
    .A0(_08391_),
    .A1(_08392_),
    .A2(_08393_),
    .A3(_08394_),
    .S1(net907),
    .X(_08395_));
 sg13g2_mux4_1 _15098_ (.S0(_08174_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(_08177_),
    .X(_08396_));
 sg13g2_mux4_1 _15099_ (.S0(net1033),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net900),
    .X(_08397_));
 sg13g2_mux4_1 _15100_ (.S0(_08056_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net1041),
    .X(_08398_));
 sg13g2_mux4_1 _15101_ (.S0(_08056_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net1041),
    .X(_08399_));
 sg13g2_mux4_1 _15102_ (.S0(_08071_),
    .A0(_08396_),
    .A1(_08397_),
    .A2(_08398_),
    .A3(_08399_),
    .S1(_08074_),
    .X(_08400_));
 sg13g2_mux2_1 _15103_ (.A0(_08395_),
    .A1(_08400_),
    .S(net1039),
    .X(_08401_));
 sg13g2_nand2b_1 _15104_ (.Y(_08402_),
    .B(_08401_),
    .A_N(net1034));
 sg13g2_buf_1 _15105_ (.A(_08402_),
    .X(_08403_));
 sg13g2_nand2_1 _15106_ (.Y(_08404_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net596));
 sg13g2_a22oi_1 _15107_ (.Y(_08405_),
    .B1(net772),
    .B2(\cpu.icache.r_tag[4][17] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[7][17] ));
 sg13g2_a22oi_1 _15108_ (.Y(_08406_),
    .B1(_08355_),
    .B2(\cpu.icache.r_tag[3][17] ),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][17] ));
 sg13g2_nor2_1 _15109_ (.A(net766),
    .B(_08406_),
    .Y(_08407_));
 sg13g2_a221oi_1 _15110_ (.B2(\cpu.icache.r_tag[6][17] ),
    .C1(_08407_),
    .B1(net544),
    .A1(\cpu.icache.r_tag[2][17] ),
    .Y(_08408_),
    .A2(net546));
 sg13g2_nand4_1 _15111_ (.B(_08404_),
    .C(_08405_),
    .A(net476),
    .Y(_08409_),
    .D(_08408_));
 sg13g2_o21ai_1 _15112_ (.B1(_08409_),
    .Y(_08410_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(net477));
 sg13g2_xor2_1 _15113_ (.B(_08410_),
    .A(net467),
    .X(_08411_));
 sg13g2_mux4_1 _15114_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net891),
    .X(_08412_));
 sg13g2_mux4_1 _15115_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net891),
    .X(_08413_));
 sg13g2_mux4_1 _15116_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net891),
    .X(_08414_));
 sg13g2_mux4_1 _15117_ (.S0(net892),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net891),
    .X(_08415_));
 sg13g2_mux4_1 _15118_ (.S0(net1040),
    .A0(_08412_),
    .A1(_08413_),
    .A2(_08414_),
    .A3(_08415_),
    .S1(net1039),
    .X(_08416_));
 sg13g2_a21oi_1 _15119_ (.A1(net1042),
    .A2(_08416_),
    .Y(_08417_),
    .B1(net1094));
 sg13g2_mux4_1 _15120_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(net889),
    .X(_08418_));
 sg13g2_mux4_1 _15121_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net889),
    .X(_08419_));
 sg13g2_mux4_1 _15122_ (.S0(_08336_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(_08337_),
    .X(_08420_));
 sg13g2_mux4_1 _15123_ (.S0(net890),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net889),
    .X(_08421_));
 sg13g2_mux4_1 _15124_ (.S0(net1040),
    .A0(_08418_),
    .A1(_08419_),
    .A2(_08420_),
    .A3(_08421_),
    .S1(net1039),
    .X(_08422_));
 sg13g2_nor3_1 _15125_ (.A(net773),
    .B(_08345_),
    .C(_08422_),
    .Y(_08423_));
 sg13g2_or2_1 _15126_ (.X(_08424_),
    .B(_08423_),
    .A(_08417_));
 sg13g2_buf_1 _15127_ (.A(_08424_),
    .X(_08425_));
 sg13g2_a22oi_1 _15128_ (.Y(_08426_),
    .B1(net700),
    .B2(\cpu.icache.r_tag[5][15] ),
    .A2(net472),
    .A1(\cpu.icache.r_tag[2][15] ));
 sg13g2_a22oi_1 _15129_ (.Y(_08427_),
    .B1(net545),
    .B2(\cpu.icache.r_tag[3][15] ),
    .A2(net702),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_mux2_1 _15130_ (.A0(\cpu.icache.r_tag[4][15] ),
    .A1(\cpu.icache.r_tag[6][15] ),
    .S(net904),
    .X(_08428_));
 sg13g2_a22oi_1 _15131_ (.Y(_08429_),
    .B1(_08428_),
    .B2(net766),
    .A2(_08236_),
    .A1(\cpu.icache.r_tag[7][15] ));
 sg13g2_or2_1 _15132_ (.X(_08430_),
    .B(_08429_),
    .A(net767));
 sg13g2_nand4_1 _15133_ (.B(_08426_),
    .C(_08427_),
    .A(net476),
    .Y(_08431_),
    .D(_08430_));
 sg13g2_o21ai_1 _15134_ (.B1(_08431_),
    .Y(_08432_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net477));
 sg13g2_xor2_1 _15135_ (.B(_08432_),
    .A(net466),
    .X(_08433_));
 sg13g2_nor3_1 _15136_ (.A(_08390_),
    .B(_08411_),
    .C(_08433_),
    .Y(_08434_));
 sg13g2_buf_1 _15137_ (.A(\cpu.ex.pc[6] ),
    .X(_08435_));
 sg13g2_nand2_1 _15138_ (.Y(_08436_),
    .A(\cpu.icache.r_tag[1][6] ),
    .B(net698));
 sg13g2_a22oi_1 _15139_ (.Y(_08437_),
    .B1(net895),
    .B2(\cpu.icache.r_tag[4][6] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[7][6] ));
 sg13g2_buf_1 _15140_ (.A(_08119_),
    .X(_08438_));
 sg13g2_a22oi_1 _15141_ (.Y(_08439_),
    .B1(_08355_),
    .B2(\cpu.icache.r_tag[3][6] ),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_nor2_1 _15142_ (.A(net894),
    .B(_08439_),
    .Y(_08440_));
 sg13g2_a221oi_1 _15143_ (.B2(\cpu.icache.r_tag[6][6] ),
    .C1(_08440_),
    .B1(net597),
    .A1(\cpu.icache.r_tag[2][6] ),
    .Y(_08441_),
    .A2(net540));
 sg13g2_nand4_1 _15144_ (.B(_08436_),
    .C(_08437_),
    .A(net548),
    .Y(_08442_),
    .D(_08441_));
 sg13g2_o21ai_1 _15145_ (.B1(_08442_),
    .Y(_08443_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net476));
 sg13g2_xor2_1 _15146_ (.B(_08443_),
    .A(_08435_),
    .X(_08444_));
 sg13g2_inv_1 _15147_ (.Y(_08445_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15148_ (.A(_08445_),
    .X(_08446_));
 sg13g2_buf_1 _15149_ (.A(_08098_),
    .X(_08447_));
 sg13g2_nand2_1 _15150_ (.Y(_08448_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(net597));
 sg13g2_a22oi_1 _15151_ (.Y(_08449_),
    .B1(net697),
    .B2(\cpu.icache.r_tag[7][11] ),
    .A2(net543),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_buf_1 _15152_ (.A(_08125_),
    .X(_08450_));
 sg13g2_a22oi_1 _15153_ (.Y(_08451_),
    .B1(_08355_),
    .B2(\cpu.icache.r_tag[3][11] ),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][11] ));
 sg13g2_nor2_1 _15154_ (.A(net894),
    .B(_08451_),
    .Y(_08452_));
 sg13g2_a221oi_1 _15155_ (.B2(\cpu.icache.r_tag[4][11] ),
    .C1(_08452_),
    .B1(net895),
    .A1(\cpu.icache.r_tag[1][11] ),
    .Y(_08453_),
    .A2(_08450_));
 sg13g2_nand4_1 _15156_ (.B(_08448_),
    .C(_08449_),
    .A(net548),
    .Y(_08454_),
    .D(_08453_));
 sg13g2_o21ai_1 _15157_ (.B1(_08454_),
    .Y(_08455_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net539));
 sg13g2_xnor2_1 _15158_ (.Y(_08456_),
    .A(net1030),
    .B(_08455_));
 sg13g2_mux4_1 _15159_ (.S0(net770),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net703),
    .X(_08457_));
 sg13g2_mux4_1 _15160_ (.S0(net770),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net703),
    .X(_08458_));
 sg13g2_mux2_1 _15161_ (.A0(_08457_),
    .A1(_08458_),
    .S(_08093_),
    .X(_08459_));
 sg13g2_buf_1 _15162_ (.A(\cpu.ex.pc[9] ),
    .X(_08460_));
 sg13g2_inv_1 _15163_ (.Y(_08461_),
    .A(_08460_));
 sg13g2_buf_1 _15164_ (.A(_08461_),
    .X(_08462_));
 sg13g2_a22oi_1 _15165_ (.Y(_08463_),
    .B1(_08199_),
    .B2(\cpu.icache.r_tag[5][9] ),
    .A2(net698),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_a22oi_1 _15166_ (.Y(_08464_),
    .B1(net895),
    .B2(\cpu.icache.r_tag[4][9] ),
    .A2(net543),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_mux2_1 _15167_ (.A0(\cpu.icache.r_tag[7][9] ),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(net1093),
    .X(_08465_));
 sg13g2_nor2_1 _15168_ (.A(net1037),
    .B(net1035),
    .Y(_08466_));
 sg13g2_a22oi_1 _15169_ (.Y(_08467_),
    .B1(_08466_),
    .B2(\cpu.icache.r_tag[6][9] ),
    .A2(_08465_),
    .A1(net1037));
 sg13g2_nand2b_1 _15170_ (.Y(_08468_),
    .B(net776),
    .A_N(_08467_));
 sg13g2_nand4_1 _15171_ (.B(_08463_),
    .C(_08464_),
    .A(net547),
    .Y(_08469_),
    .D(_08468_));
 sg13g2_o21ai_1 _15172_ (.B1(_08469_),
    .Y(_08470_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net539));
 sg13g2_xnor2_1 _15173_ (.Y(_08471_),
    .A(net888),
    .B(_08470_));
 sg13g2_nand4_1 _15174_ (.B(_08456_),
    .C(_08459_),
    .A(_08444_),
    .Y(_08472_),
    .D(_08471_));
 sg13g2_inv_1 _15175_ (.Y(_08473_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_nand2_1 _15176_ (.Y(_08474_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net702));
 sg13g2_a22oi_1 _15177_ (.Y(_08475_),
    .B1(net895),
    .B2(\cpu.icache.r_tag[4][8] ),
    .A2(net697),
    .A1(\cpu.icache.r_tag[7][8] ));
 sg13g2_a22oi_1 _15178_ (.Y(_08476_),
    .B1(_08355_),
    .B2(\cpu.icache.r_tag[3][8] ),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][8] ));
 sg13g2_nor2_1 _15179_ (.A(net894),
    .B(_08476_),
    .Y(_08477_));
 sg13g2_a221oi_1 _15180_ (.B2(\cpu.icache.r_tag[6][8] ),
    .C1(_08477_),
    .B1(net597),
    .A1(\cpu.icache.r_tag[2][8] ),
    .Y(_08478_),
    .A2(net540));
 sg13g2_nand4_1 _15181_ (.B(_08474_),
    .C(_08475_),
    .A(net548),
    .Y(_08479_),
    .D(_08478_));
 sg13g2_o21ai_1 _15182_ (.B1(_08479_),
    .Y(_08480_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net476));
 sg13g2_xnor2_1 _15183_ (.Y(_08481_),
    .A(_08473_),
    .B(_08480_));
 sg13g2_buf_2 _15184_ (.A(\cpu.ex.pc[5] ),
    .X(_08482_));
 sg13g2_a22oi_1 _15185_ (.Y(_08483_),
    .B1(_08199_),
    .B2(\cpu.icache.r_tag[5][5] ),
    .A2(net698),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_a22oi_1 _15186_ (.Y(_08484_),
    .B1(net597),
    .B2(\cpu.icache.r_tag[6][5] ),
    .A2(net543),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_mux2_1 _15187_ (.A0(\cpu.icache.r_tag[7][5] ),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net1035),
    .X(_08485_));
 sg13g2_a22oi_1 _15188_ (.Y(_08486_),
    .B1(_08485_),
    .B2(net696),
    .A2(net895),
    .A1(\cpu.icache.r_tag[4][5] ));
 sg13g2_nand4_1 _15189_ (.B(_08483_),
    .C(_08484_),
    .A(net548),
    .Y(_08487_),
    .D(_08486_));
 sg13g2_o21ai_1 _15190_ (.B1(_08487_),
    .Y(_08488_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net539));
 sg13g2_xor2_1 _15191_ (.B(_08488_),
    .A(_08482_),
    .X(_08489_));
 sg13g2_buf_1 _15192_ (.A(\cpu.ex.pc[10] ),
    .X(_08490_));
 sg13g2_a22oi_1 _15193_ (.Y(_08491_),
    .B1(net895),
    .B2(\cpu.icache.r_tag[4][10] ),
    .A2(net543),
    .A1(\cpu.icache.r_tag[2][10] ));
 sg13g2_a22oi_1 _15194_ (.Y(_08492_),
    .B1(net597),
    .B2(\cpu.icache.r_tag[6][10] ),
    .A2(net698),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_mux2_1 _15195_ (.A0(\cpu.icache.r_tag[7][10] ),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net1093),
    .X(_08493_));
 sg13g2_a22oi_1 _15196_ (.Y(_08494_),
    .B1(_08493_),
    .B2(net902),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][10] ));
 sg13g2_nand2b_1 _15197_ (.Y(_08495_),
    .B(net905),
    .A_N(_08494_));
 sg13g2_nand4_1 _15198_ (.B(_08491_),
    .C(_08492_),
    .A(net547),
    .Y(_08496_),
    .D(_08495_));
 sg13g2_o21ai_1 _15199_ (.B1(_08496_),
    .Y(_08497_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net539));
 sg13g2_xor2_1 _15200_ (.B(_08497_),
    .A(_08490_),
    .X(_08498_));
 sg13g2_inv_1 _15201_ (.Y(_08499_),
    .A(\cpu.ex.pc[7] ));
 sg13g2_buf_1 _15202_ (.A(_08499_),
    .X(_08500_));
 sg13g2_a22oi_1 _15203_ (.Y(_08501_),
    .B1(net895),
    .B2(\cpu.icache.r_tag[4][7] ),
    .A2(net597),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_a22oi_1 _15204_ (.Y(_08502_),
    .B1(net698),
    .B2(\cpu.icache.r_tag[1][7] ),
    .A2(net543),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_mux2_1 _15205_ (.A0(\cpu.icache.r_tag[7][7] ),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net1093),
    .X(_08503_));
 sg13g2_a22oi_1 _15206_ (.Y(_08504_),
    .B1(_08503_),
    .B2(net902),
    .A2(net893),
    .A1(\cpu.icache.r_tag[5][7] ));
 sg13g2_nand2b_1 _15207_ (.Y(_08505_),
    .B(net905),
    .A_N(_08504_));
 sg13g2_nand4_1 _15208_ (.B(_08501_),
    .C(_08502_),
    .A(net548),
    .Y(_08506_),
    .D(_08505_));
 sg13g2_o21ai_1 _15209_ (.B1(_08506_),
    .Y(_08507_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net539));
 sg13g2_xnor2_1 _15210_ (.Y(_08508_),
    .A(net1029),
    .B(_08507_));
 sg13g2_nand4_1 _15211_ (.B(_08489_),
    .C(_08498_),
    .A(_08481_),
    .Y(_08509_),
    .D(_08508_));
 sg13g2_nor2_1 _15212_ (.A(_08472_),
    .B(_08509_),
    .Y(_08510_));
 sg13g2_nand4_1 _15213_ (.B(_08367_),
    .C(_08434_),
    .A(_08314_),
    .Y(_08511_),
    .D(_08510_));
 sg13g2_or3_1 _15214_ (.A(_08171_),
    .B(_08287_),
    .C(_08511_),
    .X(_08512_));
 sg13g2_inv_1 _15215_ (.Y(_08513_),
    .A(_00189_));
 sg13g2_buf_2 _15216_ (.A(_00193_),
    .X(_08514_));
 sg13g2_buf_8 _15217_ (.A(\cpu.ex.ifetch ),
    .X(_08515_));
 sg13g2_buf_1 _15218_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08516_));
 sg13g2_nor2b_1 _15219_ (.A(_08515_),
    .B_N(_08516_),
    .Y(_08517_));
 sg13g2_buf_1 _15220_ (.A(_08517_),
    .X(_08518_));
 sg13g2_nor2_1 _15221_ (.A(_08514_),
    .B(_08518_),
    .Y(_08519_));
 sg13g2_buf_16 _15222_ (.X(_08520_),
    .A(\cpu.addr[13] ));
 sg13g2_buf_2 _15223_ (.A(\cpu.addr[14] ),
    .X(_08521_));
 sg13g2_buf_8 _15224_ (.A(_08521_),
    .X(_08522_));
 sg13g2_mux4_1 _15225_ (.S0(_08520_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .S1(net1028),
    .X(_08523_));
 sg13g2_mux4_1 _15226_ (.S0(_08520_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .S1(net1028),
    .X(_08524_));
 sg13g2_mux4_1 _15227_ (.S0(_08520_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(_08521_),
    .X(_08525_));
 sg13g2_mux4_1 _15228_ (.S0(_08520_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net1028),
    .X(_08526_));
 sg13g2_buf_8 _15229_ (.A(\cpu.addr[15] ),
    .X(_08527_));
 sg13g2_inv_1 _15230_ (.Y(_08528_),
    .A(_08527_));
 sg13g2_buf_4 _15231_ (.X(_08529_),
    .A(_08528_));
 sg13g2_buf_8 _15232_ (.A(\cpu.addr[12] ),
    .X(_08530_));
 sg13g2_buf_8 _15233_ (.A(_08530_),
    .X(_08531_));
 sg13g2_mux4_1 _15234_ (.S0(_08529_),
    .A0(_08523_),
    .A1(_08524_),
    .A2(_08525_),
    .A3(_08526_),
    .S1(net1027),
    .X(_08532_));
 sg13g2_nand2_1 _15235_ (.Y(_08533_),
    .A(_08519_),
    .B(_08532_));
 sg13g2_buf_2 _15236_ (.A(\cpu.ex.io_access ),
    .X(_08534_));
 sg13g2_buf_2 _15237_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08535_));
 sg13g2_nor2_2 _15238_ (.A(\cpu.ex.r_wmask[1] ),
    .B(_08535_),
    .Y(_08536_));
 sg13g2_nor3_2 _15239_ (.A(_08345_),
    .B(_08534_),
    .C(_08536_),
    .Y(_08537_));
 sg13g2_buf_8 _15240_ (.A(_08520_),
    .X(_08538_));
 sg13g2_mux4_1 _15241_ (.S0(net1026),
    .A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(net1028),
    .X(_08539_));
 sg13g2_nor2b_1 _15242_ (.A(_08539_),
    .B_N(_08530_),
    .Y(_08540_));
 sg13g2_mux2_1 _15243_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .S(_08521_),
    .X(_08541_));
 sg13g2_nor3_1 _15244_ (.A(_08530_),
    .B(net1026),
    .C(_08541_),
    .Y(_08542_));
 sg13g2_nand2b_1 _15245_ (.Y(_08543_),
    .B(net1026),
    .A_N(_08530_));
 sg13g2_mux2_1 _15246_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .S(net1028),
    .X(_08544_));
 sg13g2_nor2_1 _15247_ (.A(_08543_),
    .B(_08544_),
    .Y(_08545_));
 sg13g2_o21ai_1 _15248_ (.B1(_08529_),
    .Y(_08546_),
    .A1(_08514_),
    .A2(_08518_));
 sg13g2_or4_1 _15249_ (.A(_08540_),
    .B(_08542_),
    .C(_08545_),
    .D(_08546_),
    .X(_08547_));
 sg13g2_mux4_1 _15250_ (.S0(net1026),
    .A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(net1028),
    .X(_08548_));
 sg13g2_nor2b_1 _15251_ (.A(_08548_),
    .B_N(_08530_),
    .Y(_08549_));
 sg13g2_mux2_1 _15252_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .S(_08521_),
    .X(_08550_));
 sg13g2_nor3_1 _15253_ (.A(_08530_),
    .B(net1026),
    .C(_08550_),
    .Y(_08551_));
 sg13g2_mux2_1 _15254_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .S(net1028),
    .X(_08552_));
 sg13g2_nor2_1 _15255_ (.A(_08543_),
    .B(_08552_),
    .Y(_08553_));
 sg13g2_o21ai_1 _15256_ (.B1(_08527_),
    .Y(_08554_),
    .A1(_08514_),
    .A2(_08518_));
 sg13g2_or4_1 _15257_ (.A(_08549_),
    .B(_08551_),
    .C(_08553_),
    .D(_08554_),
    .X(_08555_));
 sg13g2_and4_1 _15258_ (.A(_08533_),
    .B(_08537_),
    .C(_08547_),
    .D(_08555_),
    .X(_08556_));
 sg13g2_buf_2 _15259_ (.A(_08556_),
    .X(_08557_));
 sg13g2_buf_1 _15260_ (.A(\cpu.ex.r_read_stall ),
    .X(_08558_));
 sg13g2_inv_1 _15261_ (.Y(_08559_),
    .A(\cpu.ex.r_wmask[1] ));
 sg13g2_inv_2 _15262_ (.Y(_08560_),
    .A(_08535_));
 sg13g2_nand2_2 _15263_ (.Y(_08561_),
    .A(_08559_),
    .B(_08560_));
 sg13g2_nor3_1 _15264_ (.A(_08513_),
    .B(_08558_),
    .C(_08561_),
    .Y(_08562_));
 sg13g2_nand3_1 _15265_ (.B(_08053_),
    .C(_08515_),
    .A(_08081_),
    .Y(_08563_));
 sg13g2_mux4_1 _15266_ (.S0(net1095),
    .A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S1(net1040),
    .X(_08564_));
 sg13g2_nor2_1 _15267_ (.A(_08055_),
    .B(_08564_),
    .Y(_08565_));
 sg13g2_mux2_1 _15268_ (.A0(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S(_08072_),
    .X(_08566_));
 sg13g2_nor3_1 _15269_ (.A(_08149_),
    .B(_08084_),
    .C(_08566_),
    .Y(_08567_));
 sg13g2_mux2_1 _15270_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(_08072_),
    .X(_08568_));
 sg13g2_nor3_1 _15271_ (.A(_08149_),
    .B(_08058_),
    .C(_08568_),
    .Y(_08569_));
 sg13g2_nor4_1 _15272_ (.A(_08070_),
    .B(_08565_),
    .C(_08567_),
    .D(_08569_),
    .Y(_08570_));
 sg13g2_nand3b_1 _15273_ (.B(_08053_),
    .C(_08515_),
    .Y(_08571_),
    .A_N(_08081_));
 sg13g2_buf_1 _15274_ (.A(_08571_),
    .X(_08572_));
 sg13g2_mux4_1 _15275_ (.S0(net1095),
    .A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S1(_08072_),
    .X(_08573_));
 sg13g2_nor4_1 _15276_ (.A(_08055_),
    .B(net1094),
    .C(_08572_),
    .D(_08573_),
    .Y(_08574_));
 sg13g2_mux4_1 _15277_ (.S0(net1095),
    .A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S1(_08072_),
    .X(_08575_));
 sg13g2_nor4_1 _15278_ (.A(_08149_),
    .B(_08069_),
    .C(_08572_),
    .D(_08575_),
    .Y(_08576_));
 sg13g2_mux4_1 _15279_ (.S0(_08055_),
    .A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S1(_08073_),
    .X(_08577_));
 sg13g2_nor3_1 _15280_ (.A(_08058_),
    .B(_08572_),
    .C(_08577_),
    .Y(_08578_));
 sg13g2_mux4_1 _15281_ (.S0(_08055_),
    .A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S1(net1040),
    .X(_08579_));
 sg13g2_nor3_1 _15282_ (.A(_08084_),
    .B(_08572_),
    .C(_08579_),
    .Y(_08580_));
 sg13g2_nor4_1 _15283_ (.A(_08574_),
    .B(_08576_),
    .C(_08578_),
    .D(_08580_),
    .Y(_08581_));
 sg13g2_o21ai_1 _15284_ (.B1(_08581_),
    .Y(_08582_),
    .A1(_08563_),
    .A2(_08570_));
 sg13g2_mux4_1 _15285_ (.S0(net1095),
    .A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S1(_08072_),
    .X(_08583_));
 sg13g2_mux4_1 _15286_ (.S0(net1095),
    .A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S1(_08072_),
    .X(_08584_));
 sg13g2_mux2_1 _15287_ (.A0(_08583_),
    .A1(_08584_),
    .S(_08149_),
    .X(_08585_));
 sg13g2_o21ai_1 _15288_ (.B1(_08070_),
    .Y(_08586_),
    .A1(_08563_),
    .A2(_08585_));
 sg13g2_or3_1 _15289_ (.A(_08574_),
    .B(_08576_),
    .C(_08586_),
    .X(_08587_));
 sg13g2_buf_2 _15290_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08588_));
 sg13g2_buf_2 _15291_ (.A(_00198_),
    .X(_08589_));
 sg13g2_a21oi_1 _15292_ (.A1(_08588_),
    .A2(\cpu.cond[0] ),
    .Y(_08590_),
    .B1(_08589_));
 sg13g2_or2_1 _15293_ (.X(_08591_),
    .B(_08590_),
    .A(net1091));
 sg13g2_buf_1 _15294_ (.A(\cpu.cond[0] ),
    .X(_08592_));
 sg13g2_nor2b_1 _15295_ (.A(_08588_),
    .B_N(net1090),
    .Y(_08593_));
 sg13g2_nand2_1 _15296_ (.Y(_08594_),
    .A(net1096),
    .B(_00197_));
 sg13g2_a21oi_1 _15297_ (.A1(_08589_),
    .A2(_08593_),
    .Y(_08595_),
    .B1(_08594_));
 sg13g2_a21oi_2 _15298_ (.B1(_08537_),
    .Y(_08596_),
    .A2(_08595_),
    .A1(_08591_));
 sg13g2_nor2_1 _15299_ (.A(_08519_),
    .B(_08596_),
    .Y(_08597_));
 sg13g2_mux4_1 _15300_ (.S0(net1027),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(_08538_),
    .X(_08598_));
 sg13g2_mux4_1 _15301_ (.S0(net1027),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(_08538_),
    .X(_08599_));
 sg13g2_mux4_1 _15302_ (.S0(_08530_),
    .A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[2] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S1(net1026),
    .X(_08600_));
 sg13g2_mux4_1 _15303_ (.S0(net1027),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(net1026),
    .X(_08601_));
 sg13g2_buf_8 _15304_ (.A(net1028),
    .X(_08602_));
 sg13g2_mux4_1 _15305_ (.S0(net887),
    .A0(_08598_),
    .A1(_08599_),
    .A2(_08600_),
    .A3(_08601_),
    .S1(_08529_),
    .X(_08603_));
 sg13g2_inv_1 _15306_ (.Y(_08604_),
    .A(_08603_));
 sg13g2_or2_1 _15307_ (.X(_08605_),
    .B(_08518_),
    .A(_08514_));
 sg13g2_buf_4 _15308_ (.X(_08606_),
    .A(_08605_));
 sg13g2_mux4_1 _15309_ (.S0(net1027),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net887),
    .X(_08607_));
 sg13g2_mux4_1 _15310_ (.S0(net1027),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(_08602_),
    .X(_08608_));
 sg13g2_mux4_1 _15311_ (.S0(_08531_),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(_08522_),
    .X(_08609_));
 sg13g2_mux4_1 _15312_ (.S0(_08531_),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(_08522_),
    .X(_08610_));
 sg13g2_buf_1 _15313_ (.A(net1026),
    .X(_08611_));
 sg13g2_mux4_1 _15314_ (.S0(_08611_),
    .A0(_08607_),
    .A1(_08608_),
    .A2(_08609_),
    .A3(_08610_),
    .S1(_08529_),
    .X(_08612_));
 sg13g2_nor3_1 _15315_ (.A(_08606_),
    .B(_08596_),
    .C(_08612_),
    .Y(_08613_));
 sg13g2_a221oi_1 _15316_ (.B2(_08604_),
    .C1(_08613_),
    .B1(_08597_),
    .A1(_08582_),
    .Y(_08614_),
    .A2(_08587_));
 sg13g2_buf_2 _15317_ (.A(_08614_),
    .X(_08615_));
 sg13g2_nor2_1 _15318_ (.A(_08562_),
    .B(_08615_),
    .Y(_08616_));
 sg13g2_buf_2 _15319_ (.A(_08616_),
    .X(_08617_));
 sg13g2_nor2_1 _15320_ (.A(_08557_),
    .B(_08617_),
    .Y(_08618_));
 sg13g2_buf_2 _15321_ (.A(_08618_),
    .X(_08619_));
 sg13g2_buf_1 _15322_ (.A(_08619_),
    .X(_08620_));
 sg13g2_nand3b_1 _15323_ (.B(_08513_),
    .C(net253),
    .Y(_08621_),
    .A_N(_08512_));
 sg13g2_buf_1 _15324_ (.A(_08621_),
    .X(_08622_));
 sg13g2_buf_1 _15325_ (.A(_08622_),
    .X(_08623_));
 sg13g2_buf_1 _15326_ (.A(net113),
    .X(_08624_));
 sg13g2_buf_1 _15327_ (.A(\cpu.ex.pc[1] ),
    .X(_08625_));
 sg13g2_buf_1 _15328_ (.A(net1089),
    .X(_08626_));
 sg13g2_buf_1 _15329_ (.A(net1025),
    .X(_08627_));
 sg13g2_nand2_1 _15330_ (.Y(_08628_),
    .A(\cpu.icache.r_data[1][16] ),
    .B(net596));
 sg13g2_a22oi_1 _15331_ (.Y(_08629_),
    .B1(net544),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net546),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_a22oi_1 _15332_ (.Y(_08630_),
    .B1(_08200_),
    .B2(\cpu.icache.r_data[5][16] ),
    .A2(net772),
    .A1(\cpu.icache.r_data[4][16] ));
 sg13g2_a22oi_1 _15333_ (.Y(_08631_),
    .B1(_08210_),
    .B2(\cpu.icache.r_data[7][16] ),
    .A2(_08132_),
    .A1(\cpu.icache.r_data[3][16] ));
 sg13g2_nand4_1 _15334_ (.B(_08629_),
    .C(_08630_),
    .A(_08628_),
    .Y(_08632_),
    .D(_08631_));
 sg13g2_a21o_1 _15335_ (.A2(net541),
    .A1(\cpu.icache.r_data[0][16] ),
    .B1(_08632_),
    .X(_08633_));
 sg13g2_a22oi_1 _15336_ (.Y(_08634_),
    .B1(net697),
    .B2(\cpu.icache.r_data[7][0] ),
    .A2(net698),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_and2_1 _15337_ (.A(\cpu.icache.r_data[4][0] ),
    .B(_08202_),
    .X(_08635_));
 sg13g2_a221oi_1 _15338_ (.B2(\cpu.icache.r_data[6][0] ),
    .C1(_08635_),
    .B1(net597),
    .A1(\cpu.icache.r_data[3][0] ),
    .Y(_08636_),
    .A2(net598));
 sg13g2_a22oi_1 _15339_ (.Y(_08637_),
    .B1(net700),
    .B2(\cpu.icache.r_data[5][0] ),
    .A2(net543),
    .A1(\cpu.icache.r_data[2][0] ));
 sg13g2_nand4_1 _15340_ (.B(_08634_),
    .C(_08636_),
    .A(_08447_),
    .Y(_08638_),
    .D(_08637_));
 sg13g2_o21ai_1 _15341_ (.B1(_08638_),
    .Y(_08639_),
    .A1(\cpu.icache.r_data[0][0] ),
    .A2(net476));
 sg13g2_nor2_1 _15342_ (.A(net1025),
    .B(_08639_),
    .Y(_08640_));
 sg13g2_a21oi_1 _15343_ (.A1(net885),
    .A2(_08633_),
    .Y(_08641_),
    .B1(_08640_));
 sg13g2_buf_2 _15344_ (.A(_08641_),
    .X(_08642_));
 sg13g2_a22oi_1 _15345_ (.Y(_08643_),
    .B1(net702),
    .B2(\cpu.icache.r_data[1][1] ),
    .A2(net546),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_a22oi_1 _15346_ (.Y(_08644_),
    .B1(net772),
    .B2(\cpu.icache.r_data[4][1] ),
    .A2(net598),
    .A1(\cpu.icache.r_data[3][1] ));
 sg13g2_mux2_1 _15347_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(\cpu.icache.r_data[7][1] ),
    .S(net1036),
    .X(_08645_));
 sg13g2_a22oi_1 _15348_ (.Y(_08646_),
    .B1(_08645_),
    .B2(net1037),
    .A2(_08117_),
    .A1(\cpu.icache.r_data[6][1] ));
 sg13g2_or2_1 _15349_ (.X(_08647_),
    .B(_08646_),
    .A(net775));
 sg13g2_nand3_1 _15350_ (.B(_08644_),
    .C(_08647_),
    .A(_08643_),
    .Y(_08648_));
 sg13g2_mux2_1 _15351_ (.A0(\cpu.icache.r_data[0][1] ),
    .A1(_08648_),
    .S(_08103_),
    .X(_08649_));
 sg13g2_buf_1 _15352_ (.A(_08383_),
    .X(_08650_));
 sg13g2_mux2_1 _15353_ (.A0(\cpu.icache.r_data[4][17] ),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(net902),
    .X(_08651_));
 sg13g2_a22oi_1 _15354_ (.Y(_08652_),
    .B1(_08651_),
    .B2(net771),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][17] ));
 sg13g2_or2_1 _15355_ (.X(_08653_),
    .B(_08652_),
    .A(net701));
 sg13g2_buf_1 _15356_ (.A(_08129_),
    .X(_08654_));
 sg13g2_and2_1 _15357_ (.A(net903),
    .B(\cpu.icache.r_data[3][17] ),
    .X(_08655_));
 sg13g2_a21oi_1 _15358_ (.A1(net906),
    .A2(\cpu.icache.r_data[7][17] ),
    .Y(_08656_),
    .B1(_08655_));
 sg13g2_a22oi_1 _15359_ (.Y(_08657_),
    .B1(_08126_),
    .B2(\cpu.icache.r_data[1][17] ),
    .A2(net546),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_o21ai_1 _15360_ (.B1(_08657_),
    .Y(_08658_),
    .A1(net765),
    .A2(_08656_));
 sg13g2_a21oi_1 _15361_ (.A1(\cpu.icache.r_data[0][17] ),
    .A2(_08362_),
    .Y(_08659_),
    .B1(_08658_));
 sg13g2_nand3_1 _15362_ (.B(_08653_),
    .C(_08659_),
    .A(net1025),
    .Y(_08660_));
 sg13g2_o21ai_1 _15363_ (.B1(_08660_),
    .Y(_08661_),
    .A1(net885),
    .A2(_08649_));
 sg13g2_buf_1 _15364_ (.A(_08661_),
    .X(_08662_));
 sg13g2_inv_1 _15365_ (.Y(_08663_),
    .A(_08662_));
 sg13g2_nor2_2 _15366_ (.A(_08642_),
    .B(_08663_),
    .Y(_08664_));
 sg13g2_nor2_1 _15367_ (.A(_00202_),
    .B(_08098_),
    .Y(_08665_));
 sg13g2_mux2_1 _15368_ (.A0(\cpu.icache.r_data[4][30] ),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(net1036),
    .X(_08666_));
 sg13g2_a22oi_1 _15369_ (.Y(_08667_),
    .B1(_08666_),
    .B2(net894),
    .A2(_08235_),
    .A1(\cpu.icache.r_data[7][30] ));
 sg13g2_nor2_1 _15370_ (.A(_08161_),
    .B(_08667_),
    .Y(_08668_));
 sg13g2_a22oi_1 _15371_ (.Y(_08669_),
    .B1(_08131_),
    .B2(\cpu.icache.r_data[3][30] ),
    .A2(_08125_),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_a22oi_1 _15372_ (.Y(_08670_),
    .B1(_08199_),
    .B2(\cpu.icache.r_data[5][30] ),
    .A2(_08119_),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_nand2_1 _15373_ (.Y(_08671_),
    .A(_08669_),
    .B(_08670_));
 sg13g2_nor3_1 _15374_ (.A(_08665_),
    .B(_08668_),
    .C(_08671_),
    .Y(_08672_));
 sg13g2_nand2_1 _15375_ (.Y(_08673_),
    .A(_00201_),
    .B(_08361_));
 sg13g2_mux4_1 _15376_ (.S0(net1037),
    .A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[5][14] ),
    .A2(\cpu.icache.r_data[6][14] ),
    .A3(\cpu.icache.r_data[7][14] ),
    .S1(_08110_),
    .X(_08674_));
 sg13g2_nand2_1 _15377_ (.Y(_08675_),
    .A(_08105_),
    .B(_08674_));
 sg13g2_nand2_1 _15378_ (.Y(_08676_),
    .A(\cpu.icache.r_data[2][14] ),
    .B(_08119_));
 sg13g2_a22oi_1 _15379_ (.Y(_08677_),
    .B1(_08131_),
    .B2(\cpu.icache.r_data[3][14] ),
    .A2(_08125_),
    .A1(\cpu.icache.r_data[1][14] ));
 sg13g2_nand4_1 _15380_ (.B(_08675_),
    .C(_08676_),
    .A(_08098_),
    .Y(_08678_),
    .D(_08677_));
 sg13g2_a21oi_1 _15381_ (.A1(_08673_),
    .A2(_08678_),
    .Y(_08679_),
    .B1(net1089));
 sg13g2_a21oi_1 _15382_ (.A1(net1089),
    .A2(_08672_),
    .Y(_08680_),
    .B1(_08679_));
 sg13g2_buf_2 _15383_ (.A(_08680_),
    .X(_08681_));
 sg13g2_nor2_1 _15384_ (.A(_00204_),
    .B(_08100_),
    .Y(_08682_));
 sg13g2_mux2_1 _15385_ (.A0(\cpu.icache.r_data[4][31] ),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(net776),
    .X(_08683_));
 sg13g2_a22oi_1 _15386_ (.Y(_08684_),
    .B1(_08683_),
    .B2(net771),
    .A2(net696),
    .A1(\cpu.icache.r_data[7][31] ));
 sg13g2_nor2_1 _15387_ (.A(net701),
    .B(_08684_),
    .Y(_08685_));
 sg13g2_a22oi_1 _15388_ (.Y(_08686_),
    .B1(net596),
    .B2(\cpu.icache.r_data[1][31] ),
    .A2(_08230_),
    .A1(\cpu.icache.r_data[2][31] ));
 sg13g2_a22oi_1 _15389_ (.Y(_08687_),
    .B1(net700),
    .B2(\cpu.icache.r_data[5][31] ),
    .A2(net545),
    .A1(\cpu.icache.r_data[3][31] ));
 sg13g2_nand2_1 _15390_ (.Y(_08688_),
    .A(_08686_),
    .B(_08687_));
 sg13g2_nor3_1 _15391_ (.A(_08682_),
    .B(_08685_),
    .C(_08688_),
    .Y(_08689_));
 sg13g2_nand2_1 _15392_ (.Y(_08690_),
    .A(_00203_),
    .B(_08362_));
 sg13g2_a22oi_1 _15393_ (.Y(_08691_),
    .B1(_08204_),
    .B2(\cpu.icache.r_data[4][15] ),
    .A2(_08230_),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_a22oi_1 _15394_ (.Y(_08692_),
    .B1(_08133_),
    .B2(\cpu.icache.r_data[3][15] ),
    .A2(_08208_),
    .A1(\cpu.icache.r_data[1][15] ));
 sg13g2_mux2_1 _15395_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(\cpu.icache.r_data[7][15] ),
    .S(net904),
    .X(_08693_));
 sg13g2_a22oi_1 _15396_ (.Y(_08694_),
    .B1(_08693_),
    .B2(net905),
    .A2(_08117_),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_or2_1 _15397_ (.X(_08695_),
    .B(_08694_),
    .A(net767));
 sg13g2_nand4_1 _15398_ (.B(_08691_),
    .C(_08692_),
    .A(_08100_),
    .Y(_08696_),
    .D(_08695_));
 sg13g2_a21oi_1 _15399_ (.A1(_08690_),
    .A2(_08696_),
    .Y(_08697_),
    .B1(net1025));
 sg13g2_a21oi_1 _15400_ (.A1(_08627_),
    .A2(_08689_),
    .Y(_08698_),
    .B1(_08697_));
 sg13g2_buf_1 _15401_ (.A(_08698_),
    .X(_08699_));
 sg13g2_mux2_1 _15402_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_08088_),
    .X(_08700_));
 sg13g2_a22oi_1 _15403_ (.Y(_08701_),
    .B1(_08700_),
    .B2(net904),
    .A2(_08279_),
    .A1(\cpu.icache.r_data[5][29] ));
 sg13g2_nand2b_1 _15404_ (.Y(_08702_),
    .B(net1037),
    .A_N(_08701_));
 sg13g2_a22oi_1 _15405_ (.Y(_08703_),
    .B1(_08203_),
    .B2(\cpu.icache.r_data[4][29] ),
    .A2(_08154_),
    .A1(\cpu.icache.r_data[6][29] ));
 sg13g2_a22oi_1 _15406_ (.Y(_08704_),
    .B1(net695),
    .B2(\cpu.icache.r_data[1][29] ),
    .A2(_08119_),
    .A1(\cpu.icache.r_data[2][29] ));
 sg13g2_nand3_1 _15407_ (.B(_08703_),
    .C(_08704_),
    .A(_08702_),
    .Y(_08705_));
 sg13g2_a21oi_1 _15408_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net541),
    .Y(_08706_),
    .B1(_08705_));
 sg13g2_nand2b_1 _15409_ (.Y(_08707_),
    .B(_08361_),
    .A_N(\cpu.icache.r_data[0][13] ));
 sg13g2_a22oi_1 _15410_ (.Y(_08708_),
    .B1(_08202_),
    .B2(\cpu.icache.r_data[4][13] ),
    .A2(_08119_),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_a22oi_1 _15411_ (.Y(_08709_),
    .B1(_08131_),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(_08125_),
    .A1(\cpu.icache.r_data[1][13] ));
 sg13g2_mux2_1 _15412_ (.A0(\cpu.icache.r_data[5][13] ),
    .A1(\cpu.icache.r_data[7][13] ),
    .S(net1092),
    .X(_08710_));
 sg13g2_a22oi_1 _15413_ (.Y(_08711_),
    .B1(_08710_),
    .B2(_08108_),
    .A2(_08117_),
    .A1(\cpu.icache.r_data[6][13] ));
 sg13g2_or2_1 _15414_ (.X(_08712_),
    .B(_08711_),
    .A(_08160_));
 sg13g2_nand4_1 _15415_ (.B(_08708_),
    .C(_08709_),
    .A(_08098_),
    .Y(_08713_),
    .D(_08712_));
 sg13g2_a21oi_1 _15416_ (.A1(_08707_),
    .A2(_08713_),
    .Y(_08714_),
    .B1(net1089));
 sg13g2_a21o_1 _15417_ (.A2(_08706_),
    .A1(_08627_),
    .B1(_08714_),
    .X(_08715_));
 sg13g2_buf_1 _15418_ (.A(_08715_),
    .X(_08716_));
 sg13g2_nand2_1 _15419_ (.Y(_08717_),
    .A(net252),
    .B(net339));
 sg13g2_nor2_1 _15420_ (.A(_08681_),
    .B(_08717_),
    .Y(_08718_));
 sg13g2_buf_1 _15421_ (.A(_08718_),
    .X(_08719_));
 sg13g2_nand2_1 _15422_ (.Y(_08720_),
    .A(_08664_),
    .B(net155));
 sg13g2_inv_1 _15423_ (.Y(_08721_),
    .A(net1089));
 sg13g2_buf_1 _15424_ (.A(_08721_),
    .X(_08722_));
 sg13g2_nand2_1 _15425_ (.Y(_08723_),
    .A(_00207_),
    .B(net541));
 sg13g2_mux4_1 _15426_ (.S0(net1037),
    .A0(\cpu.icache.r_data[4][11] ),
    .A1(\cpu.icache.r_data[5][11] ),
    .A2(\cpu.icache.r_data[6][11] ),
    .A3(\cpu.icache.r_data[7][11] ),
    .S1(net904),
    .X(_08724_));
 sg13g2_nand2_1 _15427_ (.Y(_08725_),
    .A(net906),
    .B(_08724_));
 sg13g2_nand2_1 _15428_ (.Y(_08726_),
    .A(\cpu.icache.r_data[2][11] ),
    .B(net543));
 sg13g2_a22oi_1 _15429_ (.Y(_08727_),
    .B1(_08132_),
    .B2(\cpu.icache.r_data[3][11] ),
    .A2(net695),
    .A1(\cpu.icache.r_data[1][11] ));
 sg13g2_nand4_1 _15430_ (.B(_08725_),
    .C(_08726_),
    .A(net547),
    .Y(_08728_),
    .D(_08727_));
 sg13g2_nand3_1 _15431_ (.B(_08723_),
    .C(_08728_),
    .A(_08722_),
    .Y(_08729_));
 sg13g2_nor2_1 _15432_ (.A(_00208_),
    .B(net547),
    .Y(_08730_));
 sg13g2_mux2_1 _15433_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(net1036),
    .X(_08731_));
 sg13g2_a22oi_1 _15434_ (.Y(_08732_),
    .B1(_08731_),
    .B2(net766),
    .A2(_08383_),
    .A1(\cpu.icache.r_data[5][27] ));
 sg13g2_nand2_1 _15435_ (.Y(_08733_),
    .A(net1035),
    .B(\cpu.icache.r_data[3][27] ));
 sg13g2_nand2_1 _15436_ (.Y(_08734_),
    .A(_08105_),
    .B(\cpu.icache.r_data[7][27] ));
 sg13g2_a21oi_1 _15437_ (.A1(_08733_),
    .A2(_08734_),
    .Y(_08735_),
    .B1(_08129_));
 sg13g2_a221oi_1 _15438_ (.B2(\cpu.icache.r_data[1][27] ),
    .C1(_08735_),
    .B1(net695),
    .A1(\cpu.icache.r_data[2][27] ),
    .Y(_08736_),
    .A2(net540));
 sg13g2_o21ai_1 _15439_ (.B1(_08736_),
    .Y(_08737_),
    .A1(_08161_),
    .A2(_08732_));
 sg13g2_o21ai_1 _15440_ (.B1(net1089),
    .Y(_08738_),
    .A1(_08730_),
    .A2(_08737_));
 sg13g2_and2_1 _15441_ (.A(_08729_),
    .B(_08738_),
    .X(_08739_));
 sg13g2_buf_1 _15442_ (.A(_08739_),
    .X(_08740_));
 sg13g2_inv_1 _15443_ (.Y(_08741_),
    .A(_08740_));
 sg13g2_nor2_1 _15444_ (.A(_00206_),
    .B(_08098_),
    .Y(_08742_));
 sg13g2_mux2_1 _15445_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(net904),
    .X(_08743_));
 sg13g2_a22oi_1 _15446_ (.Y(_08744_),
    .B1(_08743_),
    .B2(net766),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][26] ));
 sg13g2_nor2_1 _15447_ (.A(net767),
    .B(_08744_),
    .Y(_08745_));
 sg13g2_and2_1 _15448_ (.A(net1035),
    .B(\cpu.icache.r_data[3][26] ),
    .X(_08746_));
 sg13g2_a21oi_1 _15449_ (.A1(net906),
    .A2(\cpu.icache.r_data[7][26] ),
    .Y(_08747_),
    .B1(_08746_));
 sg13g2_a22oi_1 _15450_ (.Y(_08748_),
    .B1(net698),
    .B2(\cpu.icache.r_data[1][26] ),
    .A2(net540),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_o21ai_1 _15451_ (.B1(_08748_),
    .Y(_08749_),
    .A1(net765),
    .A2(_08747_));
 sg13g2_nor4_1 _15452_ (.A(net884),
    .B(_08742_),
    .C(_08745_),
    .D(_08749_),
    .Y(_08750_));
 sg13g2_nand2_1 _15453_ (.Y(_08751_),
    .A(_00205_),
    .B(net541));
 sg13g2_mux2_1 _15454_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(\cpu.icache.r_data[3][10] ),
    .S(net1035),
    .X(_08752_));
 sg13g2_a22oi_1 _15455_ (.Y(_08753_),
    .B1(_08752_),
    .B2(net696),
    .A2(_08203_),
    .A1(\cpu.icache.r_data[4][10] ));
 sg13g2_a22oi_1 _15456_ (.Y(_08754_),
    .B1(net695),
    .B2(\cpu.icache.r_data[1][10] ),
    .A2(net540),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_a22oi_1 _15457_ (.Y(_08755_),
    .B1(_08199_),
    .B2(\cpu.icache.r_data[5][10] ),
    .A2(net597),
    .A1(\cpu.icache.r_data[6][10] ));
 sg13g2_nand4_1 _15458_ (.B(_08753_),
    .C(_08754_),
    .A(net547),
    .Y(_08756_),
    .D(_08755_));
 sg13g2_a21oi_1 _15459_ (.A1(_08751_),
    .A2(_08756_),
    .Y(_08757_),
    .B1(net1089));
 sg13g2_or2_1 _15460_ (.X(_08758_),
    .B(_08757_),
    .A(_08750_));
 sg13g2_buf_1 _15461_ (.A(_08758_),
    .X(_08759_));
 sg13g2_buf_1 _15462_ (.A(_08759_),
    .X(_08760_));
 sg13g2_nor4_1 _15463_ (.A(net113),
    .B(_08720_),
    .C(_08741_),
    .D(net251),
    .Y(_08761_));
 sg13g2_a21o_1 _15464_ (.A2(net91),
    .A1(_08052_),
    .B1(_08761_),
    .X(_00016_));
 sg13g2_buf_1 _15465_ (.A(\cpu.dec.r_op[4] ),
    .X(_08762_));
 sg13g2_buf_1 _15466_ (.A(net1088),
    .X(_08763_));
 sg13g2_nor2_1 _15467_ (.A(_00214_),
    .B(_08098_),
    .Y(_08764_));
 sg13g2_mux2_1 _15468_ (.A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(net904),
    .X(_08765_));
 sg13g2_a22oi_1 _15469_ (.Y(_08766_),
    .B1(_08765_),
    .B2(net766),
    .A2(_08383_),
    .A1(\cpu.icache.r_data[5][28] ));
 sg13g2_nor2_1 _15470_ (.A(net767),
    .B(_08766_),
    .Y(_08767_));
 sg13g2_and2_1 _15471_ (.A(_08159_),
    .B(\cpu.icache.r_data[3][28] ),
    .X(_08768_));
 sg13g2_a21oi_1 _15472_ (.A1(net906),
    .A2(\cpu.icache.r_data[7][28] ),
    .Y(_08769_),
    .B1(_08768_));
 sg13g2_a22oi_1 _15473_ (.Y(_08770_),
    .B1(net695),
    .B2(\cpu.icache.r_data[1][28] ),
    .A2(net540),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_o21ai_1 _15474_ (.B1(_08770_),
    .Y(_08771_),
    .A1(net765),
    .A2(_08769_));
 sg13g2_nor4_1 _15475_ (.A(net884),
    .B(_08764_),
    .C(_08767_),
    .D(_08771_),
    .Y(_08772_));
 sg13g2_nand2_1 _15476_ (.Y(_08773_),
    .A(_00213_),
    .B(_08361_));
 sg13g2_a22oi_1 _15477_ (.Y(_08774_),
    .B1(_08199_),
    .B2(\cpu.icache.r_data[5][12] ),
    .A2(net540),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15478_ (.Y(_08775_),
    .B1(_08131_),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(net695),
    .A1(\cpu.icache.r_data[1][12] ));
 sg13g2_mux2_1 _15479_ (.A0(\cpu.icache.r_data[4][12] ),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_08089_),
    .X(_08776_));
 sg13g2_a22oi_1 _15480_ (.Y(_08777_),
    .B1(_08776_),
    .B2(net894),
    .A2(_08235_),
    .A1(\cpu.icache.r_data[7][12] ));
 sg13g2_or2_1 _15481_ (.X(_08778_),
    .B(_08777_),
    .A(_08160_));
 sg13g2_nand4_1 _15482_ (.B(_08774_),
    .C(_08775_),
    .A(net547),
    .Y(_08779_),
    .D(_08778_));
 sg13g2_a21oi_1 _15483_ (.A1(_08773_),
    .A2(_08779_),
    .Y(_08780_),
    .B1(_08625_));
 sg13g2_or2_1 _15484_ (.X(_08781_),
    .B(_08780_),
    .A(_08772_));
 sg13g2_buf_1 _15485_ (.A(_08781_),
    .X(_08782_));
 sg13g2_buf_1 _15486_ (.A(_08782_),
    .X(_08783_));
 sg13g2_buf_1 _15487_ (.A(net250),
    .X(_08784_));
 sg13g2_inv_1 _15488_ (.Y(_08785_),
    .A(_00211_));
 sg13g2_mux4_1 _15489_ (.S0(net1037),
    .A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[5][6] ),
    .A2(\cpu.icache.r_data[6][6] ),
    .A3(\cpu.icache.r_data[7][6] ),
    .S1(_08111_),
    .X(_08786_));
 sg13g2_nand2_1 _15490_ (.Y(_08787_),
    .A(net906),
    .B(_08786_));
 sg13g2_nand2_1 _15491_ (.Y(_08788_),
    .A(\cpu.icache.r_data[2][6] ),
    .B(net540));
 sg13g2_a22oi_1 _15492_ (.Y(_08789_),
    .B1(net598),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(net695),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_nand4_1 _15493_ (.B(_08787_),
    .C(_08788_),
    .A(_08102_),
    .Y(_08790_),
    .D(_08789_));
 sg13g2_o21ai_1 _15494_ (.B1(_08790_),
    .Y(_08791_),
    .A1(_08785_),
    .A2(net539));
 sg13g2_nor2_1 _15495_ (.A(_00212_),
    .B(net547),
    .Y(_08792_));
 sg13g2_mux2_1 _15496_ (.A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_08111_),
    .X(_08793_));
 sg13g2_a22oi_1 _15497_ (.Y(_08794_),
    .B1(_08793_),
    .B2(net766),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][22] ));
 sg13g2_nand2_1 _15498_ (.Y(_08795_),
    .A(_08159_),
    .B(\cpu.icache.r_data[3][22] ));
 sg13g2_nand2_1 _15499_ (.Y(_08796_),
    .A(_08105_),
    .B(\cpu.icache.r_data[7][22] ));
 sg13g2_a21oi_1 _15500_ (.A1(_08795_),
    .A2(_08796_),
    .Y(_08797_),
    .B1(_08129_));
 sg13g2_a221oi_1 _15501_ (.B2(\cpu.icache.r_data[1][22] ),
    .C1(_08797_),
    .B1(_08450_),
    .A1(\cpu.icache.r_data[2][22] ),
    .Y(_08798_),
    .A2(_08438_));
 sg13g2_o21ai_1 _15502_ (.B1(_08798_),
    .Y(_08799_),
    .A1(net767),
    .A2(_08794_));
 sg13g2_nor3_1 _15503_ (.A(net884),
    .B(_08792_),
    .C(_08799_),
    .Y(_08800_));
 sg13g2_a21oi_1 _15504_ (.A1(net884),
    .A2(_08791_),
    .Y(_08801_),
    .B1(_08800_));
 sg13g2_buf_2 _15505_ (.A(_08801_),
    .X(_08802_));
 sg13g2_inv_2 _15506_ (.Y(_08803_),
    .A(_08802_));
 sg13g2_nor2_1 _15507_ (.A(_00210_),
    .B(net548),
    .Y(_08804_));
 sg13g2_mux2_1 _15508_ (.A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(net902),
    .X(_08805_));
 sg13g2_a22oi_1 _15509_ (.Y(_08806_),
    .B1(_08805_),
    .B2(net766),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][21] ));
 sg13g2_nor2_1 _15510_ (.A(net767),
    .B(_08806_),
    .Y(_08807_));
 sg13g2_and2_1 _15511_ (.A(net903),
    .B(\cpu.icache.r_data[3][21] ),
    .X(_08808_));
 sg13g2_a21oi_1 _15512_ (.A1(_08106_),
    .A2(\cpu.icache.r_data[7][21] ),
    .Y(_08809_),
    .B1(_08808_));
 sg13g2_a22oi_1 _15513_ (.Y(_08810_),
    .B1(net702),
    .B2(\cpu.icache.r_data[1][21] ),
    .A2(_08229_),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_o21ai_1 _15514_ (.B1(_08810_),
    .Y(_08811_),
    .A1(net765),
    .A2(_08809_));
 sg13g2_nor3_1 _15515_ (.A(_08804_),
    .B(_08807_),
    .C(_08811_),
    .Y(_08812_));
 sg13g2_inv_1 _15516_ (.Y(_08813_),
    .A(_00209_));
 sg13g2_a22oi_1 _15517_ (.Y(_08814_),
    .B1(_08199_),
    .B2(\cpu.icache.r_data[5][5] ),
    .A2(_08438_),
    .A1(\cpu.icache.r_data[2][5] ));
 sg13g2_a22oi_1 _15518_ (.Y(_08815_),
    .B1(net598),
    .B2(\cpu.icache.r_data[3][5] ),
    .A2(net695),
    .A1(\cpu.icache.r_data[1][5] ));
 sg13g2_mux2_1 _15519_ (.A0(\cpu.icache.r_data[4][5] ),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(net1036),
    .X(_08816_));
 sg13g2_a22oi_1 _15520_ (.Y(_08817_),
    .B1(_08816_),
    .B2(_08257_),
    .A2(_08235_),
    .A1(\cpu.icache.r_data[7][5] ));
 sg13g2_or2_1 _15521_ (.X(_08818_),
    .B(_08817_),
    .A(net903));
 sg13g2_nand4_1 _15522_ (.B(_08814_),
    .C(_08815_),
    .A(_08102_),
    .Y(_08819_),
    .D(_08818_));
 sg13g2_o21ai_1 _15523_ (.B1(_08819_),
    .Y(_08820_),
    .A1(_08813_),
    .A2(net539));
 sg13g2_buf_1 _15524_ (.A(net884),
    .X(_08821_));
 sg13g2_mux2_1 _15525_ (.A0(_08812_),
    .A1(_08820_),
    .S(net764),
    .X(_08822_));
 sg13g2_buf_1 _15526_ (.A(_08822_),
    .X(_08823_));
 sg13g2_nand2_1 _15527_ (.Y(_08824_),
    .A(_08803_),
    .B(_08823_));
 sg13g2_buf_1 _15528_ (.A(_08824_),
    .X(_08825_));
 sg13g2_nor2_2 _15529_ (.A(_08740_),
    .B(_08759_),
    .Y(_08826_));
 sg13g2_a21oi_1 _15530_ (.A1(net1025),
    .A2(_08706_),
    .Y(_08827_),
    .B1(_08714_));
 sg13g2_buf_1 _15531_ (.A(_08827_),
    .X(_08828_));
 sg13g2_nor2_1 _15532_ (.A(_08681_),
    .B(_08828_),
    .Y(_08829_));
 sg13g2_buf_1 _15533_ (.A(_08829_),
    .X(_08830_));
 sg13g2_nand2_1 _15534_ (.Y(_08831_),
    .A(net252),
    .B(_08830_));
 sg13g2_buf_2 _15535_ (.A(_08831_),
    .X(_08832_));
 sg13g2_inv_1 _15536_ (.Y(_08833_),
    .A(_08642_));
 sg13g2_nand2_1 _15537_ (.Y(_08834_),
    .A(_08833_),
    .B(_08663_));
 sg13g2_buf_1 _15538_ (.A(_08834_),
    .X(_08835_));
 sg13g2_nor2_1 _15539_ (.A(_08832_),
    .B(_08835_),
    .Y(_08836_));
 sg13g2_nand2_1 _15540_ (.Y(_08837_),
    .A(_08826_),
    .B(_08836_));
 sg13g2_nor4_1 _15541_ (.A(net113),
    .B(_08784_),
    .C(_08825_),
    .D(_08837_),
    .Y(_08838_));
 sg13g2_a21o_1 _15542_ (.A2(net91),
    .A1(net1024),
    .B1(_08838_),
    .X(_00015_));
 sg13g2_buf_1 _15543_ (.A(\cpu.dec.r_op[3] ),
    .X(_08839_));
 sg13g2_inv_1 _15544_ (.Y(_08840_),
    .A(net1087));
 sg13g2_buf_1 _15545_ (.A(_08840_),
    .X(_08841_));
 sg13g2_nand4_1 _15546_ (.B(_08481_),
    .C(_08489_),
    .A(_08444_),
    .Y(_08842_),
    .D(_08498_));
 sg13g2_nand4_1 _15547_ (.B(_08508_),
    .C(_08459_),
    .A(_08456_),
    .Y(_08843_),
    .D(_08471_));
 sg13g2_nor3_1 _15548_ (.A(_08411_),
    .B(_08842_),
    .C(_08843_),
    .Y(_08844_));
 sg13g2_nand3b_1 _15549_ (.B(_08314_),
    .C(_08844_),
    .Y(_08845_),
    .A_N(_08390_));
 sg13g2_nand3_1 _15550_ (.B(_08215_),
    .C(_08240_),
    .A(_08367_),
    .Y(_08846_));
 sg13g2_inv_1 _15551_ (.Y(_08847_),
    .A(_08433_));
 sg13g2_nand3_1 _15552_ (.B(_08286_),
    .C(_08847_),
    .A(_08263_),
    .Y(_08848_));
 sg13g2_nor4_1 _15553_ (.A(_08171_),
    .B(_08845_),
    .C(_08846_),
    .D(_08848_),
    .Y(_08849_));
 sg13g2_and3_1 _15554_ (.X(_08850_),
    .A(_08513_),
    .B(net253),
    .C(_08849_));
 sg13g2_buf_1 _15555_ (.A(_08850_),
    .X(_08851_));
 sg13g2_buf_1 _15556_ (.A(net132),
    .X(_08852_));
 sg13g2_buf_1 _15557_ (.A(net132),
    .X(_08853_));
 sg13g2_nand2b_1 _15558_ (.Y(_08854_),
    .B(net884),
    .A_N(_08820_));
 sg13g2_o21ai_1 _15559_ (.B1(_08854_),
    .Y(_08855_),
    .A1(net764),
    .A2(_08812_));
 sg13g2_buf_1 _15560_ (.A(_08855_),
    .X(_08856_));
 sg13g2_nand3_1 _15561_ (.B(_08803_),
    .C(net248),
    .A(net250),
    .Y(_08857_));
 sg13g2_buf_1 _15562_ (.A(_08857_),
    .X(_08858_));
 sg13g2_nand3_1 _15563_ (.B(net155),
    .C(_08826_),
    .A(_08664_),
    .Y(_08859_));
 sg13g2_buf_1 _15564_ (.A(_08859_),
    .X(_08860_));
 sg13g2_nor2_2 _15565_ (.A(_08782_),
    .B(_08802_),
    .Y(_08861_));
 sg13g2_nor2_1 _15566_ (.A(_08823_),
    .B(_08837_),
    .Y(_08862_));
 sg13g2_inv_1 _15567_ (.Y(_08863_),
    .A(_00219_));
 sg13g2_mux4_1 _15568_ (.S0(_08109_),
    .A0(\cpu.icache.r_data[4][4] ),
    .A1(\cpu.icache.r_data[5][4] ),
    .A2(\cpu.icache.r_data[6][4] ),
    .A3(\cpu.icache.r_data[7][4] ),
    .S1(net776),
    .X(_08864_));
 sg13g2_nand2_1 _15569_ (.Y(_08865_),
    .A(net777),
    .B(_08864_));
 sg13g2_nand2_1 _15570_ (.Y(_08866_),
    .A(\cpu.icache.r_data[2][4] ),
    .B(net475));
 sg13g2_a22oi_1 _15571_ (.Y(_08867_),
    .B1(net545),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(net599),
    .A1(\cpu.icache.r_data[1][4] ));
 sg13g2_nand4_1 _15572_ (.B(_08865_),
    .C(_08866_),
    .A(net410),
    .Y(_08868_),
    .D(_08867_));
 sg13g2_o21ai_1 _15573_ (.B1(_08868_),
    .Y(_08869_),
    .A1(_08863_),
    .A2(_08101_));
 sg13g2_nor2_1 _15574_ (.A(_00220_),
    .B(_08104_),
    .Y(_08870_));
 sg13g2_mux2_1 _15575_ (.A0(\cpu.icache.r_data[4][20] ),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(net776),
    .X(_08871_));
 sg13g2_a22oi_1 _15576_ (.Y(_08872_),
    .B1(_08871_),
    .B2(net771),
    .A2(_08650_),
    .A1(\cpu.icache.r_data[5][20] ));
 sg13g2_nand2_1 _15577_ (.Y(_08873_),
    .A(_08306_),
    .B(\cpu.icache.r_data[3][20] ));
 sg13g2_nand2_1 _15578_ (.Y(_08874_),
    .A(net777),
    .B(\cpu.icache.r_data[7][20] ));
 sg13g2_a21oi_1 _15579_ (.A1(_08873_),
    .A2(_08874_),
    .Y(_08875_),
    .B1(_08654_));
 sg13g2_a221oi_1 _15580_ (.B2(\cpu.icache.r_data[1][20] ),
    .C1(_08875_),
    .B1(net599),
    .A1(\cpu.icache.r_data[2][20] ),
    .Y(_08876_),
    .A2(net472));
 sg13g2_o21ai_1 _15581_ (.B1(_08876_),
    .Y(_08877_),
    .A1(net701),
    .A2(_08872_));
 sg13g2_nor3_1 _15582_ (.A(net764),
    .B(_08870_),
    .C(_08877_),
    .Y(_08878_));
 sg13g2_a21oi_1 _15583_ (.A1(net764),
    .A2(_08869_),
    .Y(_08879_),
    .B1(_08878_));
 sg13g2_buf_1 _15584_ (.A(_08879_),
    .X(_08880_));
 sg13g2_inv_1 _15585_ (.Y(_08881_),
    .A(_08880_));
 sg13g2_nor2_1 _15586_ (.A(_00216_),
    .B(net548),
    .Y(_08882_));
 sg13g2_mux2_1 _15587_ (.A0(\cpu.icache.r_data[4][18] ),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(net902),
    .X(_08883_));
 sg13g2_a22oi_1 _15588_ (.Y(_08884_),
    .B1(_08883_),
    .B2(_08385_),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][18] ));
 sg13g2_nor2_1 _15589_ (.A(net767),
    .B(_08884_),
    .Y(_08885_));
 sg13g2_and2_1 _15590_ (.A(net903),
    .B(\cpu.icache.r_data[3][18] ),
    .X(_08886_));
 sg13g2_a21oi_1 _15591_ (.A1(_08106_),
    .A2(\cpu.icache.r_data[7][18] ),
    .Y(_08887_),
    .B1(_08886_));
 sg13g2_a22oi_1 _15592_ (.Y(_08888_),
    .B1(_08126_),
    .B2(\cpu.icache.r_data[1][18] ),
    .A2(_08120_),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_o21ai_1 _15593_ (.B1(_08888_),
    .Y(_08889_),
    .A1(net765),
    .A2(_08887_));
 sg13g2_nor4_1 _15594_ (.A(net884),
    .B(_08882_),
    .C(_08885_),
    .D(_08889_),
    .Y(_08890_));
 sg13g2_nand2_1 _15595_ (.Y(_08891_),
    .A(_00215_),
    .B(net541));
 sg13g2_a22oi_1 _15596_ (.Y(_08892_),
    .B1(net700),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(net546),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_a22oi_1 _15597_ (.Y(_08893_),
    .B1(net598),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(_08207_),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_mux2_1 _15598_ (.A0(\cpu.icache.r_data[4][2] ),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(net1036),
    .X(_08894_));
 sg13g2_a22oi_1 _15599_ (.Y(_08895_),
    .B1(_08894_),
    .B2(net894),
    .A2(_08235_),
    .A1(\cpu.icache.r_data[7][2] ));
 sg13g2_or2_1 _15600_ (.X(_08896_),
    .B(_08895_),
    .A(net775));
 sg13g2_nand4_1 _15601_ (.B(_08892_),
    .C(_08893_),
    .A(_08447_),
    .Y(_08897_),
    .D(_08896_));
 sg13g2_a21oi_1 _15602_ (.A1(_08891_),
    .A2(_08897_),
    .Y(_08898_),
    .B1(_08626_));
 sg13g2_or2_1 _15603_ (.X(_08899_),
    .B(_08898_),
    .A(_08890_));
 sg13g2_buf_2 _15604_ (.A(_08899_),
    .X(_08900_));
 sg13g2_mux4_1 _15605_ (.S0(net1037),
    .A0(\cpu.icache.r_data[4][3] ),
    .A1(\cpu.icache.r_data[5][3] ),
    .A2(\cpu.icache.r_data[6][3] ),
    .A3(\cpu.icache.r_data[7][3] ),
    .S1(_08163_),
    .X(_08901_));
 sg13g2_nand2_1 _15606_ (.Y(_08902_),
    .A(net906),
    .B(_08901_));
 sg13g2_nand2_1 _15607_ (.Y(_08903_),
    .A(\cpu.icache.r_data[2][3] ),
    .B(_08229_));
 sg13g2_a22oi_1 _15608_ (.Y(_08904_),
    .B1(net598),
    .B2(\cpu.icache.r_data[3][3] ),
    .A2(_08207_),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_and4_1 _15609_ (.A(_08099_),
    .B(_08902_),
    .C(_08903_),
    .D(_08904_),
    .X(_08905_));
 sg13g2_a21oi_1 _15610_ (.A1(_00217_),
    .A2(net541),
    .Y(_08906_),
    .B1(_08905_));
 sg13g2_nor2_1 _15611_ (.A(_00218_),
    .B(net548),
    .Y(_08907_));
 sg13g2_mux2_1 _15612_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(net903),
    .X(_08908_));
 sg13g2_a22oi_1 _15613_ (.Y(_08909_),
    .B1(_08908_),
    .B2(net776),
    .A2(_08279_),
    .A1(\cpu.icache.r_data[5][19] ));
 sg13g2_nor2_1 _15614_ (.A(net771),
    .B(_08909_),
    .Y(_08910_));
 sg13g2_a22oi_1 _15615_ (.Y(_08911_),
    .B1(net544),
    .B2(\cpu.icache.r_data[6][19] ),
    .A2(net702),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_a22oi_1 _15616_ (.Y(_08912_),
    .B1(net772),
    .B2(\cpu.icache.r_data[4][19] ),
    .A2(_08120_),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_nand2_1 _15617_ (.Y(_08913_),
    .A(_08911_),
    .B(_08912_));
 sg13g2_or4_1 _15618_ (.A(_08722_),
    .B(_08907_),
    .C(_08910_),
    .D(_08913_),
    .X(_08914_));
 sg13g2_o21ai_1 _15619_ (.B1(_08914_),
    .Y(_08915_),
    .A1(_08626_),
    .A2(_08906_));
 sg13g2_buf_1 _15620_ (.A(_08915_),
    .X(_08916_));
 sg13g2_nor2_1 _15621_ (.A(_08900_),
    .B(_08916_),
    .Y(_08917_));
 sg13g2_nand4_1 _15622_ (.B(_08862_),
    .C(_08881_),
    .A(_08861_),
    .Y(_08918_),
    .D(_08917_));
 sg13g2_o21ai_1 _15623_ (.B1(_08918_),
    .Y(_08919_),
    .A1(_08858_),
    .A2(_08860_));
 sg13g2_nand2_1 _15624_ (.Y(_08920_),
    .A(net111),
    .B(_08919_));
 sg13g2_o21ai_1 _15625_ (.B1(_08920_),
    .Y(_00014_),
    .A1(_08841_),
    .A2(net112));
 sg13g2_buf_1 _15626_ (.A(\cpu.dec.r_op[6] ),
    .X(_08921_));
 sg13g2_inv_2 _15627_ (.Y(_08922_),
    .A(net1086));
 sg13g2_nand2_1 _15628_ (.Y(_08923_),
    .A(_08900_),
    .B(_08916_));
 sg13g2_buf_2 _15629_ (.A(_08923_),
    .X(_08924_));
 sg13g2_and3_1 _15630_ (.X(_08925_),
    .A(_08861_),
    .B(_08862_),
    .C(net247));
 sg13g2_nor2b_1 _15631_ (.A(_08924_),
    .B_N(_08925_),
    .Y(_08926_));
 sg13g2_nor2_1 _15632_ (.A(_08825_),
    .B(_08860_),
    .Y(_08927_));
 sg13g2_o21ai_1 _15633_ (.B1(_08851_),
    .Y(_08928_),
    .A1(_08926_),
    .A2(_08927_));
 sg13g2_o21ai_1 _15634_ (.B1(_08928_),
    .Y(_00017_),
    .A1(_08922_),
    .A2(net112));
 sg13g2_buf_1 _15635_ (.A(\cpu.spi.r_count[7] ),
    .X(_08929_));
 sg13g2_buf_1 _15636_ (.A(\cpu.spi.r_count[3] ),
    .X(_08930_));
 sg13g2_buf_1 _15637_ (.A(\cpu.spi.r_count[0] ),
    .X(_08931_));
 sg13g2_buf_1 _15638_ (.A(\cpu.spi.r_count[1] ),
    .X(_08932_));
 sg13g2_nor2_1 _15639_ (.A(_08931_),
    .B(_08932_),
    .Y(_08933_));
 sg13g2_nand2b_1 _15640_ (.Y(_08934_),
    .B(_08933_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_buf_1 _15641_ (.A(_08934_),
    .X(_08935_));
 sg13g2_nor3_1 _15642_ (.A(_08930_),
    .B(\cpu.spi.r_count[4] ),
    .C(_08935_),
    .Y(_08936_));
 sg13g2_nor2b_1 _15643_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_08936_),
    .Y(_08937_));
 sg13g2_nor2b_1 _15644_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_08937_),
    .Y(_08938_));
 sg13g2_nand2b_1 _15645_ (.Y(_08939_),
    .B(_08938_),
    .A_N(_08929_));
 sg13g2_buf_1 _15646_ (.A(_08939_),
    .X(_08940_));
 sg13g2_buf_1 _15647_ (.A(\cpu.addr[3] ),
    .X(_08941_));
 sg13g2_buf_1 _15648_ (.A(_08941_),
    .X(_08942_));
 sg13g2_buf_1 _15649_ (.A(net1023),
    .X(_08943_));
 sg13g2_buf_1 _15650_ (.A(net882),
    .X(_08944_));
 sg13g2_buf_1 _15651_ (.A(net763),
    .X(_08945_));
 sg13g2_buf_1 _15652_ (.A(net693),
    .X(_08946_));
 sg13g2_buf_1 _15653_ (.A(net594),
    .X(_08947_));
 sg13g2_buf_1 _15654_ (.A(\cpu.addr[6] ),
    .X(_08948_));
 sg13g2_buf_1 _15655_ (.A(_08948_),
    .X(_08949_));
 sg13g2_inv_1 _15656_ (.Y(_08950_),
    .A(net1022));
 sg13g2_buf_1 _15657_ (.A(\cpu.addr[8] ),
    .X(_08951_));
 sg13g2_buf_2 _15658_ (.A(\cpu.addr[7] ),
    .X(_08952_));
 sg13g2_nand2b_1 _15659_ (.Y(_08953_),
    .B(_08952_),
    .A_N(net1085));
 sg13g2_buf_1 _15660_ (.A(_08953_),
    .X(_08954_));
 sg13g2_or2_1 _15661_ (.X(_08955_),
    .B(_08954_),
    .A(_08950_));
 sg13g2_buf_2 _15662_ (.A(_08955_),
    .X(_08956_));
 sg13g2_buf_1 _15663_ (.A(\cpu.addr[2] ),
    .X(_08957_));
 sg13g2_buf_1 _15664_ (.A(_08957_),
    .X(_08958_));
 sg13g2_buf_2 _15665_ (.A(net1021),
    .X(_08959_));
 sg13g2_buf_2 _15666_ (.A(net881),
    .X(_08960_));
 sg13g2_buf_1 _15667_ (.A(net762),
    .X(_08961_));
 sg13g2_buf_1 _15668_ (.A(\cpu.addr[1] ),
    .X(_08962_));
 sg13g2_buf_1 _15669_ (.A(_08962_),
    .X(_08963_));
 sg13g2_buf_1 _15670_ (.A(net1020),
    .X(_08964_));
 sg13g2_nor2_1 _15671_ (.A(net692),
    .B(net880),
    .Y(_08965_));
 sg13g2_buf_2 _15672_ (.A(_08965_),
    .X(_08966_));
 sg13g2_buf_2 _15673_ (.A(\cpu.dec.r_trap ),
    .X(_08967_));
 sg13g2_buf_1 _15674_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_08968_));
 sg13g2_buf_2 _15675_ (.A(ui_in[6]),
    .X(_08969_));
 sg13g2_buf_1 _15676_ (.A(\cpu.gpio.r_enable_io[7] ),
    .X(_08970_));
 sg13g2_buf_2 _15677_ (.A(uio_in[7]),
    .X(_08971_));
 sg13g2_a22oi_1 _15678_ (.Y(_08972_),
    .B1(_08970_),
    .B2(_08971_),
    .A2(_08969_),
    .A1(_08968_));
 sg13g2_buf_2 _15679_ (.A(ui_in[1]),
    .X(_08973_));
 sg13g2_buf_2 _15680_ (.A(ui_in[4]),
    .X(_08974_));
 sg13g2_a22oi_1 _15681_ (.Y(_08975_),
    .B1(\cpu.gpio.r_enable_in[4] ),
    .B2(_08974_),
    .A2(_08973_),
    .A1(\cpu.gpio.r_enable_in[1] ));
 sg13g2_buf_2 _15682_ (.A(ui_in[7]),
    .X(_08976_));
 sg13g2_buf_2 _15683_ (.A(\cpu.gpio.r_enable_io[4] ),
    .X(_08977_));
 sg13g2_buf_2 _15684_ (.A(uio_in[4]),
    .X(_08978_));
 sg13g2_a22oi_1 _15685_ (.Y(_08979_),
    .B1(_08977_),
    .B2(_08978_),
    .A2(_08976_),
    .A1(\cpu.gpio.r_enable_in[7] ));
 sg13g2_buf_2 _15686_ (.A(ui_in[0]),
    .X(_08980_));
 sg13g2_buf_2 _15687_ (.A(ui_in[5]),
    .X(_08981_));
 sg13g2_a22oi_1 _15688_ (.Y(_08982_),
    .B1(\cpu.gpio.r_enable_in[5] ),
    .B2(_08981_),
    .A2(_08980_),
    .A1(\cpu.gpio.r_enable_in[0] ));
 sg13g2_nand4_1 _15689_ (.B(_08975_),
    .C(_08979_),
    .A(_08972_),
    .Y(_08983_),
    .D(_08982_));
 sg13g2_buf_2 _15690_ (.A(ui_in[2]),
    .X(_08984_));
 sg13g2_buf_1 _15691_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_08985_));
 sg13g2_buf_1 _15692_ (.A(uio_in[5]),
    .X(_08986_));
 sg13g2_a22oi_1 _15693_ (.Y(_08987_),
    .B1(_08985_),
    .B2(_08986_),
    .A2(_08984_),
    .A1(\cpu.gpio.r_enable_in[2] ));
 sg13g2_buf_2 _15694_ (.A(ui_in[3]),
    .X(_08988_));
 sg13g2_buf_1 _15695_ (.A(uio_in[6]),
    .X(_08989_));
 sg13g2_a22oi_1 _15696_ (.Y(_08990_),
    .B1(\cpu.gpio.r_enable_io[6] ),
    .B2(_08989_),
    .A2(_08988_),
    .A1(\cpu.gpio.r_enable_in[3] ));
 sg13g2_nand2_1 _15697_ (.Y(_08991_),
    .A(_08987_),
    .B(_08990_));
 sg13g2_buf_2 _15698_ (.A(\cpu.intr.r_enable[4] ),
    .X(_08992_));
 sg13g2_o21ai_1 _15699_ (.B1(_08992_),
    .Y(_08993_),
    .A1(_08983_),
    .A2(_08991_));
 sg13g2_buf_1 _15700_ (.A(\cpu.intr.r_timer ),
    .X(_08994_));
 sg13g2_buf_1 _15701_ (.A(\cpu.intr.r_swi ),
    .X(_08995_));
 sg13g2_a22oi_1 _15702_ (.Y(_08996_),
    .B1(\cpu.intr.r_enable[3] ),
    .B2(_08995_),
    .A2(\cpu.intr.r_enable[2] ),
    .A1(_08994_));
 sg13g2_buf_1 _15703_ (.A(\cpu.intr.r_enable[1] ),
    .X(_08997_));
 sg13g2_buf_1 _15704_ (.A(\cpu.intr.spi_intr ),
    .X(_08998_));
 sg13g2_buf_1 _15705_ (.A(\cpu.intr.r_enable[5] ),
    .X(_08999_));
 sg13g2_a22oi_1 _15706_ (.Y(_09000_),
    .B1(_08998_),
    .B2(_08999_),
    .A2(_08997_),
    .A1(\cpu.intr.r_clock ));
 sg13g2_buf_1 _15707_ (.A(\cpu.uart.r_x_int ),
    .X(_09001_));
 sg13g2_buf_1 _15708_ (.A(\cpu.uart.r_r_int ),
    .X(_09002_));
 sg13g2_buf_1 _15709_ (.A(\cpu.intr.r_enable[0] ),
    .X(_09003_));
 sg13g2_o21ai_1 _15710_ (.B1(_09003_),
    .Y(_09004_),
    .A1(_09001_),
    .A2(_09002_));
 sg13g2_and3_1 _15711_ (.X(_09005_),
    .A(_08996_),
    .B(_09000_),
    .C(_09004_));
 sg13g2_buf_1 _15712_ (.A(_09005_),
    .X(_09006_));
 sg13g2_buf_1 _15713_ (.A(\cpu.ex.r_ie ),
    .X(_09007_));
 sg13g2_inv_1 _15714_ (.Y(_09008_),
    .A(_09007_));
 sg13g2_a21oi_1 _15715_ (.A1(_08993_),
    .A2(_09006_),
    .Y(_09009_),
    .B1(_09008_));
 sg13g2_and2_1 _15716_ (.A(_08081_),
    .B(_09009_),
    .X(_09010_));
 sg13g2_nor4_2 _15717_ (.A(_08967_),
    .B(_08557_),
    .C(_08617_),
    .Y(_09011_),
    .D(_09010_));
 sg13g2_nand3b_1 _15718_ (.B(_08966_),
    .C(_09011_),
    .Y(_09012_),
    .A_N(_00197_));
 sg13g2_inv_1 _15719_ (.Y(_09013_),
    .A(_08589_));
 sg13g2_nor2_1 _15720_ (.A(_08588_),
    .B(_08589_),
    .Y(_09014_));
 sg13g2_a21oi_1 _15721_ (.A1(_08588_),
    .A2(net1091),
    .Y(_09015_),
    .B1(_09014_));
 sg13g2_nand2_1 _15722_ (.Y(_09016_),
    .A(net1090),
    .B(_09015_));
 sg13g2_o21ai_1 _15723_ (.B1(_09016_),
    .Y(_09017_),
    .A1(_09013_),
    .A2(net1091));
 sg13g2_nor4_2 _15724_ (.A(net538),
    .B(_08956_),
    .C(_09012_),
    .Y(_09018_),
    .D(_09017_));
 sg13g2_buf_1 _15725_ (.A(\cpu.spi.r_state[1] ),
    .X(_09019_));
 sg13g2_inv_1 _15726_ (.Y(_09020_),
    .A(net1084));
 sg13g2_nand3_1 _15727_ (.B(_08561_),
    .C(_09011_),
    .A(_08534_),
    .Y(_09021_));
 sg13g2_buf_2 _15728_ (.A(_09021_),
    .X(_09022_));
 sg13g2_or2_1 _15729_ (.X(_09023_),
    .B(_09022_),
    .A(_08956_));
 sg13g2_buf_1 _15730_ (.A(_09023_),
    .X(_09024_));
 sg13g2_nor2_1 _15731_ (.A(net538),
    .B(_09024_),
    .Y(_09025_));
 sg13g2_buf_1 _15732_ (.A(_09025_),
    .X(_09026_));
 sg13g2_nor2_1 _15733_ (.A(_09020_),
    .B(net131),
    .Y(_09027_));
 sg13g2_a21oi_1 _15734_ (.A1(_09018_),
    .A2(_09027_),
    .Y(_09028_),
    .B1(\cpu.spi.r_state[3] ));
 sg13g2_nand2b_1 _15735_ (.Y(_09029_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_1 _15736_ (.A(_09029_),
    .X(_09030_));
 sg13g2_buf_1 _15737_ (.A(\cpu.spi.r_state[0] ),
    .X(_09031_));
 sg13g2_inv_1 _15738_ (.Y(_09032_),
    .A(_09031_));
 sg13g2_a21oi_1 _15739_ (.A1(_08966_),
    .A2(net131),
    .Y(_09033_),
    .B1(_09032_));
 sg13g2_nor2_1 _15740_ (.A(net1019),
    .B(_09033_),
    .Y(_09034_));
 sg13g2_o21ai_1 _15741_ (.B1(_09034_),
    .Y(_00029_),
    .A1(net406),
    .A2(_09028_));
 sg13g2_nor2b_1 _15742_ (.A(r_reset),
    .B_N(net1),
    .Y(_09035_));
 sg13g2_buf_1 _15743_ (.A(_09035_),
    .X(_09036_));
 sg13g2_buf_2 _15744_ (.A(net1018),
    .X(_09037_));
 sg13g2_buf_1 _15745_ (.A(net879),
    .X(_09038_));
 sg13g2_buf_2 _15746_ (.A(_09038_),
    .X(_09039_));
 sg13g2_inv_2 _15747_ (.Y(_09040_),
    .A(net1023));
 sg13g2_buf_1 _15748_ (.A(_09040_),
    .X(_09041_));
 sg13g2_nand2b_1 _15749_ (.Y(_09042_),
    .B(net760),
    .A_N(_09024_));
 sg13g2_buf_1 _15750_ (.A(_09042_),
    .X(_09043_));
 sg13g2_nand2_1 _15751_ (.Y(_09044_),
    .A(net1084),
    .B(net130));
 sg13g2_buf_1 _15752_ (.A(\cpu.spi.r_state[6] ),
    .X(_09045_));
 sg13g2_buf_1 _15753_ (.A(_09045_),
    .X(_09046_));
 sg13g2_nor2b_1 _15754_ (.A(_08929_),
    .B_N(_08938_),
    .Y(_09047_));
 sg13g2_buf_1 _15755_ (.A(_09047_),
    .X(_09048_));
 sg13g2_buf_1 _15756_ (.A(net405),
    .X(_09049_));
 sg13g2_buf_1 _15757_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09050_));
 sg13g2_buf_1 _15758_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09051_));
 sg13g2_nor3_1 _15759_ (.A(_09050_),
    .B(_09051_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09052_));
 sg13g2_buf_1 _15760_ (.A(\cpu.spi.r_timeout_count[7] ),
    .X(_09053_));
 sg13g2_buf_1 _15761_ (.A(\cpu.spi.r_timeout_count[0] ),
    .X(_09054_));
 sg13g2_buf_1 _15762_ (.A(\cpu.spi.r_timeout_count[1] ),
    .X(_09055_));
 sg13g2_or3_1 _15763_ (.A(_09054_),
    .B(_09055_),
    .C(\cpu.spi.r_timeout_count[2] ),
    .X(_09056_));
 sg13g2_buf_1 _15764_ (.A(_09056_),
    .X(_09057_));
 sg13g2_or2_1 _15765_ (.X(_09058_),
    .B(_09057_),
    .A(\cpu.spi.r_timeout_count[3] ));
 sg13g2_buf_1 _15766_ (.A(_09058_),
    .X(_09059_));
 sg13g2_or2_1 _15767_ (.X(_09060_),
    .B(_09059_),
    .A(\cpu.spi.r_timeout_count[4] ));
 sg13g2_buf_1 _15768_ (.A(_09060_),
    .X(_09061_));
 sg13g2_or2_1 _15769_ (.X(_09062_),
    .B(_09061_),
    .A(\cpu.spi.r_timeout_count[5] ));
 sg13g2_buf_1 _15770_ (.A(_09062_),
    .X(_09063_));
 sg13g2_or2_1 _15771_ (.X(_09064_),
    .B(_09063_),
    .A(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _15772_ (.A(_09064_),
    .X(_09065_));
 sg13g2_buf_1 _15773_ (.A(\cpu.spi.r_searching ),
    .X(_09066_));
 sg13g2_o21ai_1 _15774_ (.B1(_09066_),
    .Y(_09067_),
    .A1(_09053_),
    .A2(_09065_));
 sg13g2_nand2_1 _15775_ (.Y(_09068_),
    .A(_09052_),
    .B(_09067_));
 sg13g2_buf_1 _15776_ (.A(\cpu.spi.r_in[3] ),
    .X(_09069_));
 sg13g2_buf_1 _15777_ (.A(\cpu.spi.r_in[6] ),
    .X(_09070_));
 sg13g2_buf_1 _15778_ (.A(\cpu.spi.r_in[1] ),
    .X(_09071_));
 sg13g2_buf_1 _15779_ (.A(\cpu.spi.r_in[0] ),
    .X(_09072_));
 sg13g2_nand2_1 _15780_ (.Y(_09073_),
    .A(_09071_),
    .B(_09072_));
 sg13g2_nand3_1 _15781_ (.B(_09070_),
    .C(_09073_),
    .A(_09069_),
    .Y(_09074_));
 sg13g2_buf_1 _15782_ (.A(\cpu.spi.r_in[2] ),
    .X(_09075_));
 sg13g2_buf_1 _15783_ (.A(\cpu.spi.r_in[5] ),
    .X(_09076_));
 sg13g2_buf_1 _15784_ (.A(\cpu.spi.r_in[4] ),
    .X(_09077_));
 sg13g2_nand4_1 _15785_ (.B(_09076_),
    .C(_09077_),
    .A(_09075_),
    .Y(_09078_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _15786_ (.A(_09074_),
    .B(_09078_),
    .Y(_09079_));
 sg13g2_o21ai_1 _15787_ (.B1(_09066_),
    .Y(_09080_),
    .A1(_00222_),
    .A2(_09079_));
 sg13g2_nand2_2 _15788_ (.Y(_09081_),
    .A(_09068_),
    .B(_09080_));
 sg13g2_nand3_1 _15789_ (.B(net371),
    .C(_09081_),
    .A(_09046_),
    .Y(_09082_));
 sg13g2_o21ai_1 _15790_ (.B1(_09082_),
    .Y(_09083_),
    .A1(_09018_),
    .A2(_09044_));
 sg13g2_and2_1 _15791_ (.A(net691),
    .B(_09083_),
    .X(_00030_));
 sg13g2_buf_1 _15792_ (.A(net1084),
    .X(_09084_));
 sg13g2_buf_1 _15793_ (.A(net1016),
    .X(_09085_));
 sg13g2_buf_1 _15794_ (.A(net131),
    .X(_09086_));
 sg13g2_a21oi_1 _15795_ (.A1(_09085_),
    .A2(net110),
    .Y(_09087_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_buf_2 _15796_ (.A(\cpu.spi.r_state[4] ),
    .X(_09088_));
 sg13g2_inv_1 _15797_ (.Y(_09089_),
    .A(_09045_));
 sg13g2_nor2_1 _15798_ (.A(_09089_),
    .B(_09081_),
    .Y(_09090_));
 sg13g2_nor3_1 _15799_ (.A(_09088_),
    .B(net406),
    .C(_09090_),
    .Y(_09091_));
 sg13g2_buf_1 _15800_ (.A(\cpu.spi.r_state[2] ),
    .X(_09092_));
 sg13g2_buf_1 _15801_ (.A(net879),
    .X(_09093_));
 sg13g2_o21ai_1 _15802_ (.B1(net759),
    .Y(_09094_),
    .A1(net1083),
    .A2(net371));
 sg13g2_a21oi_1 _15803_ (.A1(_09087_),
    .A2(_09091_),
    .Y(_00031_),
    .B1(_09094_));
 sg13g2_buf_1 _15804_ (.A(_09030_),
    .X(_09095_));
 sg13g2_buf_1 _15805_ (.A(net877),
    .X(_09096_));
 sg13g2_buf_1 _15806_ (.A(_09096_),
    .X(_09097_));
 sg13g2_nor3_1 _15807_ (.A(net690),
    .B(net371),
    .C(_09028_),
    .Y(_00032_));
 sg13g2_nand3_1 _15808_ (.B(_08966_),
    .C(_09086_),
    .A(_09031_),
    .Y(_09098_));
 sg13g2_nand2_1 _15809_ (.Y(_09099_),
    .A(_09088_),
    .B(net406));
 sg13g2_buf_1 _15810_ (.A(_09096_),
    .X(_09100_));
 sg13g2_a21oi_1 _15811_ (.A1(_09098_),
    .A2(_09099_),
    .Y(_00033_),
    .B1(_09100_));
 sg13g2_nor3_1 _15812_ (.A(net690),
    .B(net371),
    .C(_09087_),
    .Y(_00034_));
 sg13g2_nand2_1 _15813_ (.Y(_09101_),
    .A(_09046_),
    .B(net406));
 sg13g2_nand2_1 _15814_ (.Y(_09102_),
    .A(net1083),
    .B(net371));
 sg13g2_buf_2 _15815_ (.A(net877),
    .X(_09103_));
 sg13g2_buf_1 _15816_ (.A(_09103_),
    .X(_09104_));
 sg13g2_a21oi_1 _15817_ (.A1(_09101_),
    .A2(_09102_),
    .Y(_00035_),
    .B1(_09104_));
 sg13g2_buf_1 _15818_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09105_));
 sg13g2_buf_2 _15819_ (.A(\cpu.dec.mult ),
    .X(_09106_));
 sg13g2_nand3b_1 _15820_ (.B(\cpu.dec.iready ),
    .C(_00199_),
    .Y(_09107_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_2 _15821_ (.A(_09107_),
    .X(_09108_));
 sg13g2_nor2_1 _15822_ (.A(_09029_),
    .B(_09108_),
    .Y(_09109_));
 sg13g2_buf_2 _15823_ (.A(_09109_),
    .X(_09110_));
 sg13g2_and2_1 _15824_ (.A(_09106_),
    .B(_09110_),
    .X(_09111_));
 sg13g2_buf_2 _15825_ (.A(_09111_),
    .X(_09112_));
 sg13g2_buf_1 _15826_ (.A(\cpu.dec.div ),
    .X(_09113_));
 sg13g2_and2_1 _15827_ (.A(_09113_),
    .B(_09110_),
    .X(_09114_));
 sg13g2_buf_2 _15828_ (.A(_09114_),
    .X(_09115_));
 sg13g2_nor2_2 _15829_ (.A(_09112_),
    .B(_09115_),
    .Y(_09116_));
 sg13g2_nand2_1 _15830_ (.Y(_09117_),
    .A(_09105_),
    .B(_09116_));
 sg13g2_buf_2 _15831_ (.A(_09117_),
    .X(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _15832_ (.A(\cpu.ex.r_div_running ),
    .X(_09118_));
 sg13g2_buf_1 _15833_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09119_));
 sg13g2_nor4_2 _15834_ (.A(_09119_),
    .B(\cpu.ex.r_mult_off[2] ),
    .C(\cpu.ex.r_mult_off[3] ),
    .Y(_09120_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _15835_ (.A(_09115_),
    .X(_09121_));
 sg13g2_o21ai_1 _15836_ (.B1(net1018),
    .Y(_09122_),
    .A1(_09118_),
    .A2(_09121_));
 sg13g2_a21oi_1 _15837_ (.A1(_09118_),
    .A2(_09120_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09122_));
 sg13g2_buf_1 _15838_ (.A(\cpu.ex.r_mult_running ),
    .X(_09123_));
 sg13g2_inv_2 _15839_ (.Y(_09124_),
    .A(_09123_));
 sg13g2_nand2_1 _15840_ (.Y(_09125_),
    .A(_09106_),
    .B(_09110_));
 sg13g2_buf_1 _15841_ (.A(_09125_),
    .X(_09126_));
 sg13g2_nand2_2 _15842_ (.Y(_09127_),
    .A(_09124_),
    .B(_09126_));
 sg13g2_nand2_1 _15843_ (.Y(_09128_),
    .A(net1018),
    .B(_09127_));
 sg13g2_a21oi_1 _15844_ (.A1(_09123_),
    .A2(_09120_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09128_));
 sg13g2_buf_1 _15845_ (.A(\cpu.qspi.r_state[17] ),
    .X(_09129_));
 sg13g2_buf_1 _15846_ (.A(_08515_),
    .X(_09130_));
 sg13g2_buf_1 _15847_ (.A(\cpu.dcache.flush_write ),
    .X(_09131_));
 sg13g2_inv_1 _15848_ (.Y(_09132_),
    .A(_09131_));
 sg13g2_inv_1 _15849_ (.Y(_09133_),
    .A(_00244_));
 sg13g2_buf_2 _15850_ (.A(\cpu.addr[4] ),
    .X(_09134_));
 sg13g2_or2_1 _15851_ (.X(_09135_),
    .B(net1023),
    .A(_09134_));
 sg13g2_buf_1 _15852_ (.A(_09135_),
    .X(_09136_));
 sg13g2_buf_1 _15853_ (.A(_00227_),
    .X(_09137_));
 sg13g2_and2_1 _15854_ (.A(net1021),
    .B(_09137_),
    .X(_09138_));
 sg13g2_buf_1 _15855_ (.A(_09138_),
    .X(_09139_));
 sg13g2_nor2_1 _15856_ (.A(_09136_),
    .B(_09139_),
    .Y(_09140_));
 sg13g2_buf_1 _15857_ (.A(_09140_),
    .X(_09141_));
 sg13g2_buf_1 _15858_ (.A(net593),
    .X(_09142_));
 sg13g2_nor2b_1 _15859_ (.A(_08957_),
    .B_N(_09137_),
    .Y(_09143_));
 sg13g2_and2_1 _15860_ (.A(net1023),
    .B(_09143_),
    .X(_09144_));
 sg13g2_buf_1 _15861_ (.A(_09144_),
    .X(_09145_));
 sg13g2_buf_1 _15862_ (.A(_09145_),
    .X(_09146_));
 sg13g2_buf_1 _15863_ (.A(net687),
    .X(_09147_));
 sg13g2_a22oi_1 _15864_ (.Y(_09148_),
    .B1(_09147_),
    .B2(\cpu.dcache.r_tag[2][13] ),
    .A2(net536),
    .A1(_09133_));
 sg13g2_buf_1 _15865_ (.A(_09134_),
    .X(_09149_));
 sg13g2_nor2b_1 _15866_ (.A(_08941_),
    .B_N(_08957_),
    .Y(_09150_));
 sg13g2_buf_2 _15867_ (.A(_09150_),
    .X(_09151_));
 sg13g2_and2_1 _15868_ (.A(net1014),
    .B(_09151_),
    .X(_09152_));
 sg13g2_buf_2 _15869_ (.A(_09152_),
    .X(_09153_));
 sg13g2_buf_1 _15870_ (.A(_09153_),
    .X(_09154_));
 sg13g2_buf_1 _15871_ (.A(_09137_),
    .X(_09155_));
 sg13g2_and2_1 _15872_ (.A(_08957_),
    .B(_08941_),
    .X(_09156_));
 sg13g2_buf_2 _15873_ (.A(_09156_),
    .X(_09157_));
 sg13g2_and2_1 _15874_ (.A(net1013),
    .B(_09157_),
    .X(_09158_));
 sg13g2_buf_1 _15875_ (.A(_09158_),
    .X(_09159_));
 sg13g2_buf_1 _15876_ (.A(_09159_),
    .X(_09160_));
 sg13g2_buf_1 _15877_ (.A(net590),
    .X(_09161_));
 sg13g2_a22oi_1 _15878_ (.Y(_09162_),
    .B1(net535),
    .B2(\cpu.dcache.r_tag[3][13] ),
    .A2(net591),
    .A1(\cpu.dcache.r_tag[5][13] ));
 sg13g2_inv_2 _15879_ (.Y(_09163_),
    .A(_09134_));
 sg13g2_nand2_1 _15880_ (.Y(_09164_),
    .A(net1021),
    .B(net1023));
 sg13g2_nor2_1 _15881_ (.A(_09163_),
    .B(_09164_),
    .Y(_09165_));
 sg13g2_buf_1 _15882_ (.A(_09165_),
    .X(_09166_));
 sg13g2_nand2b_1 _15883_ (.Y(_09167_),
    .B(_09134_),
    .A_N(net1021));
 sg13g2_nor2_1 _15884_ (.A(net882),
    .B(_09167_),
    .Y(_09168_));
 sg13g2_buf_1 _15885_ (.A(_09168_),
    .X(_09169_));
 sg13g2_buf_1 _15886_ (.A(net685),
    .X(_09170_));
 sg13g2_a22oi_1 _15887_ (.Y(_09171_),
    .B1(_09170_),
    .B2(\cpu.dcache.r_tag[4][13] ),
    .A2(net686),
    .A1(\cpu.dcache.r_tag[7][13] ));
 sg13g2_and2_1 _15888_ (.A(net1013),
    .B(_09151_),
    .X(_09172_));
 sg13g2_buf_1 _15889_ (.A(_09172_),
    .X(_09173_));
 sg13g2_buf_1 _15890_ (.A(_09173_),
    .X(_09174_));
 sg13g2_buf_1 _15891_ (.A(net588),
    .X(_09175_));
 sg13g2_nor2_1 _15892_ (.A(_09040_),
    .B(_09167_),
    .Y(_09176_));
 sg13g2_buf_2 _15893_ (.A(_09176_),
    .X(_09177_));
 sg13g2_buf_1 _15894_ (.A(_09177_),
    .X(_09178_));
 sg13g2_a22oi_1 _15895_ (.Y(_09179_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][13] ),
    .A2(net534),
    .A1(\cpu.dcache.r_tag[1][13] ));
 sg13g2_nand4_1 _15896_ (.B(_09162_),
    .C(_09171_),
    .A(_09148_),
    .Y(_09180_),
    .D(_09179_));
 sg13g2_buf_1 _15897_ (.A(_08606_),
    .X(_09181_));
 sg13g2_buf_8 _15898_ (.A(net1027),
    .X(_09182_));
 sg13g2_buf_1 _15899_ (.A(net876),
    .X(_09183_));
 sg13g2_buf_2 _15900_ (.A(net758),
    .X(_09184_));
 sg13g2_buf_1 _15901_ (.A(net886),
    .X(_09185_));
 sg13g2_buf_1 _15902_ (.A(net757),
    .X(_09186_));
 sg13g2_mux4_1 _15903_ (.S0(_09184_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net683),
    .X(_09187_));
 sg13g2_mux4_1 _15904_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net683),
    .X(_09188_));
 sg13g2_mux4_1 _15905_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net683),
    .X(_09189_));
 sg13g2_mux4_1 _15906_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net683),
    .X(_09190_));
 sg13g2_buf_1 _15907_ (.A(_08529_),
    .X(_09191_));
 sg13g2_buf_2 _15908_ (.A(_09191_),
    .X(_09192_));
 sg13g2_buf_2 _15909_ (.A(_08602_),
    .X(_09193_));
 sg13g2_buf_2 _15910_ (.A(net755),
    .X(_09194_));
 sg13g2_mux4_1 _15911_ (.S0(_09192_),
    .A0(_09187_),
    .A1(_09188_),
    .A2(_09189_),
    .A3(_09190_),
    .S1(_09194_),
    .X(_09195_));
 sg13g2_buf_1 _15912_ (.A(_08519_),
    .X(_09196_));
 sg13g2_mux4_1 _15913_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net757),
    .X(_09197_));
 sg13g2_mux4_1 _15914_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net757),
    .X(_09198_));
 sg13g2_mux4_1 _15915_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net757),
    .X(_09199_));
 sg13g2_mux4_1 _15916_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net757),
    .X(_09200_));
 sg13g2_mux4_1 _15917_ (.S0(net756),
    .A0(_09197_),
    .A1(_09198_),
    .A2(_09199_),
    .A3(_09200_),
    .S1(net755),
    .X(_09201_));
 sg13g2_and2_1 _15918_ (.A(net680),
    .B(_09201_),
    .X(_09202_));
 sg13g2_a21oi_1 _15919_ (.A1(net586),
    .A2(_09195_),
    .Y(_09203_),
    .B1(_09202_));
 sg13g2_nor2_1 _15920_ (.A(net1096),
    .B(net683),
    .Y(_09204_));
 sg13g2_a21oi_2 _15921_ (.B1(_09204_),
    .Y(_09205_),
    .A2(_09203_),
    .A1(_08054_));
 sg13g2_buf_1 _15922_ (.A(_09205_),
    .X(_09206_));
 sg13g2_xor2_1 _15923_ (.B(_09206_),
    .A(_09180_),
    .X(_09207_));
 sg13g2_buf_1 _15924_ (.A(net587),
    .X(_09208_));
 sg13g2_a22oi_1 _15925_ (.Y(_09209_),
    .B1(_09208_),
    .B2(\cpu.dcache.r_tag[6][12] ),
    .A2(net534),
    .A1(\cpu.dcache.r_tag[1][12] ));
 sg13g2_inv_1 _15926_ (.Y(_09210_),
    .A(_00243_));
 sg13g2_a22oi_1 _15927_ (.Y(_09211_),
    .B1(net591),
    .B2(\cpu.dcache.r_tag[5][12] ),
    .A2(net536),
    .A1(_09210_));
 sg13g2_buf_1 _15928_ (.A(net686),
    .X(_09212_));
 sg13g2_a22oi_1 _15929_ (.Y(_09213_),
    .B1(_09212_),
    .B2(\cpu.dcache.r_tag[7][12] ),
    .A2(_09161_),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_a22oi_1 _15930_ (.Y(_09214_),
    .B1(_09170_),
    .B2(\cpu.dcache.r_tag[4][12] ),
    .A2(_09147_),
    .A1(\cpu.dcache.r_tag[2][12] ));
 sg13g2_nand4_1 _15931_ (.B(_09211_),
    .C(_09213_),
    .A(_09209_),
    .Y(_09215_),
    .D(_09214_));
 sg13g2_mux4_1 _15932_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net683),
    .X(_09216_));
 sg13g2_mux4_1 _15933_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(_09186_),
    .X(_09217_));
 sg13g2_mux4_1 _15934_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(net683),
    .X(_09218_));
 sg13g2_mux4_1 _15935_ (.S0(_09184_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(_09186_),
    .X(_09219_));
 sg13g2_buf_1 _15936_ (.A(net756),
    .X(_09220_));
 sg13g2_mux4_1 _15937_ (.S0(net679),
    .A0(_09216_),
    .A1(_09217_),
    .A2(_09218_),
    .A3(_09219_),
    .S1(_09194_),
    .X(_09221_));
 sg13g2_buf_8 _15938_ (.A(_09182_),
    .X(_09222_));
 sg13g2_buf_8 _15939_ (.A(_09222_),
    .X(_09223_));
 sg13g2_buf_1 _15940_ (.A(net886),
    .X(_09224_));
 sg13g2_buf_1 _15941_ (.A(_09224_),
    .X(_09225_));
 sg13g2_mux4_1 _15942_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net677),
    .X(_09226_));
 sg13g2_mux4_1 _15943_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net677),
    .X(_09227_));
 sg13g2_mux4_1 _15944_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net757),
    .X(_09228_));
 sg13g2_mux4_1 _15945_ (.S0(net758),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net757),
    .X(_09229_));
 sg13g2_mux4_1 _15946_ (.S0(net682),
    .A0(_09226_),
    .A1(_09227_),
    .A2(_09228_),
    .A3(_09229_),
    .S1(net755),
    .X(_09230_));
 sg13g2_and2_1 _15947_ (.A(net680),
    .B(_09230_),
    .X(_09231_));
 sg13g2_a21oi_1 _15948_ (.A1(net586),
    .A2(_09221_),
    .Y(_09232_),
    .B1(_09231_));
 sg13g2_nor2_1 _15949_ (.A(_08054_),
    .B(net684),
    .Y(_09233_));
 sg13g2_a21oi_2 _15950_ (.B1(_09233_),
    .Y(_09234_),
    .A2(_09232_),
    .A1(net1042));
 sg13g2_buf_1 _15951_ (.A(_09234_),
    .X(_09235_));
 sg13g2_xor2_1 _15952_ (.B(net338),
    .A(_09215_),
    .X(_09236_));
 sg13g2_buf_8 _15953_ (.A(net758),
    .X(_09237_));
 sg13g2_buf_2 _15954_ (.A(net757),
    .X(_09238_));
 sg13g2_mux4_1 _15955_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net675),
    .X(_09239_));
 sg13g2_mux4_1 _15956_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net675),
    .X(_09240_));
 sg13g2_buf_8 _15957_ (.A(_09183_),
    .X(_09241_));
 sg13g2_buf_2 _15958_ (.A(_09185_),
    .X(_09242_));
 sg13g2_mux4_1 _15959_ (.S0(_09241_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(_09242_),
    .X(_09243_));
 sg13g2_mux4_1 _15960_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net673),
    .X(_09244_));
 sg13g2_mux4_1 _15961_ (.S0(net682),
    .A0(_09239_),
    .A1(_09240_),
    .A2(_09243_),
    .A3(_09244_),
    .S1(net681),
    .X(_09245_));
 sg13g2_nand2_1 _15962_ (.Y(_09246_),
    .A(net680),
    .B(_09245_));
 sg13g2_mux4_1 _15963_ (.S0(_09237_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(_09238_),
    .X(_09247_));
 sg13g2_mux4_1 _15964_ (.S0(_09237_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(_09238_),
    .X(_09248_));
 sg13g2_mux4_1 _15965_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net673),
    .X(_09249_));
 sg13g2_mux4_1 _15966_ (.S0(_09241_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(_09242_),
    .X(_09250_));
 sg13g2_mux4_1 _15967_ (.S0(net682),
    .A0(_09247_),
    .A1(_09248_),
    .A2(_09249_),
    .A3(_09250_),
    .S1(net681),
    .X(_09251_));
 sg13g2_nand2_1 _15968_ (.Y(_09252_),
    .A(net586),
    .B(_09251_));
 sg13g2_a21oi_2 _15969_ (.B1(_08173_),
    .Y(_09253_),
    .A2(_09252_),
    .A1(_09246_));
 sg13g2_buf_1 _15970_ (.A(_09253_),
    .X(_09254_));
 sg13g2_nand2_1 _15971_ (.Y(_09255_),
    .A(\cpu.dcache.r_tag[2][21] ),
    .B(net592));
 sg13g2_a22oi_1 _15972_ (.Y(_09256_),
    .B1(_09175_),
    .B2(\cpu.dcache.r_tag[1][21] ),
    .A2(net535),
    .A1(\cpu.dcache.r_tag[3][21] ));
 sg13g2_a22oi_1 _15973_ (.Y(_09257_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][21] ),
    .A2(_09142_),
    .A1(\cpu.dcache.r_tag[0][21] ));
 sg13g2_mux2_1 _15974_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(\cpu.dcache.r_tag[7][21] ),
    .S(net763),
    .X(_09258_));
 sg13g2_nor2_1 _15975_ (.A(net1021),
    .B(net1023),
    .Y(_09259_));
 sg13g2_buf_2 _15976_ (.A(_09259_),
    .X(_09260_));
 sg13g2_a22oi_1 _15977_ (.Y(_09261_),
    .B1(_09260_),
    .B2(\cpu.dcache.r_tag[4][21] ),
    .A2(_09258_),
    .A1(net762));
 sg13g2_buf_1 _15978_ (.A(net1014),
    .X(_09262_));
 sg13g2_nand2b_1 _15979_ (.Y(_09263_),
    .B(_09262_),
    .A_N(_09261_));
 sg13g2_nand4_1 _15980_ (.B(_09256_),
    .C(_09257_),
    .A(_09255_),
    .Y(_09264_),
    .D(_09263_));
 sg13g2_xnor2_1 _15981_ (.Y(_09265_),
    .A(net369),
    .B(_09264_));
 sg13g2_buf_8 _15982_ (.A(net876),
    .X(_09266_));
 sg13g2_buf_2 _15983_ (.A(net752),
    .X(_09267_));
 sg13g2_buf_1 _15984_ (.A(_09185_),
    .X(_09268_));
 sg13g2_mux4_1 _15985_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net671),
    .X(_09269_));
 sg13g2_mux4_1 _15986_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net671),
    .X(_09270_));
 sg13g2_buf_2 _15987_ (.A(net752),
    .X(_09271_));
 sg13g2_buf_1 _15988_ (.A(net886),
    .X(_09272_));
 sg13g2_buf_1 _15989_ (.A(net751),
    .X(_09273_));
 sg13g2_mux4_1 _15990_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net669),
    .X(_09274_));
 sg13g2_mux4_1 _15991_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net669),
    .X(_09275_));
 sg13g2_mux4_1 _15992_ (.S0(net682),
    .A0(_09269_),
    .A1(_09270_),
    .A2(_09274_),
    .A3(_09275_),
    .S1(net681),
    .X(_09276_));
 sg13g2_nand2_1 _15993_ (.Y(_09277_),
    .A(_09196_),
    .B(_09276_));
 sg13g2_mux4_1 _15994_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net671),
    .X(_09278_));
 sg13g2_mux4_1 _15995_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net671),
    .X(_09279_));
 sg13g2_mux4_1 _15996_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net677),
    .X(_09280_));
 sg13g2_mux4_1 _15997_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(net677),
    .X(_09281_));
 sg13g2_mux4_1 _15998_ (.S0(net682),
    .A0(_09278_),
    .A1(_09279_),
    .A2(_09280_),
    .A3(_09281_),
    .S1(_09193_),
    .X(_09282_));
 sg13g2_nand2_1 _15999_ (.Y(_09283_),
    .A(net586),
    .B(_09282_));
 sg13g2_a21oi_2 _16000_ (.B1(_08172_),
    .Y(_09284_),
    .A2(_09283_),
    .A1(_09277_));
 sg13g2_buf_1 _16001_ (.A(_09284_),
    .X(_09285_));
 sg13g2_a22oi_1 _16002_ (.Y(_09286_),
    .B1(_09175_),
    .B2(\cpu.dcache.r_tag[1][16] ),
    .A2(net591),
    .A1(\cpu.dcache.r_tag[5][16] ));
 sg13g2_a22oi_1 _16003_ (.Y(_09287_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][16] ),
    .A2(net590),
    .A1(\cpu.dcache.r_tag[3][16] ));
 sg13g2_inv_1 _16004_ (.Y(_09288_),
    .A(_00247_));
 sg13g2_a22oi_1 _16005_ (.Y(_09289_),
    .B1(net686),
    .B2(\cpu.dcache.r_tag[7][16] ),
    .A2(net593),
    .A1(_09288_));
 sg13g2_a22oi_1 _16006_ (.Y(_09290_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][16] ),
    .A2(net687),
    .A1(\cpu.dcache.r_tag[2][16] ));
 sg13g2_nand4_1 _16007_ (.B(_09287_),
    .C(_09289_),
    .A(_09286_),
    .Y(_09291_),
    .D(_09290_));
 sg13g2_xnor2_1 _16008_ (.Y(_09292_),
    .A(_09285_),
    .B(_09291_));
 sg13g2_mux4_1 _16009_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net669),
    .X(_09293_));
 sg13g2_mux4_1 _16010_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net669),
    .X(_09294_));
 sg13g2_mux4_1 _16011_ (.S0(_09223_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(_09225_),
    .X(_09295_));
 sg13g2_mux4_1 _16012_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net677),
    .X(_09296_));
 sg13g2_mux4_1 _16013_ (.S0(net682),
    .A0(_09293_),
    .A1(_09294_),
    .A2(_09295_),
    .A3(_09296_),
    .S1(net755),
    .X(_09297_));
 sg13g2_nand2_1 _16014_ (.Y(_09298_),
    .A(_09196_),
    .B(_09297_));
 sg13g2_mux4_1 _16015_ (.S0(_09271_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(_09273_),
    .X(_09299_));
 sg13g2_mux4_1 _16016_ (.S0(_09271_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(_09273_),
    .X(_09300_));
 sg13g2_mux4_1 _16017_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(net677),
    .X(_09301_));
 sg13g2_mux4_1 _16018_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net677),
    .X(_09302_));
 sg13g2_mux4_1 _16019_ (.S0(_09192_),
    .A0(_09299_),
    .A1(_09300_),
    .A2(_09301_),
    .A3(_09302_),
    .S1(_09193_),
    .X(_09303_));
 sg13g2_nand2_1 _16020_ (.Y(_09304_),
    .A(_09181_),
    .B(_09303_));
 sg13g2_a21oi_2 _16021_ (.B1(_08172_),
    .Y(_09305_),
    .A2(_09304_),
    .A1(_09298_));
 sg13g2_buf_1 _16022_ (.A(_09305_),
    .X(_09306_));
 sg13g2_inv_1 _16023_ (.Y(_09307_),
    .A(_00250_));
 sg13g2_a22oi_1 _16024_ (.Y(_09308_),
    .B1(net687),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(net593),
    .A1(_09307_));
 sg13g2_a22oi_1 _16025_ (.Y(_09309_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][19] ),
    .A2(_09174_),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_a22oi_1 _16026_ (.Y(_09310_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(net686),
    .A1(\cpu.dcache.r_tag[7][19] ));
 sg13g2_a22oi_1 _16027_ (.Y(_09311_),
    .B1(net590),
    .B2(\cpu.dcache.r_tag[3][19] ),
    .A2(_09153_),
    .A1(\cpu.dcache.r_tag[5][19] ));
 sg13g2_nand4_1 _16028_ (.B(_09309_),
    .C(_09310_),
    .A(_09308_),
    .Y(_09312_),
    .D(_09311_));
 sg13g2_xnor2_1 _16029_ (.Y(_09313_),
    .A(_09306_),
    .B(_09312_));
 sg13g2_buf_2 _16030_ (.A(net1027),
    .X(_09314_));
 sg13g2_buf_2 _16031_ (.A(net886),
    .X(_09315_));
 sg13g2_mux4_1 _16032_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net750),
    .X(_09316_));
 sg13g2_mux4_1 _16033_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net750),
    .X(_09317_));
 sg13g2_mux4_1 _16034_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net750),
    .X(_09318_));
 sg13g2_mux4_1 _16035_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(_09315_),
    .X(_09319_));
 sg13g2_mux4_1 _16036_ (.S0(net756),
    .A0(_09316_),
    .A1(_09317_),
    .A2(_09318_),
    .A3(_09319_),
    .S1(net887),
    .X(_09320_));
 sg13g2_nand2_1 _16037_ (.Y(_09321_),
    .A(net680),
    .B(_09320_));
 sg13g2_mux4_1 _16038_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(net750),
    .X(_09322_));
 sg13g2_mux4_1 _16039_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(_09315_),
    .X(_09323_));
 sg13g2_mux4_1 _16040_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net886),
    .X(_09324_));
 sg13g2_mux4_1 _16041_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net886),
    .X(_09325_));
 sg13g2_mux4_1 _16042_ (.S0(_08529_),
    .A0(_09322_),
    .A1(_09323_),
    .A2(_09324_),
    .A3(_09325_),
    .S1(net887),
    .X(_09326_));
 sg13g2_nand2_1 _16043_ (.Y(_09327_),
    .A(_08606_),
    .B(_09326_));
 sg13g2_a21oi_2 _16044_ (.B1(_08172_),
    .Y(_09328_),
    .A2(_09327_),
    .A1(_09321_));
 sg13g2_buf_1 _16045_ (.A(_09328_),
    .X(_09329_));
 sg13g2_inv_1 _16046_ (.Y(_09330_),
    .A(_00251_));
 sg13g2_a22oi_1 _16047_ (.Y(_09331_),
    .B1(_09153_),
    .B2(\cpu.dcache.r_tag[5][23] ),
    .A2(net593),
    .A1(_09330_));
 sg13g2_a22oi_1 _16048_ (.Y(_09332_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][23] ),
    .A2(net686),
    .A1(\cpu.dcache.r_tag[7][23] ));
 sg13g2_a22oi_1 _16049_ (.Y(_09333_),
    .B1(net588),
    .B2(\cpu.dcache.r_tag[1][23] ),
    .A2(net687),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_a22oi_1 _16050_ (.Y(_09334_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][23] ),
    .A2(net590),
    .A1(\cpu.dcache.r_tag[3][23] ));
 sg13g2_nand4_1 _16051_ (.B(_09332_),
    .C(_09333_),
    .A(_09331_),
    .Y(_09335_),
    .D(_09334_));
 sg13g2_xor2_1 _16052_ (.B(_09335_),
    .A(net404),
    .X(_09336_));
 sg13g2_mux4_1 _16053_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net753),
    .X(_09337_));
 sg13g2_mux4_1 _16054_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net753),
    .X(_09338_));
 sg13g2_mux4_1 _16055_ (.S0(_09314_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net750),
    .X(_09339_));
 sg13g2_mux4_1 _16056_ (.S0(_09314_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net750),
    .X(_09340_));
 sg13g2_mux4_1 _16057_ (.S0(net756),
    .A0(_09337_),
    .A1(_09338_),
    .A2(_09339_),
    .A3(_09340_),
    .S1(net887),
    .X(_09341_));
 sg13g2_nand2_1 _16058_ (.Y(_09342_),
    .A(net680),
    .B(_09341_));
 sg13g2_mux4_1 _16059_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(net750),
    .X(_09343_));
 sg13g2_mux4_1 _16060_ (.S0(net874),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net750),
    .X(_09344_));
 sg13g2_mux4_1 _16061_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net886),
    .X(_09345_));
 sg13g2_mux4_1 _16062_ (.S0(net876),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net886),
    .X(_09346_));
 sg13g2_mux4_1 _16063_ (.S0(_08529_),
    .A0(_09343_),
    .A1(_09344_),
    .A2(_09345_),
    .A3(_09346_),
    .S1(net887),
    .X(_09347_));
 sg13g2_nand2_1 _16064_ (.Y(_09348_),
    .A(net586),
    .B(_09347_));
 sg13g2_a21oi_2 _16065_ (.B1(_08172_),
    .Y(_09349_),
    .A2(_09348_),
    .A1(_09342_));
 sg13g2_buf_1 _16066_ (.A(_09349_),
    .X(_09350_));
 sg13g2_inv_1 _16067_ (.Y(_09351_),
    .A(_00248_));
 sg13g2_a22oi_1 _16068_ (.Y(_09352_),
    .B1(net686),
    .B2(\cpu.dcache.r_tag[7][17] ),
    .A2(_09141_),
    .A1(_09351_));
 sg13g2_a22oi_1 _16069_ (.Y(_09353_),
    .B1(net588),
    .B2(\cpu.dcache.r_tag[1][17] ),
    .A2(_09153_),
    .A1(\cpu.dcache.r_tag[5][17] ));
 sg13g2_a22oi_1 _16070_ (.Y(_09354_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][17] ),
    .A2(net687),
    .A1(\cpu.dcache.r_tag[2][17] ));
 sg13g2_a22oi_1 _16071_ (.Y(_09355_),
    .B1(_09178_),
    .B2(\cpu.dcache.r_tag[6][17] ),
    .A2(net590),
    .A1(\cpu.dcache.r_tag[3][17] ));
 sg13g2_nand4_1 _16072_ (.B(_09353_),
    .C(_09354_),
    .A(_09352_),
    .Y(_09356_),
    .D(_09355_));
 sg13g2_xor2_1 _16073_ (.B(_09356_),
    .A(_09350_),
    .X(_09357_));
 sg13g2_mux4_1 _16074_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net753),
    .X(_09358_));
 sg13g2_mux4_1 _16075_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net751),
    .X(_09359_));
 sg13g2_mux4_1 _16076_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net753),
    .X(_09360_));
 sg13g2_mux4_1 _16077_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(_09224_),
    .X(_09361_));
 sg13g2_mux4_1 _16078_ (.S0(net756),
    .A0(_09358_),
    .A1(_09359_),
    .A2(_09360_),
    .A3(_09361_),
    .S1(net887),
    .X(_09362_));
 sg13g2_nand2_1 _16079_ (.Y(_09363_),
    .A(net680),
    .B(_09362_));
 sg13g2_mux4_1 _16080_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net753),
    .X(_09364_));
 sg13g2_mux4_1 _16081_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net753),
    .X(_09365_));
 sg13g2_mux4_1 _16082_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net753),
    .X(_09366_));
 sg13g2_mux4_1 _16083_ (.S0(net754),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net753),
    .X(_09367_));
 sg13g2_mux4_1 _16084_ (.S0(net756),
    .A0(_09364_),
    .A1(_09365_),
    .A2(_09366_),
    .A3(_09367_),
    .S1(net887),
    .X(_09368_));
 sg13g2_nand2_1 _16085_ (.Y(_09369_),
    .A(net586),
    .B(_09368_));
 sg13g2_a21oi_2 _16086_ (.B1(_08172_),
    .Y(_09370_),
    .A2(_09369_),
    .A1(_09363_));
 sg13g2_buf_1 _16087_ (.A(_09370_),
    .X(_09371_));
 sg13g2_nand2_1 _16088_ (.Y(_09372_),
    .A(\cpu.dcache.r_tag[3][22] ),
    .B(net590));
 sg13g2_a22oi_1 _16089_ (.Y(_09373_),
    .B1(_09169_),
    .B2(\cpu.dcache.r_tag[4][22] ),
    .A2(net593),
    .A1(\cpu.dcache.r_tag[0][22] ));
 sg13g2_a22oi_1 _16090_ (.Y(_09374_),
    .B1(net588),
    .B2(\cpu.dcache.r_tag[1][22] ),
    .A2(net687),
    .A1(\cpu.dcache.r_tag[2][22] ));
 sg13g2_nor2b_1 _16091_ (.A(_08958_),
    .B_N(_08942_),
    .Y(_09375_));
 sg13g2_buf_1 _16092_ (.A(_09375_),
    .X(_09376_));
 sg13g2_mux2_1 _16093_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(\cpu.dcache.r_tag[7][22] ),
    .S(net882),
    .X(_09377_));
 sg13g2_a22oi_1 _16094_ (.Y(_09378_),
    .B1(_09377_),
    .B2(net881),
    .A2(net749),
    .A1(\cpu.dcache.r_tag[6][22] ));
 sg13g2_nand2b_1 _16095_ (.Y(_09379_),
    .B(net1014),
    .A_N(_09378_));
 sg13g2_nand4_1 _16096_ (.B(_09373_),
    .C(_09374_),
    .A(_09372_),
    .Y(_09380_),
    .D(_09379_));
 sg13g2_xor2_1 _16097_ (.B(_09380_),
    .A(net402),
    .X(_09381_));
 sg13g2_mux4_1 _16098_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net751),
    .X(_09382_));
 sg13g2_mux4_1 _16099_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net751),
    .X(_09383_));
 sg13g2_mux4_1 _16100_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net751),
    .X(_09384_));
 sg13g2_mux4_1 _16101_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net751),
    .X(_09385_));
 sg13g2_mux4_1 _16102_ (.S0(net756),
    .A0(_09382_),
    .A1(_09383_),
    .A2(_09384_),
    .A3(_09385_),
    .S1(net755),
    .X(_09386_));
 sg13g2_nand2_1 _16103_ (.Y(_09387_),
    .A(net680),
    .B(_09386_));
 sg13g2_mux4_1 _16104_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net751),
    .X(_09388_));
 sg13g2_mux4_1 _16105_ (.S0(net752),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net751),
    .X(_09389_));
 sg13g2_mux4_1 _16106_ (.S0(_09222_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(_09272_),
    .X(_09390_));
 sg13g2_mux4_1 _16107_ (.S0(_09266_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(_09272_),
    .X(_09391_));
 sg13g2_mux4_1 _16108_ (.S0(net756),
    .A0(_09388_),
    .A1(_09389_),
    .A2(_09390_),
    .A3(_09391_),
    .S1(net755),
    .X(_09392_));
 sg13g2_nand2_1 _16109_ (.Y(_09393_),
    .A(net586),
    .B(_09392_));
 sg13g2_a21oi_2 _16110_ (.B1(_08172_),
    .Y(_09394_),
    .A2(_09393_),
    .A1(_09387_));
 sg13g2_buf_1 _16111_ (.A(_09394_),
    .X(_09395_));
 sg13g2_mux2_1 _16112_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(\cpu.dcache.r_tag[7][20] ),
    .S(net763),
    .X(_09396_));
 sg13g2_a22oi_1 _16113_ (.Y(_09397_),
    .B1(_09396_),
    .B2(net762),
    .A2(net749),
    .A1(\cpu.dcache.r_tag[6][20] ));
 sg13g2_mux2_1 _16114_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(\cpu.dcache.r_tag[3][20] ),
    .S(net882),
    .X(_09398_));
 sg13g2_a22oi_1 _16115_ (.Y(_09399_),
    .B1(_09398_),
    .B2(net881),
    .A2(net749),
    .A1(\cpu.dcache.r_tag[2][20] ));
 sg13g2_nor2b_1 _16116_ (.A(_09399_),
    .B_N(net1013),
    .Y(_09400_));
 sg13g2_a221oi_1 _16117_ (.B2(\cpu.dcache.r_tag[4][20] ),
    .C1(_09400_),
    .B1(net685),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .Y(_09401_),
    .A2(_09141_));
 sg13g2_o21ai_1 _16118_ (.B1(_09401_),
    .Y(_09402_),
    .A1(_09163_),
    .A2(_09397_));
 sg13g2_xor2_1 _16119_ (.B(_09402_),
    .A(net401),
    .X(_09403_));
 sg13g2_nor4_1 _16120_ (.A(_09336_),
    .B(_09357_),
    .C(_09381_),
    .D(_09403_),
    .Y(_09404_));
 sg13g2_nand4_1 _16121_ (.B(_09292_),
    .C(_09313_),
    .A(_09265_),
    .Y(_09405_),
    .D(_09404_));
 sg13g2_mux2_1 _16122_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(\cpu.dcache.r_tag[7][14] ),
    .S(net763),
    .X(_09406_));
 sg13g2_a22oi_1 _16123_ (.Y(_09407_),
    .B1(_09406_),
    .B2(_08960_),
    .A2(_09260_),
    .A1(\cpu.dcache.r_tag[4][14] ));
 sg13g2_inv_1 _16124_ (.Y(_09408_),
    .A(_00245_));
 sg13g2_mux2_1 _16125_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(\cpu.dcache.r_tag[3][14] ),
    .S(net763),
    .X(_09409_));
 sg13g2_a22oi_1 _16126_ (.Y(_09410_),
    .B1(_09376_),
    .B2(\cpu.dcache.r_tag[2][14] ),
    .A2(_09409_),
    .A1(net881));
 sg13g2_nor2b_1 _16127_ (.A(_09410_),
    .B_N(net1013),
    .Y(_09411_));
 sg13g2_a221oi_1 _16128_ (.B2(\cpu.dcache.r_tag[6][14] ),
    .C1(_09411_),
    .B1(net587),
    .A1(_09408_),
    .Y(_09412_),
    .A2(net593));
 sg13g2_o21ai_1 _16129_ (.B1(_09412_),
    .Y(_09413_),
    .A1(_09163_),
    .A2(_09407_));
 sg13g2_mux4_1 _16130_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net675),
    .X(_09414_));
 sg13g2_mux4_1 _16131_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net675),
    .X(_09415_));
 sg13g2_mux4_1 _16132_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net673),
    .X(_09416_));
 sg13g2_mux4_1 _16133_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net673),
    .X(_09417_));
 sg13g2_mux4_1 _16134_ (.S0(_08606_),
    .A0(_09414_),
    .A1(_09415_),
    .A2(_09416_),
    .A3(_09417_),
    .S1(_08527_),
    .X(_09418_));
 sg13g2_nand2_1 _16135_ (.Y(_09419_),
    .A(net1096),
    .B(_09418_));
 sg13g2_mux4_1 _16136_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net675),
    .X(_09420_));
 sg13g2_mux4_1 _16137_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net675),
    .X(_09421_));
 sg13g2_mux4_1 _16138_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net675),
    .X(_09422_));
 sg13g2_mux4_1 _16139_ (.S0(net676),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(net675),
    .X(_09423_));
 sg13g2_mux4_1 _16140_ (.S0(_08606_),
    .A0(_09420_),
    .A1(_09421_),
    .A2(_09422_),
    .A3(_09423_),
    .S1(_08527_),
    .X(_09424_));
 sg13g2_o21ai_1 _16141_ (.B1(net681),
    .Y(_09425_),
    .A1(_08345_),
    .A2(_09424_));
 sg13g2_o21ai_1 _16142_ (.B1(_09425_),
    .Y(_09426_),
    .A1(net681),
    .A2(_09419_));
 sg13g2_buf_1 _16143_ (.A(_09426_),
    .X(_09427_));
 sg13g2_xnor2_1 _16144_ (.Y(_09428_),
    .A(_09413_),
    .B(net366));
 sg13g2_nand2_1 _16145_ (.Y(_09429_),
    .A(net1013),
    .B(_09151_));
 sg13g2_buf_1 _16146_ (.A(_09429_),
    .X(_09430_));
 sg13g2_inv_1 _16147_ (.Y(_09431_),
    .A(\cpu.dcache.r_tag[6][9] ));
 sg13g2_nand3b_1 _16148_ (.B(_09134_),
    .C(_08941_),
    .Y(_09432_),
    .A_N(_08957_));
 sg13g2_buf_2 _16149_ (.A(_09432_),
    .X(_09433_));
 sg13g2_nand4_1 _16150_ (.B(net882),
    .C(net1013),
    .A(net1021),
    .Y(_09434_),
    .D(\cpu.dcache.r_tag[3][9] ));
 sg13g2_o21ai_1 _16151_ (.B1(_09434_),
    .Y(_09435_),
    .A1(_09431_),
    .A2(_09433_));
 sg13g2_nor2b_1 _16152_ (.A(net1021),
    .B_N(_09134_),
    .Y(_09436_));
 sg13g2_and3_1 _16153_ (.X(_09437_),
    .A(_09040_),
    .B(\cpu.dcache.r_tag[4][9] ),
    .C(_09436_));
 sg13g2_inv_1 _16154_ (.Y(_09438_),
    .A(\cpu.dcache.r_tag[2][9] ));
 sg13g2_nand3b_1 _16155_ (.B(net1023),
    .C(_09137_),
    .Y(_09439_),
    .A_N(net1021));
 sg13g2_buf_1 _16156_ (.A(_09439_),
    .X(_09440_));
 sg13g2_nor2_1 _16157_ (.A(_09438_),
    .B(_09440_),
    .Y(_09441_));
 sg13g2_inv_1 _16158_ (.Y(_09442_),
    .A(\cpu.dcache.r_tag[5][9] ));
 sg13g2_nand3b_1 _16159_ (.B(_09134_),
    .C(_08958_),
    .Y(_09443_),
    .A_N(_08942_));
 sg13g2_buf_1 _16160_ (.A(_09443_),
    .X(_09444_));
 sg13g2_nand4_1 _16161_ (.B(net1014),
    .C(net882),
    .A(net881),
    .Y(_09445_),
    .D(\cpu.dcache.r_tag[7][9] ));
 sg13g2_o21ai_1 _16162_ (.B1(_09445_),
    .Y(_09446_),
    .A1(_09442_),
    .A2(net748));
 sg13g2_nor4_1 _16163_ (.A(_09435_),
    .B(_09437_),
    .C(_09441_),
    .D(_09446_),
    .Y(_09447_));
 sg13g2_mux2_1 _16164_ (.A0(_00238_),
    .A1(_09447_),
    .S(_09136_),
    .X(_09448_));
 sg13g2_nor2_1 _16165_ (.A(\cpu.dcache.r_tag[1][9] ),
    .B(net668),
    .Y(_09449_));
 sg13g2_a22oi_1 _16166_ (.Y(_09450_),
    .B1(_09449_),
    .B2(_09447_),
    .A2(_09448_),
    .A1(net668));
 sg13g2_xnor2_1 _16167_ (.Y(_09451_),
    .A(_00237_),
    .B(_09450_));
 sg13g2_inv_1 _16168_ (.Y(_09452_),
    .A(_00234_));
 sg13g2_nor2_1 _16169_ (.A(_09134_),
    .B(net1023),
    .Y(_09453_));
 sg13g2_buf_2 _16170_ (.A(_09453_),
    .X(_09454_));
 sg13g2_nand2b_1 _16171_ (.Y(_09455_),
    .B(_09454_),
    .A_N(_09139_));
 sg13g2_buf_1 _16172_ (.A(_09455_),
    .X(_09456_));
 sg13g2_buf_1 _16173_ (.A(_09456_),
    .X(_09457_));
 sg13g2_a22oi_1 _16174_ (.Y(_09458_),
    .B1(_09177_),
    .B2(\cpu.dcache.r_tag[6][7] ),
    .A2(_09146_),
    .A1(\cpu.dcache.r_tag[2][7] ));
 sg13g2_a22oi_1 _16175_ (.Y(_09459_),
    .B1(net588),
    .B2(\cpu.dcache.r_tag[1][7] ),
    .A2(_09159_),
    .A1(\cpu.dcache.r_tag[3][7] ));
 sg13g2_mux2_1 _16176_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(\cpu.dcache.r_tag[7][7] ),
    .S(net882),
    .X(_09460_));
 sg13g2_a22oi_1 _16177_ (.Y(_09461_),
    .B1(_09460_),
    .B2(net881),
    .A2(_09260_),
    .A1(\cpu.dcache.r_tag[4][7] ));
 sg13g2_nand2b_1 _16178_ (.Y(_09462_),
    .B(net1014),
    .A_N(_09461_));
 sg13g2_nand4_1 _16179_ (.B(_09458_),
    .C(_09459_),
    .A(_09456_),
    .Y(_09463_),
    .D(_09462_));
 sg13g2_o21ai_1 _16180_ (.B1(_09463_),
    .Y(_09464_),
    .A1(_09452_),
    .A2(net532));
 sg13g2_xor2_1 _16181_ (.B(_09464_),
    .A(_00233_),
    .X(_09465_));
 sg13g2_inv_1 _16182_ (.Y(_09466_),
    .A(_00242_));
 sg13g2_a22oi_1 _16183_ (.Y(_09467_),
    .B1(_09166_),
    .B2(\cpu.dcache.r_tag[7][11] ),
    .A2(_09146_),
    .A1(\cpu.dcache.r_tag[2][11] ));
 sg13g2_a22oi_1 _16184_ (.Y(_09468_),
    .B1(_09174_),
    .B2(\cpu.dcache.r_tag[1][11] ),
    .A2(_09160_),
    .A1(\cpu.dcache.r_tag[3][11] ));
 sg13g2_mux2_1 _16185_ (.A0(\cpu.dcache.r_tag[4][11] ),
    .A1(\cpu.dcache.r_tag[6][11] ),
    .S(_08943_),
    .X(_09469_));
 sg13g2_inv_2 _16186_ (.Y(_09470_),
    .A(_08959_));
 sg13g2_a22oi_1 _16187_ (.Y(_09471_),
    .B1(_09469_),
    .B2(_09470_),
    .A2(_09151_),
    .A1(\cpu.dcache.r_tag[5][11] ));
 sg13g2_nand2b_1 _16188_ (.Y(_09472_),
    .B(net1014),
    .A_N(_09471_));
 sg13g2_nand4_1 _16189_ (.B(_09467_),
    .C(_09468_),
    .A(_09457_),
    .Y(_09473_),
    .D(_09472_));
 sg13g2_o21ai_1 _16190_ (.B1(_09473_),
    .Y(_09474_),
    .A1(_09466_),
    .A2(_09457_));
 sg13g2_xor2_1 _16191_ (.B(_09474_),
    .A(_00241_),
    .X(_09475_));
 sg13g2_buf_1 _16192_ (.A(_00229_),
    .X(_09476_));
 sg13g2_a22oi_1 _16193_ (.Y(_09477_),
    .B1(\cpu.dcache.r_tag[1][5] ),
    .B2(net1013),
    .A2(\cpu.dcache.r_tag[5][5] ),
    .A1(net1014));
 sg13g2_nand3_1 _16194_ (.B(_09155_),
    .C(\cpu.dcache.r_tag[3][5] ),
    .A(net882),
    .Y(_09478_));
 sg13g2_o21ai_1 _16195_ (.B1(_09478_),
    .Y(_09479_),
    .A1(net763),
    .A2(_09477_));
 sg13g2_nand2_1 _16196_ (.Y(_09480_),
    .A(net881),
    .B(_09479_));
 sg13g2_a22oi_1 _16197_ (.Y(_09481_),
    .B1(_09260_),
    .B2(\cpu.dcache.r_tag[4][5] ),
    .A2(_09157_),
    .A1(\cpu.dcache.r_tag[7][5] ));
 sg13g2_nand2b_1 _16198_ (.Y(_09482_),
    .B(net1014),
    .A_N(_09481_));
 sg13g2_nand2b_1 _16199_ (.Y(_09483_),
    .B(net593),
    .A_N(_00230_));
 sg13g2_a22oi_1 _16200_ (.Y(_09484_),
    .B1(_09177_),
    .B2(\cpu.dcache.r_tag[6][5] ),
    .A2(_09145_),
    .A1(\cpu.dcache.r_tag[2][5] ));
 sg13g2_and4_1 _16201_ (.A(_09480_),
    .B(_09482_),
    .C(_09483_),
    .D(_09484_),
    .X(_09485_));
 sg13g2_xnor2_1 _16202_ (.Y(_09486_),
    .A(_09476_),
    .B(_09485_));
 sg13g2_nor2_1 _16203_ (.A(_00240_),
    .B(_09456_),
    .Y(_09487_));
 sg13g2_mux2_1 _16204_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(\cpu.dcache.r_tag[7][10] ),
    .S(_08943_),
    .X(_09488_));
 sg13g2_a22oi_1 _16205_ (.Y(_09489_),
    .B1(_09488_),
    .B2(net881),
    .A2(_09260_),
    .A1(\cpu.dcache.r_tag[4][10] ));
 sg13g2_nor2_1 _16206_ (.A(_09163_),
    .B(_09489_),
    .Y(_09490_));
 sg13g2_a22oi_1 _16207_ (.Y(_09491_),
    .B1(_09436_),
    .B2(\cpu.dcache.r_tag[6][10] ),
    .A2(_09139_),
    .A1(\cpu.dcache.r_tag[3][10] ));
 sg13g2_nor2_1 _16208_ (.A(_09040_),
    .B(_09491_),
    .Y(_09492_));
 sg13g2_a22oi_1 _16209_ (.Y(_09493_),
    .B1(_09376_),
    .B2(\cpu.dcache.r_tag[2][10] ),
    .A2(_09151_),
    .A1(\cpu.dcache.r_tag[1][10] ));
 sg13g2_nor2b_1 _16210_ (.A(_09493_),
    .B_N(_09155_),
    .Y(_09494_));
 sg13g2_nor4_2 _16211_ (.A(_09487_),
    .B(_09490_),
    .C(_09492_),
    .Y(_09495_),
    .D(_09494_));
 sg13g2_xnor2_1 _16212_ (.Y(_09496_),
    .A(_00239_),
    .B(_09495_));
 sg13g2_buf_1 _16213_ (.A(_00235_),
    .X(_09497_));
 sg13g2_inv_1 _16214_ (.Y(_09498_),
    .A(_00236_));
 sg13g2_a22oi_1 _16215_ (.Y(_09499_),
    .B1(_09153_),
    .B2(\cpu.dcache.r_tag[5][8] ),
    .A2(_09140_),
    .A1(_09498_));
 sg13g2_a22oi_1 _16216_ (.Y(_09500_),
    .B1(_09177_),
    .B2(\cpu.dcache.r_tag[6][8] ),
    .A2(_09173_),
    .A1(\cpu.dcache.r_tag[1][8] ));
 sg13g2_a22oi_1 _16217_ (.Y(_09501_),
    .B1(_09160_),
    .B2(\cpu.dcache.r_tag[3][8] ),
    .A2(_09145_),
    .A1(\cpu.dcache.r_tag[2][8] ));
 sg13g2_a22oi_1 _16218_ (.Y(_09502_),
    .B1(_09169_),
    .B2(\cpu.dcache.r_tag[4][8] ),
    .A2(_09166_),
    .A1(\cpu.dcache.r_tag[7][8] ));
 sg13g2_and4_1 _16219_ (.A(_09499_),
    .B(_09500_),
    .C(_09501_),
    .D(_09502_),
    .X(_09503_));
 sg13g2_xnor2_1 _16220_ (.Y(_09504_),
    .A(_09497_),
    .B(_09503_));
 sg13g2_a22oi_1 _16221_ (.Y(_09505_),
    .B1(_09177_),
    .B2(\cpu.dcache.r_tag[6][6] ),
    .A2(_09159_),
    .A1(\cpu.dcache.r_tag[3][6] ));
 sg13g2_a22oi_1 _16222_ (.Y(_09506_),
    .B1(net588),
    .B2(\cpu.dcache.r_tag[1][6] ),
    .A2(_09145_),
    .A1(\cpu.dcache.r_tag[2][6] ));
 sg13g2_a22oi_1 _16223_ (.Y(_09507_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][6] ),
    .A2(_09165_),
    .A1(\cpu.dcache.r_tag[7][6] ));
 sg13g2_inv_1 _16224_ (.Y(_09508_),
    .A(_00232_));
 sg13g2_a22oi_1 _16225_ (.Y(_09509_),
    .B1(_09153_),
    .B2(\cpu.dcache.r_tag[5][6] ),
    .A2(_09140_),
    .A1(_09508_));
 sg13g2_and4_1 _16226_ (.A(_09505_),
    .B(_09506_),
    .C(_09507_),
    .D(_09509_),
    .X(_09510_));
 sg13g2_xnor2_1 _16227_ (.Y(_09511_),
    .A(_00231_),
    .B(_09510_));
 sg13g2_nand4_1 _16228_ (.B(_09496_),
    .C(_09504_),
    .A(_09486_),
    .Y(_09512_),
    .D(_09511_));
 sg13g2_nor4_1 _16229_ (.A(_09451_),
    .B(_09465_),
    .C(_09475_),
    .D(_09512_),
    .Y(_09513_));
 sg13g2_mux4_1 _16230_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net673),
    .X(_09514_));
 sg13g2_mux4_1 _16231_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net673),
    .X(_09515_));
 sg13g2_mux4_1 _16232_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net671),
    .X(_09516_));
 sg13g2_mux4_1 _16233_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net671),
    .X(_09517_));
 sg13g2_mux4_1 _16234_ (.S0(net682),
    .A0(_09514_),
    .A1(_09515_),
    .A2(_09516_),
    .A3(_09517_),
    .S1(net681),
    .X(_09518_));
 sg13g2_nand2_1 _16235_ (.Y(_09519_),
    .A(net680),
    .B(_09518_));
 sg13g2_mux4_1 _16236_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net673),
    .X(_09520_));
 sg13g2_mux4_1 _16237_ (.S0(net674),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(net673),
    .X(_09521_));
 sg13g2_mux4_1 _16238_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(net671),
    .X(_09522_));
 sg13g2_mux4_1 _16239_ (.S0(net672),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(net671),
    .X(_09523_));
 sg13g2_mux4_1 _16240_ (.S0(net682),
    .A0(_09520_),
    .A1(_09521_),
    .A2(_09522_),
    .A3(_09523_),
    .S1(net681),
    .X(_09524_));
 sg13g2_nand2_1 _16241_ (.Y(_09525_),
    .A(net586),
    .B(_09524_));
 sg13g2_a21oi_2 _16242_ (.B1(_08173_),
    .Y(_09526_),
    .A2(_09525_),
    .A1(_09519_));
 sg13g2_buf_1 _16243_ (.A(_09526_),
    .X(_09527_));
 sg13g2_inv_1 _16244_ (.Y(_09528_),
    .A(_00249_));
 sg13g2_a22oi_1 _16245_ (.Y(_09529_),
    .B1(net687),
    .B2(\cpu.dcache.r_tag[2][18] ),
    .A2(_09142_),
    .A1(_09528_));
 sg13g2_a22oi_1 _16246_ (.Y(_09530_),
    .B1(net590),
    .B2(\cpu.dcache.r_tag[3][18] ),
    .A2(_09154_),
    .A1(\cpu.dcache.r_tag[5][18] ));
 sg13g2_a22oi_1 _16247_ (.Y(_09531_),
    .B1(net589),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(net686),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_a22oi_1 _16248_ (.Y(_09532_),
    .B1(net587),
    .B2(\cpu.dcache.r_tag[6][18] ),
    .A2(net588),
    .A1(\cpu.dcache.r_tag[1][18] ));
 sg13g2_nand4_1 _16249_ (.B(_09530_),
    .C(_09531_),
    .A(_09529_),
    .Y(_09533_),
    .D(_09532_));
 sg13g2_xnor2_1 _16250_ (.Y(_09534_),
    .A(_09527_),
    .B(_09533_));
 sg13g2_inv_1 _16251_ (.Y(_09535_),
    .A(_00246_));
 sg13g2_a22oi_1 _16252_ (.Y(_09536_),
    .B1(_09154_),
    .B2(\cpu.dcache.r_tag[5][15] ),
    .A2(net593),
    .A1(_09535_));
 sg13g2_a22oi_1 _16253_ (.Y(_09537_),
    .B1(net685),
    .B2(\cpu.dcache.r_tag[4][15] ),
    .A2(net686),
    .A1(\cpu.dcache.r_tag[7][15] ));
 sg13g2_a22oi_1 _16254_ (.Y(_09538_),
    .B1(net590),
    .B2(\cpu.dcache.r_tag[3][15] ),
    .A2(net687),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_a22oi_1 _16255_ (.Y(_09539_),
    .B1(_09178_),
    .B2(\cpu.dcache.r_tag[6][15] ),
    .A2(net588),
    .A1(\cpu.dcache.r_tag[1][15] ));
 sg13g2_nand4_1 _16256_ (.B(_09537_),
    .C(_09538_),
    .A(_09536_),
    .Y(_09540_),
    .D(_09539_));
 sg13g2_mux4_1 _16257_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net669),
    .X(_09541_));
 sg13g2_mux4_1 _16258_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net669),
    .X(_09542_));
 sg13g2_mux4_1 _16259_ (.S0(net678),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net677),
    .X(_09543_));
 sg13g2_mux4_1 _16260_ (.S0(_09223_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(_09225_),
    .X(_09544_));
 sg13g2_mux4_1 _16261_ (.S0(_08606_),
    .A0(_09541_),
    .A1(_09542_),
    .A2(_09543_),
    .A3(_09544_),
    .S1(net755),
    .X(_09545_));
 sg13g2_nand2_1 _16262_ (.Y(_09546_),
    .A(net1096),
    .B(_09545_));
 sg13g2_mux4_1 _16263_ (.S0(_09267_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(_09268_),
    .X(_09547_));
 sg13g2_mux4_1 _16264_ (.S0(_09267_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(_09268_),
    .X(_09548_));
 sg13g2_mux4_1 _16265_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net669),
    .X(_09549_));
 sg13g2_mux4_1 _16266_ (.S0(net670),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net669),
    .X(_09550_));
 sg13g2_mux4_1 _16267_ (.S0(_08606_),
    .A0(_09547_),
    .A1(_09548_),
    .A2(_09549_),
    .A3(_09550_),
    .S1(net755),
    .X(_09551_));
 sg13g2_o21ai_1 _16268_ (.B1(_08527_),
    .Y(_09552_),
    .A1(_08345_),
    .A2(_09551_));
 sg13g2_o21ai_1 _16269_ (.B1(_09552_),
    .Y(_09553_),
    .A1(_08527_),
    .A2(_09546_));
 sg13g2_buf_1 _16270_ (.A(_09553_),
    .X(_09554_));
 sg13g2_xnor2_1 _16271_ (.Y(_09555_),
    .A(_09540_),
    .B(_09554_));
 sg13g2_nand4_1 _16272_ (.B(_09513_),
    .C(_09534_),
    .A(_09428_),
    .Y(_09556_),
    .D(_09555_));
 sg13g2_nor4_1 _16273_ (.A(_09207_),
    .B(_09236_),
    .C(_09405_),
    .D(_09556_),
    .Y(_09557_));
 sg13g2_mux4_1 _16274_ (.S0(_08960_),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net763),
    .X(_09558_));
 sg13g2_mux4_1 _16275_ (.S0(net762),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net763),
    .X(_09559_));
 sg13g2_mux2_1 _16276_ (.A0(_09558_),
    .A1(_09559_),
    .S(_09163_),
    .X(_09560_));
 sg13g2_mux4_1 _16277_ (.S0(net762),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(_08945_),
    .X(_09561_));
 sg13g2_mux4_1 _16278_ (.S0(net762),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(_08945_),
    .X(_09562_));
 sg13g2_mux2_1 _16279_ (.A0(_09561_),
    .A1(_09562_),
    .S(_09163_),
    .X(_09563_));
 sg13g2_nand3_1 _16280_ (.B(_09560_),
    .C(_09563_),
    .A(_09011_),
    .Y(_09564_));
 sg13g2_a21o_1 _16281_ (.A2(_09557_),
    .A1(_09132_),
    .B1(_09564_),
    .X(_09565_));
 sg13g2_buf_1 _16282_ (.A(_09565_),
    .X(_09566_));
 sg13g2_and2_1 _16283_ (.A(_09560_),
    .B(_09557_),
    .X(_09567_));
 sg13g2_buf_1 _16284_ (.A(_09567_),
    .X(_09568_));
 sg13g2_and2_1 _16285_ (.A(_09132_),
    .B(_09564_),
    .X(_09569_));
 sg13g2_nand2b_1 _16286_ (.Y(_09570_),
    .B(_09569_),
    .A_N(_09568_));
 sg13g2_buf_1 _16287_ (.A(_09570_),
    .X(_09571_));
 sg13g2_nand2b_1 _16288_ (.Y(_09572_),
    .B(_09011_),
    .A_N(_08534_));
 sg13g2_a221oi_1 _16289_ (.B2(_09571_),
    .C1(_09572_),
    .B1(_09566_),
    .A1(_08536_),
    .Y(_09573_),
    .A2(_09017_));
 sg13g2_a21o_1 _16290_ (.A2(_08512_),
    .A1(net1015),
    .B1(_09573_),
    .X(_09574_));
 sg13g2_inv_1 _16291_ (.Y(_09575_),
    .A(_09574_));
 sg13g2_nand2_1 _16292_ (.Y(_09576_),
    .A(_09129_),
    .B(_09575_));
 sg13g2_buf_1 _16293_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09577_));
 sg13g2_buf_2 _16294_ (.A(\cpu.qspi.r_ind ),
    .X(_09578_));
 sg13g2_buf_1 _16295_ (.A(_00252_),
    .X(_09579_));
 sg13g2_buf_1 _16296_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09580_));
 sg13g2_buf_2 _16297_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09581_));
 sg13g2_buf_1 _16298_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09582_));
 sg13g2_nor3_1 _16299_ (.A(_09580_),
    .B(_09581_),
    .C(_09582_),
    .Y(_09583_));
 sg13g2_nor2b_1 _16300_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09583_),
    .Y(_09584_));
 sg13g2_buf_1 _16301_ (.A(_09584_),
    .X(_09585_));
 sg13g2_and2_1 _16302_ (.A(_09579_),
    .B(_09585_),
    .X(_09586_));
 sg13g2_buf_1 _16303_ (.A(_09586_),
    .X(_09587_));
 sg13g2_buf_1 _16304_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09588_));
 sg13g2_buf_1 _16305_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09589_));
 sg13g2_a221oi_1 _16306_ (.B2(_09588_),
    .C1(_09589_),
    .B1(_09587_),
    .A1(_09577_),
    .Y(_09590_),
    .A2(_09578_));
 sg13g2_a21oi_1 _16307_ (.A1(_09576_),
    .A2(_09590_),
    .Y(_00026_),
    .B1(net688));
 sg13g2_buf_1 _16308_ (.A(net877),
    .X(_09591_));
 sg13g2_buf_2 _16309_ (.A(net747),
    .X(_09592_));
 sg13g2_buf_1 _16310_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09593_));
 sg13g2_nand2_1 _16311_ (.Y(_09594_),
    .A(_09579_),
    .B(_09585_));
 sg13g2_buf_1 _16312_ (.A(_09594_),
    .X(_09595_));
 sg13g2_nor2_1 _16313_ (.A(_08515_),
    .B(_09566_),
    .Y(_09596_));
 sg13g2_buf_1 _16314_ (.A(_09596_),
    .X(_09597_));
 sg13g2_buf_2 _16315_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09598_));
 sg13g2_a22oi_1 _16316_ (.Y(_09599_),
    .B1(net128),
    .B2(_09598_),
    .A2(net584),
    .A1(_09593_));
 sg13g2_nor2_1 _16317_ (.A(net667),
    .B(_09599_),
    .Y(_00025_));
 sg13g2_buf_1 _16318_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09600_));
 sg13g2_buf_1 _16319_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09601_));
 sg13g2_a21oi_1 _16320_ (.A1(_09600_),
    .A2(_09587_),
    .Y(_09602_),
    .B1(_09601_));
 sg13g2_nor2_1 _16321_ (.A(net667),
    .B(_09602_),
    .Y(_00022_));
 sg13g2_buf_1 _16322_ (.A(_00277_),
    .X(_09603_));
 sg13g2_buf_1 _16323_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09604_));
 sg13g2_nand2_1 _16324_ (.Y(_09605_),
    .A(net1082),
    .B(net584));
 sg13g2_a21oi_1 _16325_ (.A1(_09603_),
    .A2(_09605_),
    .Y(_00023_),
    .B1(net688));
 sg13g2_buf_1 _16326_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09606_));
 sg13g2_buf_1 _16327_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09607_));
 sg13g2_inv_1 _16328_ (.Y(_09608_),
    .A(_09607_));
 sg13g2_inv_2 _16329_ (.Y(_09609_),
    .A(_08515_));
 sg13g2_nor2_1 _16330_ (.A(_09609_),
    .B(_08326_),
    .Y(_09610_));
 sg13g2_a21oi_1 _16331_ (.A1(_09609_),
    .A2(_09329_),
    .Y(_09611_),
    .B1(_09610_));
 sg13g2_or2_1 _16332_ (.X(_09612_),
    .B(_09611_),
    .A(_09607_));
 sg13g2_o21ai_1 _16333_ (.B1(_09612_),
    .Y(_09613_),
    .A1(_09608_),
    .A2(net128));
 sg13g2_and2_1 _16334_ (.A(_09606_),
    .B(_09613_),
    .X(_09614_));
 sg13g2_buf_2 _16335_ (.A(_09614_),
    .X(_09615_));
 sg13g2_nor3_1 _16336_ (.A(_09607_),
    .B(_09606_),
    .C(_09611_),
    .Y(_09616_));
 sg13g2_buf_2 _16337_ (.A(_09616_),
    .X(_09617_));
 sg13g2_nor2_1 _16338_ (.A(_09617_),
    .B(_09615_),
    .Y(_09618_));
 sg13g2_buf_2 _16339_ (.A(_09618_),
    .X(_09619_));
 sg13g2_and2_1 _16340_ (.A(\cpu.qspi.r_quad[2] ),
    .B(_09617_),
    .X(_09620_));
 sg13g2_a221oi_1 _16341_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09620_),
    .B1(_09619_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09621_),
    .A2(_09615_));
 sg13g2_buf_2 _16342_ (.A(_09621_),
    .X(_09622_));
 sg13g2_inv_1 _16343_ (.Y(_09623_),
    .A(_09622_));
 sg13g2_nand3_1 _16344_ (.B(net879),
    .C(_09574_),
    .A(_09129_),
    .Y(_09624_));
 sg13g2_nand3_1 _16345_ (.B(net759),
    .C(net584),
    .A(_09600_),
    .Y(_09625_));
 sg13g2_o21ai_1 _16346_ (.B1(_09625_),
    .Y(_00028_),
    .A1(_09623_),
    .A2(_09624_));
 sg13g2_nand2_1 _16347_ (.Y(_09626_),
    .A(_09588_),
    .B(net584));
 sg13g2_buf_2 _16348_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09627_));
 sg13g2_nand2_1 _16349_ (.Y(_09628_),
    .A(_09627_),
    .B(_09587_));
 sg13g2_a21oi_1 _16350_ (.A1(_09626_),
    .A2(_09628_),
    .Y(_00027_),
    .B1(_09104_));
 sg13g2_inv_1 _16351_ (.Y(_09629_),
    .A(_09578_));
 sg13g2_a21o_1 _16352_ (.A2(_09629_),
    .A1(_09577_),
    .B1(_09097_),
    .X(_00021_));
 sg13g2_buf_1 _16353_ (.A(net113),
    .X(_09630_));
 sg13g2_buf_1 _16354_ (.A(net155),
    .X(_09631_));
 sg13g2_inv_1 _16355_ (.Y(_09632_),
    .A(net251));
 sg13g2_nor2_1 _16356_ (.A(_08741_),
    .B(net213),
    .Y(_09633_));
 sg13g2_nand3_1 _16357_ (.B(net127),
    .C(_09633_),
    .A(_08664_),
    .Y(_09634_));
 sg13g2_buf_1 _16358_ (.A(\cpu.dec.r_op[10] ),
    .X(_09635_));
 sg13g2_buf_1 _16359_ (.A(_08622_),
    .X(_09636_));
 sg13g2_nand2_1 _16360_ (.Y(_09637_),
    .A(_09635_),
    .B(net109));
 sg13g2_o21ai_1 _16361_ (.B1(_09637_),
    .Y(_00011_),
    .A1(net90),
    .A2(_09634_));
 sg13g2_buf_1 _16362_ (.A(_08900_),
    .X(_09638_));
 sg13g2_inv_1 _16363_ (.Y(_09639_),
    .A(_08916_));
 sg13g2_nand3_1 _16364_ (.B(_08826_),
    .C(_08861_),
    .A(_08856_),
    .Y(_09640_));
 sg13g2_nand2b_1 _16365_ (.Y(_09641_),
    .B(_08881_),
    .A_N(_09640_));
 sg13g2_buf_1 _16366_ (.A(_09641_),
    .X(_09642_));
 sg13g2_nor4_1 _16367_ (.A(_08835_),
    .B(net246),
    .C(_09639_),
    .D(_09642_),
    .Y(_09643_));
 sg13g2_nand2_1 _16368_ (.Y(_09644_),
    .A(_08741_),
    .B(net213));
 sg13g2_buf_1 _16369_ (.A(_08835_),
    .X(_09645_));
 sg13g2_buf_1 _16370_ (.A(_08823_),
    .X(_09646_));
 sg13g2_inv_2 _16371_ (.Y(_09647_),
    .A(net250));
 sg13g2_nor2_1 _16372_ (.A(_09647_),
    .B(_08803_),
    .Y(_09648_));
 sg13g2_nand2_1 _16373_ (.Y(_09649_),
    .A(net245),
    .B(_09648_));
 sg13g2_nor3_1 _16374_ (.A(_09644_),
    .B(net126),
    .C(_09649_),
    .Y(_09650_));
 sg13g2_o21ai_1 _16375_ (.B1(net127),
    .Y(_09651_),
    .A1(_09643_),
    .A2(_09650_));
 sg13g2_buf_2 _16376_ (.A(\cpu.dec.r_op[1] ),
    .X(_09652_));
 sg13g2_nand2_1 _16377_ (.Y(_09653_),
    .A(_09652_),
    .B(net109));
 sg13g2_o21ai_1 _16378_ (.B1(_09653_),
    .Y(_00012_),
    .A1(net90),
    .A2(_09651_));
 sg13g2_buf_1 _16379_ (.A(\cpu.dec.r_op[9] ),
    .X(_09654_));
 sg13g2_buf_1 _16380_ (.A(_09654_),
    .X(_09655_));
 sg13g2_buf_1 _16381_ (.A(_08622_),
    .X(_09656_));
 sg13g2_buf_1 _16382_ (.A(_08740_),
    .X(_09657_));
 sg13g2_nor3_1 _16383_ (.A(_08720_),
    .B(net251),
    .C(_09649_),
    .Y(_09658_));
 sg13g2_a21oi_1 _16384_ (.A1(net251),
    .A2(_08836_),
    .Y(_09659_),
    .B1(_09658_));
 sg13g2_nor3_1 _16385_ (.A(net108),
    .B(net244),
    .C(_09659_),
    .Y(_09660_));
 sg13g2_a21o_1 _16386_ (.A2(net91),
    .A1(net1012),
    .B1(_09660_),
    .X(_00020_));
 sg13g2_buf_1 _16387_ (.A(\cpu.dec.r_op[8] ),
    .X(_09661_));
 sg13g2_inv_2 _16388_ (.Y(_09662_),
    .A(_09661_));
 sg13g2_inv_1 _16389_ (.Y(_09663_),
    .A(net252));
 sg13g2_nand2_2 _16390_ (.Y(_09664_),
    .A(net212),
    .B(net249));
 sg13g2_nand2_1 _16391_ (.Y(_09665_),
    .A(_08642_),
    .B(_08663_));
 sg13g2_buf_2 _16392_ (.A(_09665_),
    .X(_09666_));
 sg13g2_nor2_1 _16393_ (.A(_09664_),
    .B(_09666_),
    .Y(_09667_));
 sg13g2_nand2_1 _16394_ (.Y(_09668_),
    .A(net111),
    .B(_09667_));
 sg13g2_o21ai_1 _16395_ (.B1(_09668_),
    .Y(_00019_),
    .A1(_09662_),
    .A2(net112));
 sg13g2_buf_1 _16396_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09669_));
 sg13g2_inv_1 _16397_ (.Y(_09670_),
    .A(_09669_));
 sg13g2_nand2_1 _16398_ (.Y(_09671_),
    .A(_09627_),
    .B(_09595_));
 sg13g2_a21oi_1 _16399_ (.A1(_09670_),
    .A2(_09671_),
    .Y(_00024_),
    .B1(net688));
 sg13g2_buf_1 _16400_ (.A(\cpu.dec.r_op[2] ),
    .X(_09672_));
 sg13g2_buf_1 _16401_ (.A(net1079),
    .X(_09673_));
 sg13g2_a21oi_1 _16402_ (.A1(net248),
    .A2(_09648_),
    .Y(_09674_),
    .B1(net251));
 sg13g2_nor4_1 _16403_ (.A(net113),
    .B(_08720_),
    .C(net244),
    .D(_09674_),
    .Y(_09675_));
 sg13g2_a21o_1 _16404_ (.A2(net91),
    .A1(net1011),
    .B1(_09675_),
    .X(_00013_));
 sg13g2_buf_1 _16405_ (.A(\cpu.dec.r_op[7] ),
    .X(_09676_));
 sg13g2_buf_1 _16406_ (.A(net113),
    .X(_09677_));
 sg13g2_inv_2 _16407_ (.Y(_09678_),
    .A(_08900_));
 sg13g2_buf_1 _16408_ (.A(net247),
    .X(_09679_));
 sg13g2_buf_1 _16409_ (.A(_08916_),
    .X(_09680_));
 sg13g2_nor3_1 _16410_ (.A(_09678_),
    .B(net211),
    .C(net243),
    .Y(_09681_));
 sg13g2_a21oi_1 _16411_ (.A1(_08861_),
    .A2(_09681_),
    .Y(_09682_),
    .B1(_09648_));
 sg13g2_nor4_1 _16412_ (.A(net113),
    .B(net245),
    .C(_08837_),
    .D(_09682_),
    .Y(_09683_));
 sg13g2_a21o_1 _16413_ (.A2(net89),
    .A1(_09676_),
    .B1(_09683_),
    .X(_00018_));
 sg13g2_buf_1 _16414_ (.A(\cpu.uart.r_div[11] ),
    .X(_09684_));
 sg13g2_nor3_1 _16415_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09685_));
 sg13g2_nor2b_1 _16416_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09685_),
    .Y(_09686_));
 sg13g2_nor2b_1 _16417_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09686_),
    .Y(_09687_));
 sg13g2_nor2b_1 _16418_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09687_),
    .Y(_09688_));
 sg13g2_nor2b_1 _16419_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09688_),
    .Y(_09689_));
 sg13g2_nand2b_1 _16420_ (.Y(_09690_),
    .B(_09689_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16421_ (.A(\cpu.uart.r_div[8] ),
    .B(_09690_),
    .Y(_09691_));
 sg13g2_nand2b_1 _16422_ (.Y(_09692_),
    .B(_09691_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16423_ (.A(_09692_),
    .X(_09693_));
 sg13g2_nor3_1 _16424_ (.A(_09684_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09693_),
    .Y(_09694_));
 sg13g2_buf_1 _16425_ (.A(_09694_),
    .X(_09695_));
 sg13g2_nor2_1 _16426_ (.A(net1019),
    .B(net337),
    .Y(_09696_));
 sg13g2_buf_1 _16427_ (.A(_09696_),
    .X(_09697_));
 sg13g2_buf_1 _16428_ (.A(net242),
    .X(_09698_));
 sg13g2_mux2_1 _16429_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00279_),
    .S(net210),
    .X(_00079_));
 sg13g2_xnor2_1 _16430_ (.Y(_09699_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16431_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09699_),
    .S(net210),
    .X(_00082_));
 sg13g2_o21ai_1 _16432_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09700_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16433_ (.A(_09685_),
    .B_N(_09700_),
    .Y(_09701_));
 sg13g2_nor2_1 _16434_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net242),
    .Y(_09702_));
 sg13g2_a21oi_1 _16435_ (.A1(net210),
    .A2(_09701_),
    .Y(_00083_),
    .B1(_09702_));
 sg13g2_xnor2_1 _16436_ (.Y(_09703_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09685_));
 sg13g2_nor2_1 _16437_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net242),
    .Y(_09704_));
 sg13g2_a21oi_1 _16438_ (.A1(net210),
    .A2(_09703_),
    .Y(_00084_),
    .B1(_09704_));
 sg13g2_xnor2_1 _16439_ (.Y(_09705_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09686_));
 sg13g2_nor2_1 _16440_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net242),
    .Y(_09706_));
 sg13g2_a21oi_1 _16441_ (.A1(net210),
    .A2(_09705_),
    .Y(_00085_),
    .B1(_09706_));
 sg13g2_xnor2_1 _16442_ (.Y(_09707_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09687_));
 sg13g2_nor2_1 _16443_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net242),
    .Y(_09708_));
 sg13g2_a21oi_1 _16444_ (.A1(net210),
    .A2(_09707_),
    .Y(_00086_),
    .B1(_09708_));
 sg13g2_xnor2_1 _16445_ (.Y(_09709_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09688_));
 sg13g2_nor2_1 _16446_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net242),
    .Y(_09710_));
 sg13g2_a21oi_1 _16447_ (.A1(_09698_),
    .A2(_09709_),
    .Y(_00087_),
    .B1(_09710_));
 sg13g2_xnor2_1 _16448_ (.Y(_09711_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09689_));
 sg13g2_nor2_1 _16449_ (.A(\cpu.uart.r_div_value[7] ),
    .B(_09697_),
    .Y(_09712_));
 sg13g2_a21oi_1 _16450_ (.A1(_09698_),
    .A2(_09711_),
    .Y(_00088_),
    .B1(_09712_));
 sg13g2_xor2_1 _16451_ (.B(_09690_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09713_));
 sg13g2_nor2_1 _16452_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net242),
    .Y(_09714_));
 sg13g2_a21oi_1 _16453_ (.A1(net210),
    .A2(_09713_),
    .Y(_00089_),
    .B1(_09714_));
 sg13g2_xnor2_1 _16454_ (.Y(_09715_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09691_));
 sg13g2_nor2_1 _16455_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net242),
    .Y(_09716_));
 sg13g2_a21oi_1 _16456_ (.A1(net210),
    .A2(_09715_),
    .Y(_00090_),
    .B1(_09716_));
 sg13g2_buf_1 _16457_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09717_));
 sg13g2_inv_1 _16458_ (.Y(_09718_),
    .A(_09717_));
 sg13g2_nand2_1 _16459_ (.Y(_09719_),
    .A(net879),
    .B(_09693_));
 sg13g2_o21ai_1 _16460_ (.B1(_09719_),
    .Y(_09720_),
    .A1(_09684_),
    .A2(_09717_));
 sg13g2_inv_1 _16461_ (.Y(_09721_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16462_ (.A(_09721_),
    .B(_09096_),
    .C(_09693_),
    .Y(_09722_));
 sg13g2_a221oi_1 _16463_ (.B2(_09721_),
    .C1(_09722_),
    .B1(_09720_),
    .A1(_09718_),
    .Y(_00080_),
    .A2(net747));
 sg13g2_nor2_1 _16464_ (.A(\cpu.uart.r_div[10] ),
    .B(_09693_),
    .Y(_09723_));
 sg13g2_nand2_1 _16465_ (.Y(_09724_),
    .A(_09684_),
    .B(net761));
 sg13g2_o21ai_1 _16466_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09725_),
    .A1(_09096_),
    .A2(net337));
 sg13g2_o21ai_1 _16467_ (.B1(_09725_),
    .Y(_00081_),
    .A1(_09723_),
    .A2(_09724_));
 sg13g2_inv_1 _16468_ (.Y(_09726_),
    .A(_08962_));
 sg13g2_buf_1 _16469_ (.A(_09726_),
    .X(_09727_));
 sg13g2_buf_1 _16470_ (.A(net873),
    .X(_09728_));
 sg13g2_buf_1 _16471_ (.A(_09728_),
    .X(_09729_));
 sg13g2_nand2_1 _16472_ (.Y(_09730_),
    .A(net875),
    .B(_09157_));
 sg13g2_buf_1 _16473_ (.A(_09730_),
    .X(_09731_));
 sg13g2_buf_1 _16474_ (.A(\cpu.addr[5] ),
    .X(_09732_));
 sg13g2_buf_1 _16475_ (.A(_09732_),
    .X(_09733_));
 sg13g2_nor3_1 _16476_ (.A(_09733_),
    .B(net1085),
    .C(_08952_),
    .Y(_09734_));
 sg13g2_nand2_1 _16477_ (.Y(_09735_),
    .A(net1022),
    .B(_09734_));
 sg13g2_buf_1 _16478_ (.A(_09735_),
    .X(_09736_));
 sg13g2_buf_1 _16479_ (.A(_09736_),
    .X(_09737_));
 sg13g2_nor4_1 _16480_ (.A(net666),
    .B(_09022_),
    .C(_09731_),
    .D(net583),
    .Y(_09738_));
 sg13g2_buf_1 _16481_ (.A(_09738_),
    .X(_09739_));
 sg13g2_buf_1 _16482_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09740_));
 sg13g2_buf_1 _16483_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09741_));
 sg13g2_buf_1 _16484_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09742_));
 sg13g2_buf_1 _16485_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09743_));
 sg13g2_buf_1 _16486_ (.A(\cpu.intr.r_timer_count[11] ),
    .X(_09744_));
 sg13g2_buf_1 _16487_ (.A(\cpu.intr.r_timer_count[8] ),
    .X(_09745_));
 sg13g2_buf_2 _16488_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09746_));
 sg13g2_nor3_2 _16489_ (.A(_09746_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09747_));
 sg13g2_nor2b_1 _16490_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09747_),
    .Y(_09748_));
 sg13g2_nor2b_1 _16491_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09748_),
    .Y(_09749_));
 sg13g2_nor2b_1 _16492_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09749_),
    .Y(_09750_));
 sg13g2_nor2b_1 _16493_ (.A(\cpu.intr.r_timer_count[6] ),
    .B_N(_09750_),
    .Y(_09751_));
 sg13g2_nand2b_1 _16494_ (.Y(_09752_),
    .B(_09751_),
    .A_N(\cpu.intr.r_timer_count[7] ));
 sg13g2_nor3_2 _16495_ (.A(\cpu.intr.r_timer_count[9] ),
    .B(_09745_),
    .C(_09752_),
    .Y(_09753_));
 sg13g2_nand2b_1 _16496_ (.Y(_09754_),
    .B(_09753_),
    .A_N(\cpu.intr.r_timer_count[10] ));
 sg13g2_nor3_2 _16497_ (.A(_09744_),
    .B(\cpu.intr.r_timer_count[12] ),
    .C(_09754_),
    .Y(_09755_));
 sg13g2_nand2b_1 _16498_ (.Y(_09756_),
    .B(_09755_),
    .A_N(\cpu.intr.r_timer_count[13] ));
 sg13g2_nor2_1 _16499_ (.A(\cpu.intr.r_timer_count[14] ),
    .B(_09756_),
    .Y(_09757_));
 sg13g2_nand2b_1 _16500_ (.Y(_09758_),
    .B(_09757_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_nor3_1 _16501_ (.A(_09742_),
    .B(_09743_),
    .C(_09758_),
    .Y(_09759_));
 sg13g2_nor2b_1 _16502_ (.A(_09741_),
    .B_N(_09759_),
    .Y(_09760_));
 sg13g2_nand2b_1 _16503_ (.Y(_09761_),
    .B(_09760_),
    .A_N(_09740_));
 sg13g2_buf_2 _16504_ (.A(_09761_),
    .X(_09762_));
 sg13g2_buf_1 _16505_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09763_));
 sg13g2_buf_1 _16506_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09764_));
 sg13g2_buf_1 _16507_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09765_));
 sg13g2_buf_1 _16508_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09766_));
 sg13g2_nor4_2 _16509_ (.A(_09763_),
    .B(_09764_),
    .C(_09765_),
    .Y(_09767_),
    .D(_09766_));
 sg13g2_nand2b_1 _16510_ (.Y(_09768_),
    .B(_09767_),
    .A_N(_09762_));
 sg13g2_buf_2 _16511_ (.A(_09768_),
    .X(_09769_));
 sg13g2_nand2b_1 _16512_ (.Y(_09770_),
    .B(_09769_),
    .A_N(_09739_));
 sg13g2_buf_2 _16513_ (.A(_09770_),
    .X(_09771_));
 sg13g2_buf_8 _16514_ (.A(_09771_),
    .X(_09772_));
 sg13g2_mux2_1 _16515_ (.A0(_00285_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net70),
    .X(_00055_));
 sg13g2_buf_1 _16516_ (.A(_09771_),
    .X(_09773_));
 sg13g2_xor2_1 _16517_ (.B(\cpu.intr.r_timer_count[0] ),
    .A(_09746_),
    .X(_09774_));
 sg13g2_nand2_1 _16518_ (.Y(_09775_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net70));
 sg13g2_o21ai_1 _16519_ (.B1(_09775_),
    .Y(_00066_),
    .A1(net69),
    .A2(_09774_));
 sg13g2_o21ai_1 _16520_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_09776_),
    .A1(_09746_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16521_ (.A(_09747_),
    .B_N(_09776_),
    .Y(_09777_));
 sg13g2_nand2_1 _16522_ (.Y(_09778_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net70));
 sg13g2_o21ai_1 _16523_ (.B1(_09778_),
    .Y(_00071_),
    .A1(net69),
    .A2(_09777_));
 sg13g2_xnor2_1 _16524_ (.Y(_09779_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09747_));
 sg13g2_nand2_1 _16525_ (.Y(_09780_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(net70));
 sg13g2_o21ai_1 _16526_ (.B1(_09780_),
    .Y(_00072_),
    .A1(net69),
    .A2(_09779_));
 sg13g2_xnor2_1 _16527_ (.Y(_09781_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09748_));
 sg13g2_nand2_1 _16528_ (.Y(_09782_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_09772_));
 sg13g2_o21ai_1 _16529_ (.B1(_09782_),
    .Y(_00073_),
    .A1(_09773_),
    .A2(_09781_));
 sg13g2_xnor2_1 _16530_ (.Y(_09783_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09749_));
 sg13g2_buf_8 _16531_ (.A(_09771_),
    .X(_09784_));
 sg13g2_nand2_1 _16532_ (.Y(_09785_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(net68));
 sg13g2_o21ai_1 _16533_ (.B1(_09785_),
    .Y(_00074_),
    .A1(_09773_),
    .A2(_09783_));
 sg13g2_xnor2_1 _16534_ (.Y(_09786_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09750_));
 sg13g2_nand2_1 _16535_ (.Y(_09787_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(_09784_));
 sg13g2_o21ai_1 _16536_ (.B1(_09787_),
    .Y(_00075_),
    .A1(net69),
    .A2(_09786_));
 sg13g2_xnor2_1 _16537_ (.Y(_09788_),
    .A(\cpu.intr.r_timer_count[7] ),
    .B(_09751_));
 sg13g2_nand2_1 _16538_ (.Y(_09789_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_09784_));
 sg13g2_o21ai_1 _16539_ (.B1(_09789_),
    .Y(_00076_),
    .A1(net69),
    .A2(_09788_));
 sg13g2_xor2_1 _16540_ (.B(_09752_),
    .A(_09745_),
    .X(_09790_));
 sg13g2_nand2_1 _16541_ (.Y(_09791_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(net68));
 sg13g2_o21ai_1 _16542_ (.B1(_09791_),
    .Y(_00077_),
    .A1(net69),
    .A2(_09790_));
 sg13g2_o21ai_1 _16543_ (.B1(\cpu.intr.r_timer_count[9] ),
    .Y(_09792_),
    .A1(_09745_),
    .A2(_09752_));
 sg13g2_nor2b_1 _16544_ (.A(_09753_),
    .B_N(_09792_),
    .Y(_09793_));
 sg13g2_nand2_1 _16545_ (.Y(_09794_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net68));
 sg13g2_o21ai_1 _16546_ (.B1(_09794_),
    .Y(_00078_),
    .A1(net69),
    .A2(_09793_));
 sg13g2_xnor2_1 _16547_ (.Y(_09795_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(_09753_));
 sg13g2_nand2_1 _16548_ (.Y(_09796_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net68));
 sg13g2_o21ai_1 _16549_ (.B1(_09796_),
    .Y(_00056_),
    .A1(net69),
    .A2(_09795_));
 sg13g2_xor2_1 _16550_ (.B(_09754_),
    .A(_09744_),
    .X(_09797_));
 sg13g2_nand2_1 _16551_ (.Y(_09798_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net68));
 sg13g2_o21ai_1 _16552_ (.B1(_09798_),
    .Y(_00057_),
    .A1(net70),
    .A2(_09797_));
 sg13g2_o21ai_1 _16553_ (.B1(\cpu.intr.r_timer_count[12] ),
    .Y(_09799_),
    .A1(_09744_),
    .A2(_09754_));
 sg13g2_nor2b_1 _16554_ (.A(_09755_),
    .B_N(_09799_),
    .Y(_09800_));
 sg13g2_nand2_1 _16555_ (.Y(_09801_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net68));
 sg13g2_o21ai_1 _16556_ (.B1(_09801_),
    .Y(_00058_),
    .A1(net70),
    .A2(_09800_));
 sg13g2_xnor2_1 _16557_ (.Y(_09802_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_09755_));
 sg13g2_nand2_1 _16558_ (.Y(_09803_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net68));
 sg13g2_o21ai_1 _16559_ (.B1(_09803_),
    .Y(_00059_),
    .A1(net70),
    .A2(_09802_));
 sg13g2_xor2_1 _16560_ (.B(_09756_),
    .A(\cpu.intr.r_timer_count[14] ),
    .X(_09804_));
 sg13g2_nand2_1 _16561_ (.Y(_09805_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net68));
 sg13g2_o21ai_1 _16562_ (.B1(_09805_),
    .Y(_00060_),
    .A1(net70),
    .A2(_09804_));
 sg13g2_xnor2_1 _16563_ (.Y(_09806_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_09757_));
 sg13g2_nand2_1 _16564_ (.Y(_09807_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_09771_));
 sg13g2_o21ai_1 _16565_ (.B1(_09807_),
    .Y(_00061_),
    .A1(_09772_),
    .A2(_09806_));
 sg13g2_buf_1 _16566_ (.A(\cpu.dcache.wdata[0] ),
    .X(_09808_));
 sg13g2_inv_1 _16567_ (.Y(_09809_),
    .A(_09808_));
 sg13g2_buf_1 _16568_ (.A(_09809_),
    .X(_09810_));
 sg13g2_buf_1 _16569_ (.A(net872),
    .X(_09811_));
 sg13g2_buf_1 _16570_ (.A(_09739_),
    .X(_09812_));
 sg13g2_buf_1 _16571_ (.A(_09739_),
    .X(_09813_));
 sg13g2_nor4_1 _16572_ (.A(_09742_),
    .B(_09741_),
    .C(_09740_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_09814_));
 sg13g2_a21oi_1 _16573_ (.A1(_09767_),
    .A2(_09814_),
    .Y(_09815_),
    .B1(_09743_));
 sg13g2_mux2_1 _16574_ (.A0(_09815_),
    .A1(_09743_),
    .S(_09758_),
    .X(_09816_));
 sg13g2_nor2_1 _16575_ (.A(net153),
    .B(_09816_),
    .Y(_09817_));
 sg13g2_a21oi_1 _16576_ (.A1(net745),
    .A2(net154),
    .Y(_00062_),
    .B1(_09817_));
 sg13g2_buf_2 _16577_ (.A(\cpu.dcache.wdata[1] ),
    .X(_09818_));
 sg13g2_buf_1 _16578_ (.A(_09818_),
    .X(_09819_));
 sg13g2_buf_1 _16579_ (.A(net1009),
    .X(_09820_));
 sg13g2_nor2_1 _16580_ (.A(\cpu.intr.r_timer_reload[17] ),
    .B(_09769_),
    .Y(_09821_));
 sg13g2_o21ai_1 _16581_ (.B1(_09742_),
    .Y(_09822_),
    .A1(_09743_),
    .A2(_09758_));
 sg13g2_nor2b_1 _16582_ (.A(_09759_),
    .B_N(_09822_),
    .Y(_09823_));
 sg13g2_nor3_1 _16583_ (.A(_09739_),
    .B(_09821_),
    .C(_09823_),
    .Y(_09824_));
 sg13g2_a21o_1 _16584_ (.A2(net154),
    .A1(net871),
    .B1(_09824_),
    .X(_00063_));
 sg13g2_buf_1 _16585_ (.A(\cpu.dcache.wdata[2] ),
    .X(_09825_));
 sg13g2_buf_1 _16586_ (.A(_09825_),
    .X(_09826_));
 sg13g2_buf_1 _16587_ (.A(net1008),
    .X(_09827_));
 sg13g2_nor2_1 _16588_ (.A(\cpu.intr.r_timer_reload[18] ),
    .B(_09769_),
    .Y(_09828_));
 sg13g2_xnor2_1 _16589_ (.Y(_09829_),
    .A(_09741_),
    .B(_09759_));
 sg13g2_nor3_1 _16590_ (.A(_09739_),
    .B(_09828_),
    .C(_09829_),
    .Y(_09830_));
 sg13g2_a21o_1 _16591_ (.A2(net153),
    .A1(net870),
    .B1(_09830_),
    .X(_00064_));
 sg13g2_xor2_1 _16592_ (.B(_09760_),
    .A(_09740_),
    .X(_09831_));
 sg13g2_o21ai_1 _16593_ (.B1(_09831_),
    .Y(_09832_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09769_));
 sg13g2_buf_1 _16594_ (.A(\cpu.dcache.wdata[3] ),
    .X(_09833_));
 sg13g2_nand2_1 _16595_ (.Y(_09834_),
    .A(net1078),
    .B(net153));
 sg13g2_o21ai_1 _16596_ (.B1(_09834_),
    .Y(_00065_),
    .A1(net154),
    .A2(_09832_));
 sg13g2_inv_1 _16597_ (.Y(_09835_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_a21oi_1 _16598_ (.A1(_09835_),
    .A2(_09767_),
    .Y(_09836_),
    .B1(_09763_));
 sg13g2_nor2b_1 _16599_ (.A(_09762_),
    .B_N(_09836_),
    .Y(_09837_));
 sg13g2_a21oi_1 _16600_ (.A1(_09763_),
    .A2(_09762_),
    .Y(_09838_),
    .B1(_09837_));
 sg13g2_buf_2 _16601_ (.A(\cpu.dcache.wdata[4] ),
    .X(_09839_));
 sg13g2_buf_1 _16602_ (.A(_09839_),
    .X(_09840_));
 sg13g2_nand2_1 _16603_ (.Y(_09841_),
    .A(net1007),
    .B(net153));
 sg13g2_o21ai_1 _16604_ (.B1(_09841_),
    .Y(_00067_),
    .A1(_09812_),
    .A2(_09838_));
 sg13g2_nor2_1 _16605_ (.A(_09763_),
    .B(_09762_),
    .Y(_09842_));
 sg13g2_xor2_1 _16606_ (.B(_09842_),
    .A(_09764_),
    .X(_09843_));
 sg13g2_o21ai_1 _16607_ (.B1(_09843_),
    .Y(_09844_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09769_));
 sg13g2_buf_2 _16608_ (.A(\cpu.dcache.wdata[5] ),
    .X(_09845_));
 sg13g2_buf_1 _16609_ (.A(_09845_),
    .X(_09846_));
 sg13g2_nand2_1 _16610_ (.Y(_09847_),
    .A(net1006),
    .B(net153));
 sg13g2_o21ai_1 _16611_ (.B1(_09847_),
    .Y(_00068_),
    .A1(net154),
    .A2(_09844_));
 sg13g2_nor3_1 _16612_ (.A(_09763_),
    .B(_09764_),
    .C(_09762_),
    .Y(_09848_));
 sg13g2_xor2_1 _16613_ (.B(_09848_),
    .A(_09765_),
    .X(_09849_));
 sg13g2_o21ai_1 _16614_ (.B1(_09849_),
    .Y(_09850_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09769_));
 sg13g2_buf_2 _16615_ (.A(\cpu.dcache.wdata[6] ),
    .X(_09851_));
 sg13g2_nand2_1 _16616_ (.Y(_09852_),
    .A(_09851_),
    .B(_09739_));
 sg13g2_o21ai_1 _16617_ (.B1(_09852_),
    .Y(_00069_),
    .A1(net154),
    .A2(_09850_));
 sg13g2_nor2b_1 _16618_ (.A(_09766_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_09853_));
 sg13g2_nor2b_1 _16619_ (.A(_09765_),
    .B_N(_09848_),
    .Y(_09854_));
 sg13g2_mux2_1 _16620_ (.A0(_09766_),
    .A1(_09853_),
    .S(_09854_),
    .X(_09855_));
 sg13g2_buf_2 _16621_ (.A(\cpu.dcache.wdata[7] ),
    .X(_09856_));
 sg13g2_buf_1 _16622_ (.A(_09856_),
    .X(_09857_));
 sg13g2_mux2_1 _16623_ (.A0(_09855_),
    .A1(net1005),
    .S(_09813_),
    .X(_00070_));
 sg13g2_buf_1 _16624_ (.A(net589),
    .X(_09858_));
 sg13g2_buf_1 _16625_ (.A(net531),
    .X(_09859_));
 sg13g2_buf_1 _16626_ (.A(net465),
    .X(_09860_));
 sg13g2_nor2_1 _16627_ (.A(_09022_),
    .B(_09736_),
    .Y(_09861_));
 sg13g2_buf_1 _16628_ (.A(_09861_),
    .X(_09862_));
 sg13g2_nand2_1 _16629_ (.Y(_09863_),
    .A(net400),
    .B(_09862_));
 sg13g2_buf_1 _16630_ (.A(_09863_),
    .X(_09864_));
 sg13g2_buf_1 _16631_ (.A(net125),
    .X(_09865_));
 sg13g2_buf_1 _16632_ (.A(net880),
    .X(_09866_));
 sg13g2_buf_1 _16633_ (.A(net744),
    .X(_09867_));
 sg13g2_buf_1 _16634_ (.A(net665),
    .X(_09868_));
 sg13g2_buf_2 _16635_ (.A(net582),
    .X(_09869_));
 sg13g2_nor3_1 _16636_ (.A(net530),
    .B(net872),
    .C(net107),
    .Y(_09870_));
 sg13g2_a21o_1 _16637_ (.A2(net107),
    .A1(_00286_),
    .B1(_09870_),
    .X(_00036_));
 sg13g2_nand2_1 _16638_ (.Y(_09871_),
    .A(_09040_),
    .B(_09436_));
 sg13g2_nor3_1 _16639_ (.A(_09022_),
    .B(_09871_),
    .C(net583),
    .Y(_09872_));
 sg13g2_buf_2 _16640_ (.A(_09872_),
    .X(_09873_));
 sg13g2_buf_1 _16641_ (.A(_09873_),
    .X(_09874_));
 sg13g2_buf_1 _16642_ (.A(net152),
    .X(_09875_));
 sg13g2_buf_2 _16643_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_09876_));
 sg13g2_buf_2 _16644_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_09877_));
 sg13g2_xnor2_1 _16645_ (.Y(_09878_),
    .A(_09876_),
    .B(_09877_));
 sg13g2_buf_1 _16646_ (.A(net666),
    .X(_09879_));
 sg13g2_buf_2 _16647_ (.A(net581),
    .X(_09880_));
 sg13g2_buf_1 _16648_ (.A(net529),
    .X(_09881_));
 sg13g2_buf_1 _16649_ (.A(net464),
    .X(_09882_));
 sg13g2_buf_1 _16650_ (.A(_09818_),
    .X(_09883_));
 sg13g2_buf_1 _16651_ (.A(net152),
    .X(_09884_));
 sg13g2_nand3_1 _16652_ (.B(net1004),
    .C(net123),
    .A(net399),
    .Y(_09885_));
 sg13g2_o21ai_1 _16653_ (.B1(_09885_),
    .Y(_00043_),
    .A1(net124),
    .A2(_09878_));
 sg13g2_buf_2 _16654_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_09886_));
 sg13g2_nand2_1 _16655_ (.Y(_09887_),
    .A(_09876_),
    .B(_09877_));
 sg13g2_xor2_1 _16656_ (.B(_09887_),
    .A(_09886_),
    .X(_09888_));
 sg13g2_buf_1 _16657_ (.A(net1008),
    .X(_09889_));
 sg13g2_nand3_1 _16658_ (.B(net869),
    .C(net123),
    .A(net399),
    .Y(_09890_));
 sg13g2_o21ai_1 _16659_ (.B1(_09890_),
    .Y(_00044_),
    .A1(net124),
    .A2(_09888_));
 sg13g2_buf_1 _16660_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_09891_));
 sg13g2_nand2_1 _16661_ (.Y(_09892_),
    .A(_09877_),
    .B(_09886_));
 sg13g2_nor2_1 _16662_ (.A(_00286_),
    .B(_09892_),
    .Y(_09893_));
 sg13g2_xnor2_1 _16663_ (.Y(_09894_),
    .A(_09891_),
    .B(_09893_));
 sg13g2_nand3_1 _16664_ (.B(net1078),
    .C(net123),
    .A(net399),
    .Y(_09895_));
 sg13g2_o21ai_1 _16665_ (.B1(_09895_),
    .Y(_00045_),
    .A1(net124),
    .A2(_09894_));
 sg13g2_buf_2 _16666_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_09896_));
 sg13g2_and4_1 _16667_ (.A(_09876_),
    .B(_09877_),
    .C(_09886_),
    .D(_09891_),
    .X(_09897_));
 sg13g2_buf_1 _16668_ (.A(_09897_),
    .X(_09898_));
 sg13g2_xnor2_1 _16669_ (.Y(_09899_),
    .A(_09896_),
    .B(_09898_));
 sg13g2_nand3_1 _16670_ (.B(net1007),
    .C(_09884_),
    .A(net399),
    .Y(_09900_));
 sg13g2_o21ai_1 _16671_ (.B1(_09900_),
    .Y(_00046_),
    .A1(_09875_),
    .A2(_09899_));
 sg13g2_buf_2 _16672_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_09901_));
 sg13g2_nand3_1 _16673_ (.B(_09896_),
    .C(_09893_),
    .A(_09891_),
    .Y(_09902_));
 sg13g2_buf_1 _16674_ (.A(_09902_),
    .X(_09903_));
 sg13g2_xor2_1 _16675_ (.B(_09903_),
    .A(_09901_),
    .X(_09904_));
 sg13g2_nand3_1 _16676_ (.B(net1006),
    .C(_09884_),
    .A(_09882_),
    .Y(_09905_));
 sg13g2_o21ai_1 _16677_ (.B1(_09905_),
    .Y(_00047_),
    .A1(_09875_),
    .A2(_09904_));
 sg13g2_buf_2 _16678_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_09906_));
 sg13g2_nand3_1 _16679_ (.B(_09901_),
    .C(_09898_),
    .A(_09896_),
    .Y(_09907_));
 sg13g2_xor2_1 _16680_ (.B(_09907_),
    .A(_09906_),
    .X(_09908_));
 sg13g2_buf_1 _16681_ (.A(net152),
    .X(_09909_));
 sg13g2_nand3_1 _16682_ (.B(_09851_),
    .C(net122),
    .A(net399),
    .Y(_09910_));
 sg13g2_o21ai_1 _16683_ (.B1(_09910_),
    .Y(_00048_),
    .A1(net124),
    .A2(_09908_));
 sg13g2_buf_1 _16684_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_09911_));
 sg13g2_nand2_1 _16685_ (.Y(_09912_),
    .A(_09901_),
    .B(_09906_));
 sg13g2_nor2_1 _16686_ (.A(_09903_),
    .B(_09912_),
    .Y(_09913_));
 sg13g2_xnor2_1 _16687_ (.Y(_09914_),
    .A(_09911_),
    .B(_09913_));
 sg13g2_nand3_1 _16688_ (.B(_09856_),
    .C(_09909_),
    .A(net399),
    .Y(_09915_));
 sg13g2_o21ai_1 _16689_ (.B1(_09915_),
    .Y(_00049_),
    .A1(net124),
    .A2(_09914_));
 sg13g2_buf_2 _16690_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_09916_));
 sg13g2_nand2_1 _16691_ (.Y(_09917_),
    .A(_09896_),
    .B(_09898_));
 sg13g2_nand3_1 _16692_ (.B(_09906_),
    .C(_09911_),
    .A(_09901_),
    .Y(_09918_));
 sg13g2_nor2_1 _16693_ (.A(_09917_),
    .B(_09918_),
    .Y(_09919_));
 sg13g2_xnor2_1 _16694_ (.Y(_09920_),
    .A(_09916_),
    .B(_09919_));
 sg13g2_buf_1 _16695_ (.A(\cpu.dcache.wdata[8] ),
    .X(_09921_));
 sg13g2_nand3_1 _16696_ (.B(_09921_),
    .C(net122),
    .A(net399),
    .Y(_09922_));
 sg13g2_o21ai_1 _16697_ (.B1(_09922_),
    .Y(_00050_),
    .A1(net124),
    .A2(_09920_));
 sg13g2_buf_1 _16698_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_09923_));
 sg13g2_nand2_1 _16699_ (.Y(_09924_),
    .A(_09916_),
    .B(_09919_));
 sg13g2_xor2_1 _16700_ (.B(_09924_),
    .A(_09923_),
    .X(_09925_));
 sg13g2_buf_2 _16701_ (.A(\cpu.dcache.wdata[9] ),
    .X(_09926_));
 sg13g2_nand3_1 _16702_ (.B(_09926_),
    .C(net122),
    .A(net399),
    .Y(_09927_));
 sg13g2_o21ai_1 _16703_ (.B1(_09927_),
    .Y(_00051_),
    .A1(net124),
    .A2(_09925_));
 sg13g2_buf_1 _16704_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_09928_));
 sg13g2_nand3_1 _16705_ (.B(_09923_),
    .C(_09919_),
    .A(_09916_),
    .Y(_09929_));
 sg13g2_xor2_1 _16706_ (.B(_09929_),
    .A(_09928_),
    .X(_09930_));
 sg13g2_nand3_1 _16707_ (.B(\cpu.dcache.wdata[10] ),
    .C(net122),
    .A(net464),
    .Y(_09931_));
 sg13g2_o21ai_1 _16708_ (.B1(_09931_),
    .Y(_00037_),
    .A1(net124),
    .A2(_09930_));
 sg13g2_buf_1 _16709_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_09932_));
 sg13g2_nand3_1 _16710_ (.B(_09923_),
    .C(_09928_),
    .A(_09916_),
    .Y(_09933_));
 sg13g2_nor2_1 _16711_ (.A(_09918_),
    .B(_09933_),
    .Y(_09934_));
 sg13g2_nor2b_1 _16712_ (.A(_09903_),
    .B_N(_09934_),
    .Y(_09935_));
 sg13g2_xnor2_1 _16713_ (.Y(_09936_),
    .A(_09932_),
    .B(_09935_));
 sg13g2_buf_2 _16714_ (.A(\cpu.dcache.wdata[11] ),
    .X(_09937_));
 sg13g2_nand3_1 _16715_ (.B(_09937_),
    .C(net122),
    .A(net464),
    .Y(_09938_));
 sg13g2_o21ai_1 _16716_ (.B1(_09938_),
    .Y(_00038_),
    .A1(net123),
    .A2(_09936_));
 sg13g2_buf_1 _16717_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_09939_));
 sg13g2_nand4_1 _16718_ (.B(_09932_),
    .C(_09898_),
    .A(_09896_),
    .Y(_09940_),
    .D(_09934_));
 sg13g2_xor2_1 _16719_ (.B(_09940_),
    .A(_09939_),
    .X(_09941_));
 sg13g2_buf_2 _16720_ (.A(\cpu.dcache.wdata[12] ),
    .X(_09942_));
 sg13g2_nand3_1 _16721_ (.B(_09942_),
    .C(net122),
    .A(net464),
    .Y(_09943_));
 sg13g2_o21ai_1 _16722_ (.B1(_09943_),
    .Y(_00039_),
    .A1(net123),
    .A2(_09941_));
 sg13g2_buf_2 _16723_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_09944_));
 sg13g2_nand3_1 _16724_ (.B(_09939_),
    .C(_09934_),
    .A(_09932_),
    .Y(_09945_));
 sg13g2_buf_1 _16725_ (.A(_09945_),
    .X(_09946_));
 sg13g2_nor2_1 _16726_ (.A(_09903_),
    .B(_09946_),
    .Y(_09947_));
 sg13g2_xnor2_1 _16727_ (.Y(_09948_),
    .A(_09944_),
    .B(_09947_));
 sg13g2_nand3_1 _16728_ (.B(\cpu.dcache.wdata[13] ),
    .C(net122),
    .A(net464),
    .Y(_09949_));
 sg13g2_o21ai_1 _16729_ (.B1(_09949_),
    .Y(_00040_),
    .A1(net123),
    .A2(_09948_));
 sg13g2_buf_2 _16730_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_09950_));
 sg13g2_nor2_1 _16731_ (.A(_09917_),
    .B(_09946_),
    .Y(_09951_));
 sg13g2_nand2_1 _16732_ (.Y(_09952_),
    .A(_09944_),
    .B(_09951_));
 sg13g2_xor2_1 _16733_ (.B(_09952_),
    .A(_09950_),
    .X(_09953_));
 sg13g2_nand3_1 _16734_ (.B(\cpu.dcache.wdata[14] ),
    .C(_09909_),
    .A(net464),
    .Y(_09954_));
 sg13g2_o21ai_1 _16735_ (.B1(_09954_),
    .Y(_00041_),
    .A1(net123),
    .A2(_09953_));
 sg13g2_buf_2 _16736_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_09955_));
 sg13g2_nand3_1 _16737_ (.B(_09950_),
    .C(_09947_),
    .A(_09944_),
    .Y(_09956_));
 sg13g2_xor2_1 _16738_ (.B(_09956_),
    .A(_09955_),
    .X(_09957_));
 sg13g2_buf_2 _16739_ (.A(\cpu.dcache.wdata[15] ),
    .X(_09958_));
 sg13g2_nand3_1 _16740_ (.B(_09958_),
    .C(net122),
    .A(net464),
    .Y(_09959_));
 sg13g2_o21ai_1 _16741_ (.B1(_09959_),
    .Y(_00042_),
    .A1(net123),
    .A2(_09957_));
 sg13g2_buf_2 _16742_ (.A(\cpu.ex.r_wb_valid ),
    .X(_09960_));
 sg13g2_inv_1 _16743_ (.Y(_09961_),
    .A(_09960_));
 sg13g2_buf_1 _16744_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_09962_));
 sg13g2_buf_2 _16745_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_09963_));
 sg13g2_buf_8 _16746_ (.A(_09963_),
    .X(_09964_));
 sg13g2_nand2_1 _16747_ (.Y(_09965_),
    .A(net1077),
    .B(net1003));
 sg13g2_buf_1 _16748_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_09966_));
 sg13g2_buf_2 _16749_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_09967_));
 sg13g2_inv_1 _16750_ (.Y(_09968_),
    .A(_09967_));
 sg13g2_nor2_1 _16751_ (.A(net1076),
    .B(_09968_),
    .Y(_09969_));
 sg13g2_inv_1 _16752_ (.Y(_09970_),
    .A(_09969_));
 sg13g2_nor3_1 _16753_ (.A(_09961_),
    .B(_09965_),
    .C(_09970_),
    .Y(_09971_));
 sg13g2_nand2_2 _16754_ (.Y(_09972_),
    .A(_09960_),
    .B(\cpu.ex.r_set_cc ));
 sg13g2_nor2b_1 _16755_ (.A(_09971_),
    .B_N(_09972_),
    .Y(_09973_));
 sg13g2_buf_2 _16756_ (.A(_09973_),
    .X(_09974_));
 sg13g2_buf_1 _16757_ (.A(_09974_),
    .X(_09975_));
 sg13g2_buf_1 _16758_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_09976_));
 sg13g2_buf_1 _16759_ (.A(_09976_),
    .X(_09977_));
 sg13g2_buf_1 _16760_ (.A(net1002),
    .X(_09978_));
 sg13g2_buf_2 _16761_ (.A(\cpu.dec.r_rs2_inv ),
    .X(_09979_));
 sg13g2_nor2_1 _16762_ (.A(_09976_),
    .B(_09979_),
    .Y(_09980_));
 sg13g2_buf_1 _16763_ (.A(_09980_),
    .X(_09981_));
 sg13g2_buf_1 _16764_ (.A(\cpu.dec.needs_rs2 ),
    .X(_09982_));
 sg13g2_buf_1 _16765_ (.A(_09982_),
    .X(_09983_));
 sg13g2_buf_1 _16766_ (.A(net1001),
    .X(_09984_));
 sg13g2_buf_2 _16767_ (.A(\cpu.addr[9] ),
    .X(_09985_));
 sg13g2_nor2_1 _16768_ (.A(net1077),
    .B(net1003),
    .Y(_09986_));
 sg13g2_nor2_1 _16769_ (.A(net1076),
    .B(_09967_),
    .Y(_09987_));
 sg13g2_a21oi_2 _16770_ (.B1(_09961_),
    .Y(_09988_),
    .A2(_09987_),
    .A1(_09986_));
 sg13g2_buf_2 _16771_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_09989_));
 sg13g2_xor2_1 _16772_ (.B(_09989_),
    .A(_09967_),
    .X(_09990_));
 sg13g2_buf_2 _16773_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_09991_));
 sg13g2_xor2_1 _16774_ (.B(_09991_),
    .A(_09964_),
    .X(_09992_));
 sg13g2_buf_2 _16775_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_09993_));
 sg13g2_xor2_1 _16776_ (.B(_09993_),
    .A(_09966_),
    .X(_09994_));
 sg13g2_buf_2 _16777_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_09995_));
 sg13g2_buf_8 _16778_ (.A(_09995_),
    .X(_09996_));
 sg13g2_xor2_1 _16779_ (.B(_09996_),
    .A(_09962_),
    .X(_09997_));
 sg13g2_nor4_2 _16780_ (.A(_09990_),
    .B(_09992_),
    .C(_09994_),
    .Y(_09998_),
    .D(_09997_));
 sg13g2_and2_1 _16781_ (.A(_09988_),
    .B(_09998_),
    .X(_09999_));
 sg13g2_buf_1 _16782_ (.A(_09999_),
    .X(_10000_));
 sg13g2_buf_1 _16783_ (.A(net580),
    .X(_10001_));
 sg13g2_nor2_1 _16784_ (.A(_09993_),
    .B(_09989_),
    .Y(_10002_));
 sg13g2_buf_1 _16785_ (.A(_10002_),
    .X(_10003_));
 sg13g2_nor2_1 _16786_ (.A(_09991_),
    .B(_09995_),
    .Y(_10004_));
 sg13g2_buf_1 _16787_ (.A(_10004_),
    .X(_10005_));
 sg13g2_and2_1 _16788_ (.A(net866),
    .B(_10005_),
    .X(_10006_));
 sg13g2_a21oi_1 _16789_ (.A1(_09988_),
    .A2(_09998_),
    .Y(_10007_),
    .B1(_10006_));
 sg13g2_buf_2 _16790_ (.A(_10007_),
    .X(_10008_));
 sg13g2_buf_1 _16791_ (.A(_10008_),
    .X(_10009_));
 sg13g2_buf_8 _16792_ (.A(net1000),
    .X(_10010_));
 sg13g2_inv_2 _16793_ (.Y(_10011_),
    .A(_10010_));
 sg13g2_buf_1 _16794_ (.A(_10011_),
    .X(_10012_));
 sg13g2_buf_1 _16795_ (.A(_09989_),
    .X(_10013_));
 sg13g2_buf_8 _16796_ (.A(_09993_),
    .X(_10014_));
 sg13g2_nor2b_1 _16797_ (.A(net999),
    .B_N(net998),
    .Y(_10015_));
 sg13g2_buf_1 _16798_ (.A(_10015_),
    .X(_10016_));
 sg13g2_nand3_1 _16799_ (.B(net664),
    .C(net743),
    .A(\cpu.ex.r_9[9] ),
    .Y(_10017_));
 sg13g2_nor2b_1 _16800_ (.A(_10014_),
    .B_N(_09996_),
    .Y(_10018_));
 sg13g2_buf_2 _16801_ (.A(_10018_),
    .X(_10019_));
 sg13g2_buf_1 _16802_ (.A(_10019_),
    .X(_10020_));
 sg13g2_buf_1 _16803_ (.A(_09989_),
    .X(_10021_));
 sg13g2_buf_8 _16804_ (.A(net997),
    .X(_10022_));
 sg13g2_mux2_1 _16805_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(\cpu.ex.r_mult[25] ),
    .S(net864),
    .X(_10023_));
 sg13g2_nand2_1 _16806_ (.Y(_10024_),
    .A(net663),
    .B(_10023_));
 sg13g2_buf_8 _16807_ (.A(_09991_),
    .X(_10025_));
 sg13g2_inv_1 _16808_ (.Y(_10026_),
    .A(net996));
 sg13g2_buf_1 _16809_ (.A(_10026_),
    .X(_10027_));
 sg13g2_buf_1 _16810_ (.A(_10027_),
    .X(_10028_));
 sg13g2_a21o_1 _16811_ (.A2(_10024_),
    .A1(_10017_),
    .B1(net662),
    .X(_10029_));
 sg13g2_buf_1 _16812_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10030_));
 sg13g2_nor2_1 _16813_ (.A(net996),
    .B(net999),
    .Y(_10031_));
 sg13g2_buf_2 _16814_ (.A(_10031_),
    .X(_10032_));
 sg13g2_and2_1 _16815_ (.A(net663),
    .B(_10032_),
    .X(_10033_));
 sg13g2_buf_8 _16816_ (.A(net1000),
    .X(_10034_));
 sg13g2_buf_8 _16817_ (.A(net863),
    .X(_10035_));
 sg13g2_mux2_1 _16818_ (.A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_10[9] ),
    .S(net741),
    .X(_10036_));
 sg13g2_buf_8 _16819_ (.A(net996),
    .X(_10037_));
 sg13g2_buf_1 _16820_ (.A(net862),
    .X(_10038_));
 sg13g2_and3_1 _16821_ (.X(_10039_),
    .A(\cpu.ex.r_11[9] ),
    .B(net740),
    .C(net741));
 sg13g2_a21o_1 _16822_ (.A2(_10036_),
    .A1(net662),
    .B1(_10039_),
    .X(_10040_));
 sg13g2_a22oi_1 _16823_ (.Y(_10041_),
    .B1(_10040_),
    .B2(net743),
    .A2(_10033_),
    .A1(_10030_));
 sg13g2_and2_1 _16824_ (.A(_09993_),
    .B(_09989_),
    .X(_10042_));
 sg13g2_buf_1 _16825_ (.A(_10042_),
    .X(_10043_));
 sg13g2_buf_1 _16826_ (.A(_10043_),
    .X(_10044_));
 sg13g2_inv_1 _16827_ (.Y(_10045_),
    .A(_00267_));
 sg13g2_mux4_1 _16828_ (.S0(net742),
    .A0(_10045_),
    .A1(\cpu.ex.r_14[9] ),
    .A2(\cpu.ex.r_13[9] ),
    .A3(\cpu.ex.r_12[9] ),
    .S1(net664),
    .X(_10046_));
 sg13g2_nand2_1 _16829_ (.Y(_10047_),
    .A(net739),
    .B(_10046_));
 sg13g2_inv_1 _16830_ (.Y(_10048_),
    .A(\cpu.ex.r_stmp[9] ));
 sg13g2_buf_8 _16831_ (.A(net740),
    .X(_10049_));
 sg13g2_nand2_2 _16832_ (.Y(_10050_),
    .A(net741),
    .B(net864));
 sg13g2_nor3_1 _16833_ (.A(_10048_),
    .B(net661),
    .C(_10050_),
    .Y(_10051_));
 sg13g2_inv_1 _16834_ (.Y(_10052_),
    .A(net997));
 sg13g2_buf_1 _16835_ (.A(_10052_),
    .X(_10053_));
 sg13g2_nor2b_1 _16836_ (.A(_09995_),
    .B_N(_09991_),
    .Y(_10054_));
 sg13g2_buf_1 _16837_ (.A(_10054_),
    .X(_10055_));
 sg13g2_and3_1 _16838_ (.X(_10056_),
    .A(\cpu.ex.r_lr[9] ),
    .B(net738),
    .C(net861));
 sg13g2_inv_1 _16839_ (.Y(_10057_),
    .A(_09993_));
 sg13g2_buf_1 _16840_ (.A(_10057_),
    .X(_10058_));
 sg13g2_o21ai_1 _16841_ (.B1(net860),
    .Y(_10059_),
    .A1(_10051_),
    .A2(_10056_));
 sg13g2_nand4_1 _16842_ (.B(_10041_),
    .C(_10047_),
    .A(_10029_),
    .Y(_10060_),
    .D(_10059_));
 sg13g2_a22oi_1 _16843_ (.Y(_10061_),
    .B1(net527),
    .B2(_10060_),
    .A2(net528),
    .A1(_09985_));
 sg13g2_nor2_1 _16844_ (.A(net1001),
    .B(\cpu.dec.imm[9] ),
    .Y(_10062_));
 sg13g2_a21o_1 _16845_ (.A2(_10061_),
    .A1(_09984_),
    .B1(_10062_),
    .X(_10063_));
 sg13g2_a22oi_1 _16846_ (.Y(_10064_),
    .B1(_09981_),
    .B2(_10063_),
    .A2(_09978_),
    .A1(_08461_));
 sg13g2_buf_1 _16847_ (.A(_10064_),
    .X(_10065_));
 sg13g2_nor2b_1 _16848_ (.A(\cpu.ex.pc[8] ),
    .B_N(net868),
    .Y(_10066_));
 sg13g2_buf_2 _16849_ (.A(_10066_),
    .X(_10067_));
 sg13g2_nand2_1 _16850_ (.Y(_10068_),
    .A(net1085),
    .B(net580));
 sg13g2_nor2b_1 _16851_ (.A(net996),
    .B_N(net999),
    .Y(_10069_));
 sg13g2_buf_1 _16852_ (.A(_10069_),
    .X(_10070_));
 sg13g2_nor2b_1 _16853_ (.A(net999),
    .B_N(net996),
    .Y(_10071_));
 sg13g2_buf_2 _16854_ (.A(_10071_),
    .X(_10072_));
 sg13g2_a22oi_1 _16855_ (.Y(_10073_),
    .B1(_10072_),
    .B2(\cpu.ex.r_9[8] ),
    .A2(net737),
    .A1(\cpu.ex.r_12[8] ));
 sg13g2_and2_1 _16856_ (.A(net996),
    .B(net999),
    .X(_10074_));
 sg13g2_buf_2 _16857_ (.A(_10074_),
    .X(_10075_));
 sg13g2_a22oi_1 _16858_ (.Y(_10076_),
    .B1(_10032_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(_10075_),
    .A1(\cpu.ex.r_13[8] ));
 sg13g2_buf_8 _16859_ (.A(net998),
    .X(_10077_));
 sg13g2_nand2b_1 _16860_ (.Y(_10078_),
    .B(net859),
    .A_N(net863));
 sg13g2_a21oi_1 _16861_ (.A1(_10073_),
    .A2(_10076_),
    .Y(_10079_),
    .B1(_10078_));
 sg13g2_and2_1 _16862_ (.A(_10003_),
    .B(_10055_),
    .X(_10080_));
 sg13g2_nor2b_1 _16863_ (.A(net996),
    .B_N(net1000),
    .Y(_10081_));
 sg13g2_buf_1 _16864_ (.A(_10081_),
    .X(_10082_));
 sg13g2_buf_1 _16865_ (.A(_10082_),
    .X(_10083_));
 sg13g2_and2_1 _16866_ (.A(net660),
    .B(net739),
    .X(_10084_));
 sg13g2_buf_1 _16867_ (.A(_10084_),
    .X(_10085_));
 sg13g2_a22oi_1 _16868_ (.Y(_10086_),
    .B1(_10085_),
    .B2(\cpu.ex.r_14[8] ),
    .A2(_10080_),
    .A1(\cpu.ex.r_lr[8] ));
 sg13g2_nand2b_1 _16869_ (.Y(_10087_),
    .B(_10086_),
    .A_N(_10079_));
 sg13g2_inv_1 _16870_ (.Y(_10088_),
    .A(_00266_));
 sg13g2_mux2_1 _16871_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(\cpu.ex.r_mult[24] ),
    .S(net864),
    .X(_10089_));
 sg13g2_a22oi_1 _16872_ (.Y(_10090_),
    .B1(_10089_),
    .B2(net860),
    .A2(net739),
    .A1(_10088_));
 sg13g2_buf_1 _16873_ (.A(net661),
    .X(_10091_));
 sg13g2_nand2b_1 _16874_ (.Y(_10092_),
    .B(_10091_),
    .A_N(_10090_));
 sg13g2_nor2b_1 _16875_ (.A(net998),
    .B_N(net999),
    .Y(_10093_));
 sg13g2_buf_1 _16876_ (.A(_10093_),
    .X(_10094_));
 sg13g2_nor2b_1 _16877_ (.A(net661),
    .B_N(\cpu.ex.r_stmp[8] ),
    .Y(_10095_));
 sg13g2_buf_1 _16878_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10096_));
 sg13g2_buf_8 _16879_ (.A(net859),
    .X(_10097_));
 sg13g2_mux2_1 _16880_ (.A0(_10096_),
    .A1(\cpu.ex.r_10[8] ),
    .S(net736),
    .X(_10098_));
 sg13g2_and3_1 _16881_ (.X(_10099_),
    .A(\cpu.ex.r_11[8] ),
    .B(net740),
    .C(net743));
 sg13g2_a221oi_1 _16882_ (.B2(_10032_),
    .C1(_10099_),
    .B1(_10098_),
    .A1(_10094_),
    .Y(_10100_),
    .A2(_10095_));
 sg13g2_a21oi_1 _16883_ (.A1(_10092_),
    .A2(_10100_),
    .Y(_10101_),
    .B1(net664));
 sg13g2_o21ai_1 _16884_ (.B1(net527),
    .Y(_10102_),
    .A1(_10087_),
    .A2(_10101_));
 sg13g2_nand3_1 _16885_ (.B(_10068_),
    .C(_10102_),
    .A(net1001),
    .Y(_10103_));
 sg13g2_or2_1 _16886_ (.X(_10104_),
    .B(\cpu.dec.imm[8] ),
    .A(net1001));
 sg13g2_or2_1 _16887_ (.X(_10105_),
    .B(_09979_),
    .A(_09976_));
 sg13g2_buf_1 _16888_ (.A(_10105_),
    .X(_10106_));
 sg13g2_a21oi_1 _16889_ (.A1(_10103_),
    .A2(_10104_),
    .Y(_10107_),
    .B1(_10106_));
 sg13g2_buf_2 _16890_ (.A(_10107_),
    .X(_10108_));
 sg13g2_buf_2 _16891_ (.A(_00303_),
    .X(_10109_));
 sg13g2_inv_1 _16892_ (.Y(_10110_),
    .A(_10109_));
 sg13g2_o21ai_1 _16893_ (.B1(_10110_),
    .Y(_10111_),
    .A1(_10067_),
    .A2(_10108_));
 sg13g2_buf_2 _16894_ (.A(_00302_),
    .X(_10112_));
 sg13g2_a21o_1 _16895_ (.A2(_10111_),
    .A1(net296),
    .B1(_10112_),
    .X(_10113_));
 sg13g2_inv_1 _16896_ (.Y(_10114_),
    .A(net296));
 sg13g2_or2_1 _16897_ (.X(_10115_),
    .B(_10108_),
    .A(_10067_));
 sg13g2_buf_1 _16898_ (.A(_10115_),
    .X(_10116_));
 sg13g2_nand3_1 _16899_ (.B(_10114_),
    .C(net182),
    .A(_10110_),
    .Y(_10117_));
 sg13g2_a21oi_1 _16900_ (.A1(_10113_),
    .A2(_10117_),
    .Y(_10118_),
    .B1(net537));
 sg13g2_buf_2 _16901_ (.A(_10118_),
    .X(_10119_));
 sg13g2_buf_1 _16902_ (.A(_09981_),
    .X(_10120_));
 sg13g2_inv_1 _16903_ (.Y(_10121_),
    .A(_09982_));
 sg13g2_buf_1 _16904_ (.A(_10121_),
    .X(_10122_));
 sg13g2_a21o_1 _16905_ (.A2(_09998_),
    .A1(_09988_),
    .B1(_10006_),
    .X(_10123_));
 sg13g2_buf_1 _16906_ (.A(_10123_),
    .X(_10124_));
 sg13g2_buf_1 _16907_ (.A(net864),
    .X(_10125_));
 sg13g2_buf_1 _16908_ (.A(net734),
    .X(_10126_));
 sg13g2_nand3_1 _16909_ (.B(net579),
    .C(net663),
    .A(\cpu.ex.r_mult[27] ),
    .Y(_10127_));
 sg13g2_nor2b_1 _16910_ (.A(net1000),
    .B_N(_09993_),
    .Y(_10128_));
 sg13g2_buf_1 _16911_ (.A(_10128_),
    .X(_10129_));
 sg13g2_buf_1 _16912_ (.A(_10129_),
    .X(_10130_));
 sg13g2_nand3_1 _16913_ (.B(net662),
    .C(net658),
    .A(\cpu.ex.r_12[11] ),
    .Y(_10131_));
 sg13g2_nand3_1 _16914_ (.B(net662),
    .C(net663),
    .A(\cpu.ex.r_stmp[11] ),
    .Y(_10132_));
 sg13g2_nand3_1 _16915_ (.B(net579),
    .C(net658),
    .A(\cpu.ex.r_13[11] ),
    .Y(_10133_));
 sg13g2_nand4_1 _16916_ (.B(_10131_),
    .C(_10132_),
    .A(_10127_),
    .Y(_10134_),
    .D(_10133_));
 sg13g2_buf_1 _16917_ (.A(_10035_),
    .X(_10135_));
 sg13g2_buf_1 _16918_ (.A(net736),
    .X(_10136_));
 sg13g2_nand3_1 _16919_ (.B(_10136_),
    .C(net734),
    .A(net657),
    .Y(_10137_));
 sg13g2_nand3_1 _16920_ (.B(net664),
    .C(net866),
    .A(\cpu.ex.r_lr[11] ),
    .Y(_10138_));
 sg13g2_o21ai_1 _16921_ (.B1(_10138_),
    .Y(_10139_),
    .A1(_00269_),
    .A2(_10137_));
 sg13g2_nand3_1 _16922_ (.B(net660),
    .C(net739),
    .A(\cpu.ex.r_14[11] ),
    .Y(_10140_));
 sg13g2_mux2_1 _16923_ (.A0(\cpu.ex.r_sp[11] ),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net661),
    .X(_10141_));
 sg13g2_nand3_1 _16924_ (.B(net663),
    .C(_10141_),
    .A(_10053_),
    .Y(_10142_));
 sg13g2_mux4_1 _16925_ (.S0(net661),
    .A0(\cpu.ex.r_8[11] ),
    .A1(\cpu.ex.r_9[11] ),
    .A2(\cpu.ex.r_10[11] ),
    .A3(\cpu.ex.r_11[11] ),
    .S1(net657),
    .X(_10143_));
 sg13g2_nand2_1 _16926_ (.Y(_10144_),
    .A(net743),
    .B(_10143_));
 sg13g2_nand3_1 _16927_ (.B(_10142_),
    .C(_10144_),
    .A(_10140_),
    .Y(_10145_));
 sg13g2_a221oi_1 _16928_ (.B2(net579),
    .C1(_10145_),
    .B1(_10139_),
    .A1(net659),
    .Y(_10146_),
    .A2(_10134_));
 sg13g2_buf_2 _16929_ (.A(\cpu.addr[11] ),
    .X(_10147_));
 sg13g2_nand2_1 _16930_ (.Y(_10148_),
    .A(_10147_),
    .B(net528));
 sg13g2_o21ai_1 _16931_ (.B1(_10148_),
    .Y(_10149_),
    .A1(_10124_),
    .A2(_10146_));
 sg13g2_or2_1 _16932_ (.X(_10150_),
    .B(\cpu.dec.imm[11] ),
    .A(net867));
 sg13g2_o21ai_1 _16933_ (.B1(_10150_),
    .Y(_10151_),
    .A1(net858),
    .A2(_10149_));
 sg13g2_a22oi_1 _16934_ (.Y(_10152_),
    .B1(net735),
    .B2(_10151_),
    .A2(net868),
    .A1(_08445_));
 sg13g2_buf_2 _16935_ (.A(_10152_),
    .X(_10153_));
 sg13g2_buf_1 _16936_ (.A(_10153_),
    .X(_10154_));
 sg13g2_nand2b_1 _16937_ (.Y(_10155_),
    .B(net868),
    .A_N(_08490_));
 sg13g2_buf_1 _16938_ (.A(\cpu.addr[10] ),
    .X(_10156_));
 sg13g2_nor2b_1 _16939_ (.A(net657),
    .B_N(\cpu.ex.r_9[10] ),
    .Y(_10157_));
 sg13g2_buf_1 _16940_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10158_));
 sg13g2_and2_1 _16941_ (.A(_10158_),
    .B(net657),
    .X(_10159_));
 sg13g2_a22oi_1 _16942_ (.Y(_10160_),
    .B1(_10159_),
    .B2(_10094_),
    .A2(_10157_),
    .A1(net743));
 sg13g2_buf_1 _16943_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10161_));
 sg13g2_and2_1 _16944_ (.A(_10161_),
    .B(_10135_),
    .X(_10162_));
 sg13g2_nor2b_1 _16945_ (.A(_10135_),
    .B_N(\cpu.ex.r_12[10] ),
    .Y(_10163_));
 sg13g2_a221oi_1 _16946_ (.B2(_10044_),
    .C1(net579),
    .B1(_10163_),
    .A1(net866),
    .Y(_10164_),
    .A2(_10162_));
 sg13g2_a21o_1 _16947_ (.A2(_10160_),
    .A1(net579),
    .B1(_10164_),
    .X(_10165_));
 sg13g2_a22oi_1 _16948_ (.Y(_10166_),
    .B1(_10032_),
    .B2(\cpu.ex.r_8[10] ),
    .A2(_10075_),
    .A1(\cpu.ex.r_13[10] ));
 sg13g2_nand2b_1 _16949_ (.Y(_10167_),
    .B(_10130_),
    .A_N(_10166_));
 sg13g2_a22oi_1 _16950_ (.Y(_10168_),
    .B1(_10072_),
    .B2(\cpu.ex.r_epc[10] ),
    .A2(net737),
    .A1(\cpu.ex.r_stmp[10] ));
 sg13g2_nand2b_1 _16951_ (.Y(_10169_),
    .B(_10020_),
    .A_N(_10168_));
 sg13g2_mux2_1 _16952_ (.A0(\cpu.ex.r_10[10] ),
    .A1(\cpu.ex.r_11[10] ),
    .S(net661),
    .X(_10170_));
 sg13g2_nand2b_1 _16953_ (.Y(_10171_),
    .B(_10014_),
    .A_N(_09989_));
 sg13g2_buf_1 _16954_ (.A(_10171_),
    .X(_10172_));
 sg13g2_nor2_1 _16955_ (.A(_10012_),
    .B(_10172_),
    .Y(_10173_));
 sg13g2_nand2b_1 _16956_ (.Y(_10174_),
    .B(_10049_),
    .A_N(_00268_));
 sg13g2_nand2b_1 _16957_ (.Y(_10175_),
    .B(\cpu.ex.r_14[10] ),
    .A_N(_10049_));
 sg13g2_a21oi_1 _16958_ (.A1(_10174_),
    .A2(_10175_),
    .Y(_10176_),
    .B1(_10137_));
 sg13g2_a221oi_1 _16959_ (.B2(_10173_),
    .C1(_10176_),
    .B1(_10170_),
    .A1(\cpu.ex.r_lr[10] ),
    .Y(_10177_),
    .A2(_10080_));
 sg13g2_nand4_1 _16960_ (.B(_10167_),
    .C(_10169_),
    .A(_10165_),
    .Y(_10178_),
    .D(_10177_));
 sg13g2_a221oi_1 _16961_ (.B2(_10178_),
    .C1(net858),
    .B1(net527),
    .A1(net1075),
    .Y(_10179_),
    .A2(net528));
 sg13g2_nor2_1 _16962_ (.A(net867),
    .B(\cpu.dec.imm[10] ),
    .Y(_10180_));
 sg13g2_o21ai_1 _16963_ (.B1(net735),
    .Y(_10181_),
    .A1(_10179_),
    .A2(_10180_));
 sg13g2_and2_1 _16964_ (.A(_10155_),
    .B(_10181_),
    .X(_10182_));
 sg13g2_buf_2 _16965_ (.A(_10182_),
    .X(_10183_));
 sg13g2_buf_1 _16966_ (.A(_10183_),
    .X(_10184_));
 sg13g2_nor2_1 _16967_ (.A(net209),
    .B(net208),
    .Y(_10185_));
 sg13g2_nand2_1 _16968_ (.Y(_10186_),
    .A(_10155_),
    .B(_10181_));
 sg13g2_buf_2 _16969_ (.A(_10186_),
    .X(_10187_));
 sg13g2_buf_1 _16970_ (.A(_10187_),
    .X(_10188_));
 sg13g2_inv_2 _16971_ (.Y(_10189_),
    .A(_10158_));
 sg13g2_buf_2 _16972_ (.A(_00301_),
    .X(_10190_));
 sg13g2_a21oi_1 _16973_ (.A1(_10189_),
    .A2(net209),
    .Y(_10191_),
    .B1(_10190_));
 sg13g2_o21ai_1 _16974_ (.B1(_10191_),
    .Y(_10192_),
    .A1(net207),
    .A2(_10119_));
 sg13g2_inv_2 _16975_ (.Y(_10193_),
    .A(_10153_));
 sg13g2_a221oi_1 _16976_ (.B2(_10117_),
    .C1(net208),
    .B1(_10113_),
    .A1(_09113_),
    .Y(_10194_),
    .A2(_09110_));
 sg13g2_buf_1 _16977_ (.A(_10158_),
    .X(_10195_));
 sg13g2_o21ai_1 _16978_ (.B1(net995),
    .Y(_10196_),
    .A1(_10193_),
    .A2(_10194_));
 sg13g2_buf_1 _16979_ (.A(net537),
    .X(_10197_));
 sg13g2_a21oi_1 _16980_ (.A1(_10192_),
    .A2(_10196_),
    .Y(_10198_),
    .B1(_10197_));
 sg13g2_a21o_1 _16981_ (.A2(_10185_),
    .A1(_10119_),
    .B1(_10198_),
    .X(_10199_));
 sg13g2_buf_1 _16982_ (.A(_08527_),
    .X(_10200_));
 sg13g2_nor2_1 _16983_ (.A(net742),
    .B(_10078_),
    .Y(_10201_));
 sg13g2_nand2b_1 _16984_ (.Y(_10202_),
    .B(net865),
    .A_N(net859));
 sg13g2_nor2_2 _16985_ (.A(net740),
    .B(_10202_),
    .Y(_10203_));
 sg13g2_a22oi_1 _16986_ (.Y(_10204_),
    .B1(_10203_),
    .B2(\cpu.ex.r_stmp[15] ),
    .A2(_10201_),
    .A1(\cpu.ex.r_13[15] ));
 sg13g2_nor2_1 _16987_ (.A(net742),
    .B(_10202_),
    .Y(_10205_));
 sg13g2_nor2_1 _16988_ (.A(net740),
    .B(_10078_),
    .Y(_10206_));
 sg13g2_a221oi_1 _16989_ (.B2(\cpu.ex.r_8[15] ),
    .C1(net659),
    .B1(_10206_),
    .A1(\cpu.ex.r_epc[15] ),
    .Y(_10207_),
    .A2(_10205_));
 sg13g2_a21oi_1 _16990_ (.A1(net659),
    .A2(_10204_),
    .Y(_10208_),
    .B1(_10207_));
 sg13g2_buf_1 _16991_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10209_));
 sg13g2_a22oi_1 _16992_ (.Y(_10210_),
    .B1(net660),
    .B2(_10209_),
    .A2(net861),
    .A1(\cpu.ex.r_lr[15] ));
 sg13g2_nor2b_1 _16993_ (.A(_10210_),
    .B_N(net866),
    .Y(_10211_));
 sg13g2_a21o_1 _16994_ (.A2(_10085_),
    .A1(\cpu.ex.r_14[15] ),
    .B1(_10211_),
    .X(_10212_));
 sg13g2_a22oi_1 _16995_ (.Y(_10213_),
    .B1(net660),
    .B2(\cpu.ex.r_10[15] ),
    .A2(net861),
    .A1(\cpu.ex.r_9[15] ));
 sg13g2_and2_1 _16996_ (.A(_09991_),
    .B(_09995_),
    .X(_10214_));
 sg13g2_buf_2 _16997_ (.A(_10214_),
    .X(_10215_));
 sg13g2_a22oi_1 _16998_ (.Y(_10216_),
    .B1(_10215_),
    .B2(\cpu.ex.r_15[15] ),
    .A2(_10005_),
    .A1(\cpu.ex.r_12[15] ));
 sg13g2_nand2b_1 _16999_ (.Y(_10217_),
    .B(net739),
    .A_N(_10216_));
 sg13g2_o21ai_1 _17000_ (.B1(_10217_),
    .Y(_10218_),
    .A1(_10172_),
    .A2(_10213_));
 sg13g2_a22oi_1 _17001_ (.Y(_10219_),
    .B1(_10094_),
    .B2(\cpu.ex.r_mult[31] ),
    .A2(_10016_),
    .A1(\cpu.ex.r_11[15] ));
 sg13g2_buf_2 _17002_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10220_));
 sg13g2_nand3_1 _17003_ (.B(net664),
    .C(_10094_),
    .A(_10220_),
    .Y(_10221_));
 sg13g2_o21ai_1 _17004_ (.B1(_10221_),
    .Y(_10222_),
    .A1(net664),
    .A2(_10219_));
 sg13g2_and2_1 _17005_ (.A(net579),
    .B(_10222_),
    .X(_10223_));
 sg13g2_or4_1 _17006_ (.A(_10208_),
    .B(_10212_),
    .C(_10218_),
    .D(_10223_),
    .X(_10224_));
 sg13g2_a22oi_1 _17007_ (.Y(_10225_),
    .B1(net527),
    .B2(_10224_),
    .A2(net528),
    .A1(net994));
 sg13g2_nor2_1 _17008_ (.A(net867),
    .B(\cpu.dec.imm[15] ),
    .Y(_10226_));
 sg13g2_a21o_1 _17009_ (.A2(_10225_),
    .A1(net867),
    .B1(_10226_),
    .X(_10227_));
 sg13g2_nor2b_1 _17010_ (.A(net1094),
    .B_N(net868),
    .Y(_10228_));
 sg13g2_a21oi_1 _17011_ (.A1(_10227_),
    .A2(net735),
    .Y(_10229_),
    .B1(_10228_));
 sg13g2_buf_1 _17012_ (.A(_10229_),
    .X(_10230_));
 sg13g2_buf_1 _17013_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10231_));
 sg13g2_buf_2 _17014_ (.A(_00299_),
    .X(_10232_));
 sg13g2_a22oi_1 _17015_ (.Y(_10233_),
    .B1(_10215_),
    .B2(\cpu.ex.r_11[14] ),
    .A2(net861),
    .A1(\cpu.ex.r_9[14] ));
 sg13g2_nor2_1 _17016_ (.A(_10172_),
    .B(_10233_),
    .Y(_10234_));
 sg13g2_nor2b_1 _17017_ (.A(net862),
    .B_N(net998),
    .Y(_10235_));
 sg13g2_buf_1 _17018_ (.A(_10235_),
    .X(_10236_));
 sg13g2_mux2_1 _17019_ (.A0(\cpu.ex.r_8[14] ),
    .A1(\cpu.ex.r_12[14] ),
    .S(net659),
    .X(_10237_));
 sg13g2_nor2b_1 _17020_ (.A(net859),
    .B_N(_10025_),
    .Y(_10238_));
 sg13g2_buf_1 _17021_ (.A(_10238_),
    .X(_10239_));
 sg13g2_buf_1 _17022_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10240_));
 sg13g2_inv_1 _17023_ (.Y(_10241_),
    .A(net1073));
 sg13g2_nor2_1 _17024_ (.A(\cpu.ex.r_lr[14] ),
    .B(_10126_),
    .Y(_10242_));
 sg13g2_a21oi_1 _17025_ (.A1(_10241_),
    .A2(_10126_),
    .Y(_10243_),
    .B1(_10242_));
 sg13g2_a22oi_1 _17026_ (.Y(_10244_),
    .B1(_10239_),
    .B2(_10243_),
    .A2(_10237_),
    .A1(_10236_));
 sg13g2_nor2_1 _17027_ (.A(net657),
    .B(_10244_),
    .Y(_10245_));
 sg13g2_a22oi_1 _17028_ (.Y(_10246_),
    .B1(_10239_),
    .B2(\cpu.ex.r_mult[30] ),
    .A2(_10236_),
    .A1(\cpu.ex.r_14[14] ));
 sg13g2_a22oi_1 _17029_ (.Y(_10247_),
    .B1(_10072_),
    .B2(\cpu.ex.r_epc[14] ),
    .A2(net737),
    .A1(\cpu.ex.r_stmp[14] ));
 sg13g2_nand2b_1 _17030_ (.Y(_10248_),
    .B(_10020_),
    .A_N(_10247_));
 sg13g2_o21ai_1 _17031_ (.B1(_10248_),
    .Y(_10249_),
    .A1(_10246_),
    .A2(_10050_));
 sg13g2_buf_1 _17032_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10250_));
 sg13g2_nor3_1 _17033_ (.A(net579),
    .B(_10136_),
    .C(net659),
    .Y(_10251_));
 sg13g2_nor2_1 _17034_ (.A(_00272_),
    .B(net662),
    .Y(_10252_));
 sg13g2_a22oi_1 _17035_ (.Y(_10253_),
    .B1(net739),
    .B2(_10252_),
    .A2(_10251_),
    .A1(_10250_));
 sg13g2_nor2b_2 _17036_ (.A(net863),
    .B_N(net999),
    .Y(_10254_));
 sg13g2_nand3_1 _17037_ (.B(net579),
    .C(_10254_),
    .A(\cpu.ex.r_13[14] ),
    .Y(_10255_));
 sg13g2_nor2b_1 _17038_ (.A(net999),
    .B_N(net1000),
    .Y(_10256_));
 sg13g2_buf_2 _17039_ (.A(_10256_),
    .X(_10257_));
 sg13g2_nand3_1 _17040_ (.B(net662),
    .C(_10257_),
    .A(\cpu.ex.r_10[14] ),
    .Y(_10258_));
 sg13g2_a21o_1 _17041_ (.A2(_10258_),
    .A1(_10255_),
    .B1(net860),
    .X(_10259_));
 sg13g2_o21ai_1 _17042_ (.B1(_10259_),
    .Y(_10260_),
    .A1(_10012_),
    .A2(_10253_));
 sg13g2_nor4_1 _17043_ (.A(_10234_),
    .B(_10245_),
    .C(_10249_),
    .D(_10260_),
    .Y(_10261_));
 sg13g2_buf_1 _17044_ (.A(net681),
    .X(_10262_));
 sg13g2_nand2_1 _17045_ (.Y(_10263_),
    .A(net578),
    .B(_10001_));
 sg13g2_o21ai_1 _17046_ (.B1(_10263_),
    .Y(_10264_),
    .A1(_10124_),
    .A2(_10261_));
 sg13g2_inv_1 _17047_ (.Y(_10265_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_nand2_1 _17048_ (.Y(_10266_),
    .A(net858),
    .B(_10265_));
 sg13g2_o21ai_1 _17049_ (.B1(_10266_),
    .Y(_10267_),
    .A1(net858),
    .A2(_10264_));
 sg13g2_a22oi_1 _17050_ (.Y(_10268_),
    .B1(net735),
    .B2(_10267_),
    .A2(net868),
    .A1(_08344_));
 sg13g2_buf_1 _17051_ (.A(_10268_),
    .X(_10269_));
 sg13g2_nor3_1 _17052_ (.A(net1074),
    .B(_10232_),
    .C(net206),
    .Y(_10270_));
 sg13g2_inv_1 _17053_ (.Y(_10271_),
    .A(net1074));
 sg13g2_inv_1 _17054_ (.Y(_10272_),
    .A(net206));
 sg13g2_nor2_1 _17055_ (.A(_10271_),
    .B(_10272_),
    .Y(_10273_));
 sg13g2_a21o_1 _17056_ (.A2(net735),
    .A1(_10227_),
    .B1(_10228_),
    .X(_10274_));
 sg13g2_buf_2 _17057_ (.A(_10274_),
    .X(_10275_));
 sg13g2_xnor2_1 _17058_ (.Y(_10276_),
    .A(_10232_),
    .B(_10275_));
 sg13g2_a22oi_1 _17059_ (.Y(_10277_),
    .B1(_10273_),
    .B2(_10276_),
    .A2(_10270_),
    .A1(net241));
 sg13g2_nor2_1 _17060_ (.A(_10229_),
    .B(net206),
    .Y(_10278_));
 sg13g2_inv_1 _17061_ (.Y(_10279_),
    .A(_10232_));
 sg13g2_nand2_1 _17062_ (.Y(_10280_),
    .A(_09113_),
    .B(_09110_));
 sg13g2_buf_1 _17063_ (.A(_10280_),
    .X(_10281_));
 sg13g2_buf_1 _17064_ (.A(_10281_),
    .X(_10282_));
 sg13g2_o21ai_1 _17065_ (.B1(net526),
    .Y(_10283_),
    .A1(net1074),
    .A2(_10279_));
 sg13g2_nand2_1 _17066_ (.Y(_10284_),
    .A(_10278_),
    .B(_10283_));
 sg13g2_o21ai_1 _17067_ (.B1(_10284_),
    .Y(_10285_),
    .A1(net537),
    .A2(_10277_));
 sg13g2_buf_1 _17068_ (.A(net683),
    .X(_10286_));
 sg13g2_buf_1 _17069_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10287_));
 sg13g2_mux2_1 _17070_ (.A0(_10287_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(_10125_),
    .X(_10288_));
 sg13g2_a22oi_1 _17071_ (.Y(_10289_),
    .B1(_10288_),
    .B2(_10028_),
    .A2(_10075_),
    .A1(_10231_));
 sg13g2_nor2_1 _17072_ (.A(_10202_),
    .B(_10289_),
    .Y(_10290_));
 sg13g2_nand3_1 _17073_ (.B(_10058_),
    .C(net861),
    .A(\cpu.ex.r_lr[13] ),
    .Y(_10291_));
 sg13g2_nand3_1 _17074_ (.B(net656),
    .C(net660),
    .A(\cpu.ex.r_10[13] ),
    .Y(_10292_));
 sg13g2_a21oi_1 _17075_ (.A1(_10291_),
    .A2(_10292_),
    .Y(_10293_),
    .B1(net659));
 sg13g2_nand3_1 _17076_ (.B(_10053_),
    .C(net663),
    .A(\cpu.ex.r_epc[13] ),
    .Y(_10294_));
 sg13g2_nand3_1 _17077_ (.B(net659),
    .C(net658),
    .A(\cpu.ex.r_13[13] ),
    .Y(_10295_));
 sg13g2_a21oi_1 _17078_ (.A1(_10294_),
    .A2(_10295_),
    .Y(_10296_),
    .B1(net662));
 sg13g2_nor3_1 _17079_ (.A(_10290_),
    .B(_10293_),
    .C(_10296_),
    .Y(_10297_));
 sg13g2_a22oi_1 _17080_ (.Y(_10298_),
    .B1(_10215_),
    .B2(\cpu.ex.r_11[13] ),
    .A2(_10005_),
    .A1(\cpu.ex.r_8[13] ));
 sg13g2_nand2b_1 _17081_ (.Y(_10299_),
    .B(net743),
    .A_N(_10298_));
 sg13g2_a22oi_1 _17082_ (.Y(_10300_),
    .B1(_10072_),
    .B2(\cpu.ex.r_9[13] ),
    .A2(net737),
    .A1(\cpu.ex.r_12[13] ));
 sg13g2_nand2b_1 _17083_ (.Y(_10301_),
    .B(net658),
    .A_N(_10300_));
 sg13g2_buf_1 _17084_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10302_));
 sg13g2_nor2_1 _17085_ (.A(net657),
    .B(net656),
    .Y(_10303_));
 sg13g2_and2_1 _17086_ (.A(net1000),
    .B(net998),
    .X(_10304_));
 sg13g2_buf_1 _17087_ (.A(_10304_),
    .X(_10305_));
 sg13g2_nor2b_1 _17088_ (.A(_00271_),
    .B_N(_10305_),
    .Y(_10306_));
 sg13g2_a21o_1 _17089_ (.A2(_10303_),
    .A1(_10302_),
    .B1(_10306_),
    .X(_10307_));
 sg13g2_a22oi_1 _17090_ (.Y(_10308_),
    .B1(_10075_),
    .B2(_10307_),
    .A2(_10085_),
    .A1(\cpu.ex.r_14[13] ));
 sg13g2_nand4_1 _17091_ (.B(_10299_),
    .C(_10301_),
    .A(_10297_),
    .Y(_10309_),
    .D(_10308_));
 sg13g2_a22oi_1 _17092_ (.Y(_10310_),
    .B1(_10009_),
    .B2(_10309_),
    .A2(net528),
    .A1(net577));
 sg13g2_nor2_1 _17093_ (.A(net867),
    .B(\cpu.dec.imm[13] ),
    .Y(_10311_));
 sg13g2_a21o_1 _17094_ (.A2(_10310_),
    .A1(net867),
    .B1(_10311_),
    .X(_10312_));
 sg13g2_nor2b_1 _17095_ (.A(net768),
    .B_N(net868),
    .Y(_10313_));
 sg13g2_a21oi_1 _17096_ (.A1(net735),
    .A2(_10312_),
    .Y(_10314_),
    .B1(_10313_));
 sg13g2_buf_2 _17097_ (.A(_10314_),
    .X(_10315_));
 sg13g2_buf_1 _17098_ (.A(net684),
    .X(_10316_));
 sg13g2_buf_2 _17099_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10317_));
 sg13g2_inv_1 _17100_ (.Y(_10318_),
    .A(_00270_));
 sg13g2_a22oi_1 _17101_ (.Y(_10319_),
    .B1(_10305_),
    .B2(_10318_),
    .A2(_10303_),
    .A1(_10317_));
 sg13g2_nand2b_1 _17102_ (.Y(_10320_),
    .B(_10075_),
    .A_N(_10319_));
 sg13g2_buf_1 _17103_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10321_));
 sg13g2_mux2_1 _17104_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(_10321_),
    .S(net734),
    .X(_10322_));
 sg13g2_a22oi_1 _17105_ (.Y(_10323_),
    .B1(_10322_),
    .B2(net860),
    .A2(_10016_),
    .A1(\cpu.ex.r_11[12] ));
 sg13g2_nand2b_1 _17106_ (.Y(_10324_),
    .B(_10215_),
    .A_N(_10323_));
 sg13g2_mux2_1 _17107_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_12[12] ),
    .S(_10125_),
    .X(_10325_));
 sg13g2_nand3_1 _17108_ (.B(_10130_),
    .C(_10325_),
    .A(net662),
    .Y(_10326_));
 sg13g2_nand3_1 _17109_ (.B(_10083_),
    .C(_10044_),
    .A(\cpu.ex.r_14[12] ),
    .Y(_10327_));
 sg13g2_mux2_1 _17110_ (.A0(\cpu.ex.r_9[12] ),
    .A1(\cpu.ex.r_13[12] ),
    .S(net734),
    .X(_10328_));
 sg13g2_nand3_1 _17111_ (.B(net658),
    .C(_10328_),
    .A(_10091_),
    .Y(_10329_));
 sg13g2_nand3_1 _17112_ (.B(_10003_),
    .C(net861),
    .A(\cpu.ex.r_lr[12] ),
    .Y(_10330_));
 sg13g2_and4_1 _17113_ (.A(_10326_),
    .B(_10327_),
    .C(_10329_),
    .D(_10330_),
    .X(_10331_));
 sg13g2_buf_1 _17114_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10332_));
 sg13g2_inv_1 _17115_ (.Y(_10333_),
    .A(\cpu.ex.r_10[12] ));
 sg13g2_nand3b_1 _17116_ (.B(net659),
    .C(\cpu.ex.r_stmp[12] ),
    .Y(_10334_),
    .A_N(net656));
 sg13g2_o21ai_1 _17117_ (.B1(_10334_),
    .Y(_10335_),
    .A1(_10333_),
    .A2(_10172_));
 sg13g2_a22oi_1 _17118_ (.Y(_10336_),
    .B1(_10335_),
    .B2(_10083_),
    .A2(_10033_),
    .A1(_10332_));
 sg13g2_nand4_1 _17119_ (.B(_10324_),
    .C(_10331_),
    .A(_10320_),
    .Y(_10337_),
    .D(_10336_));
 sg13g2_a22oi_1 _17120_ (.Y(_10338_),
    .B1(_10009_),
    .B2(_10337_),
    .A2(net528),
    .A1(net576));
 sg13g2_nor2_1 _17121_ (.A(net867),
    .B(\cpu.dec.imm[12] ),
    .Y(_10339_));
 sg13g2_a21o_1 _17122_ (.A2(_10338_),
    .A1(net867),
    .B1(_10339_),
    .X(_10340_));
 sg13g2_a22oi_1 _17123_ (.Y(_10341_),
    .B1(net735),
    .B2(_10340_),
    .A2(net868),
    .A1(_08149_));
 sg13g2_buf_2 _17124_ (.A(_10341_),
    .X(_10342_));
 sg13g2_inv_1 _17125_ (.Y(_10343_),
    .A(net1071));
 sg13g2_buf_8 _17126_ (.A(_00300_),
    .X(_10344_));
 sg13g2_a21oi_1 _17127_ (.A1(_10343_),
    .A2(_10344_),
    .Y(_10345_),
    .B1(net537));
 sg13g2_nor3_1 _17128_ (.A(_10315_),
    .B(_10342_),
    .C(_10345_),
    .Y(_10346_));
 sg13g2_inv_2 _17129_ (.Y(_10347_),
    .A(_10344_));
 sg13g2_a21o_1 _17130_ (.A2(_10312_),
    .A1(net735),
    .B1(_10313_),
    .X(_10348_));
 sg13g2_buf_2 _17131_ (.A(_10348_),
    .X(_10349_));
 sg13g2_nand4_1 _17132_ (.B(_10347_),
    .C(_10349_),
    .A(_10343_),
    .Y(_10350_),
    .D(_10342_));
 sg13g2_xnor2_1 _17133_ (.Y(_10351_),
    .A(_10347_),
    .B(_10342_));
 sg13g2_nand3_1 _17134_ (.B(_10315_),
    .C(_10351_),
    .A(_10321_),
    .Y(_10352_));
 sg13g2_a21oi_1 _17135_ (.A1(_10350_),
    .A2(_10352_),
    .Y(_10353_),
    .B1(net537));
 sg13g2_or2_1 _17136_ (.X(_10354_),
    .B(_10353_),
    .A(_10346_));
 sg13g2_buf_1 _17137_ (.A(_10354_),
    .X(_10355_));
 sg13g2_and2_1 _17138_ (.A(_10285_),
    .B(_10355_),
    .X(_10356_));
 sg13g2_nor4_1 _17139_ (.A(_10158_),
    .B(_10190_),
    .C(_10153_),
    .D(_10187_),
    .Y(_10357_));
 sg13g2_xnor2_1 _17140_ (.Y(_10358_),
    .A(_10190_),
    .B(_10187_));
 sg13g2_nand3_1 _17141_ (.B(_10153_),
    .C(_10358_),
    .A(_10195_),
    .Y(_10359_));
 sg13g2_nand2b_1 _17142_ (.Y(_10360_),
    .B(_10359_),
    .A_N(_10357_));
 sg13g2_inv_1 _17143_ (.Y(_10361_),
    .A(_10190_));
 sg13g2_o21ai_1 _17144_ (.B1(net526),
    .Y(_10362_),
    .A1(_10195_),
    .A2(_10361_));
 sg13g2_a22oi_1 _17145_ (.Y(_10363_),
    .B1(_10362_),
    .B2(_10185_),
    .A2(_10360_),
    .A1(net526));
 sg13g2_inv_1 _17146_ (.Y(_10364_),
    .A(_10363_));
 sg13g2_buf_1 _17147_ (.A(_10114_),
    .X(_10365_));
 sg13g2_nor2_1 _17148_ (.A(_10109_),
    .B(net537),
    .Y(_10366_));
 sg13g2_nor2_1 _17149_ (.A(_10067_),
    .B(_10108_),
    .Y(_10367_));
 sg13g2_buf_1 _17150_ (.A(_10367_),
    .X(_10368_));
 sg13g2_mux2_1 _17151_ (.A0(_10109_),
    .A1(_10366_),
    .S(net181),
    .X(_10369_));
 sg13g2_a22oi_1 _17152_ (.Y(_10370_),
    .B1(_10369_),
    .B2(_10112_),
    .A2(net182),
    .A1(net537));
 sg13g2_xnor2_1 _17153_ (.Y(_10371_),
    .A(_10109_),
    .B(net182));
 sg13g2_nor2_1 _17154_ (.A(_10112_),
    .B(net537),
    .Y(_10372_));
 sg13g2_a21oi_1 _17155_ (.A1(_10371_),
    .A2(_10372_),
    .Y(_10373_),
    .B1(net205));
 sg13g2_a21oi_1 _17156_ (.A1(net205),
    .A2(_10370_),
    .Y(_10374_),
    .B1(_10373_));
 sg13g2_buf_1 _17157_ (.A(_10374_),
    .X(_10375_));
 sg13g2_and4_1 _17158_ (.A(_10285_),
    .B(_10355_),
    .C(_10364_),
    .D(_10375_),
    .X(_10376_));
 sg13g2_inv_1 _17159_ (.Y(_10377_),
    .A(_00265_));
 sg13g2_mux4_1 _17160_ (.S0(net738),
    .A0(_10377_),
    .A1(\cpu.ex.r_11[7] ),
    .A2(\cpu.ex.r_mult[23] ),
    .A3(\cpu.ex.r_epc[7] ),
    .S1(net860),
    .X(_10378_));
 sg13g2_nand2_1 _17161_ (.Y(_10379_),
    .A(_10215_),
    .B(_10378_));
 sg13g2_a22oi_1 _17162_ (.Y(_10380_),
    .B1(net663),
    .B2(\cpu.ex.r_stmp[7] ),
    .A2(net658),
    .A1(\cpu.ex.r_12[7] ));
 sg13g2_nand2b_1 _17163_ (.Y(_10381_),
    .B(net737),
    .A_N(_10380_));
 sg13g2_a22oi_1 _17164_ (.Y(_10382_),
    .B1(_10032_),
    .B2(\cpu.ex.r_8[7] ),
    .A2(_10075_),
    .A1(\cpu.ex.r_13[7] ));
 sg13g2_nand2b_1 _17165_ (.Y(_10383_),
    .B(net658),
    .A_N(_10382_));
 sg13g2_or2_1 _17166_ (.X(_10384_),
    .B(net997),
    .A(net865));
 sg13g2_nor2_1 _17167_ (.A(net742),
    .B(_10384_),
    .Y(_10385_));
 sg13g2_mux2_1 _17168_ (.A0(\cpu.ex.r_lr[7] ),
    .A1(\cpu.ex.r_9[7] ),
    .S(net736),
    .X(_10386_));
 sg13g2_nor2_1 _17169_ (.A(net862),
    .B(net859),
    .Y(_10387_));
 sg13g2_buf_1 _17170_ (.A(\cpu.dec.user_io ),
    .X(_10388_));
 sg13g2_nand3b_1 _17171_ (.B(net734),
    .C(_10388_),
    .Y(_10389_),
    .A_N(net741));
 sg13g2_buf_1 _17172_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10390_));
 sg13g2_nand3b_1 _17173_ (.B(net741),
    .C(_10390_),
    .Y(_10391_),
    .A_N(_10022_));
 sg13g2_nand2_1 _17174_ (.Y(_10392_),
    .A(_10389_),
    .B(_10391_));
 sg13g2_mux2_1 _17175_ (.A0(\cpu.ex.r_10[7] ),
    .A1(\cpu.ex.r_14[7] ),
    .S(net864),
    .X(_10393_));
 sg13g2_and3_1 _17176_ (.X(_10394_),
    .A(net736),
    .B(net660),
    .C(_10393_));
 sg13g2_a221oi_1 _17177_ (.B2(_10392_),
    .C1(_10394_),
    .B1(_10387_),
    .A1(_10385_),
    .Y(_10395_),
    .A2(_10386_));
 sg13g2_nand4_1 _17178_ (.B(_10381_),
    .C(_10383_),
    .A(_10379_),
    .Y(_10396_),
    .D(_10395_));
 sg13g2_a22oi_1 _17179_ (.Y(_10397_),
    .B1(net527),
    .B2(_10396_),
    .A2(_10001_),
    .A1(_08952_));
 sg13g2_nor2_1 _17180_ (.A(net1001),
    .B(\cpu.dec.imm[7] ),
    .Y(_10398_));
 sg13g2_a21o_1 _17181_ (.A2(_10397_),
    .A1(_09984_),
    .B1(_10398_),
    .X(_10399_));
 sg13g2_a22oi_1 _17182_ (.Y(_10400_),
    .B1(_10120_),
    .B2(_10399_),
    .A2(net868),
    .A1(_08499_));
 sg13g2_buf_2 _17183_ (.A(_10400_),
    .X(_10401_));
 sg13g2_buf_1 _17184_ (.A(_10401_),
    .X(_10402_));
 sg13g2_nor2b_1 _17185_ (.A(_08435_),
    .B_N(net1002),
    .Y(_10403_));
 sg13g2_inv_1 _17186_ (.Y(_10404_),
    .A(_00264_));
 sg13g2_and3_1 _17187_ (.X(_10405_),
    .A(_10037_),
    .B(net863),
    .C(net997));
 sg13g2_nor2b_1 _17188_ (.A(net661),
    .B_N(\cpu.ex.r_8[6] ),
    .Y(_10406_));
 sg13g2_nor2_2 _17189_ (.A(net1000),
    .B(_10013_),
    .Y(_10407_));
 sg13g2_a22oi_1 _17190_ (.Y(_10408_),
    .B1(_10406_),
    .B2(_10407_),
    .A2(_10405_),
    .A1(_10404_));
 sg13g2_nor2_1 _17191_ (.A(_10038_),
    .B(_10050_),
    .Y(_10409_));
 sg13g2_a221oi_1 _17192_ (.B2(\cpu.ex.r_lr[6] ),
    .C1(net656),
    .B1(_10385_),
    .A1(\cpu.ex.r_stmp[6] ),
    .Y(_10410_),
    .A2(_10409_));
 sg13g2_a21oi_1 _17193_ (.A1(net656),
    .A2(_10408_),
    .Y(_10411_),
    .B1(_10410_));
 sg13g2_nand3_1 _17194_ (.B(net738),
    .C(_10019_),
    .A(\cpu.ex.r_epc[6] ),
    .Y(_10412_));
 sg13g2_nand3_1 _17195_ (.B(_10022_),
    .C(net658),
    .A(\cpu.ex.r_13[6] ),
    .Y(_10413_));
 sg13g2_a21oi_1 _17196_ (.A1(_10412_),
    .A2(_10413_),
    .Y(_10414_),
    .B1(net742));
 sg13g2_buf_2 _17197_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10415_));
 sg13g2_a22oi_1 _17198_ (.Y(_10416_),
    .B1(_10239_),
    .B2(_10415_),
    .A2(_10236_),
    .A1(\cpu.ex.r_14[6] ));
 sg13g2_nor2_1 _17199_ (.A(_10050_),
    .B(_10416_),
    .Y(_10417_));
 sg13g2_nand3_1 _17200_ (.B(net861),
    .C(net743),
    .A(\cpu.ex.r_9[6] ),
    .Y(_10418_));
 sg13g2_nand3_1 _17201_ (.B(_10236_),
    .C(_10254_),
    .A(\cpu.ex.r_12[6] ),
    .Y(_10419_));
 sg13g2_nand2_1 _17202_ (.Y(_10420_),
    .A(_10418_),
    .B(_10419_));
 sg13g2_buf_1 _17203_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10421_));
 sg13g2_and2_1 _17204_ (.A(_10025_),
    .B(net998),
    .X(_10422_));
 sg13g2_buf_1 _17205_ (.A(_10422_),
    .X(_10423_));
 sg13g2_a22oi_1 _17206_ (.Y(_10424_),
    .B1(_10423_),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10387_),
    .A1(_10421_));
 sg13g2_nand2_1 _17207_ (.Y(_10425_),
    .A(\cpu.ex.r_10[6] ),
    .B(_10236_));
 sg13g2_nand2_1 _17208_ (.Y(_10426_),
    .A(net657),
    .B(net738));
 sg13g2_a21oi_1 _17209_ (.A1(_10424_),
    .A2(_10425_),
    .Y(_10427_),
    .B1(_10426_));
 sg13g2_or4_1 _17210_ (.A(_10414_),
    .B(_10417_),
    .C(_10420_),
    .D(_10427_),
    .X(_10428_));
 sg13g2_o21ai_1 _17211_ (.B1(net527),
    .Y(_10429_),
    .A1(_10411_),
    .A2(_10428_));
 sg13g2_nand2_1 _17212_ (.Y(_10430_),
    .A(_08948_),
    .B(net580));
 sg13g2_nand3_1 _17213_ (.B(_10429_),
    .C(_10430_),
    .A(net1001),
    .Y(_10431_));
 sg13g2_or2_1 _17214_ (.X(_10432_),
    .B(\cpu.dec.imm[6] ),
    .A(_09983_));
 sg13g2_a21oi_1 _17215_ (.A1(_10431_),
    .A2(_10432_),
    .Y(_10433_),
    .B1(_10106_));
 sg13g2_nor2_1 _17216_ (.A(_10403_),
    .B(_10433_),
    .Y(_10434_));
 sg13g2_buf_2 _17217_ (.A(_10434_),
    .X(_10435_));
 sg13g2_buf_1 _17218_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10436_));
 sg13g2_a22oi_1 _17219_ (.Y(_10437_),
    .B1(_10203_),
    .B2(_10436_),
    .A2(_10201_),
    .A1(\cpu.ex.r_9[5] ));
 sg13g2_a221oi_1 _17220_ (.B2(\cpu.ex.r_12[5] ),
    .C1(net738),
    .B1(_10206_),
    .A1(\cpu.ex.r_mult[21] ),
    .Y(_10438_),
    .A2(_10205_));
 sg13g2_a21oi_1 _17221_ (.A1(net738),
    .A2(_10437_),
    .Y(_10439_),
    .B1(_10438_));
 sg13g2_nand2_1 _17222_ (.Y(_10440_),
    .A(net862),
    .B(net736));
 sg13g2_a22oi_1 _17223_ (.Y(_10441_),
    .B1(_10257_),
    .B2(\cpu.ex.r_11[5] ),
    .A2(_10254_),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_nand4_1 _17224_ (.B(net736),
    .C(_10052_),
    .A(\cpu.ex.r_10[5] ),
    .Y(_10442_),
    .D(_10082_));
 sg13g2_o21ai_1 _17225_ (.B1(_10442_),
    .Y(_10443_),
    .A1(_10440_),
    .A2(_10441_));
 sg13g2_inv_1 _17226_ (.Y(_10444_),
    .A(_00263_));
 sg13g2_a22oi_1 _17227_ (.Y(_10445_),
    .B1(_10423_),
    .B2(_10444_),
    .A2(_10387_),
    .A1(\cpu.ex.r_stmp[5] ));
 sg13g2_nor2_1 _17228_ (.A(_10050_),
    .B(_10445_),
    .Y(_10446_));
 sg13g2_a22oi_1 _17229_ (.Y(_10447_),
    .B1(_10239_),
    .B2(\cpu.ex.r_lr[5] ),
    .A2(_10236_),
    .A1(\cpu.ex.r_8[5] ));
 sg13g2_nor2_1 _17230_ (.A(_10384_),
    .B(_10447_),
    .Y(_10448_));
 sg13g2_nand3_1 _17231_ (.B(net742),
    .C(net739),
    .A(\cpu.ex.r_14[5] ),
    .Y(_10449_));
 sg13g2_nand3_1 _17232_ (.B(net740),
    .C(net866),
    .A(\cpu.ex.r_epc[5] ),
    .Y(_10450_));
 sg13g2_a21oi_1 _17233_ (.A1(_10449_),
    .A2(_10450_),
    .Y(_10451_),
    .B1(net664));
 sg13g2_or4_1 _17234_ (.A(_10443_),
    .B(_10446_),
    .C(_10448_),
    .D(_10451_),
    .X(_10452_));
 sg13g2_o21ai_1 _17235_ (.B1(_10008_),
    .Y(_10453_),
    .A1(_10439_),
    .A2(_10452_));
 sg13g2_nand2_1 _17236_ (.Y(_10454_),
    .A(_09732_),
    .B(net580));
 sg13g2_nand3_1 _17237_ (.B(_10453_),
    .C(_10454_),
    .A(net1001),
    .Y(_10455_));
 sg13g2_inv_1 _17238_ (.Y(_10456_),
    .A(\cpu.dec.imm[5] ));
 sg13g2_a21oi_1 _17239_ (.A1(net858),
    .A2(_10456_),
    .Y(_10457_),
    .B1(_09977_));
 sg13g2_mux2_1 _17240_ (.A0(_09979_),
    .A1(_08482_),
    .S(net1002),
    .X(_10458_));
 sg13g2_a21o_1 _17241_ (.A2(_10457_),
    .A1(_10455_),
    .B1(_10458_),
    .X(_10459_));
 sg13g2_buf_1 _17242_ (.A(_10459_),
    .X(_10460_));
 sg13g2_buf_1 _17243_ (.A(_00306_),
    .X(_10461_));
 sg13g2_inv_1 _17244_ (.Y(_10462_),
    .A(_00262_));
 sg13g2_mux2_1 _17245_ (.A0(_10462_),
    .A1(\cpu.ex.r_mult[20] ),
    .S(net860),
    .X(_10463_));
 sg13g2_mux2_1 _17246_ (.A0(_08516_),
    .A1(\cpu.ex.r_12[4] ),
    .S(net998),
    .X(_10464_));
 sg13g2_and2_1 _17247_ (.A(_10005_),
    .B(_10464_),
    .X(_10465_));
 sg13g2_a21o_1 _17248_ (.A2(_10463_),
    .A1(_10215_),
    .B1(_10465_),
    .X(_10466_));
 sg13g2_a22oi_1 _17249_ (.Y(_10467_),
    .B1(_10032_),
    .B2(\cpu.ex.r_8[4] ),
    .A2(_10075_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_nand3b_1 _17250_ (.B(net862),
    .C(\cpu.ex.r_9[4] ),
    .Y(_10468_),
    .A_N(net865));
 sg13g2_nand3b_1 _17251_ (.B(net865),
    .C(\cpu.ex.r_10[4] ),
    .Y(_10469_),
    .A_N(net862));
 sg13g2_a21o_1 _17252_ (.A2(_10469_),
    .A1(_10468_),
    .B1(net864),
    .X(_10470_));
 sg13g2_o21ai_1 _17253_ (.B1(_10470_),
    .Y(_10471_),
    .A1(net741),
    .A2(_10467_));
 sg13g2_nand3_1 _17254_ (.B(net743),
    .C(_10215_),
    .A(\cpu.ex.r_11[4] ),
    .Y(_10472_));
 sg13g2_nand3_1 _17255_ (.B(net660),
    .C(net739),
    .A(\cpu.ex.r_14[4] ),
    .Y(_10473_));
 sg13g2_buf_1 _17256_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10474_));
 sg13g2_mux2_1 _17257_ (.A0(_10474_),
    .A1(\cpu.ex.r_stmp[4] ),
    .S(net997),
    .X(_10475_));
 sg13g2_nand3_1 _17258_ (.B(_10019_),
    .C(_10475_),
    .A(net742),
    .Y(_10476_));
 sg13g2_mux2_1 _17259_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_epc[4] ),
    .S(net863),
    .X(_10477_));
 sg13g2_nand3_1 _17260_ (.B(net866),
    .C(_10477_),
    .A(net740),
    .Y(_10478_));
 sg13g2_nand4_1 _17261_ (.B(_10473_),
    .C(_10476_),
    .A(_10472_),
    .Y(_10479_),
    .D(_10478_));
 sg13g2_a221oi_1 _17262_ (.B2(net656),
    .C1(_10479_),
    .B1(_10471_),
    .A1(net734),
    .Y(_10480_),
    .A2(_10466_));
 sg13g2_nand2_1 _17263_ (.Y(_10481_),
    .A(_09149_),
    .B(net580));
 sg13g2_o21ai_1 _17264_ (.B1(_10481_),
    .Y(_10482_),
    .A1(_10124_),
    .A2(_10480_));
 sg13g2_or2_1 _17265_ (.X(_10483_),
    .B(\cpu.dec.imm[4] ),
    .A(net1001));
 sg13g2_o21ai_1 _17266_ (.B1(_10483_),
    .Y(_10484_),
    .A1(net858),
    .A2(_10482_));
 sg13g2_nor2b_1 _17267_ (.A(net1038),
    .B_N(_09977_),
    .Y(_10485_));
 sg13g2_a21o_1 _17268_ (.A2(_10484_),
    .A1(_09981_),
    .B1(_10485_),
    .X(_10486_));
 sg13g2_buf_1 _17269_ (.A(_10486_),
    .X(_10487_));
 sg13g2_nand2b_1 _17270_ (.Y(_10488_),
    .B(_10487_),
    .A_N(_10461_));
 sg13g2_buf_2 _17271_ (.A(_00305_),
    .X(_10489_));
 sg13g2_a21oi_1 _17272_ (.A1(net295),
    .A2(_10488_),
    .Y(_10490_),
    .B1(_10489_));
 sg13g2_nor2_1 _17273_ (.A(net295),
    .B(_10488_),
    .Y(_10491_));
 sg13g2_o21ai_1 _17274_ (.B1(_10282_),
    .Y(_10492_),
    .A1(_10490_),
    .A2(_10491_));
 sg13g2_buf_1 _17275_ (.A(_10492_),
    .X(_10493_));
 sg13g2_nand3_1 _17276_ (.B(_10435_),
    .C(_10493_),
    .A(net240),
    .Y(_10494_));
 sg13g2_nand2b_1 _17277_ (.Y(_10495_),
    .B(_10281_),
    .A_N(_00304_));
 sg13g2_buf_1 _17278_ (.A(_10495_),
    .X(_10496_));
 sg13g2_nand2_1 _17279_ (.Y(_10497_),
    .A(net240),
    .B(_10496_));
 sg13g2_nand2b_1 _17280_ (.Y(_10498_),
    .B(_10493_),
    .A_N(_10497_));
 sg13g2_xor2_1 _17281_ (.B(_09119_),
    .A(_09105_),
    .X(_10499_));
 sg13g2_and3_1 _17282_ (.X(_10500_),
    .A(_09126_),
    .B(_10281_),
    .C(_10499_));
 sg13g2_buf_2 _17283_ (.A(_10500_),
    .X(_10501_));
 sg13g2_nor2_1 _17284_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_10501_),
    .Y(_10502_));
 sg13g2_buf_1 _17285_ (.A(_00273_),
    .X(_10503_));
 sg13g2_buf_8 _17286_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10504_));
 sg13g2_buf_8 _17287_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10505_));
 sg13g2_buf_2 _17288_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10506_));
 sg13g2_buf_1 _17289_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10507_));
 sg13g2_nor4_2 _17290_ (.A(_10504_),
    .B(_10505_),
    .C(_10506_),
    .Y(_10508_),
    .D(_10507_));
 sg13g2_nor2_1 _17291_ (.A(_10503_),
    .B(_10508_),
    .Y(_10509_));
 sg13g2_inv_1 _17292_ (.Y(_10510_),
    .A(_10509_));
 sg13g2_nor4_1 _17293_ (.A(_08967_),
    .B(_08557_),
    .C(_09009_),
    .D(_10510_),
    .Y(_10511_));
 sg13g2_inv_1 _17294_ (.Y(_10512_),
    .A(net1091));
 sg13g2_nand3_1 _17295_ (.B(_10512_),
    .C(_08536_),
    .A(_00189_),
    .Y(_10513_));
 sg13g2_nor2_1 _17296_ (.A(_08983_),
    .B(_08991_),
    .Y(_10514_));
 sg13g2_inv_1 _17297_ (.Y(_10515_),
    .A(_08967_));
 sg13g2_and3_1 _17298_ (.X(_10516_),
    .A(_10515_),
    .B(_09006_),
    .C(_10509_));
 sg13g2_nor4_1 _17299_ (.A(_08967_),
    .B(_08992_),
    .C(_10503_),
    .D(_10508_),
    .Y(_10517_));
 sg13g2_nor4_1 _17300_ (.A(_08967_),
    .B(_09007_),
    .C(_10503_),
    .D(_10508_),
    .Y(_10518_));
 sg13g2_a221oi_1 _17301_ (.B2(_09006_),
    .C1(_10518_),
    .B1(_10517_),
    .A1(_10514_),
    .Y(_10519_),
    .A2(_10516_));
 sg13g2_buf_1 _17302_ (.A(_10519_),
    .X(_10520_));
 sg13g2_buf_1 _17303_ (.A(\cpu.br ),
    .X(_10521_));
 sg13g2_o21ai_1 _17304_ (.B1(_10521_),
    .Y(_10522_),
    .A1(_10513_),
    .A2(_10520_));
 sg13g2_a21o_1 _17305_ (.A2(_10511_),
    .A1(_08615_),
    .B1(_10522_),
    .X(_10523_));
 sg13g2_buf_8 _17306_ (.A(_10523_),
    .X(_10524_));
 sg13g2_buf_8 _17307_ (.A(_10524_),
    .X(_10525_));
 sg13g2_buf_8 _17308_ (.A(_10525_),
    .X(_10526_));
 sg13g2_inv_1 _17309_ (.Y(_10527_),
    .A(_00291_));
 sg13g2_inv_1 _17310_ (.Y(_10528_),
    .A(_00297_));
 sg13g2_or3_1 _17311_ (.A(_09105_),
    .B(_09119_),
    .C(\cpu.ex.r_mult_off[2] ),
    .X(_10529_));
 sg13g2_xor2_1 _17312_ (.B(_10529_),
    .A(\cpu.ex.r_mult_off[3] ),
    .X(_10530_));
 sg13g2_and2_1 _17313_ (.A(_09116_),
    .B(_10530_),
    .X(_10531_));
 sg13g2_buf_2 _17314_ (.A(_10531_),
    .X(_10532_));
 sg13g2_mux2_1 _17315_ (.A0(_10527_),
    .A1(_10528_),
    .S(_10532_),
    .X(_10533_));
 sg13g2_xor2_1 _17316_ (.B(_10506_),
    .A(net1076),
    .X(_10534_));
 sg13g2_buf_1 _17317_ (.A(_10504_),
    .X(_10535_));
 sg13g2_xor2_1 _17318_ (.B(_10535_),
    .A(_09963_),
    .X(_10536_));
 sg13g2_buf_8 _17319_ (.A(_10507_),
    .X(_10537_));
 sg13g2_xor2_1 _17320_ (.B(_10537_),
    .A(_09967_),
    .X(_10538_));
 sg13g2_xor2_1 _17321_ (.B(_10505_),
    .A(net1077),
    .X(_10539_));
 sg13g2_nor4_1 _17322_ (.A(_10534_),
    .B(_10536_),
    .C(_10538_),
    .D(_10539_),
    .Y(_10540_));
 sg13g2_nand3_1 _17323_ (.B(_09988_),
    .C(_10540_),
    .A(_09470_),
    .Y(_10541_));
 sg13g2_nand2_1 _17324_ (.Y(_10542_),
    .A(_09988_),
    .B(_10540_));
 sg13g2_buf_1 _17325_ (.A(_10542_),
    .X(_10543_));
 sg13g2_buf_1 _17326_ (.A(_10506_),
    .X(_10544_));
 sg13g2_buf_1 _17327_ (.A(net991),
    .X(_10545_));
 sg13g2_buf_1 _17328_ (.A(net857),
    .X(_10546_));
 sg13g2_buf_1 _17329_ (.A(net733),
    .X(_10547_));
 sg13g2_buf_2 _17330_ (.A(net993),
    .X(_10548_));
 sg13g2_buf_8 _17331_ (.A(_10548_),
    .X(_10549_));
 sg13g2_nor2b_1 _17332_ (.A(_10505_),
    .B_N(net992),
    .Y(_10550_));
 sg13g2_buf_1 _17333_ (.A(_10550_),
    .X(_10551_));
 sg13g2_nor2b_1 _17334_ (.A(_10537_),
    .B_N(_10505_),
    .Y(_10552_));
 sg13g2_buf_2 _17335_ (.A(_10552_),
    .X(_10553_));
 sg13g2_buf_1 _17336_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10554_));
 sg13g2_buf_1 _17337_ (.A(_10505_),
    .X(_10555_));
 sg13g2_buf_1 _17338_ (.A(net992),
    .X(_10556_));
 sg13g2_and3_1 _17339_ (.X(_10557_),
    .A(net990),
    .B(net855),
    .C(\cpu.ex.r_stmp[2] ));
 sg13g2_a221oi_1 _17340_ (.B2(_10554_),
    .C1(_10557_),
    .B1(_10553_),
    .A1(_08081_),
    .Y(_10558_),
    .A2(_10551_));
 sg13g2_inv_1 _17341_ (.Y(_10559_),
    .A(net992));
 sg13g2_buf_1 _17342_ (.A(_10559_),
    .X(_10560_));
 sg13g2_and2_1 _17343_ (.A(net993),
    .B(_10505_),
    .X(_10561_));
 sg13g2_buf_2 _17344_ (.A(_10561_),
    .X(_10562_));
 sg13g2_nand3_1 _17345_ (.B(\cpu.ex.r_epc[2] ),
    .C(_10562_),
    .A(net731),
    .Y(_10563_));
 sg13g2_o21ai_1 _17346_ (.B1(_10563_),
    .Y(_10564_),
    .A1(net732),
    .A2(_10558_));
 sg13g2_nor3_1 _17347_ (.A(net993),
    .B(net990),
    .C(net855),
    .Y(_10565_));
 sg13g2_nand2_1 _17348_ (.Y(_10566_),
    .A(\cpu.ex.r_8[2] ),
    .B(_10565_));
 sg13g2_buf_8 _17349_ (.A(net855),
    .X(_10567_));
 sg13g2_inv_1 _17350_ (.Y(_10568_),
    .A(_00260_));
 sg13g2_nand3_1 _17351_ (.B(_10568_),
    .C(_10562_),
    .A(net730),
    .Y(_10569_));
 sg13g2_nand3_1 _17352_ (.B(_10566_),
    .C(_10569_),
    .A(_10546_),
    .Y(_10570_));
 sg13g2_o21ai_1 _17353_ (.B1(_10570_),
    .Y(_10571_),
    .A1(net655),
    .A2(_10564_));
 sg13g2_nor2b_1 _17354_ (.A(_10535_),
    .B_N(_10505_),
    .Y(_10572_));
 sg13g2_buf_1 _17355_ (.A(_10572_),
    .X(_10573_));
 sg13g2_nand3_1 _17356_ (.B(\cpu.ex.r_14[2] ),
    .C(_10573_),
    .A(net857),
    .Y(_10574_));
 sg13g2_inv_2 _17357_ (.Y(_10575_),
    .A(net991));
 sg13g2_buf_2 _17358_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10576_));
 sg13g2_nor2b_1 _17359_ (.A(_10505_),
    .B_N(_10504_),
    .Y(_10577_));
 sg13g2_buf_2 _17360_ (.A(_10577_),
    .X(_10578_));
 sg13g2_nand3_1 _17361_ (.B(_10576_),
    .C(_10578_),
    .A(_10575_),
    .Y(_10579_));
 sg13g2_a21oi_1 _17362_ (.A1(_10574_),
    .A2(_10579_),
    .Y(_10580_),
    .B1(net731));
 sg13g2_nor2b_1 _17363_ (.A(net993),
    .B_N(net992),
    .Y(_10581_));
 sg13g2_buf_2 _17364_ (.A(_10581_),
    .X(_10582_));
 sg13g2_nor2b_1 _17365_ (.A(net992),
    .B_N(net993),
    .Y(_10583_));
 sg13g2_buf_1 _17366_ (.A(_10583_),
    .X(_10584_));
 sg13g2_a22oi_1 _17367_ (.Y(_10585_),
    .B1(_10584_),
    .B2(\cpu.ex.r_9[2] ),
    .A2(_10582_),
    .A1(\cpu.ex.r_12[2] ));
 sg13g2_nor2b_1 _17368_ (.A(net990),
    .B_N(net991),
    .Y(_10586_));
 sg13g2_buf_1 _17369_ (.A(_10586_),
    .X(_10587_));
 sg13g2_nor2b_1 _17370_ (.A(_10585_),
    .B_N(_10587_),
    .Y(_10588_));
 sg13g2_nand2_1 _17371_ (.Y(_10589_),
    .A(net856),
    .B(net731));
 sg13g2_nor2_1 _17372_ (.A(net990),
    .B(net991),
    .Y(_10590_));
 sg13g2_and2_1 _17373_ (.A(net990),
    .B(net991),
    .X(_10591_));
 sg13g2_buf_1 _17374_ (.A(_10591_),
    .X(_10592_));
 sg13g2_a22oi_1 _17375_ (.Y(_10593_),
    .B1(_10592_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10590_),
    .A1(\cpu.ex.r_lr[2] ));
 sg13g2_nand4_1 _17376_ (.B(net730),
    .C(\cpu.ex.r_13[2] ),
    .A(net857),
    .Y(_10594_),
    .D(_10578_));
 sg13g2_o21ai_1 _17377_ (.B1(_10594_),
    .Y(_10595_),
    .A1(_10589_),
    .A2(_10593_));
 sg13g2_nor3_1 _17378_ (.A(_10580_),
    .B(_10588_),
    .C(_10595_),
    .Y(_10596_));
 sg13g2_nor2b_1 _17379_ (.A(_10504_),
    .B_N(_10506_),
    .Y(_10597_));
 sg13g2_buf_2 _17380_ (.A(_10597_),
    .X(_10598_));
 sg13g2_and2_1 _17381_ (.A(net731),
    .B(_10598_),
    .X(_10599_));
 sg13g2_buf_2 _17382_ (.A(_10599_),
    .X(_10600_));
 sg13g2_nand2b_1 _17383_ (.Y(_10601_),
    .B(_10504_),
    .A_N(_10506_));
 sg13g2_buf_2 _17384_ (.A(_10601_),
    .X(_10602_));
 sg13g2_nor2_1 _17385_ (.A(net731),
    .B(_10602_),
    .Y(_10603_));
 sg13g2_buf_2 _17386_ (.A(_10603_),
    .X(_10604_));
 sg13g2_a22oi_1 _17387_ (.Y(_10605_),
    .B1(_10604_),
    .B2(\cpu.ex.r_mult[18] ),
    .A2(_10600_),
    .A1(\cpu.ex.r_10[2] ));
 sg13g2_buf_1 _17388_ (.A(_10555_),
    .X(_10606_));
 sg13g2_buf_8 _17389_ (.A(net854),
    .X(_10607_));
 sg13g2_buf_1 _17390_ (.A(_10607_),
    .X(_10608_));
 sg13g2_nand2b_1 _17391_ (.Y(_10609_),
    .B(net654),
    .A_N(_10605_));
 sg13g2_nand4_1 _17392_ (.B(_10571_),
    .C(_10596_),
    .A(net575),
    .Y(_10610_),
    .D(_10609_));
 sg13g2_buf_1 _17393_ (.A(_10610_),
    .X(_10611_));
 sg13g2_nand3_1 _17394_ (.B(_10541_),
    .C(_10611_),
    .A(_10532_),
    .Y(_10612_));
 sg13g2_inv_1 _17395_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(_10532_));
 sg13g2_a22oi_1 _17396_ (.Y(_10613_),
    .B1(_10592_),
    .B2(\cpu.ex.r_11[10] ),
    .A2(_10590_),
    .A1(\cpu.ex.r_lr[10] ));
 sg13g2_nand2b_1 _17397_ (.Y(_10614_),
    .B(_10584_),
    .A_N(_10613_));
 sg13g2_nor2b_1 _17398_ (.A(net992),
    .B_N(_10544_),
    .Y(_10615_));
 sg13g2_buf_2 _17399_ (.A(_10615_),
    .X(_10616_));
 sg13g2_and2_1 _17400_ (.A(_10616_),
    .B(_10578_),
    .X(_10617_));
 sg13g2_buf_1 _17401_ (.A(_10617_),
    .X(_10618_));
 sg13g2_nor2b_1 _17402_ (.A(_10506_),
    .B_N(net992),
    .Y(_10619_));
 sg13g2_buf_2 _17403_ (.A(_10619_),
    .X(_10620_));
 sg13g2_and2_1 _17404_ (.A(_10573_),
    .B(_10620_),
    .X(_10621_));
 sg13g2_buf_1 _17405_ (.A(_10621_),
    .X(_10622_));
 sg13g2_a22oi_1 _17406_ (.Y(_10623_),
    .B1(_10622_),
    .B2(\cpu.ex.r_stmp[10] ),
    .A2(_10618_),
    .A1(\cpu.ex.r_9[10] ));
 sg13g2_buf_1 _17407_ (.A(net730),
    .X(_10624_));
 sg13g2_mux2_1 _17408_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(_10158_),
    .S(_10624_),
    .X(_10625_));
 sg13g2_buf_1 _17409_ (.A(_10562_),
    .X(_10626_));
 sg13g2_and2_1 _17410_ (.A(_10575_),
    .B(_10626_),
    .X(_10627_));
 sg13g2_mux2_1 _17411_ (.A0(_10161_),
    .A1(\cpu.ex.r_10[10] ),
    .S(_10547_),
    .X(_10628_));
 sg13g2_buf_1 _17412_ (.A(_10624_),
    .X(_10629_));
 sg13g2_nand2b_1 _17413_ (.Y(_10630_),
    .B(_10555_),
    .A_N(net993));
 sg13g2_buf_1 _17414_ (.A(_10630_),
    .X(_10631_));
 sg13g2_nor2_1 _17415_ (.A(_10629_),
    .B(_10631_),
    .Y(_10632_));
 sg13g2_a22oi_1 _17416_ (.Y(_10633_),
    .B1(_10628_),
    .B2(_10632_),
    .A2(_10627_),
    .A1(_10625_));
 sg13g2_buf_1 _17417_ (.A(_10587_),
    .X(_10634_));
 sg13g2_buf_1 _17418_ (.A(net855),
    .X(_10635_));
 sg13g2_nor2_1 _17419_ (.A(net732),
    .B(net728),
    .Y(_10636_));
 sg13g2_and3_1 _17420_ (.X(_10637_),
    .A(net732),
    .B(_10635_),
    .C(\cpu.ex.r_13[10] ));
 sg13g2_a21o_1 _17421_ (.A2(_10636_),
    .A1(\cpu.ex.r_8[10] ),
    .B1(_10637_),
    .X(_10638_));
 sg13g2_nand2_1 _17422_ (.Y(_10639_),
    .A(_10545_),
    .B(net855));
 sg13g2_nor2_1 _17423_ (.A(_00268_),
    .B(_10639_),
    .Y(_10640_));
 sg13g2_mux2_1 _17424_ (.A0(\cpu.ex.r_12[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net729),
    .X(_10641_));
 sg13g2_and3_1 _17425_ (.X(_10642_),
    .A(_10629_),
    .B(_10598_),
    .C(_10641_));
 sg13g2_a221oi_1 _17426_ (.B2(_10626_),
    .C1(_10642_),
    .B1(_10640_),
    .A1(_10634_),
    .Y(_10643_),
    .A2(_10638_));
 sg13g2_nand4_1 _17427_ (.B(_10623_),
    .C(_10633_),
    .A(_10614_),
    .Y(_10644_),
    .D(_10643_));
 sg13g2_buf_1 _17428_ (.A(net575),
    .X(_10645_));
 sg13g2_mux2_1 _17429_ (.A0(net1075),
    .A1(_10644_),
    .S(_10645_),
    .X(_10646_));
 sg13g2_nand2_1 _17430_ (.Y(_10647_),
    .A(\cpu.ex.c_mult_off[3] ),
    .B(_10646_));
 sg13g2_nand3_1 _17431_ (.B(_10612_),
    .C(_10647_),
    .A(_10526_),
    .Y(_10648_));
 sg13g2_o21ai_1 _17432_ (.B1(_10648_),
    .Y(_10649_),
    .A1(net294),
    .A2(_10533_));
 sg13g2_nand2b_1 _17433_ (.Y(_10650_),
    .B(_10521_),
    .A_N(_08514_));
 sg13g2_or3_1 _17434_ (.A(_08562_),
    .B(_08615_),
    .C(_10650_),
    .X(_10651_));
 sg13g2_buf_1 _17435_ (.A(_10651_),
    .X(_10652_));
 sg13g2_nand4_1 _17436_ (.B(_08537_),
    .C(_08547_),
    .A(_08533_),
    .Y(_10653_),
    .D(_08555_));
 sg13g2_nor2_1 _17437_ (.A(_08967_),
    .B(_09009_),
    .Y(_10654_));
 sg13g2_a21o_1 _17438_ (.A2(_10654_),
    .A1(_10653_),
    .B1(_10650_),
    .X(_10655_));
 sg13g2_buf_1 _17439_ (.A(_10655_),
    .X(_10656_));
 sg13g2_nor2_1 _17440_ (.A(_08588_),
    .B(net575),
    .Y(_10657_));
 sg13g2_mux2_1 _17441_ (.A0(\cpu.ex.r_9[0] ),
    .A1(\cpu.ex.r_13[0] ),
    .S(net855),
    .X(_10658_));
 sg13g2_buf_1 _17442_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10659_));
 sg13g2_mux4_1 _17443_ (.S0(net991),
    .A0(_10659_),
    .A1(\cpu.ex.r_11[0] ),
    .A2(\cpu.ex.r_mult[16] ),
    .A3(\cpu.ex.r_15[0] ),
    .S1(net730),
    .X(_10660_));
 sg13g2_a22oi_1 _17444_ (.Y(_10661_),
    .B1(_10660_),
    .B2(net729),
    .A2(_10658_),
    .A1(net651));
 sg13g2_buf_1 _17445_ (.A(_10549_),
    .X(_10662_));
 sg13g2_nand2b_1 _17446_ (.Y(_10663_),
    .B(net650),
    .A_N(_10661_));
 sg13g2_nor2b_1 _17447_ (.A(net991),
    .B_N(net990),
    .Y(_10664_));
 sg13g2_buf_1 _17448_ (.A(_10664_),
    .X(_10665_));
 sg13g2_nand3_1 _17449_ (.B(\cpu.ex.r_stmp[0] ),
    .C(_10665_),
    .A(net728),
    .Y(_10666_));
 sg13g2_nand3_1 _17450_ (.B(\cpu.ex.r_8[0] ),
    .C(_10587_),
    .A(net731),
    .Y(_10667_));
 sg13g2_a21o_1 _17451_ (.A2(_10667_),
    .A1(_10666_),
    .B1(net650),
    .X(_10668_));
 sg13g2_and3_1 _17452_ (.X(_10669_),
    .A(_10606_),
    .B(net857),
    .C(\cpu.ex.r_14[0] ));
 sg13g2_a21o_1 _17453_ (.A2(_10590_),
    .A1(_09007_),
    .B1(_10669_),
    .X(_10670_));
 sg13g2_nand3b_1 _17454_ (.B(_10567_),
    .C(\cpu.ex.r_12[0] ),
    .Y(_10671_),
    .A_N(net854));
 sg13g2_nand3b_1 _17455_ (.B(\cpu.ex.r_10[0] ),
    .C(_10606_),
    .Y(_10672_),
    .A_N(_10567_));
 sg13g2_nand2_1 _17456_ (.Y(_10673_),
    .A(_10671_),
    .B(_10672_));
 sg13g2_a22oi_1 _17457_ (.Y(_10674_),
    .B1(_10673_),
    .B2(_10598_),
    .A2(_10670_),
    .A1(_10582_));
 sg13g2_and4_1 _17458_ (.A(net575),
    .B(_10663_),
    .C(_10668_),
    .D(_10674_),
    .X(_10675_));
 sg13g2_nor2_1 _17459_ (.A(_10657_),
    .B(_10675_),
    .Y(_10676_));
 sg13g2_nor4_1 _17460_ (.A(_08557_),
    .B(_10520_),
    .C(_10657_),
    .D(_10675_),
    .Y(_10677_));
 sg13g2_a22oi_1 _17461_ (.Y(_10678_),
    .B1(_10677_),
    .B2(_08615_),
    .A2(_10676_),
    .A1(_10522_));
 sg13g2_and3_1 _17462_ (.X(_10679_),
    .A(_10652_),
    .B(_10656_),
    .C(_10678_));
 sg13g2_buf_1 _17463_ (.A(_10679_),
    .X(_10680_));
 sg13g2_inv_1 _17464_ (.Y(_10681_),
    .A(_00293_));
 sg13g2_nor2_1 _17465_ (.A(net991),
    .B(net992),
    .Y(_10682_));
 sg13g2_buf_2 _17466_ (.A(_10682_),
    .X(_10683_));
 sg13g2_buf_1 _17467_ (.A(_10683_),
    .X(_10684_));
 sg13g2_buf_1 _17468_ (.A(_10573_),
    .X(_10685_));
 sg13g2_nand3_1 _17469_ (.B(net649),
    .C(net648),
    .A(_10096_),
    .Y(_10686_));
 sg13g2_buf_1 _17470_ (.A(_10578_),
    .X(_10687_));
 sg13g2_mux2_1 _17471_ (.A0(\cpu.ex.r_9[8] ),
    .A1(\cpu.ex.r_13[8] ),
    .S(net730),
    .X(_10688_));
 sg13g2_nand3_1 _17472_ (.B(net727),
    .C(_10688_),
    .A(net655),
    .Y(_10689_));
 sg13g2_nor2_1 _17473_ (.A(net993),
    .B(net990),
    .Y(_10690_));
 sg13g2_buf_1 _17474_ (.A(_10690_),
    .X(_10691_));
 sg13g2_nand4_1 _17475_ (.B(net653),
    .C(\cpu.ex.r_12[8] ),
    .A(net655),
    .Y(_10692_),
    .D(_10691_));
 sg13g2_nor2b_1 _17476_ (.A(_00266_),
    .B_N(net730),
    .Y(_10693_));
 sg13g2_nor2b_1 _17477_ (.A(net728),
    .B_N(\cpu.ex.r_11[8] ),
    .Y(_10694_));
 sg13g2_and3_1 _17478_ (.X(_10695_),
    .A(net732),
    .B(net854),
    .C(net857));
 sg13g2_o21ai_1 _17479_ (.B1(_10695_),
    .Y(_10696_),
    .A1(_10693_),
    .A2(_10694_));
 sg13g2_nand4_1 _17480_ (.B(_10689_),
    .C(_10692_),
    .A(_10686_),
    .Y(_10697_),
    .D(_10696_));
 sg13g2_a22oi_1 _17481_ (.Y(_10698_),
    .B1(_10620_),
    .B2(\cpu.ex.r_stmp[8] ),
    .A2(_10616_),
    .A1(\cpu.ex.r_10[8] ));
 sg13g2_nand3_1 _17482_ (.B(net649),
    .C(net652),
    .A(\cpu.ex.r_epc[8] ),
    .Y(_10699_));
 sg13g2_o21ai_1 _17483_ (.B1(_10699_),
    .Y(_10700_),
    .A1(_10631_),
    .A2(_10698_));
 sg13g2_and2_1 _17484_ (.A(net854),
    .B(net730),
    .X(_10701_));
 sg13g2_buf_1 _17485_ (.A(_10701_),
    .X(_10702_));
 sg13g2_nor2_2 _17486_ (.A(net729),
    .B(net728),
    .Y(_10703_));
 sg13g2_a22oi_1 _17487_ (.Y(_10704_),
    .B1(_10703_),
    .B2(\cpu.ex.r_lr[8] ),
    .A2(_10702_),
    .A1(\cpu.ex.r_mult[24] ));
 sg13g2_nor2_1 _17488_ (.A(_10602_),
    .B(_10704_),
    .Y(_10705_));
 sg13g2_a22oi_1 _17489_ (.Y(_10706_),
    .B1(_10703_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(_10702_),
    .A1(\cpu.ex.r_14[8] ));
 sg13g2_nor2b_1 _17490_ (.A(_10706_),
    .B_N(_10598_),
    .Y(_10707_));
 sg13g2_nor4_1 _17491_ (.A(_10697_),
    .B(_10700_),
    .C(_10705_),
    .D(_10707_),
    .Y(_10708_));
 sg13g2_buf_1 _17492_ (.A(net575),
    .X(_10709_));
 sg13g2_nor2_1 _17493_ (.A(\cpu.addr[8] ),
    .B(net524),
    .Y(_10710_));
 sg13g2_a21oi_1 _17494_ (.A1(net525),
    .A2(_10708_),
    .Y(_10711_),
    .B1(_10710_));
 sg13g2_mux2_1 _17495_ (.A0(_10681_),
    .A1(_10711_),
    .S(_10524_),
    .X(_10712_));
 sg13g2_buf_2 _17496_ (.A(_10712_),
    .X(_10713_));
 sg13g2_inv_1 _17497_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_10501_));
 sg13g2_nor2_1 _17498_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(\cpu.ex.c_mult_off[1] ),
    .Y(_10714_));
 sg13g2_inv_1 _17499_ (.Y(_10715_),
    .A(_10714_));
 sg13g2_a21oi_1 _17500_ (.A1(\cpu.ex.c_mult_off[3] ),
    .A2(_10713_),
    .Y(_10716_),
    .B1(_10715_));
 sg13g2_inv_1 _17501_ (.Y(_10717_),
    .A(\cpu.ex.c_mult_off[0] ));
 sg13g2_inv_1 _17502_ (.Y(_10718_),
    .A(_00292_));
 sg13g2_nor2_1 _17503_ (.A(_00290_),
    .B(_10501_),
    .Y(_10719_));
 sg13g2_a21oi_1 _17504_ (.A1(_10718_),
    .A2(_10501_),
    .Y(_10720_),
    .B1(_10719_));
 sg13g2_nor3_1 _17505_ (.A(_10532_),
    .B(net294),
    .C(_10720_),
    .Y(_10721_));
 sg13g2_mux2_1 _17506_ (.A0(\cpu.ex.r_12[9] ),
    .A1(\cpu.ex.r_14[9] ),
    .S(net854),
    .X(_10722_));
 sg13g2_nand3_1 _17507_ (.B(_10598_),
    .C(_10722_),
    .A(net653),
    .Y(_10723_));
 sg13g2_nand3_1 _17508_ (.B(_10616_),
    .C(net727),
    .A(\cpu.ex.r_9[9] ),
    .Y(_10724_));
 sg13g2_nor2b_1 _17509_ (.A(_00267_),
    .B_N(net728),
    .Y(_10725_));
 sg13g2_nor2b_1 _17510_ (.A(net728),
    .B_N(\cpu.ex.r_11[9] ),
    .Y(_10726_));
 sg13g2_o21ai_1 _17511_ (.B1(_10695_),
    .Y(_10727_),
    .A1(_10725_),
    .A2(_10726_));
 sg13g2_mux2_1 _17512_ (.A0(_10030_),
    .A1(\cpu.ex.r_epc[9] ),
    .S(net856),
    .X(_10728_));
 sg13g2_nand3_1 _17513_ (.B(net649),
    .C(_10728_),
    .A(net654),
    .Y(_10729_));
 sg13g2_nand4_1 _17514_ (.B(_10724_),
    .C(_10727_),
    .A(_10723_),
    .Y(_10730_),
    .D(_10729_));
 sg13g2_a22oi_1 _17515_ (.Y(_10731_),
    .B1(_10703_),
    .B2(\cpu.ex.r_lr[9] ),
    .A2(_10702_),
    .A1(\cpu.ex.r_mult[25] ));
 sg13g2_nor2_1 _17516_ (.A(_10602_),
    .B(_10731_),
    .Y(_10732_));
 sg13g2_buf_1 _17517_ (.A(_10560_),
    .X(_10733_));
 sg13g2_nand3_1 _17518_ (.B(\cpu.ex.r_10[9] ),
    .C(net648),
    .A(net647),
    .Y(_10734_));
 sg13g2_nand3_1 _17519_ (.B(\cpu.ex.r_13[9] ),
    .C(net727),
    .A(net653),
    .Y(_10735_));
 sg13g2_a21oi_1 _17520_ (.A1(_10734_),
    .A2(_10735_),
    .Y(_10736_),
    .B1(_10575_));
 sg13g2_nand3_1 _17521_ (.B(\cpu.ex.r_8[9] ),
    .C(net651),
    .A(net647),
    .Y(_10737_));
 sg13g2_nand3_1 _17522_ (.B(\cpu.ex.r_stmp[9] ),
    .C(_10665_),
    .A(net574),
    .Y(_10738_));
 sg13g2_a21oi_1 _17523_ (.A1(_10737_),
    .A2(_10738_),
    .Y(_10739_),
    .B1(net650));
 sg13g2_nor4_1 _17524_ (.A(_10730_),
    .B(_10732_),
    .C(_10736_),
    .D(_10739_),
    .Y(_10740_));
 sg13g2_nor2_1 _17525_ (.A(_09985_),
    .B(_10709_),
    .Y(_10741_));
 sg13g2_a21oi_2 _17526_ (.B1(_10741_),
    .Y(_10742_),
    .A2(_10740_),
    .A1(net525));
 sg13g2_nand2_1 _17527_ (.Y(_10743_),
    .A(_10501_),
    .B(_10742_));
 sg13g2_a22oi_1 _17528_ (.Y(_10744_),
    .B1(_10620_),
    .B2(\cpu.ex.r_mult[27] ),
    .A2(_10616_),
    .A1(\cpu.ex.r_11[11] ));
 sg13g2_inv_1 _17529_ (.Y(_10745_),
    .A(_10744_));
 sg13g2_inv_2 _17530_ (.Y(_10746_),
    .A(_10607_));
 sg13g2_inv_1 _17531_ (.Y(_10747_),
    .A(_00269_));
 sg13g2_and2_1 _17532_ (.A(net856),
    .B(net855),
    .X(_10748_));
 sg13g2_mux2_1 _17533_ (.A0(\cpu.ex.r_10[11] ),
    .A1(\cpu.ex.r_14[11] ),
    .S(_10556_),
    .X(_10749_));
 sg13g2_inv_1 _17534_ (.Y(_10750_),
    .A(net856));
 sg13g2_a22oi_1 _17535_ (.Y(_10751_),
    .B1(_10749_),
    .B2(_10750_),
    .A2(_10748_),
    .A1(_10747_));
 sg13g2_nand3_1 _17536_ (.B(\cpu.ex.r_13[11] ),
    .C(_10687_),
    .A(_10635_),
    .Y(_10752_));
 sg13g2_o21ai_1 _17537_ (.B1(_10752_),
    .Y(_10753_),
    .A1(_10746_),
    .A2(_10751_));
 sg13g2_mux2_1 _17538_ (.A0(\cpu.ex.r_8[11] ),
    .A1(\cpu.ex.r_12[11] ),
    .S(_10556_),
    .X(_10754_));
 sg13g2_nand3_1 _17539_ (.B(_10691_),
    .C(_10754_),
    .A(net733),
    .Y(_10755_));
 sg13g2_nand3_1 _17540_ (.B(net648),
    .C(_10620_),
    .A(\cpu.ex.r_stmp[11] ),
    .Y(_10756_));
 sg13g2_mux2_1 _17541_ (.A0(\cpu.ex.r_sp[11] ),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net856),
    .X(_10757_));
 sg13g2_nand3_1 _17542_ (.B(_10683_),
    .C(_10757_),
    .A(net729),
    .Y(_10758_));
 sg13g2_mux2_1 _17543_ (.A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_9[11] ),
    .S(net857),
    .X(_10759_));
 sg13g2_nand3_1 _17544_ (.B(net727),
    .C(_10759_),
    .A(net647),
    .Y(_10760_));
 sg13g2_nand4_1 _17545_ (.B(_10756_),
    .C(_10758_),
    .A(_10755_),
    .Y(_10761_),
    .D(_10760_));
 sg13g2_a221oi_1 _17546_ (.B2(_10547_),
    .C1(_10761_),
    .B1(_10753_),
    .A1(net652),
    .Y(_10762_),
    .A2(_10745_));
 sg13g2_nor2_1 _17547_ (.A(_10147_),
    .B(net575),
    .Y(_10763_));
 sg13g2_a21o_1 _17548_ (.A2(_10762_),
    .A1(net575),
    .B1(_10763_),
    .X(_10764_));
 sg13g2_buf_1 _17549_ (.A(_10764_),
    .X(_10765_));
 sg13g2_nand2b_1 _17550_ (.Y(_10766_),
    .B(\cpu.ex.c_mult_off[1] ),
    .A_N(_10765_));
 sg13g2_a21oi_1 _17551_ (.A1(_08615_),
    .A2(_10511_),
    .Y(_10767_),
    .B1(_10522_));
 sg13g2_buf_1 _17552_ (.A(_10767_),
    .X(_10768_));
 sg13g2_a221oi_1 _17553_ (.B2(_10766_),
    .C1(net363),
    .B1(_10743_),
    .A1(_09116_),
    .Y(_10769_),
    .A2(_10530_));
 sg13g2_inv_1 _17554_ (.Y(_10770_),
    .A(_00191_));
 sg13g2_buf_1 _17555_ (.A(_00200_),
    .X(_10771_));
 sg13g2_inv_1 _17556_ (.Y(_10772_),
    .A(_10771_));
 sg13g2_mux2_1 _17557_ (.A0(\cpu.ex.r_stmp[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net733),
    .X(_10773_));
 sg13g2_a22oi_1 _17558_ (.Y(_10774_),
    .B1(_10773_),
    .B2(net654),
    .A2(_10590_),
    .A1(net1096));
 sg13g2_nor2b_1 _17559_ (.A(_10774_),
    .B_N(_10582_),
    .Y(_10775_));
 sg13g2_inv_1 _17560_ (.Y(_10776_),
    .A(_00261_));
 sg13g2_a22oi_1 _17561_ (.Y(_10777_),
    .B1(net652),
    .B2(_10776_),
    .A2(_10691_),
    .A1(\cpu.ex.r_12[3] ));
 sg13g2_or2_1 _17562_ (.X(_10778_),
    .B(_10777_),
    .A(_10639_));
 sg13g2_a22oi_1 _17563_ (.Y(_10779_),
    .B1(_10553_),
    .B2(\cpu.ex.r_epc[3] ),
    .A2(_10551_),
    .A1(\cpu.ex.mmu_read[3] ));
 sg13g2_or2_1 _17564_ (.X(_10780_),
    .B(_10779_),
    .A(_10602_));
 sg13g2_buf_2 _17565_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10781_));
 sg13g2_a22oi_1 _17566_ (.Y(_10782_),
    .B1(_10685_),
    .B2(_10781_),
    .A2(_10578_),
    .A1(\cpu.ex.r_lr[3] ));
 sg13g2_nand2b_1 _17567_ (.Y(_10783_),
    .B(_10684_),
    .A_N(_10782_));
 sg13g2_nand3_1 _17568_ (.B(_10780_),
    .C(_10783_),
    .A(_10778_),
    .Y(_10784_));
 sg13g2_a22oi_1 _17569_ (.Y(_10785_),
    .B1(_10604_),
    .B2(\cpu.ex.r_mult[19] ),
    .A2(_10600_),
    .A1(\cpu.ex.r_10[3] ));
 sg13g2_nor2_1 _17570_ (.A(_10746_),
    .B(_10785_),
    .Y(_10786_));
 sg13g2_and2_1 _17571_ (.A(net857),
    .B(_10578_),
    .X(_10787_));
 sg13g2_buf_2 _17572_ (.A(_10787_),
    .X(_10788_));
 sg13g2_mux2_1 _17573_ (.A0(\cpu.ex.r_9[3] ),
    .A1(\cpu.ex.r_13[3] ),
    .S(net728),
    .X(_10789_));
 sg13g2_a22oi_1 _17574_ (.Y(_10790_),
    .B1(net652),
    .B2(\cpu.ex.r_11[3] ),
    .A2(_10691_),
    .A1(\cpu.ex.r_8[3] ));
 sg13g2_nor2b_1 _17575_ (.A(_10790_),
    .B_N(_10616_),
    .Y(_10791_));
 sg13g2_a21o_1 _17576_ (.A2(_10789_),
    .A1(_10788_),
    .B1(_10791_),
    .X(_10792_));
 sg13g2_nor4_2 _17577_ (.A(_10775_),
    .B(_10784_),
    .C(_10786_),
    .Y(_10793_),
    .D(_10792_));
 sg13g2_nor2_1 _17578_ (.A(_08944_),
    .B(net524),
    .Y(_10794_));
 sg13g2_a21oi_1 _17579_ (.A1(net525),
    .A2(_10793_),
    .Y(_10795_),
    .B1(_10794_));
 sg13g2_buf_1 _17580_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10796_));
 sg13g2_a22oi_1 _17581_ (.Y(_10797_),
    .B1(_10584_),
    .B2(\cpu.ex.r_lr[1] ),
    .A2(_10582_),
    .A1(_10796_));
 sg13g2_a22oi_1 _17582_ (.Y(_10798_),
    .B1(net648),
    .B2(\cpu.ex.r_stmp[1] ),
    .A2(net727),
    .A1(\cpu.ex.mmu_read[1] ));
 sg13g2_nand2b_1 _17583_ (.Y(_10799_),
    .B(net574),
    .A_N(_10798_));
 sg13g2_o21ai_1 _17584_ (.B1(_10799_),
    .Y(_10800_),
    .A1(net654),
    .A2(_10797_));
 sg13g2_nand2_1 _17585_ (.Y(_10801_),
    .A(\cpu.ex.r_9[1] ),
    .B(_10788_));
 sg13g2_mux2_1 _17586_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(net733),
    .X(_10802_));
 sg13g2_a21oi_1 _17587_ (.A1(net652),
    .A2(_10802_),
    .Y(_10803_),
    .B1(net574));
 sg13g2_nand2_1 _17588_ (.Y(_10804_),
    .A(_10801_),
    .B(_10803_));
 sg13g2_a21oi_1 _17589_ (.A1(\cpu.ex.r_mult[17] ),
    .A2(_10627_),
    .Y(_10805_),
    .B1(net647));
 sg13g2_and2_1 _17590_ (.A(net857),
    .B(_10691_),
    .X(_10806_));
 sg13g2_buf_1 _17591_ (.A(_10806_),
    .X(_10807_));
 sg13g2_nand2_1 _17592_ (.Y(_10808_),
    .A(\cpu.ex.r_12[1] ),
    .B(_10807_));
 sg13g2_nand2_1 _17593_ (.Y(_10809_),
    .A(_10805_),
    .B(_10808_));
 sg13g2_buf_1 _17594_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10810_));
 sg13g2_nand3_1 _17595_ (.B(net649),
    .C(net648),
    .A(_10810_),
    .Y(_10811_));
 sg13g2_nand3_1 _17596_ (.B(\cpu.ex.r_13[1] ),
    .C(_10788_),
    .A(net574),
    .Y(_10812_));
 sg13g2_mux2_1 _17597_ (.A0(\cpu.ex.r_8[1] ),
    .A1(\cpu.ex.r_10[1] ),
    .S(net729),
    .X(_10813_));
 sg13g2_and3_1 _17598_ (.X(_10814_),
    .A(net990),
    .B(_10544_),
    .C(net855));
 sg13g2_buf_2 _17599_ (.A(_10814_),
    .X(_10815_));
 sg13g2_inv_1 _17600_ (.Y(_10816_),
    .A(_00259_));
 sg13g2_mux2_1 _17601_ (.A0(\cpu.ex.r_14[1] ),
    .A1(_10816_),
    .S(net732),
    .X(_10817_));
 sg13g2_a22oi_1 _17602_ (.Y(_10818_),
    .B1(_10815_),
    .B2(_10817_),
    .A2(_10813_),
    .A1(_10600_));
 sg13g2_nand3_1 _17603_ (.B(_10812_),
    .C(_10818_),
    .A(_10811_),
    .Y(_10819_));
 sg13g2_a221oi_1 _17604_ (.B2(_10809_),
    .C1(_10819_),
    .B1(_10804_),
    .A1(_10575_),
    .Y(_10820_),
    .A2(_10800_));
 sg13g2_nor2_1 _17605_ (.A(_08962_),
    .B(net524),
    .Y(_10821_));
 sg13g2_a21oi_2 _17606_ (.B1(_10821_),
    .Y(_10822_),
    .A2(_10820_),
    .A1(net525));
 sg13g2_mux4_1 _17607_ (.S0(_10501_),
    .A0(_10770_),
    .A1(_10772_),
    .A2(_10795_),
    .A3(_10822_),
    .S1(net294),
    .X(_10823_));
 sg13g2_nor4_1 _17608_ (.A(_10717_),
    .B(_10721_),
    .C(_10769_),
    .D(_10823_),
    .Y(_10824_));
 sg13g2_a221oi_1 _17609_ (.B2(_10716_),
    .C1(_10824_),
    .B1(net293),
    .A1(_10502_),
    .Y(_10825_),
    .A2(_10649_));
 sg13g2_nor4_1 _17610_ (.A(_10717_),
    .B(_10532_),
    .C(_10721_),
    .D(_10769_),
    .Y(_10826_));
 sg13g2_nor3_1 _17611_ (.A(_10532_),
    .B(_10715_),
    .C(_10713_),
    .Y(_10827_));
 sg13g2_o21ai_1 _17612_ (.B1(\cpu.ex.r_mult_off[2] ),
    .Y(_10828_),
    .A1(_09105_),
    .A2(_09119_));
 sg13g2_nand3_1 _17613_ (.B(_10529_),
    .C(_10828_),
    .A(_09116_),
    .Y(_10829_));
 sg13g2_buf_1 _17614_ (.A(_10829_),
    .X(\cpu.ex.c_mult_off[2] ));
 sg13g2_nor3_1 _17615_ (.A(_10826_),
    .B(_10827_),
    .C(\cpu.ex.c_mult_off[2] ),
    .Y(_10830_));
 sg13g2_inv_1 _17616_ (.Y(_10831_),
    .A(_00195_));
 sg13g2_nand3_1 _17617_ (.B(\cpu.ex.r_14[14] ),
    .C(_10598_),
    .A(net574),
    .Y(_10832_));
 sg13g2_nand3_1 _17618_ (.B(\cpu.ex.r_epc[14] ),
    .C(_10684_),
    .A(net650),
    .Y(_10833_));
 sg13g2_a21oi_1 _17619_ (.A1(_10832_),
    .A2(_10833_),
    .Y(_10834_),
    .B1(_10746_));
 sg13g2_nor2_1 _17620_ (.A(net647),
    .B(_00272_),
    .Y(_10835_));
 sg13g2_a22oi_1 _17621_ (.Y(_10836_),
    .B1(_10835_),
    .B2(net652),
    .A2(_10565_),
    .A1(\cpu.ex.r_8[14] ));
 sg13g2_and2_1 _17622_ (.A(_10560_),
    .B(_10578_),
    .X(_10837_));
 sg13g2_nor2_1 _17623_ (.A(net731),
    .B(_10631_),
    .Y(_10838_));
 sg13g2_a221oi_1 _17624_ (.B2(\cpu.ex.r_stmp[14] ),
    .C1(net655),
    .B1(_10838_),
    .A1(\cpu.ex.r_lr[14] ),
    .Y(_10839_),
    .A2(_10837_));
 sg13g2_a21oi_1 _17625_ (.A1(net655),
    .A2(_10836_),
    .Y(_10840_),
    .B1(_10839_));
 sg13g2_and2_1 _17626_ (.A(_10616_),
    .B(_10573_),
    .X(_10841_));
 sg13g2_buf_1 _17627_ (.A(_10841_),
    .X(_10842_));
 sg13g2_nand2_1 _17628_ (.Y(_10843_),
    .A(\cpu.ex.r_10[14] ),
    .B(_10842_));
 sg13g2_mux2_1 _17629_ (.A0(\cpu.ex.r_12[14] ),
    .A1(\cpu.ex.r_13[14] ),
    .S(net732),
    .X(_10844_));
 sg13g2_nand3_1 _17630_ (.B(net651),
    .C(_10844_),
    .A(net574),
    .Y(_10845_));
 sg13g2_nand2_1 _17631_ (.Y(_10846_),
    .A(net729),
    .B(\cpu.ex.r_mult[30] ));
 sg13g2_o21ai_1 _17632_ (.B1(_10846_),
    .Y(_10847_),
    .A1(net654),
    .A2(_10241_));
 sg13g2_a22oi_1 _17633_ (.Y(_10848_),
    .B1(_10604_),
    .B2(_10847_),
    .A2(_10618_),
    .A1(\cpu.ex.r_9[14] ));
 sg13g2_and2_1 _17634_ (.A(net993),
    .B(_10545_),
    .X(_10849_));
 sg13g2_buf_1 _17635_ (.A(_10849_),
    .X(_10850_));
 sg13g2_nor2_2 _17636_ (.A(_10548_),
    .B(_10546_),
    .Y(_10851_));
 sg13g2_a22oi_1 _17637_ (.Y(_10852_),
    .B1(_10851_),
    .B2(_10250_),
    .A2(_10850_),
    .A1(\cpu.ex.r_11[14] ));
 sg13g2_nand2b_1 _17638_ (.Y(_10853_),
    .B(_10553_),
    .A_N(_10852_));
 sg13g2_nand4_1 _17639_ (.B(_10845_),
    .C(_10848_),
    .A(_10843_),
    .Y(_10854_),
    .D(_10853_));
 sg13g2_nor3_1 _17640_ (.A(_10834_),
    .B(_10840_),
    .C(_10854_),
    .Y(_10855_));
 sg13g2_nor2_1 _17641_ (.A(net578),
    .B(_10709_),
    .Y(_10856_));
 sg13g2_a21oi_1 _17642_ (.A1(net525),
    .A2(_10855_),
    .Y(_10857_),
    .B1(_10856_));
 sg13g2_mux2_1 _17643_ (.A0(_10831_),
    .A1(_10857_),
    .S(net336),
    .X(_10858_));
 sg13g2_buf_2 _17644_ (.A(_10858_),
    .X(_10859_));
 sg13g2_mux4_1 _17645_ (.S0(net647),
    .A0(\cpu.ex.r_14[12] ),
    .A1(\cpu.ex.r_10[12] ),
    .A2(_10318_),
    .A3(\cpu.ex.r_11[12] ),
    .S1(net650),
    .X(_10860_));
 sg13g2_nor2b_1 _17646_ (.A(net655),
    .B_N(\cpu.ex.r_stmp[12] ),
    .Y(_10861_));
 sg13g2_a22oi_1 _17647_ (.Y(_10862_),
    .B1(_10861_),
    .B2(_10582_),
    .A2(_10860_),
    .A1(net655));
 sg13g2_a22oi_1 _17648_ (.Y(_10863_),
    .B1(net651),
    .B2(\cpu.ex.r_8[12] ),
    .A2(_10665_),
    .A1(_10332_));
 sg13g2_mux2_1 _17649_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_epc[12] ),
    .S(net854),
    .X(_10864_));
 sg13g2_nand2b_1 _17650_ (.Y(_10865_),
    .B(_10864_),
    .A_N(_10602_));
 sg13g2_o21ai_1 _17651_ (.B1(_10865_),
    .Y(_10866_),
    .A1(net650),
    .A2(_10863_));
 sg13g2_a22oi_1 _17652_ (.Y(_10867_),
    .B1(net651),
    .B2(\cpu.ex.r_13[12] ),
    .A2(_10665_),
    .A1(\cpu.ex.r_mult[28] ));
 sg13g2_a22oi_1 _17653_ (.Y(_10868_),
    .B1(_10620_),
    .B2(_10317_),
    .A2(_10616_),
    .A1(\cpu.ex.r_9[12] ));
 sg13g2_or2_1 _17654_ (.X(_10869_),
    .B(_10868_),
    .A(net729));
 sg13g2_o21ai_1 _17655_ (.B1(_10869_),
    .Y(_10870_),
    .A1(net647),
    .A2(_10867_));
 sg13g2_and3_1 _17656_ (.X(_10871_),
    .A(\cpu.ex.r_12[12] ),
    .B(net651),
    .C(_10582_));
 sg13g2_a221oi_1 _17657_ (.B2(net650),
    .C1(_10871_),
    .B1(_10870_),
    .A1(_10733_),
    .Y(_10872_),
    .A2(_10866_));
 sg13g2_o21ai_1 _17658_ (.B1(_10872_),
    .Y(_10873_),
    .A1(_10746_),
    .A2(_10862_));
 sg13g2_mux2_1 _17659_ (.A0(net576),
    .A1(_10873_),
    .S(_10645_),
    .X(_10874_));
 sg13g2_nor2_1 _17660_ (.A(_00289_),
    .B(_10524_),
    .Y(_10875_));
 sg13g2_a21o_1 _17661_ (.A2(_10874_),
    .A1(net336),
    .B1(_10875_),
    .X(_10876_));
 sg13g2_buf_2 _17662_ (.A(_10876_),
    .X(_10877_));
 sg13g2_a22oi_1 _17663_ (.Y(_10878_),
    .B1(_10851_),
    .B2(_10209_),
    .A2(_10850_),
    .A1(\cpu.ex.r_11[15] ));
 sg13g2_nor2b_1 _17664_ (.A(_10878_),
    .B_N(_10553_),
    .Y(_10879_));
 sg13g2_a22oi_1 _17665_ (.Y(_10880_),
    .B1(_10634_),
    .B2(\cpu.ex.r_12[15] ),
    .A2(_10665_),
    .A1(\cpu.ex.r_stmp[15] ));
 sg13g2_nor2b_1 _17666_ (.A(_10880_),
    .B_N(_10582_),
    .Y(_10881_));
 sg13g2_nand3_1 _17667_ (.B(\cpu.ex.r_15[15] ),
    .C(_10815_),
    .A(_10549_),
    .Y(_10882_));
 sg13g2_nand3_1 _17668_ (.B(_10683_),
    .C(_10687_),
    .A(\cpu.ex.r_lr[15] ),
    .Y(_10883_));
 sg13g2_a22oi_1 _17669_ (.Y(_10884_),
    .B1(_10685_),
    .B2(\cpu.ex.r_14[15] ),
    .A2(_10578_),
    .A1(\cpu.ex.r_13[15] ));
 sg13g2_or2_1 _17670_ (.X(_10885_),
    .B(_10884_),
    .A(_10639_));
 sg13g2_nand4_1 _17671_ (.B(_10882_),
    .C(_10883_),
    .A(_10543_),
    .Y(_10886_),
    .D(_10885_));
 sg13g2_and2_1 _17672_ (.A(_10683_),
    .B(_10562_),
    .X(_10887_));
 sg13g2_buf_1 _17673_ (.A(_10887_),
    .X(_10888_));
 sg13g2_a22oi_1 _17674_ (.Y(_10889_),
    .B1(_10842_),
    .B2(\cpu.ex.r_10[15] ),
    .A2(_10888_),
    .A1(\cpu.ex.r_epc[15] ));
 sg13g2_and2_1 _17675_ (.A(net731),
    .B(_10587_),
    .X(_10890_));
 sg13g2_mux2_1 _17676_ (.A0(\cpu.ex.r_8[15] ),
    .A1(\cpu.ex.r_9[15] ),
    .S(net856),
    .X(_10891_));
 sg13g2_inv_2 _17677_ (.Y(_10892_),
    .A(_10220_));
 sg13g2_nand2_1 _17678_ (.Y(_10893_),
    .A(net854),
    .B(\cpu.ex.r_mult[31] ));
 sg13g2_o21ai_1 _17679_ (.B1(_10893_),
    .Y(_10894_),
    .A1(net729),
    .A2(_10892_));
 sg13g2_a22oi_1 _17680_ (.Y(_10895_),
    .B1(_10894_),
    .B2(_10604_),
    .A2(_10891_),
    .A1(_10890_));
 sg13g2_nand2_1 _17681_ (.Y(_10896_),
    .A(_10889_),
    .B(_10895_));
 sg13g2_or4_1 _17682_ (.A(_10879_),
    .B(_10881_),
    .C(_10886_),
    .D(_10896_),
    .X(_10897_));
 sg13g2_o21ai_1 _17683_ (.B1(_10897_),
    .Y(_10898_),
    .A1(net994),
    .A2(net524));
 sg13g2_nor2_1 _17684_ (.A(net363),
    .B(_10898_),
    .Y(_10899_));
 sg13g2_inv_1 _17685_ (.Y(_10900_),
    .A(_00194_));
 sg13g2_nand2_1 _17686_ (.Y(_10901_),
    .A(_10900_),
    .B(net363));
 sg13g2_nand2b_1 _17687_ (.Y(_10902_),
    .B(_10901_),
    .A_N(_10899_));
 sg13g2_buf_1 _17688_ (.A(_10902_),
    .X(_10903_));
 sg13g2_nand3_1 _17689_ (.B(\cpu.ex.r_epc[13] ),
    .C(_10683_),
    .A(net654),
    .Y(_10904_));
 sg13g2_nand3_1 _17690_ (.B(\cpu.ex.r_13[13] ),
    .C(net651),
    .A(net653),
    .Y(_10905_));
 sg13g2_nand2b_1 _17691_ (.Y(_10906_),
    .B(_10815_),
    .A_N(_00271_));
 sg13g2_nand3_1 _17692_ (.B(\cpu.ex.r_lr[13] ),
    .C(_10683_),
    .A(_10746_),
    .Y(_10907_));
 sg13g2_nand4_1 _17693_ (.B(_10905_),
    .C(_10906_),
    .A(_10904_),
    .Y(_10908_),
    .D(_10907_));
 sg13g2_and2_1 _17694_ (.A(net650),
    .B(_10908_),
    .X(_10909_));
 sg13g2_nand3_1 _17695_ (.B(_10287_),
    .C(net649),
    .A(net654),
    .Y(_10910_));
 sg13g2_nand3_1 _17696_ (.B(\cpu.ex.r_12[13] ),
    .C(net651),
    .A(net574),
    .Y(_10911_));
 sg13g2_a21oi_1 _17697_ (.A1(_10910_),
    .A2(_10911_),
    .Y(_10912_),
    .B1(_10662_));
 sg13g2_a22oi_1 _17698_ (.Y(_10913_),
    .B1(_10584_),
    .B2(\cpu.ex.r_11[13] ),
    .A2(_10582_),
    .A1(\cpu.ex.r_14[13] ));
 sg13g2_nand2b_1 _17699_ (.Y(_10914_),
    .B(_10592_),
    .A_N(_10913_));
 sg13g2_a22oi_1 _17700_ (.Y(_10915_),
    .B1(_10622_),
    .B2(\cpu.ex.r_stmp[13] ),
    .A2(_10618_),
    .A1(\cpu.ex.r_9[13] ));
 sg13g2_nand2_1 _17701_ (.Y(_10916_),
    .A(_10914_),
    .B(_10915_));
 sg13g2_a22oi_1 _17702_ (.Y(_10917_),
    .B1(_10604_),
    .B2(\cpu.ex.r_mult[29] ),
    .A2(_10600_),
    .A1(\cpu.ex.r_10[13] ));
 sg13g2_a221oi_1 _17703_ (.B2(\cpu.ex.mmu_read[13] ),
    .C1(_10608_),
    .B1(_10604_),
    .A1(\cpu.ex.r_8[13] ),
    .Y(_10918_),
    .A2(_10600_));
 sg13g2_a21oi_1 _17704_ (.A1(_10608_),
    .A2(_10917_),
    .Y(_10919_),
    .B1(_10918_));
 sg13g2_nor4_1 _17705_ (.A(_10909_),
    .B(_10912_),
    .C(_10916_),
    .D(_10919_),
    .Y(_10920_));
 sg13g2_nor2_1 _17706_ (.A(net577),
    .B(net525),
    .Y(_10921_));
 sg13g2_a21oi_1 _17707_ (.A1(net525),
    .A2(_10920_),
    .Y(_10922_),
    .B1(_10921_));
 sg13g2_nor2_1 _17708_ (.A(_00196_),
    .B(net336),
    .Y(_10923_));
 sg13g2_a21o_1 _17709_ (.A2(_10922_),
    .A1(net336),
    .B1(_10923_),
    .X(_10924_));
 sg13g2_buf_1 _17710_ (.A(_10924_),
    .X(_10925_));
 sg13g2_mux4_1 _17711_ (.S0(_10501_),
    .A0(_10859_),
    .A1(_10877_),
    .A2(net239),
    .A3(_10925_),
    .S1(\cpu.ex.c_mult_off[0] ),
    .X(_10926_));
 sg13g2_and2_1 _17712_ (.A(\cpu.ex.c_mult_off[3] ),
    .B(\cpu.ex.c_mult_off[2] ),
    .X(_10927_));
 sg13g2_and2_1 _17713_ (.A(_10532_),
    .B(\cpu.ex.c_mult_off[2] ),
    .X(_10928_));
 sg13g2_inv_1 _17714_ (.Y(_10929_),
    .A(_00296_));
 sg13g2_a22oi_1 _17715_ (.Y(_10930_),
    .B1(net648),
    .B2(_10436_),
    .A2(net727),
    .A1(\cpu.ex.r_lr[5] ));
 sg13g2_nand2b_1 _17716_ (.Y(_10931_),
    .B(net649),
    .A_N(_10930_));
 sg13g2_a22oi_1 _17717_ (.Y(_10932_),
    .B1(_10553_),
    .B2(\cpu.ex.r_11[5] ),
    .A2(_10551_),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_nor2b_1 _17718_ (.A(_10932_),
    .B_N(_10850_),
    .Y(_10933_));
 sg13g2_a221oi_1 _17719_ (.B2(\cpu.ex.r_epc[5] ),
    .C1(_10933_),
    .B1(_10888_),
    .A1(\cpu.ex.r_stmp[5] ),
    .Y(_10934_),
    .A2(_10622_));
 sg13g2_a22oi_1 _17720_ (.Y(_10935_),
    .B1(_10838_),
    .B2(\cpu.ex.r_14[5] ),
    .A2(_10837_),
    .A1(\cpu.ex.r_9[5] ));
 sg13g2_nand2b_1 _17721_ (.Y(_10936_),
    .B(net655),
    .A_N(_10935_));
 sg13g2_mux2_1 _17722_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_12[5] ),
    .S(net728),
    .X(_10937_));
 sg13g2_mux2_1 _17723_ (.A0(_10444_),
    .A1(\cpu.ex.r_mult[21] ),
    .S(_10575_),
    .X(_10938_));
 sg13g2_and3_1 _17724_ (.X(_10939_),
    .A(net653),
    .B(net652),
    .C(_10938_));
 sg13g2_a221oi_1 _17725_ (.B2(_10807_),
    .C1(_10939_),
    .B1(_10937_),
    .A1(\cpu.ex.r_10[5] ),
    .Y(_10940_),
    .A2(_10842_));
 sg13g2_nand4_1 _17726_ (.B(_10934_),
    .C(_10936_),
    .A(_10931_),
    .Y(_10941_),
    .D(_10940_));
 sg13g2_mux2_1 _17727_ (.A0(_09732_),
    .A1(_10941_),
    .S(net524),
    .X(_10942_));
 sg13g2_mux2_1 _17728_ (.A0(_10929_),
    .A1(_10942_),
    .S(net336),
    .X(_10943_));
 sg13g2_buf_1 _17729_ (.A(_10943_),
    .X(_10944_));
 sg13g2_inv_1 _17730_ (.Y(_10945_),
    .A(_00294_));
 sg13g2_mux2_1 _17731_ (.A0(\cpu.ex.r_stmp[7] ),
    .A1(\cpu.ex.r_mult[23] ),
    .S(net732),
    .X(_10946_));
 sg13g2_and2_1 _17732_ (.A(net654),
    .B(_10620_),
    .X(_10947_));
 sg13g2_a22oi_1 _17733_ (.Y(_10948_),
    .B1(_10946_),
    .B2(_10947_),
    .A2(_10842_),
    .A1(\cpu.ex.r_10[7] ));
 sg13g2_and2_1 _17734_ (.A(net647),
    .B(net652),
    .X(_10949_));
 sg13g2_mux2_1 _17735_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(\cpu.ex.r_11[7] ),
    .S(net733),
    .X(_10950_));
 sg13g2_mux2_1 _17736_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_12[7] ),
    .S(net653),
    .X(_10951_));
 sg13g2_a22oi_1 _17737_ (.Y(_10952_),
    .B1(_10951_),
    .B2(_10807_),
    .A2(_10950_),
    .A1(_10949_));
 sg13g2_a22oi_1 _17738_ (.Y(_10953_),
    .B1(_10851_),
    .B2(_10388_),
    .A2(_10850_),
    .A1(\cpu.ex.r_13[7] ));
 sg13g2_nand2b_1 _17739_ (.Y(_10954_),
    .B(_10551_),
    .A_N(_10953_));
 sg13g2_mux2_1 _17740_ (.A0(\cpu.ex.r_14[7] ),
    .A1(_10377_),
    .S(net732),
    .X(_10955_));
 sg13g2_a22oi_1 _17741_ (.Y(_10956_),
    .B1(net648),
    .B2(_10390_),
    .A2(net727),
    .A1(\cpu.ex.r_lr[7] ));
 sg13g2_nor2b_1 _17742_ (.A(_10956_),
    .B_N(net649),
    .Y(_10957_));
 sg13g2_a221oi_1 _17743_ (.B2(_10955_),
    .C1(_10957_),
    .B1(_10815_),
    .A1(\cpu.ex.r_9[7] ),
    .Y(_10958_),
    .A2(_10618_));
 sg13g2_nand4_1 _17744_ (.B(_10952_),
    .C(_10954_),
    .A(_10948_),
    .Y(_10959_),
    .D(_10958_));
 sg13g2_mux2_1 _17745_ (.A0(_08952_),
    .A1(_10959_),
    .S(net524),
    .X(_10960_));
 sg13g2_mux2_1 _17746_ (.A0(_10945_),
    .A1(_10960_),
    .S(_10524_),
    .X(_10961_));
 sg13g2_buf_2 _17747_ (.A(_10961_),
    .X(_10962_));
 sg13g2_a22oi_1 _17748_ (.Y(_10963_),
    .B1(_10703_),
    .B2(\cpu.ex.r_lr[4] ),
    .A2(_10702_),
    .A1(\cpu.ex.r_mult[20] ));
 sg13g2_nor2_1 _17749_ (.A(_10602_),
    .B(_10963_),
    .Y(_10964_));
 sg13g2_mux2_1 _17750_ (.A0(_08516_),
    .A1(\cpu.ex.r_12[4] ),
    .S(net733),
    .X(_10965_));
 sg13g2_nand3_1 _17751_ (.B(_10691_),
    .C(_10965_),
    .A(net653),
    .Y(_10966_));
 sg13g2_mux2_1 _17752_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(\cpu.ex.r_11[4] ),
    .S(net733),
    .X(_10967_));
 sg13g2_nand2_1 _17753_ (.Y(_10968_),
    .A(_10949_),
    .B(_10967_));
 sg13g2_mux2_1 _17754_ (.A0(\cpu.ex.r_14[4] ),
    .A1(_10462_),
    .S(net856),
    .X(_10969_));
 sg13g2_mux2_1 _17755_ (.A0(\cpu.ex.r_8[4] ),
    .A1(\cpu.ex.r_10[4] ),
    .S(net854),
    .X(_10970_));
 sg13g2_a22oi_1 _17756_ (.Y(_10971_),
    .B1(_10970_),
    .B2(_10600_),
    .A2(_10969_),
    .A1(_10815_));
 sg13g2_nand3_1 _17757_ (.B(_10968_),
    .C(_10971_),
    .A(_10966_),
    .Y(_10972_));
 sg13g2_nor2_1 _17758_ (.A(net733),
    .B(_10631_),
    .Y(_10973_));
 sg13g2_a22oi_1 _17759_ (.Y(_10974_),
    .B1(_10973_),
    .B2(\cpu.ex.r_stmp[4] ),
    .A2(_10788_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_a221oi_1 _17760_ (.B2(_10474_),
    .C1(net653),
    .B1(_10973_),
    .A1(\cpu.ex.r_9[4] ),
    .Y(_10975_),
    .A2(_10788_));
 sg13g2_a21oi_1 _17761_ (.A1(net574),
    .A2(_10974_),
    .Y(_10976_),
    .B1(_10975_));
 sg13g2_nor3_1 _17762_ (.A(_10964_),
    .B(_10972_),
    .C(_10976_),
    .Y(_10977_));
 sg13g2_nor2_1 _17763_ (.A(_09149_),
    .B(net575),
    .Y(_10978_));
 sg13g2_a21oi_1 _17764_ (.A1(net524),
    .A2(_10977_),
    .Y(_10979_),
    .B1(_10978_));
 sg13g2_mux2_1 _17765_ (.A0(_08105_),
    .A1(_10979_),
    .S(_10524_),
    .X(_10980_));
 sg13g2_buf_2 _17766_ (.A(_10980_),
    .X(_10981_));
 sg13g2_inv_1 _17767_ (.Y(_10982_),
    .A(_00295_));
 sg13g2_nand2_1 _17768_ (.Y(_10983_),
    .A(\cpu.ex.r_10[6] ),
    .B(_10842_));
 sg13g2_mux2_1 _17769_ (.A0(\cpu.ex.r_14[6] ),
    .A1(_10404_),
    .S(net856),
    .X(_10984_));
 sg13g2_nand2_1 _17770_ (.Y(_10985_),
    .A(_10815_),
    .B(_10984_));
 sg13g2_and2_1 _17771_ (.A(_10562_),
    .B(_10620_),
    .X(_10986_));
 sg13g2_a22oi_1 _17772_ (.Y(_10987_),
    .B1(_10986_),
    .B2(_10415_),
    .A2(_10622_),
    .A1(\cpu.ex.r_stmp[6] ));
 sg13g2_mux2_1 _17773_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_12[6] ),
    .S(net730),
    .X(_10988_));
 sg13g2_nand2_1 _17774_ (.Y(_10989_),
    .A(_10807_),
    .B(_10988_));
 sg13g2_and4_1 _17775_ (.A(_10983_),
    .B(_10985_),
    .C(_10987_),
    .D(_10989_),
    .X(_10990_));
 sg13g2_a22oi_1 _17776_ (.Y(_10991_),
    .B1(net648),
    .B2(_10421_),
    .A2(net727),
    .A1(\cpu.ex.r_lr[6] ));
 sg13g2_nand2b_1 _17777_ (.Y(_10992_),
    .B(net649),
    .A_N(_10991_));
 sg13g2_a22oi_1 _17778_ (.Y(_10993_),
    .B1(_10888_),
    .B2(\cpu.ex.r_epc[6] ),
    .A2(_10618_),
    .A1(\cpu.ex.r_9[6] ));
 sg13g2_a22oi_1 _17779_ (.Y(_10994_),
    .B1(_10553_),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10551_),
    .A1(\cpu.ex.r_13[6] ));
 sg13g2_nand2b_1 _17780_ (.Y(_10995_),
    .B(_10850_),
    .A_N(_10994_));
 sg13g2_nand4_1 _17781_ (.B(_10992_),
    .C(_10993_),
    .A(_10990_),
    .Y(_10996_),
    .D(_10995_));
 sg13g2_mux2_1 _17782_ (.A0(_08948_),
    .A1(_10996_),
    .S(net524),
    .X(_10997_));
 sg13g2_mux2_1 _17783_ (.A0(_10982_),
    .A1(_10997_),
    .S(_10524_),
    .X(_10998_));
 sg13g2_buf_2 _17784_ (.A(_10998_),
    .X(_10999_));
 sg13g2_mux4_1 _17785_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(_10944_),
    .A1(_10962_),
    .A2(_10981_),
    .A3(_10999_),
    .S1(_10717_),
    .X(_11000_));
 sg13g2_and2_1 _17786_ (.A(_10928_),
    .B(_11000_),
    .X(_11001_));
 sg13g2_a221oi_1 _17787_ (.B2(_10927_),
    .C1(_11001_),
    .B1(_10926_),
    .A1(_10825_),
    .Y(_11002_),
    .A2(_10830_));
 sg13g2_buf_8 _17788_ (.A(_11002_),
    .X(_11003_));
 sg13g2_nand2_1 _17789_ (.Y(_11004_),
    .A(\cpu.ex.r_9[0] ),
    .B(_10407_));
 sg13g2_nand3_1 _17790_ (.B(net865),
    .C(net997),
    .A(\cpu.ex.r_15[0] ),
    .Y(_11005_));
 sg13g2_a21oi_1 _17791_ (.A1(_11004_),
    .A2(_11005_),
    .Y(_11006_),
    .B1(_10440_));
 sg13g2_a22oi_1 _17792_ (.Y(_11007_),
    .B1(_10019_),
    .B2(\cpu.ex.r_stmp[0] ),
    .A2(_10129_),
    .A1(\cpu.ex.r_12[0] ));
 sg13g2_nor2b_1 _17793_ (.A(_11007_),
    .B_N(net737),
    .Y(_11008_));
 sg13g2_a221oi_1 _17794_ (.B2(\cpu.ex.r_mult[16] ),
    .C1(net859),
    .B1(_10215_),
    .A1(_09007_),
    .Y(_11009_),
    .A2(_10005_));
 sg13g2_a221oi_1 _17795_ (.B2(\cpu.ex.r_14[0] ),
    .C1(net860),
    .B1(_10082_),
    .A1(\cpu.ex.r_13[0] ),
    .Y(_11010_),
    .A2(net861));
 sg13g2_nor3_1 _17796_ (.A(_10052_),
    .B(_11009_),
    .C(_11010_),
    .Y(_11011_));
 sg13g2_mux2_1 _17797_ (.A0(_10659_),
    .A1(\cpu.ex.r_11[0] ),
    .S(net998),
    .X(_11012_));
 sg13g2_nand3_1 _17798_ (.B(net865),
    .C(_11012_),
    .A(_10037_),
    .Y(_11013_));
 sg13g2_mux2_1 _17799_ (.A0(\cpu.ex.r_8[0] ),
    .A1(\cpu.ex.r_10[0] ),
    .S(net1000),
    .X(_11014_));
 sg13g2_nand3_1 _17800_ (.B(_10097_),
    .C(_11014_),
    .A(_10026_),
    .Y(_11015_));
 sg13g2_a21oi_1 _17801_ (.A1(_11013_),
    .A2(_11015_),
    .Y(_11016_),
    .B1(net864));
 sg13g2_or4_1 _17802_ (.A(_11006_),
    .B(_11008_),
    .C(_11011_),
    .D(_11016_),
    .X(_11017_));
 sg13g2_a22oi_1 _17803_ (.Y(_11018_),
    .B1(_10008_),
    .B2(_11017_),
    .A2(net580),
    .A1(_08588_));
 sg13g2_buf_1 _17804_ (.A(_11018_),
    .X(_11019_));
 sg13g2_nor2_1 _17805_ (.A(_10122_),
    .B(_09979_),
    .Y(_11020_));
 sg13g2_buf_1 _17806_ (.A(\cpu.dec.imm[0] ),
    .X(_11021_));
 sg13g2_nor3_1 _17807_ (.A(_11021_),
    .B(_09982_),
    .C(_09979_),
    .Y(_11022_));
 sg13g2_or2_1 _17808_ (.X(_11023_),
    .B(_11022_),
    .A(net1002));
 sg13g2_a21o_1 _17809_ (.A2(_11020_),
    .A1(_11019_),
    .B1(_11023_),
    .X(_11024_));
 sg13g2_buf_1 _17810_ (.A(_11024_),
    .X(_11025_));
 sg13g2_inv_1 _17811_ (.Y(_11026_),
    .A(_00309_));
 sg13g2_a22oi_1 _17812_ (.Y(_11027_),
    .B1(_10423_),
    .B2(_10816_),
    .A2(_10387_),
    .A1(\cpu.ex.r_stmp[1] ));
 sg13g2_nand2b_1 _17813_ (.Y(_11028_),
    .B(net657),
    .A_N(_11027_));
 sg13g2_mux2_1 _17814_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(_10034_),
    .X(_11029_));
 sg13g2_a22oi_1 _17815_ (.Y(_11030_),
    .B1(_11029_),
    .B2(_10038_),
    .A2(_10005_),
    .A1(_10796_));
 sg13g2_or2_1 _17816_ (.X(_11031_),
    .B(_11030_),
    .A(net736));
 sg13g2_a21oi_1 _17817_ (.A1(_11028_),
    .A2(_11031_),
    .Y(_11032_),
    .B1(net738));
 sg13g2_nand3_1 _17818_ (.B(_10026_),
    .C(_10043_),
    .A(\cpu.ex.r_14[1] ),
    .Y(_11033_));
 sg13g2_nand3_1 _17819_ (.B(net862),
    .C(net866),
    .A(\cpu.ex.r_epc[1] ),
    .Y(_11034_));
 sg13g2_a21oi_1 _17820_ (.A1(_11033_),
    .A2(_11034_),
    .Y(_11035_),
    .B1(_10011_));
 sg13g2_nand3_1 _17821_ (.B(net740),
    .C(net866),
    .A(\cpu.ex.r_lr[1] ),
    .Y(_11036_));
 sg13g2_nand3_1 _17822_ (.B(_10026_),
    .C(_10043_),
    .A(\cpu.ex.r_12[1] ),
    .Y(_11037_));
 sg13g2_a21oi_1 _17823_ (.A1(_11036_),
    .A2(_11037_),
    .Y(_11038_),
    .B1(_10035_));
 sg13g2_a22oi_1 _17824_ (.Y(_11039_),
    .B1(_10257_),
    .B2(\cpu.ex.r_11[1] ),
    .A2(_10254_),
    .A1(\cpu.ex.r_13[1] ));
 sg13g2_nor2_1 _17825_ (.A(_10440_),
    .B(_11039_),
    .Y(_11040_));
 sg13g2_mux2_1 _17826_ (.A0(\cpu.ex.r_8[1] ),
    .A1(\cpu.ex.r_9[1] ),
    .S(net996),
    .X(_11041_));
 sg13g2_mux2_1 _17827_ (.A0(_10810_),
    .A1(\cpu.ex.r_10[1] ),
    .S(net859),
    .X(_11042_));
 sg13g2_a22oi_1 _17828_ (.Y(_11043_),
    .B1(_11042_),
    .B2(_10082_),
    .A2(_11041_),
    .A1(_10129_));
 sg13g2_nor2_1 _17829_ (.A(net734),
    .B(_11043_),
    .Y(_11044_));
 sg13g2_or4_1 _17830_ (.A(_11035_),
    .B(_11038_),
    .C(_11040_),
    .D(_11044_),
    .X(_11045_));
 sg13g2_nor2_1 _17831_ (.A(net858),
    .B(_10124_),
    .Y(_11046_));
 sg13g2_o21ai_1 _17832_ (.B1(_11046_),
    .Y(_11047_),
    .A1(_11032_),
    .A2(_11045_));
 sg13g2_buf_1 _17833_ (.A(\cpu.dec.imm[1] ),
    .X(_11048_));
 sg13g2_nor2_1 _17834_ (.A(_09727_),
    .B(_10121_),
    .Y(_11049_));
 sg13g2_a221oi_1 _17835_ (.B2(_11049_),
    .C1(_10106_),
    .B1(_10000_),
    .A1(_11048_),
    .Y(_11050_),
    .A2(_10122_));
 sg13g2_buf_1 _17836_ (.A(_11050_),
    .X(_11051_));
 sg13g2_nor2b_1 _17837_ (.A(net1089),
    .B_N(net1002),
    .Y(_11052_));
 sg13g2_a21o_1 _17838_ (.A2(_11051_),
    .A1(_11047_),
    .B1(_11052_),
    .X(_11053_));
 sg13g2_buf_1 _17839_ (.A(_11053_),
    .X(_11054_));
 sg13g2_buf_1 _17840_ (.A(_11054_),
    .X(_11055_));
 sg13g2_mux2_1 _17841_ (.A0(\cpu.ex.r_12[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net863),
    .X(_11056_));
 sg13g2_a22oi_1 _17842_ (.Y(_11057_),
    .B1(_11056_),
    .B2(net737),
    .A2(_10405_),
    .A1(_10568_));
 sg13g2_nand3_1 _17843_ (.B(_10027_),
    .C(_10407_),
    .A(\cpu.ex.r_8[2] ),
    .Y(_11058_));
 sg13g2_a21oi_1 _17844_ (.A1(_11057_),
    .A2(_11058_),
    .Y(_11059_),
    .B1(net860));
 sg13g2_inv_1 _17845_ (.Y(_11060_),
    .A(\cpu.ex.r_10[2] ));
 sg13g2_nand3b_1 _17846_ (.B(_10021_),
    .C(\cpu.ex.r_stmp[2] ),
    .Y(_11061_),
    .A_N(_10077_));
 sg13g2_o21ai_1 _17847_ (.B1(_11061_),
    .Y(_11062_),
    .A1(_11060_),
    .A2(_10172_));
 sg13g2_nand3b_1 _17848_ (.B(net865),
    .C(_10554_),
    .Y(_11063_),
    .A_N(net997));
 sg13g2_nand3b_1 _17849_ (.B(_10021_),
    .C(_08081_),
    .Y(_11064_),
    .A_N(_10034_));
 sg13g2_or2_1 _17850_ (.X(_11065_),
    .B(net859),
    .A(net862));
 sg13g2_a21oi_1 _17851_ (.A1(_11063_),
    .A2(_11064_),
    .Y(_11066_),
    .B1(_11065_));
 sg13g2_a21o_1 _17852_ (.A2(_11062_),
    .A1(net660),
    .B1(_11066_),
    .X(_11067_));
 sg13g2_o21ai_1 _17853_ (.B1(_10008_),
    .Y(_11068_),
    .A1(_11059_),
    .A2(_11067_));
 sg13g2_mux4_1 _17854_ (.S0(net863),
    .A0(\cpu.ex.r_lr[2] ),
    .A1(\cpu.ex.r_epc[2] ),
    .A2(_10576_),
    .A3(\cpu.ex.r_mult[18] ),
    .S1(net997),
    .X(_11069_));
 sg13g2_nor2_1 _17855_ (.A(net736),
    .B(_11069_),
    .Y(_11070_));
 sg13g2_mux2_1 _17856_ (.A0(\cpu.ex.r_9[2] ),
    .A1(\cpu.ex.r_13[2] ),
    .S(_10013_),
    .X(_11071_));
 sg13g2_a221oi_1 _17857_ (.B2(_10011_),
    .C1(_10058_),
    .B1(_11071_),
    .A1(\cpu.ex.r_11[2] ),
    .Y(_11072_),
    .A2(_10257_));
 sg13g2_nor3_1 _17858_ (.A(net742),
    .B(_11070_),
    .C(_11072_),
    .Y(_11073_));
 sg13g2_a22oi_1 _17859_ (.Y(_11074_),
    .B1(_10008_),
    .B2(_11073_),
    .A2(net580),
    .A1(_08959_));
 sg13g2_nor3_2 _17860_ (.A(_10121_),
    .B(_09976_),
    .C(_09979_),
    .Y(_11075_));
 sg13g2_nand3_1 _17861_ (.B(_11074_),
    .C(_11075_),
    .A(_11068_),
    .Y(_11076_));
 sg13g2_buf_1 _17862_ (.A(_11076_),
    .X(_11077_));
 sg13g2_buf_1 _17863_ (.A(\cpu.dec.imm[2] ),
    .X(_11078_));
 sg13g2_nor2_1 _17864_ (.A(_11078_),
    .B(_09982_),
    .Y(_11079_));
 sg13g2_a22oi_1 _17865_ (.Y(_11080_),
    .B1(_09981_),
    .B2(_11079_),
    .A2(net1002),
    .A1(_08123_));
 sg13g2_buf_1 _17866_ (.A(_11080_),
    .X(_11081_));
 sg13g2_nand2_1 _17867_ (.Y(_11082_),
    .A(_11077_),
    .B(_11081_));
 sg13g2_buf_1 _17868_ (.A(_11082_),
    .X(_11083_));
 sg13g2_inv_1 _17869_ (.Y(_11084_),
    .A(_00308_));
 sg13g2_a22oi_1 _17870_ (.Y(_11085_),
    .B1(net333),
    .B2(_11084_),
    .A2(net334),
    .A1(_11026_));
 sg13g2_nor2_1 _17871_ (.A(_09115_),
    .B(_11085_),
    .Y(_11086_));
 sg13g2_a22oi_1 _17872_ (.Y(_11087_),
    .B1(_10072_),
    .B2(\cpu.ex.r_epc[3] ),
    .A2(_10070_),
    .A1(\cpu.ex.r_stmp[3] ));
 sg13g2_inv_1 _17873_ (.Y(_11088_),
    .A(_11087_));
 sg13g2_nor2_1 _17874_ (.A(\cpu.ex.r_13[3] ),
    .B(net865),
    .Y(_11089_));
 sg13g2_a21oi_1 _17875_ (.A1(_00261_),
    .A2(_10010_),
    .Y(_11090_),
    .B1(_11089_));
 sg13g2_mux2_1 _17876_ (.A0(\cpu.ex.r_8[3] ),
    .A1(\cpu.ex.r_10[3] ),
    .S(net863),
    .X(_11091_));
 sg13g2_and2_1 _17877_ (.A(_10032_),
    .B(_11091_),
    .X(_11092_));
 sg13g2_a21o_1 _17878_ (.A2(_11090_),
    .A1(_10075_),
    .B1(_11092_),
    .X(_11093_));
 sg13g2_a22oi_1 _17879_ (.Y(_11094_),
    .B1(_11093_),
    .B2(net656),
    .A2(_11088_),
    .A1(net663));
 sg13g2_inv_2 _17880_ (.Y(_11095_),
    .A(\cpu.ex.mmu_read[3] ));
 sg13g2_nand2_1 _17881_ (.Y(_11096_),
    .A(_10011_),
    .B(_10094_));
 sg13g2_nand3_1 _17882_ (.B(net741),
    .C(_10015_),
    .A(\cpu.ex.r_11[3] ),
    .Y(_11097_));
 sg13g2_o21ai_1 _17883_ (.B1(_11097_),
    .Y(_11098_),
    .A1(_11095_),
    .A2(_11096_));
 sg13g2_nand2_1 _17884_ (.Y(_11099_),
    .A(\cpu.ex.r_lr[3] ),
    .B(_10407_));
 sg13g2_nand3_1 _17885_ (.B(net741),
    .C(net864),
    .A(\cpu.ex.r_mult[19] ),
    .Y(_11100_));
 sg13g2_a21oi_1 _17886_ (.A1(_11099_),
    .A2(_11100_),
    .Y(_11101_),
    .B1(_10097_));
 sg13g2_o21ai_1 _17887_ (.B1(net661),
    .Y(_11102_),
    .A1(_11098_),
    .A2(_11101_));
 sg13g2_a21oi_1 _17888_ (.A1(_11094_),
    .A2(_11102_),
    .Y(_11103_),
    .B1(_10124_));
 sg13g2_a22oi_1 _17889_ (.Y(_11104_),
    .B1(_10203_),
    .B2(_10781_),
    .A2(_10201_),
    .A1(\cpu.ex.r_9[3] ));
 sg13g2_mux2_1 _17890_ (.A0(net1096),
    .A1(\cpu.ex.r_12[3] ),
    .S(_10077_),
    .X(_11105_));
 sg13g2_a22oi_1 _17891_ (.Y(_11106_),
    .B1(_11105_),
    .B2(_10011_),
    .A2(_10305_),
    .A1(\cpu.ex.r_14[3] ));
 sg13g2_nand2b_1 _17892_ (.Y(_11107_),
    .B(net737),
    .A_N(_11106_));
 sg13g2_o21ai_1 _17893_ (.B1(_11107_),
    .Y(_11108_),
    .A1(net734),
    .A2(_11104_));
 sg13g2_a22oi_1 _17894_ (.Y(_11109_),
    .B1(_10008_),
    .B2(_11108_),
    .A2(net580),
    .A1(_08944_));
 sg13g2_nand3b_1 _17895_ (.B(_11109_),
    .C(_11075_),
    .Y(_11110_),
    .A_N(_11103_));
 sg13g2_buf_2 _17896_ (.A(_11110_),
    .X(_11111_));
 sg13g2_buf_1 _17897_ (.A(\cpu.dec.imm[3] ),
    .X(_11112_));
 sg13g2_nor2_1 _17898_ (.A(_11112_),
    .B(_09983_),
    .Y(_11113_));
 sg13g2_a22oi_1 _17899_ (.Y(_11114_),
    .B1(_09981_),
    .B2(_11113_),
    .A2(net1002),
    .A1(_08090_));
 sg13g2_buf_1 _17900_ (.A(_11114_),
    .X(_11115_));
 sg13g2_and2_1 _17901_ (.A(_11111_),
    .B(_11115_),
    .X(_11116_));
 sg13g2_buf_1 _17902_ (.A(_11116_),
    .X(_11117_));
 sg13g2_buf_2 _17903_ (.A(_00307_),
    .X(_11118_));
 sg13g2_nand2b_1 _17904_ (.Y(_11119_),
    .B(_10281_),
    .A_N(_11118_));
 sg13g2_nor2_1 _17905_ (.A(_11117_),
    .B(_11119_),
    .Y(_11120_));
 sg13g2_nor3_1 _17906_ (.A(net335),
    .B(_11086_),
    .C(_11120_),
    .Y(_11121_));
 sg13g2_a21oi_1 _17907_ (.A1(_10120_),
    .A2(_10484_),
    .Y(_11122_),
    .B1(_10485_));
 sg13g2_buf_2 _17908_ (.A(_11122_),
    .X(_11123_));
 sg13g2_nand2b_1 _17909_ (.Y(_11124_),
    .B(_10281_),
    .A_N(_10461_));
 sg13g2_a22oi_1 _17910_ (.Y(_11125_),
    .B1(net295),
    .B2(_10489_),
    .A2(_11124_),
    .A1(_11123_));
 sg13g2_a21oi_1 _17911_ (.A1(_10455_),
    .A2(_10457_),
    .Y(_11126_),
    .B1(_10458_));
 sg13g2_buf_2 _17912_ (.A(_11126_),
    .X(_11127_));
 sg13g2_nand2b_1 _17913_ (.Y(_11128_),
    .B(_11127_),
    .A_N(_10489_));
 sg13g2_a21o_1 _17914_ (.A2(_11128_),
    .A1(_10488_),
    .B1(_09115_),
    .X(_11129_));
 sg13g2_a21o_1 _17915_ (.A2(_11117_),
    .A1(_11118_),
    .B1(_09115_),
    .X(_11130_));
 sg13g2_o21ai_1 _17916_ (.B1(_11130_),
    .Y(_11131_),
    .A1(_11117_),
    .A2(_10460_));
 sg13g2_nand2_1 _17917_ (.Y(_11132_),
    .A(_11054_),
    .B(net333));
 sg13g2_o21ai_1 _17918_ (.B1(net333),
    .Y(_11133_),
    .A1(_11026_),
    .A2(_11054_));
 sg13g2_nor3_1 _17919_ (.A(_11026_),
    .B(net334),
    .C(net333),
    .Y(_11134_));
 sg13g2_a221oi_1 _17920_ (.B2(_00308_),
    .C1(_11134_),
    .B1(_11133_),
    .A1(_09115_),
    .Y(_11135_),
    .A2(_11132_));
 sg13g2_buf_1 _17921_ (.A(_11135_),
    .X(_11136_));
 sg13g2_or2_1 _17922_ (.X(_11137_),
    .B(_11136_),
    .A(_11120_));
 sg13g2_nand4_1 _17923_ (.B(_11129_),
    .C(_11131_),
    .A(_11125_),
    .Y(_11138_),
    .D(_11137_));
 sg13g2_a21oi_2 _17924_ (.B1(_11138_),
    .Y(_11139_),
    .A2(_11121_),
    .A1(_11003_));
 sg13g2_a21o_1 _17925_ (.A2(_10498_),
    .A1(_10494_),
    .B1(_11139_),
    .X(_11140_));
 sg13g2_buf_1 _17926_ (.A(_11140_),
    .X(_11141_));
 sg13g2_nand2_2 _17927_ (.Y(_11142_),
    .A(_10415_),
    .B(_10282_));
 sg13g2_nand3_1 _17928_ (.B(_10435_),
    .C(_10493_),
    .A(_11142_),
    .Y(_11143_));
 sg13g2_nand2_1 _17929_ (.Y(_11144_),
    .A(_11142_),
    .B(_10496_));
 sg13g2_nand2b_1 _17930_ (.Y(_11145_),
    .B(_10493_),
    .A_N(_11144_));
 sg13g2_a21o_1 _17931_ (.A2(_11145_),
    .A1(_11143_),
    .B1(_11139_),
    .X(_11146_));
 sg13g2_buf_1 _17932_ (.A(_11146_),
    .X(_11147_));
 sg13g2_or2_1 _17933_ (.X(_11148_),
    .B(_10433_),
    .A(_10403_));
 sg13g2_buf_1 _17934_ (.A(_11148_),
    .X(_11149_));
 sg13g2_buf_1 _17935_ (.A(_11149_),
    .X(_11150_));
 sg13g2_a21oi_1 _17936_ (.A1(_10497_),
    .A2(_11144_),
    .Y(_11151_),
    .B1(net204));
 sg13g2_a21oi_2 _17937_ (.B1(_11151_),
    .Y(_11152_),
    .A2(_11142_),
    .A1(net240));
 sg13g2_and3_1 _17938_ (.X(_11153_),
    .A(_11141_),
    .B(_11147_),
    .C(_11152_));
 sg13g2_nor2_1 _17939_ (.A(_10344_),
    .B(_10342_),
    .Y(_11154_));
 sg13g2_nand2_1 _17940_ (.Y(_11155_),
    .A(_10349_),
    .B(_11154_));
 sg13g2_o21ai_1 _17941_ (.B1(net1071),
    .Y(_11156_),
    .A1(_10349_),
    .A2(_11154_));
 sg13g2_nand3_1 _17942_ (.B(_11155_),
    .C(_11156_),
    .A(net206),
    .Y(_11157_));
 sg13g2_a21oi_1 _17943_ (.A1(_11155_),
    .A2(_11156_),
    .Y(_11158_),
    .B1(net206));
 sg13g2_a21oi_1 _17944_ (.A1(net1074),
    .A2(_11157_),
    .Y(_11159_),
    .B1(_11158_));
 sg13g2_a21o_1 _17945_ (.A2(net241),
    .A1(_10232_),
    .B1(_11159_),
    .X(_11160_));
 sg13g2_nand2_1 _17946_ (.Y(_11161_),
    .A(_10279_),
    .B(_10275_));
 sg13g2_a21oi_1 _17947_ (.A1(_11160_),
    .A2(_11161_),
    .Y(_11162_),
    .B1(net462));
 sg13g2_a221oi_1 _17948_ (.B2(_11153_),
    .C1(_11162_),
    .B1(_10376_),
    .A1(_10199_),
    .Y(_11163_),
    .A2(_10356_));
 sg13g2_buf_1 _17949_ (.A(_11163_),
    .X(_11164_));
 sg13g2_nor2_1 _17950_ (.A(_09118_),
    .B(_09121_),
    .Y(_11165_));
 sg13g2_inv_2 _17951_ (.Y(_11166_),
    .A(net240));
 sg13g2_buf_1 _17952_ (.A(_11123_),
    .X(_11167_));
 sg13g2_nor4_1 _17953_ (.A(_10342_),
    .B(net209),
    .C(_10183_),
    .D(net238),
    .Y(_11168_));
 sg13g2_nand3_1 _17954_ (.B(_11166_),
    .C(_11168_),
    .A(_10278_),
    .Y(_11169_));
 sg13g2_a21oi_1 _17955_ (.A1(_11019_),
    .A2(_11020_),
    .Y(_11170_),
    .B1(_11023_));
 sg13g2_buf_2 _17956_ (.A(_11170_),
    .X(_11171_));
 sg13g2_a21oi_1 _17957_ (.A1(_11047_),
    .A2(_11051_),
    .Y(_11172_),
    .B1(_11052_));
 sg13g2_buf_1 _17958_ (.A(_11172_),
    .X(_11173_));
 sg13g2_nor2_1 _17959_ (.A(_11171_),
    .B(net362),
    .Y(_11174_));
 sg13g2_buf_2 _17960_ (.A(_11174_),
    .X(_11175_));
 sg13g2_and3_1 _17961_ (.X(_11176_),
    .A(_11068_),
    .B(_11074_),
    .C(_11075_));
 sg13g2_buf_1 _17962_ (.A(_11176_),
    .X(_11177_));
 sg13g2_inv_1 _17963_ (.Y(_11178_),
    .A(_11081_));
 sg13g2_nor2_1 _17964_ (.A(_11177_),
    .B(_11178_),
    .Y(_11179_));
 sg13g2_buf_1 _17965_ (.A(_11179_),
    .X(_11180_));
 sg13g2_buf_1 _17966_ (.A(_11117_),
    .X(_11181_));
 sg13g2_nor2_2 _17967_ (.A(_11180_),
    .B(_11181_),
    .Y(_11182_));
 sg13g2_nand2_2 _17968_ (.Y(_11183_),
    .A(_11175_),
    .B(_11182_));
 sg13g2_buf_1 _17969_ (.A(_10349_),
    .X(_11184_));
 sg13g2_nor2_1 _17970_ (.A(net296),
    .B(net181),
    .Y(_11185_));
 sg13g2_buf_1 _17971_ (.A(_11127_),
    .X(_11186_));
 sg13g2_nand4_1 _17972_ (.B(_11185_),
    .C(net204),
    .A(net203),
    .Y(_11187_),
    .D(_11186_));
 sg13g2_nor3_1 _17973_ (.A(_11169_),
    .B(_11183_),
    .C(_11187_),
    .Y(_11188_));
 sg13g2_or3_1 _17974_ (.A(_11165_),
    .B(_09127_),
    .C(_11188_),
    .X(_11189_));
 sg13g2_buf_1 _17975_ (.A(_11189_),
    .X(_11190_));
 sg13g2_inv_1 _17976_ (.Y(_11191_),
    .A(_11003_));
 sg13g2_buf_1 _17977_ (.A(_11191_),
    .X(_11192_));
 sg13g2_buf_1 _17978_ (.A(_11171_),
    .X(_11193_));
 sg13g2_nand3_1 _17979_ (.B(net88),
    .C(net292),
    .A(_09127_),
    .Y(_11194_));
 sg13g2_o21ai_1 _17980_ (.B1(_11194_),
    .Y(_11195_),
    .A1(net33),
    .A2(_11190_));
 sg13g2_buf_1 _17981_ (.A(_09123_),
    .X(_11196_));
 sg13g2_nor2_1 _17982_ (.A(_09118_),
    .B(net989),
    .Y(_11197_));
 sg13g2_and2_1 _17983_ (.A(_09116_),
    .B(_11197_),
    .X(_11198_));
 sg13g2_buf_2 _17984_ (.A(_11198_),
    .X(_11199_));
 sg13g2_nand2b_1 _17985_ (.Y(_11200_),
    .B(_09974_),
    .A_N(_11199_));
 sg13g2_buf_2 _17986_ (.A(_11200_),
    .X(_11201_));
 sg13g2_buf_1 _17987_ (.A(_11201_),
    .X(_11202_));
 sg13g2_buf_1 _17988_ (.A(\cpu.ex.r_mult[0] ),
    .X(_11203_));
 sg13g2_a22oi_1 _17989_ (.Y(_11204_),
    .B1(net291),
    .B2(_11203_),
    .A2(_11195_),
    .A1(net463));
 sg13g2_inv_1 _17990_ (.Y(\cpu.ex.c_mult[0] ),
    .A(_11204_));
 sg13g2_buf_1 _17991_ (.A(\cpu.dec.load ),
    .X(_11205_));
 sg13g2_o21ai_1 _17992_ (.B1(_08515_),
    .Y(_11206_),
    .A1(_08557_),
    .A2(_08617_));
 sg13g2_buf_1 _17993_ (.A(_11206_),
    .X(_11207_));
 sg13g2_nand2b_1 _17994_ (.Y(_11208_),
    .B(net1018),
    .A_N(_09120_));
 sg13g2_nand2b_1 _17995_ (.Y(_11209_),
    .B(_11208_),
    .A_N(_11197_));
 sg13g2_nor2_1 _17996_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11210_));
 sg13g2_nand2_1 _17997_ (.Y(_11211_),
    .A(_10659_),
    .B(\cpu.dec.r_swapsp ));
 sg13g2_nor3_1 _17998_ (.A(net1091),
    .B(net1019),
    .C(_09108_),
    .Y(_11212_));
 sg13g2_nand2_1 _17999_ (.Y(_11213_),
    .A(_10521_),
    .B(\cpu.cond[2] ));
 sg13g2_nand2_1 _18000_ (.Y(_11214_),
    .A(_00258_),
    .B(_11213_));
 sg13g2_nand2_1 _18001_ (.Y(_11215_),
    .A(_08592_),
    .B(_11214_));
 sg13g2_buf_2 _18002_ (.A(_11215_),
    .X(_11216_));
 sg13g2_o21ai_1 _18003_ (.B1(_11216_),
    .Y(_11217_),
    .A1(_10521_),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand4_1 _18004_ (.B(_11211_),
    .C(_11212_),
    .A(_11210_),
    .Y(_11218_),
    .D(_11217_));
 sg13g2_nand3_1 _18005_ (.B(_11209_),
    .C(_11218_),
    .A(_11207_),
    .Y(_11219_));
 sg13g2_buf_1 _18006_ (.A(_11219_),
    .X(_11220_));
 sg13g2_and2_1 _18007_ (.A(net1018),
    .B(_11220_),
    .X(_11221_));
 sg13g2_buf_1 _18008_ (.A(_11221_),
    .X(_11222_));
 sg13g2_buf_1 _18009_ (.A(_11222_),
    .X(_11223_));
 sg13g2_nand2_1 _18010_ (.Y(_11224_),
    .A(_00310_),
    .B(net106));
 sg13g2_nand2_1 _18011_ (.Y(_11225_),
    .A(net1018),
    .B(_11220_));
 sg13g2_buf_1 _18012_ (.A(_11225_),
    .X(_11226_));
 sg13g2_nor2b_1 _18013_ (.A(_08534_),
    .B_N(_09011_),
    .Y(_11227_));
 sg13g2_nand2_1 _18014_ (.Y(_11228_),
    .A(_09566_),
    .B(_09568_));
 sg13g2_a21oi_1 _18015_ (.A1(_11227_),
    .A2(_11228_),
    .Y(_11229_),
    .B1(_09017_));
 sg13g2_nand2_1 _18016_ (.Y(_11230_),
    .A(_11226_),
    .B(_11229_));
 sg13g2_a21o_1 _18017_ (.A2(_11230_),
    .A1(_11224_),
    .B1(_10512_),
    .X(_11231_));
 sg13g2_o21ai_1 _18018_ (.B1(_11231_),
    .Y(_00054_),
    .A1(_11205_),
    .A2(_11224_));
 sg13g2_nand2b_1 _18019_ (.Y(_11232_),
    .B(_09972_),
    .A_N(_09971_));
 sg13g2_buf_1 _18020_ (.A(_11232_),
    .X(_11233_));
 sg13g2_nor3_1 _18021_ (.A(_11165_),
    .B(_09127_),
    .C(_11188_),
    .Y(_11234_));
 sg13g2_buf_1 _18022_ (.A(_11234_),
    .X(_11235_));
 sg13g2_nor2_1 _18023_ (.A(_11003_),
    .B(net334),
    .Y(_11236_));
 sg13g2_buf_1 _18024_ (.A(_09112_),
    .X(_11237_));
 sg13g2_buf_1 _18025_ (.A(net522),
    .X(_11238_));
 sg13g2_buf_1 _18026_ (.A(net461),
    .X(_11239_));
 sg13g2_buf_1 _18027_ (.A(net398),
    .X(_11240_));
 sg13g2_buf_1 _18028_ (.A(_09126_),
    .X(_11241_));
 sg13g2_nand2_1 _18029_ (.Y(_11242_),
    .A(_11203_),
    .B(net521));
 sg13g2_mux2_1 _18030_ (.A0(_11242_),
    .A1(_11203_),
    .S(_11236_),
    .X(_11243_));
 sg13g2_nor2_1 _18031_ (.A(_09124_),
    .B(_11243_),
    .Y(_11244_));
 sg13g2_a221oi_1 _18032_ (.B2(net361),
    .C1(_11244_),
    .B1(_11236_),
    .A1(_11203_),
    .Y(_11245_),
    .A2(net81));
 sg13g2_buf_1 _18033_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11246_));
 sg13g2_nand2_1 _18034_ (.Y(_11247_),
    .A(_11246_),
    .B(_11201_));
 sg13g2_o21ai_1 _18035_ (.B1(_11247_),
    .Y(\cpu.ex.c_mult[1] ),
    .A1(net523),
    .A2(_11245_));
 sg13g2_buf_1 _18036_ (.A(_11241_),
    .X(_11248_));
 sg13g2_inv_1 _18037_ (.Y(_11249_),
    .A(_11203_));
 sg13g2_a221oi_1 _18038_ (.B2(_11051_),
    .C1(_11249_),
    .B1(_11047_),
    .A1(_08721_),
    .Y(_11250_),
    .A2(net1002));
 sg13g2_buf_1 _18039_ (.A(_11250_),
    .X(_11251_));
 sg13g2_inv_1 _18040_ (.Y(_11252_),
    .A(_11246_));
 sg13g2_nand3b_1 _18041_ (.B(net989),
    .C(_11252_),
    .Y(_11253_),
    .A_N(_11251_));
 sg13g2_buf_1 _18042_ (.A(_11083_),
    .X(_11254_));
 sg13g2_a21oi_1 _18043_ (.A1(net460),
    .A2(_11253_),
    .Y(_11255_),
    .B1(_11254_));
 sg13g2_buf_1 _18044_ (.A(_11003_),
    .X(_11256_));
 sg13g2_buf_1 _18045_ (.A(net105),
    .X(_11257_));
 sg13g2_buf_1 _18046_ (.A(_11180_),
    .X(_11258_));
 sg13g2_nor2_1 _18047_ (.A(net289),
    .B(_11251_),
    .Y(_11259_));
 sg13g2_o21ai_1 _18048_ (.B1(_11246_),
    .Y(_11260_),
    .A1(_11257_),
    .A2(_11259_));
 sg13g2_o21ai_1 _18049_ (.B1(_11252_),
    .Y(_11261_),
    .A1(_11177_),
    .A2(_11178_));
 sg13g2_nor2_1 _18050_ (.A(net105),
    .B(_11261_),
    .Y(_11262_));
 sg13g2_nor3_1 _18051_ (.A(_11252_),
    .B(_11177_),
    .C(_11178_),
    .Y(_11263_));
 sg13g2_o21ai_1 _18052_ (.B1(_11251_),
    .Y(_11264_),
    .A1(_11262_),
    .A2(_11263_));
 sg13g2_nand2_2 _18053_ (.Y(_11265_),
    .A(_11196_),
    .B(net460));
 sg13g2_a21oi_1 _18054_ (.A1(_11260_),
    .A2(_11264_),
    .Y(_11266_),
    .B1(_11265_));
 sg13g2_a221oi_1 _18055_ (.B2(_11192_),
    .C1(_11266_),
    .B1(_11255_),
    .A1(_11246_),
    .Y(_11267_),
    .A2(net81));
 sg13g2_nand2_1 _18056_ (.Y(_11268_),
    .A(\cpu.ex.r_mult[2] ),
    .B(_11201_));
 sg13g2_o21ai_1 _18057_ (.B1(_11268_),
    .Y(\cpu.ex.c_mult[2] ),
    .A1(_11233_),
    .A2(_11267_));
 sg13g2_buf_1 _18058_ (.A(_00120_),
    .X(_11269_));
 sg13g2_nand2_1 _18059_ (.Y(_11270_),
    .A(_11111_),
    .B(_11115_));
 sg13g2_buf_2 _18060_ (.A(_11270_),
    .X(_11271_));
 sg13g2_buf_1 _18061_ (.A(_11271_),
    .X(_11272_));
 sg13g2_buf_1 _18062_ (.A(net235),
    .X(_11273_));
 sg13g2_nand2_1 _18063_ (.Y(_11274_),
    .A(_11269_),
    .B(net202));
 sg13g2_inv_1 _18064_ (.Y(_11275_),
    .A(_11269_));
 sg13g2_nand3_1 _18065_ (.B(_11111_),
    .C(_11115_),
    .A(_11275_),
    .Y(_11276_));
 sg13g2_o21ai_1 _18066_ (.B1(_11276_),
    .Y(_11277_),
    .A1(net87),
    .A2(_11274_));
 sg13g2_a21oi_1 _18067_ (.A1(_11251_),
    .A2(_11261_),
    .Y(_11278_),
    .B1(_11263_));
 sg13g2_nor2_1 _18068_ (.A(_11239_),
    .B(_11278_),
    .Y(_11279_));
 sg13g2_a21o_1 _18069_ (.A2(_11278_),
    .A1(net202),
    .B1(net87),
    .X(_11280_));
 sg13g2_nor2_1 _18070_ (.A(_11269_),
    .B(net361),
    .Y(_11281_));
 sg13g2_buf_1 _18071_ (.A(_11181_),
    .X(_11282_));
 sg13g2_and4_1 _18072_ (.A(_11269_),
    .B(_11192_),
    .C(_11282_),
    .D(_11278_),
    .X(_11283_));
 sg13g2_a221oi_1 _18073_ (.B2(_11281_),
    .C1(_11283_),
    .B1(_11280_),
    .A1(_11277_),
    .Y(_11284_),
    .A2(_11279_));
 sg13g2_nor2_1 _18074_ (.A(net460),
    .B(net87),
    .Y(_11285_));
 sg13g2_a22oi_1 _18075_ (.Y(_11286_),
    .B1(_11285_),
    .B2(_11282_),
    .A2(net81),
    .A1(_11275_));
 sg13g2_o21ai_1 _18076_ (.B1(_11286_),
    .Y(_11287_),
    .A1(_09124_),
    .A2(_11284_));
 sg13g2_a22oi_1 _18077_ (.Y(_11288_),
    .B1(_11287_),
    .B2(_09974_),
    .A2(_11201_),
    .A1(\cpu.ex.r_mult[3] ));
 sg13g2_inv_1 _18078_ (.Y(\cpu.ex.c_mult[3] ),
    .A(_11288_));
 sg13g2_buf_1 _18079_ (.A(_11257_),
    .X(_11289_));
 sg13g2_buf_1 _18080_ (.A(_00127_),
    .X(_11290_));
 sg13g2_nor2_1 _18081_ (.A(_11290_),
    .B(net398),
    .Y(_11291_));
 sg13g2_nand2_1 _18082_ (.Y(_11292_),
    .A(_11290_),
    .B(_10487_));
 sg13g2_inv_1 _18083_ (.Y(_11293_),
    .A(_11290_));
 sg13g2_nand2_1 _18084_ (.Y(_11294_),
    .A(_11293_),
    .B(net238));
 sg13g2_o21ai_1 _18085_ (.B1(_11294_),
    .Y(_11295_),
    .A1(net87),
    .A2(_11292_));
 sg13g2_a21oi_1 _18086_ (.A1(_11111_),
    .A2(_11115_),
    .Y(_11296_),
    .B1(_11275_));
 sg13g2_a21oi_1 _18087_ (.A1(_11278_),
    .A2(_11276_),
    .Y(_11297_),
    .B1(_11296_));
 sg13g2_buf_1 _18088_ (.A(_11297_),
    .X(_11298_));
 sg13g2_and2_1 _18089_ (.A(net460),
    .B(_11298_),
    .X(_11299_));
 sg13g2_nand3b_1 _18090_ (.B(net238),
    .C(_11290_),
    .Y(_11300_),
    .A_N(net105));
 sg13g2_nand2_1 _18091_ (.Y(_11301_),
    .A(_10487_),
    .B(_11291_));
 sg13g2_a21oi_1 _18092_ (.A1(_11300_),
    .A2(_11301_),
    .Y(_11302_),
    .B1(_11298_));
 sg13g2_a221oi_1 _18093_ (.B2(_11299_),
    .C1(_11302_),
    .B1(_11295_),
    .A1(net80),
    .Y(_11303_),
    .A2(_11291_));
 sg13g2_a22oi_1 _18094_ (.Y(_11304_),
    .B1(_11285_),
    .B2(net238),
    .A2(net81),
    .A1(_11293_));
 sg13g2_o21ai_1 _18095_ (.B1(_11304_),
    .Y(_11305_),
    .A1(_09124_),
    .A2(_11303_));
 sg13g2_a22oi_1 _18096_ (.Y(_11306_),
    .B1(_11305_),
    .B2(net463),
    .A2(net291),
    .A1(\cpu.ex.r_mult[4] ));
 sg13g2_inv_1 _18097_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11306_));
 sg13g2_buf_1 _18098_ (.A(_00139_),
    .X(_11307_));
 sg13g2_inv_1 _18099_ (.Y(_11308_),
    .A(_11307_));
 sg13g2_nand2_1 _18100_ (.Y(_11309_),
    .A(net238),
    .B(_11298_));
 sg13g2_o21ai_1 _18101_ (.B1(_11293_),
    .Y(_11310_),
    .A1(net238),
    .A2(_11298_));
 sg13g2_nand2_1 _18102_ (.Y(_11311_),
    .A(_11309_),
    .B(_11310_));
 sg13g2_nand2_1 _18103_ (.Y(_11312_),
    .A(_11307_),
    .B(_11127_));
 sg13g2_nor2_1 _18104_ (.A(_11307_),
    .B(net236),
    .Y(_11313_));
 sg13g2_inv_1 _18105_ (.Y(_11314_),
    .A(_11313_));
 sg13g2_o21ai_1 _18106_ (.B1(_11314_),
    .Y(_11315_),
    .A1(net105),
    .A2(_11312_));
 sg13g2_a22oi_1 _18107_ (.Y(_11316_),
    .B1(_11311_),
    .B2(_11315_),
    .A2(net87),
    .A1(_11308_));
 sg13g2_nand2_1 _18108_ (.Y(_11317_),
    .A(_11307_),
    .B(net295));
 sg13g2_nand3_1 _18109_ (.B(net521),
    .C(net236),
    .A(_11308_),
    .Y(_11318_));
 sg13g2_o21ai_1 _18110_ (.B1(_11318_),
    .Y(_11319_),
    .A1(net105),
    .A2(_11317_));
 sg13g2_nand2b_1 _18111_ (.Y(_11320_),
    .B(_11319_),
    .A_N(_11311_));
 sg13g2_o21ai_1 _18112_ (.B1(_11320_),
    .Y(_11321_),
    .A1(net361),
    .A2(_11316_));
 sg13g2_nor3_1 _18113_ (.A(_11248_),
    .B(_11289_),
    .C(net236),
    .Y(_11322_));
 sg13g2_a221oi_1 _18114_ (.B2(net989),
    .C1(_11322_),
    .B1(_11321_),
    .A1(_11308_),
    .Y(_11323_),
    .A2(net81));
 sg13g2_nand2_1 _18115_ (.Y(_11324_),
    .A(\cpu.ex.r_mult[5] ),
    .B(_11201_));
 sg13g2_o21ai_1 _18116_ (.B1(_11324_),
    .Y(\cpu.ex.c_mult[5] ),
    .A1(net523),
    .A2(_11323_));
 sg13g2_buf_2 _18117_ (.A(_00151_),
    .X(_11325_));
 sg13g2_inv_1 _18118_ (.Y(_11326_),
    .A(_11325_));
 sg13g2_nor2_1 _18119_ (.A(_11325_),
    .B(net398),
    .Y(_11327_));
 sg13g2_a22oi_1 _18120_ (.Y(_11328_),
    .B1(net295),
    .B2(_11308_),
    .A2(_11123_),
    .A1(_11293_));
 sg13g2_nand2_1 _18121_ (.Y(_11329_),
    .A(_11298_),
    .B(_11292_));
 sg13g2_a221oi_1 _18122_ (.B2(_11329_),
    .C1(net522),
    .B1(_11328_),
    .A1(_11307_),
    .Y(_11330_),
    .A2(_11127_));
 sg13g2_buf_1 _18123_ (.A(_11330_),
    .X(_11331_));
 sg13g2_xnor2_1 _18124_ (.Y(_11332_),
    .A(_10435_),
    .B(_11331_));
 sg13g2_nor2_1 _18125_ (.A(net105),
    .B(_11332_),
    .Y(_11333_));
 sg13g2_mux2_1 _18126_ (.A0(_11327_),
    .A1(_11325_),
    .S(_11333_),
    .X(_11334_));
 sg13g2_nor3_1 _18127_ (.A(_11248_),
    .B(net204),
    .C(_11289_),
    .Y(_11335_));
 sg13g2_a221oi_1 _18128_ (.B2(net989),
    .C1(_11335_),
    .B1(_11334_),
    .A1(_11326_),
    .Y(_11336_),
    .A2(net81));
 sg13g2_nand2_1 _18129_ (.Y(_11337_),
    .A(\cpu.ex.r_mult[6] ),
    .B(_11201_));
 sg13g2_o21ai_1 _18130_ (.B1(_11337_),
    .Y(\cpu.ex.c_mult[6] ),
    .A1(net523),
    .A2(_11336_));
 sg13g2_inv_2 _18131_ (.Y(_11338_),
    .A(_00163_));
 sg13g2_nand2_1 _18132_ (.Y(_11339_),
    .A(_11338_),
    .B(_09126_));
 sg13g2_o21ai_1 _18133_ (.B1(_11325_),
    .Y(_11340_),
    .A1(_10403_),
    .A2(_10433_));
 sg13g2_and4_1 _18134_ (.A(_11298_),
    .B(_11292_),
    .C(_11312_),
    .D(_11340_),
    .X(_11341_));
 sg13g2_nor2_1 _18135_ (.A(_11325_),
    .B(net204),
    .Y(_11342_));
 sg13g2_a221oi_1 _18136_ (.B2(_11307_),
    .C1(_11328_),
    .B1(net236),
    .A1(_11325_),
    .Y(_11343_),
    .A2(_11149_));
 sg13g2_or3_1 _18137_ (.A(_11341_),
    .B(_11342_),
    .C(_11343_),
    .X(_11344_));
 sg13g2_buf_1 _18138_ (.A(_11344_),
    .X(_11345_));
 sg13g2_a21o_1 _18139_ (.A2(_11345_),
    .A1(net521),
    .B1(_11166_),
    .X(_11346_));
 sg13g2_nand3_1 _18140_ (.B(_11166_),
    .C(_11345_),
    .A(net521),
    .Y(_11347_));
 sg13g2_a21oi_1 _18141_ (.A1(_11346_),
    .A2(_11347_),
    .Y(_11348_),
    .B1(net105));
 sg13g2_mux2_1 _18142_ (.A0(_11339_),
    .A1(_11338_),
    .S(_11348_),
    .X(_11349_));
 sg13g2_a22oi_1 _18143_ (.Y(_11350_),
    .B1(_11348_),
    .B2(net361),
    .A2(net81),
    .A1(_11338_));
 sg13g2_o21ai_1 _18144_ (.B1(_11350_),
    .Y(_11351_),
    .A1(_09124_),
    .A2(_11349_));
 sg13g2_and2_1 _18145_ (.A(\cpu.ex.r_mult[7] ),
    .B(_11201_),
    .X(_11352_));
 sg13g2_a21o_1 _18146_ (.A2(_11351_),
    .A1(_09974_),
    .B1(_11352_),
    .X(\cpu.ex.c_mult[7] ));
 sg13g2_o21ai_1 _18147_ (.B1(_11326_),
    .Y(_11353_),
    .A1(_11338_),
    .A2(_10401_));
 sg13g2_nand2_1 _18148_ (.Y(_11354_),
    .A(_11338_),
    .B(_10401_));
 sg13g2_o21ai_1 _18149_ (.B1(_11354_),
    .Y(_11355_),
    .A1(_11149_),
    .A2(_11353_));
 sg13g2_mux2_1 _18150_ (.A0(_11339_),
    .A1(_11338_),
    .S(_10401_),
    .X(_11356_));
 sg13g2_nor3_1 _18151_ (.A(_11326_),
    .B(net204),
    .C(_11356_),
    .Y(_11357_));
 sg13g2_xnor2_1 _18152_ (.Y(_11358_),
    .A(_11338_),
    .B(_10401_));
 sg13g2_nor4_1 _18153_ (.A(_11325_),
    .B(net522),
    .C(_10435_),
    .D(_11358_),
    .Y(_11359_));
 sg13g2_or2_1 _18154_ (.X(_11360_),
    .B(_11359_),
    .A(_11357_));
 sg13g2_a22oi_1 _18155_ (.Y(_11361_),
    .B1(_11360_),
    .B2(_11331_),
    .A2(_11355_),
    .A1(net521));
 sg13g2_xnor2_1 _18156_ (.Y(_11362_),
    .A(_10116_),
    .B(_11361_));
 sg13g2_nor2_1 _18157_ (.A(net87),
    .B(_11362_),
    .Y(_11363_));
 sg13g2_buf_2 _18158_ (.A(_00164_),
    .X(_11364_));
 sg13g2_nor2_1 _18159_ (.A(_11364_),
    .B(net522),
    .Y(_11365_));
 sg13g2_mux2_1 _18160_ (.A0(_11365_),
    .A1(_11364_),
    .S(_11363_),
    .X(_11366_));
 sg13g2_nor2_1 _18161_ (.A(_11364_),
    .B(_11190_),
    .Y(_11367_));
 sg13g2_a221oi_1 _18162_ (.B2(net989),
    .C1(_11367_),
    .B1(_11366_),
    .A1(net361),
    .Y(_11368_),
    .A2(_11363_));
 sg13g2_nand2_1 _18163_ (.Y(_11369_),
    .A(\cpu.ex.r_mult[8] ),
    .B(net291));
 sg13g2_o21ai_1 _18164_ (.B1(_11369_),
    .Y(\cpu.ex.c_mult[8] ),
    .A1(net523),
    .A2(_11368_));
 sg13g2_buf_1 _18165_ (.A(_00165_),
    .X(_11370_));
 sg13g2_inv_1 _18166_ (.Y(_11371_),
    .A(net1070));
 sg13g2_buf_1 _18167_ (.A(_11235_),
    .X(_11372_));
 sg13g2_buf_1 _18168_ (.A(net296),
    .X(_11373_));
 sg13g2_nor3_1 _18169_ (.A(_11364_),
    .B(_10067_),
    .C(_10108_),
    .Y(_11374_));
 sg13g2_o21ai_1 _18170_ (.B1(_11364_),
    .Y(_11375_),
    .A1(_10067_),
    .A2(_10108_));
 sg13g2_nand2b_1 _18171_ (.Y(_11376_),
    .B(_11375_),
    .A_N(_11374_));
 sg13g2_nor3_1 _18172_ (.A(net461),
    .B(_11358_),
    .C(_11376_),
    .Y(_11377_));
 sg13g2_and2_1 _18173_ (.A(_11338_),
    .B(net240),
    .X(_11378_));
 sg13g2_a21oi_2 _18174_ (.B1(_11374_),
    .Y(_11379_),
    .A2(_11375_),
    .A1(_11378_));
 sg13g2_nor2_1 _18175_ (.A(net398),
    .B(_11379_),
    .Y(_11380_));
 sg13g2_a21oi_1 _18176_ (.A1(_11345_),
    .A2(_11377_),
    .Y(_11381_),
    .B1(_11380_));
 sg13g2_xnor2_1 _18177_ (.Y(_11382_),
    .A(net234),
    .B(_11381_));
 sg13g2_and2_1 _18178_ (.A(net88),
    .B(_11382_),
    .X(_11383_));
 sg13g2_a22oi_1 _18179_ (.Y(_11384_),
    .B1(_11383_),
    .B2(net361),
    .A2(_11372_),
    .A1(_11371_));
 sg13g2_buf_1 _18180_ (.A(_09110_),
    .X(_11385_));
 sg13g2_a221oi_1 _18181_ (.B2(_11382_),
    .C1(net1070),
    .B1(net88),
    .A1(_09106_),
    .Y(_11386_),
    .A2(net646));
 sg13g2_and3_1 _18182_ (.X(_11387_),
    .A(_11370_),
    .B(net88),
    .C(_11382_));
 sg13g2_o21ai_1 _18183_ (.B1(net989),
    .Y(_11388_),
    .A1(_11386_),
    .A2(_11387_));
 sg13g2_a21oi_1 _18184_ (.A1(_11384_),
    .A2(_11388_),
    .Y(_11389_),
    .B1(net523));
 sg13g2_a21oi_1 _18185_ (.A1(\cpu.ex.r_mult[9] ),
    .A2(net291),
    .Y(_11390_),
    .B1(_11389_));
 sg13g2_inv_1 _18186_ (.Y(\cpu.ex.c_mult[9] ),
    .A(_11390_));
 sg13g2_nor2_1 _18187_ (.A(net1070),
    .B(_09112_),
    .Y(_11391_));
 sg13g2_mux2_1 _18188_ (.A0(_11391_),
    .A1(net1070),
    .S(net296),
    .X(_11392_));
 sg13g2_a22oi_1 _18189_ (.Y(_11393_),
    .B1(_11392_),
    .B2(_11364_),
    .A2(net296),
    .A1(_11237_));
 sg13g2_nand3_1 _18190_ (.B(_10065_),
    .C(_11365_),
    .A(net1070),
    .Y(_11394_));
 sg13g2_mux2_1 _18191_ (.A0(_11393_),
    .A1(_11394_),
    .S(net182),
    .X(_11395_));
 sg13g2_nor3_1 _18192_ (.A(_11364_),
    .B(net1070),
    .C(_11237_),
    .Y(_11396_));
 sg13g2_o21ai_1 _18193_ (.B1(_11396_),
    .Y(_11397_),
    .A1(_11185_),
    .A2(_11003_));
 sg13g2_nand2_1 _18194_ (.Y(_11398_),
    .A(_11331_),
    .B(_11360_));
 sg13g2_a21o_1 _18195_ (.A2(_11397_),
    .A1(_11395_),
    .B1(_11398_),
    .X(_11399_));
 sg13g2_buf_1 _18196_ (.A(_11399_),
    .X(_11400_));
 sg13g2_nand3_1 _18197_ (.B(net181),
    .C(_11355_),
    .A(_09126_),
    .Y(_11401_));
 sg13g2_nor2_1 _18198_ (.A(net205),
    .B(_11401_),
    .Y(_11402_));
 sg13g2_a221oi_1 _18199_ (.B2(_11401_),
    .C1(net1070),
    .B1(_10114_),
    .A1(_09106_),
    .Y(_11403_),
    .A2(net646));
 sg13g2_a21oi_1 _18200_ (.A1(_09126_),
    .A2(_11355_),
    .Y(_11404_),
    .B1(net181));
 sg13g2_nor2_1 _18201_ (.A(_11371_),
    .B(net234),
    .Y(_11405_));
 sg13g2_nor4_1 _18202_ (.A(_11364_),
    .B(net461),
    .C(_11404_),
    .D(_11405_),
    .Y(_11406_));
 sg13g2_nor3_2 _18203_ (.A(_11402_),
    .B(_11403_),
    .C(_11406_),
    .Y(_11407_));
 sg13g2_and3_1 _18204_ (.X(_11408_),
    .A(net207),
    .B(_11400_),
    .C(_11407_));
 sg13g2_a21oi_1 _18205_ (.A1(_11400_),
    .A2(_11407_),
    .Y(_11409_),
    .B1(net207));
 sg13g2_nor3_1 _18206_ (.A(net87),
    .B(_11408_),
    .C(_11409_),
    .Y(_11410_));
 sg13g2_nand3_1 _18207_ (.B(net460),
    .C(_09974_),
    .A(net989),
    .Y(_11411_));
 sg13g2_buf_1 _18208_ (.A(_11411_),
    .X(_11412_));
 sg13g2_nand2_2 _18209_ (.Y(_11413_),
    .A(_09974_),
    .B(net81));
 sg13g2_o21ai_1 _18210_ (.B1(_11413_),
    .Y(_11414_),
    .A1(_11410_),
    .A2(_11412_));
 sg13g2_buf_1 _18211_ (.A(_00166_),
    .X(_11415_));
 sg13g2_inv_1 _18212_ (.Y(_11416_),
    .A(_11415_));
 sg13g2_nand2_1 _18213_ (.Y(_11417_),
    .A(_09127_),
    .B(_09974_));
 sg13g2_buf_2 _18214_ (.A(_11417_),
    .X(_11418_));
 sg13g2_nor2_1 _18215_ (.A(_11415_),
    .B(_09112_),
    .Y(_11419_));
 sg13g2_nor2_1 _18216_ (.A(_11418_),
    .B(_11419_),
    .Y(_11420_));
 sg13g2_and2_1 _18217_ (.A(_11410_),
    .B(_11420_),
    .X(_11421_));
 sg13g2_a221oi_1 _18218_ (.B2(_11416_),
    .C1(_11421_),
    .B1(_11414_),
    .A1(\cpu.ex.r_mult[10] ),
    .Y(_11422_),
    .A2(net291));
 sg13g2_buf_1 _18219_ (.A(_11422_),
    .X(_11423_));
 sg13g2_inv_1 _18220_ (.Y(\cpu.ex.c_mult[10] ),
    .A(_11423_));
 sg13g2_buf_1 _18221_ (.A(_00167_),
    .X(_11424_));
 sg13g2_inv_1 _18222_ (.Y(_11425_),
    .A(_11424_));
 sg13g2_buf_1 _18223_ (.A(_10154_),
    .X(_11426_));
 sg13g2_mux2_1 _18224_ (.A0(_11415_),
    .A1(_11419_),
    .S(_10187_),
    .X(_11427_));
 sg13g2_a22oi_1 _18225_ (.Y(_11428_),
    .B1(_11427_),
    .B2(net1070),
    .A2(_10183_),
    .A1(net461));
 sg13g2_xnor2_1 _18226_ (.Y(_11429_),
    .A(_11416_),
    .B(_10187_));
 sg13g2_nand3_1 _18227_ (.B(_11391_),
    .C(_11429_),
    .A(_10114_),
    .Y(_11430_));
 sg13g2_o21ai_1 _18228_ (.B1(_11430_),
    .Y(_11431_),
    .A1(net205),
    .A2(_11428_));
 sg13g2_nand3_1 _18229_ (.B(_11377_),
    .C(_11431_),
    .A(_11345_),
    .Y(_11432_));
 sg13g2_buf_1 _18230_ (.A(_11432_),
    .X(_11433_));
 sg13g2_nor4_1 _18231_ (.A(net461),
    .B(_10188_),
    .C(net205),
    .D(_11379_),
    .Y(_11434_));
 sg13g2_o21ai_1 _18232_ (.B1(_11371_),
    .Y(_11435_),
    .A1(_11416_),
    .A2(_10183_));
 sg13g2_nor3_1 _18233_ (.A(net398),
    .B(_11379_),
    .C(_11435_),
    .Y(_11436_));
 sg13g2_nor4_1 _18234_ (.A(_11415_),
    .B(net461),
    .C(net205),
    .D(_11379_),
    .Y(_11437_));
 sg13g2_nand2_1 _18235_ (.Y(_11438_),
    .A(net521),
    .B(net234));
 sg13g2_nand2_1 _18236_ (.Y(_11439_),
    .A(net208),
    .B(_11419_));
 sg13g2_o21ai_1 _18237_ (.B1(_11439_),
    .Y(_11440_),
    .A1(_11435_),
    .A2(_11438_));
 sg13g2_nor4_2 _18238_ (.A(_11434_),
    .B(_11436_),
    .C(_11437_),
    .Y(_11441_),
    .D(_11440_));
 sg13g2_nand2_1 _18239_ (.Y(_11442_),
    .A(_11433_),
    .B(_11441_));
 sg13g2_xnor2_1 _18240_ (.Y(_11443_),
    .A(net180),
    .B(_11442_));
 sg13g2_nor2_1 _18241_ (.A(net80),
    .B(_11443_),
    .Y(_11444_));
 sg13g2_o21ai_1 _18242_ (.B1(_11190_),
    .Y(_11445_),
    .A1(_11265_),
    .A2(_11444_));
 sg13g2_nand3_1 _18243_ (.B(net463),
    .C(_11445_),
    .A(_11425_),
    .Y(_11446_));
 sg13g2_nor2_1 _18244_ (.A(_11424_),
    .B(_09112_),
    .Y(_11447_));
 sg13g2_nor2_1 _18245_ (.A(_11418_),
    .B(_11447_),
    .Y(_11448_));
 sg13g2_a22oi_1 _18246_ (.Y(_11449_),
    .B1(_11444_),
    .B2(_11448_),
    .A2(net291),
    .A1(\cpu.ex.r_mult[11] ));
 sg13g2_nand2_1 _18247_ (.Y(\cpu.ex.c_mult[11] ),
    .A(_11446_),
    .B(_11449_));
 sg13g2_buf_1 _18248_ (.A(_10342_),
    .X(_11450_));
 sg13g2_and3_1 _18249_ (.X(_11451_),
    .A(_11416_),
    .B(_10155_),
    .C(_10181_));
 sg13g2_o21ai_1 _18250_ (.B1(_11451_),
    .Y(_11452_),
    .A1(_11425_),
    .A2(_10153_));
 sg13g2_nand2_1 _18251_ (.Y(_11453_),
    .A(_11425_),
    .B(_10153_));
 sg13g2_a21oi_1 _18252_ (.A1(_11452_),
    .A2(_11453_),
    .Y(_11454_),
    .B1(net461));
 sg13g2_nand2_1 _18253_ (.Y(_11455_),
    .A(_10187_),
    .B(_11419_));
 sg13g2_a21oi_1 _18254_ (.A1(_11424_),
    .A2(_10193_),
    .Y(_11456_),
    .B1(_11455_));
 sg13g2_mux2_1 _18255_ (.A0(_11447_),
    .A1(_11424_),
    .S(_10153_),
    .X(_11457_));
 sg13g2_a22oi_1 _18256_ (.Y(_11458_),
    .B1(_11457_),
    .B2(_11415_),
    .A2(_10153_),
    .A1(net522));
 sg13g2_nor2_1 _18257_ (.A(_10187_),
    .B(_11458_),
    .Y(_11459_));
 sg13g2_a21oi_1 _18258_ (.A1(_11453_),
    .A2(_11456_),
    .Y(_11460_),
    .B1(_11459_));
 sg13g2_a21oi_1 _18259_ (.A1(_11400_),
    .A2(_11407_),
    .Y(_11461_),
    .B1(_11460_));
 sg13g2_nor2_1 _18260_ (.A(_11454_),
    .B(_11461_),
    .Y(_11462_));
 sg13g2_xnor2_1 _18261_ (.Y(_11463_),
    .A(net200),
    .B(_11462_));
 sg13g2_buf_1 _18262_ (.A(_00168_),
    .X(_11464_));
 sg13g2_nor2_1 _18263_ (.A(_11464_),
    .B(net522),
    .Y(_11465_));
 sg13g2_nor2_1 _18264_ (.A(_11418_),
    .B(_11465_),
    .Y(_11466_));
 sg13g2_and3_1 _18265_ (.X(_11467_),
    .A(net88),
    .B(_11463_),
    .C(_11466_));
 sg13g2_or2_1 _18266_ (.X(_11468_),
    .B(_11412_),
    .A(_11464_));
 sg13g2_a21oi_1 _18267_ (.A1(net88),
    .A2(_11463_),
    .Y(_11469_),
    .B1(_11468_));
 sg13g2_nand2_1 _18268_ (.Y(_11470_),
    .A(\cpu.ex.r_mult[12] ),
    .B(_11201_));
 sg13g2_o21ai_1 _18269_ (.B1(_11470_),
    .Y(_11471_),
    .A1(_11464_),
    .A2(_11413_));
 sg13g2_or3_1 _18270_ (.A(_11467_),
    .B(_11469_),
    .C(_11471_),
    .X(\cpu.ex.c_mult[12] ));
 sg13g2_buf_1 _18271_ (.A(_10315_),
    .X(_11472_));
 sg13g2_nand2_1 _18272_ (.Y(_11473_),
    .A(_10928_),
    .B(_11000_));
 sg13g2_a22oi_1 _18273_ (.Y(_11474_),
    .B1(_10926_),
    .B2(_10927_),
    .A2(_10830_),
    .A1(_10825_));
 sg13g2_inv_1 _18274_ (.Y(_11475_),
    .A(_10342_));
 sg13g2_buf_1 _18275_ (.A(_11475_),
    .X(_11476_));
 sg13g2_a21oi_1 _18276_ (.A1(_11464_),
    .A2(net179),
    .Y(_11477_),
    .B1(_11424_));
 sg13g2_nand2_1 _18277_ (.Y(_11478_),
    .A(net521),
    .B(_11477_));
 sg13g2_a221oi_1 _18278_ (.B2(_11441_),
    .C1(_11478_),
    .B1(_11433_),
    .A1(_11473_),
    .Y(_11479_),
    .A2(_11474_));
 sg13g2_nand2_1 _18279_ (.Y(_11480_),
    .A(net209),
    .B(_11465_));
 sg13g2_a221oi_1 _18280_ (.B2(_11441_),
    .C1(_11480_),
    .B1(_11433_),
    .A1(_11473_),
    .Y(_11481_),
    .A2(_11474_));
 sg13g2_nand2_1 _18281_ (.Y(_11482_),
    .A(net200),
    .B(net209));
 sg13g2_a221oi_1 _18282_ (.B2(_11441_),
    .C1(_11482_),
    .B1(_11433_),
    .A1(_11473_),
    .Y(_11483_),
    .A2(_11474_));
 sg13g2_nand2_1 _18283_ (.Y(_11484_),
    .A(net200),
    .B(_11465_));
 sg13g2_nand3_1 _18284_ (.B(net180),
    .C(_11477_),
    .A(net521),
    .Y(_11485_));
 sg13g2_nand2_1 _18285_ (.Y(_11486_),
    .A(_11484_),
    .B(_11485_));
 sg13g2_or4_1 _18286_ (.A(_11479_),
    .B(_11481_),
    .C(_11483_),
    .D(_11486_),
    .X(_11487_));
 sg13g2_xnor2_1 _18287_ (.Y(_11488_),
    .A(net199),
    .B(_11487_));
 sg13g2_nor2_1 _18288_ (.A(net80),
    .B(_11488_),
    .Y(_11489_));
 sg13g2_buf_2 _18289_ (.A(_00169_),
    .X(_11490_));
 sg13g2_nor2_1 _18290_ (.A(_11490_),
    .B(net522),
    .Y(_11491_));
 sg13g2_xnor2_1 _18291_ (.Y(_11492_),
    .A(_11489_),
    .B(_11491_));
 sg13g2_nor2_1 _18292_ (.A(_11232_),
    .B(_11190_),
    .Y(_11493_));
 sg13g2_buf_2 _18293_ (.A(_11493_),
    .X(_11494_));
 sg13g2_inv_1 _18294_ (.Y(_11495_),
    .A(_11490_));
 sg13g2_a22oi_1 _18295_ (.Y(_11496_),
    .B1(_11494_),
    .B2(_11495_),
    .A2(net291),
    .A1(\cpu.ex.r_mult[13] ));
 sg13g2_o21ai_1 _18296_ (.B1(_11496_),
    .Y(\cpu.ex.c_mult[13] ),
    .A1(_11418_),
    .A2(_11492_));
 sg13g2_buf_1 _18297_ (.A(net206),
    .X(_11497_));
 sg13g2_a21oi_1 _18298_ (.A1(_11490_),
    .A2(net203),
    .Y(_11498_),
    .B1(_11464_));
 sg13g2_o21ai_1 _18299_ (.B1(_11498_),
    .Y(_11499_),
    .A1(net200),
    .A2(_11454_));
 sg13g2_a221oi_1 _18300_ (.B2(_11453_),
    .C1(_11475_),
    .B1(_11452_),
    .A1(_09106_),
    .Y(_11500_),
    .A2(_09110_));
 sg13g2_o21ai_1 _18301_ (.B1(_11495_),
    .Y(_11501_),
    .A1(_10315_),
    .A2(_11500_));
 sg13g2_a21oi_1 _18302_ (.A1(_11499_),
    .A2(_11501_),
    .Y(_11502_),
    .B1(net398));
 sg13g2_and2_1 _18303_ (.A(_10315_),
    .B(_11500_),
    .X(_11503_));
 sg13g2_or2_1 _18304_ (.X(_11504_),
    .B(_11503_),
    .A(_11502_));
 sg13g2_buf_1 _18305_ (.A(_11504_),
    .X(_11505_));
 sg13g2_mux2_1 _18306_ (.A0(_11490_),
    .A1(_11491_),
    .S(_10349_),
    .X(_11506_));
 sg13g2_a22oi_1 _18307_ (.Y(_11507_),
    .B1(_11506_),
    .B2(_11464_),
    .A2(_10315_),
    .A1(net461));
 sg13g2_xnor2_1 _18308_ (.Y(_11508_),
    .A(_11495_),
    .B(_10349_));
 sg13g2_nand2_1 _18309_ (.Y(_11509_),
    .A(_11465_),
    .B(_11508_));
 sg13g2_mux2_1 _18310_ (.A0(_11507_),
    .A1(_11509_),
    .S(net179),
    .X(_11510_));
 sg13g2_or3_1 _18311_ (.A(_11003_),
    .B(_11460_),
    .C(_11510_),
    .X(_11511_));
 sg13g2_a21oi_1 _18312_ (.A1(_11400_),
    .A2(_11407_),
    .Y(_11512_),
    .B1(_11511_));
 sg13g2_a21oi_1 _18313_ (.A1(net88),
    .A2(_11505_),
    .Y(_11513_),
    .B1(_11512_));
 sg13g2_buf_1 _18314_ (.A(_10272_),
    .X(_11514_));
 sg13g2_or4_1 _18315_ (.A(net151),
    .B(net80),
    .C(_11512_),
    .D(_11505_),
    .X(_11515_));
 sg13g2_o21ai_1 _18316_ (.B1(_11515_),
    .Y(_11516_),
    .A1(net178),
    .A2(_11513_));
 sg13g2_buf_2 _18317_ (.A(_00170_),
    .X(_11517_));
 sg13g2_nor2_1 _18318_ (.A(_11517_),
    .B(_11238_),
    .Y(_11518_));
 sg13g2_xnor2_1 _18319_ (.Y(_11519_),
    .A(_11516_),
    .B(_11518_));
 sg13g2_inv_1 _18320_ (.Y(_11520_),
    .A(_11517_));
 sg13g2_a22oi_1 _18321_ (.Y(_11521_),
    .B1(_11494_),
    .B2(_11520_),
    .A2(_11202_),
    .A1(\cpu.ex.r_mult[14] ));
 sg13g2_o21ai_1 _18322_ (.B1(_11521_),
    .Y(_11522_),
    .A1(_11418_),
    .A2(_11519_));
 sg13g2_buf_1 _18323_ (.A(_11522_),
    .X(\cpu.ex.c_mult[14] ));
 sg13g2_and2_1 _18324_ (.A(net203),
    .B(_11491_),
    .X(_11523_));
 sg13g2_and2_1 _18325_ (.A(_11517_),
    .B(net206),
    .X(_11524_));
 sg13g2_nor2b_1 _18326_ (.A(_10269_),
    .B_N(_11518_),
    .Y(_11525_));
 sg13g2_o21ai_1 _18327_ (.B1(_11490_),
    .Y(_11526_),
    .A1(_11524_),
    .A2(_11525_));
 sg13g2_o21ai_1 _18328_ (.B1(_11526_),
    .Y(_11527_),
    .A1(_11241_),
    .A2(net151));
 sg13g2_a22oi_1 _18329_ (.Y(_11528_),
    .B1(_11527_),
    .B2(net199),
    .A2(_11524_),
    .A1(_11523_));
 sg13g2_nor2_1 _18330_ (.A(net206),
    .B(net199),
    .Y(_11529_));
 sg13g2_nor3_1 _18331_ (.A(_11490_),
    .B(_11517_),
    .C(net398),
    .Y(_11530_));
 sg13g2_o21ai_1 _18332_ (.B1(_11530_),
    .Y(_11531_),
    .A1(net105),
    .A2(_11529_));
 sg13g2_o21ai_1 _18333_ (.B1(_11531_),
    .Y(_11532_),
    .A1(net87),
    .A2(_11528_));
 sg13g2_a21oi_1 _18334_ (.A1(_11517_),
    .A2(net151),
    .Y(_11533_),
    .B1(_11490_));
 sg13g2_nor2_1 _18335_ (.A(_11517_),
    .B(net151),
    .Y(_11534_));
 sg13g2_a21o_1 _18336_ (.A2(_11533_),
    .A1(net199),
    .B1(_11534_),
    .X(_11535_));
 sg13g2_a22oi_1 _18337_ (.Y(_11536_),
    .B1(_11535_),
    .B2(net460),
    .A2(_11532_),
    .A1(_11487_));
 sg13g2_or4_1 _18338_ (.A(net241),
    .B(net80),
    .C(_11494_),
    .D(_11536_),
    .X(_11537_));
 sg13g2_nand4_1 _18339_ (.B(net88),
    .C(_11413_),
    .A(net241),
    .Y(_11538_),
    .D(_11536_));
 sg13g2_buf_1 _18340_ (.A(_00171_),
    .X(_11539_));
 sg13g2_a21oi_1 _18341_ (.A1(_11413_),
    .A2(_11412_),
    .Y(_11540_),
    .B1(_11539_));
 sg13g2_nand3_1 _18342_ (.B(_11538_),
    .C(_11540_),
    .A(_11537_),
    .Y(_11541_));
 sg13g2_xnor2_1 _18343_ (.Y(_11542_),
    .A(_10275_),
    .B(_11536_));
 sg13g2_nor2_1 _18344_ (.A(_11539_),
    .B(net522),
    .Y(_11543_));
 sg13g2_or4_1 _18345_ (.A(net80),
    .B(_11418_),
    .C(_11542_),
    .D(_11543_),
    .X(_11544_));
 sg13g2_buf_1 _18346_ (.A(\cpu.ex.r_mult[15] ),
    .X(_11545_));
 sg13g2_nand2_1 _18347_ (.Y(_11546_),
    .A(_11545_),
    .B(_11202_));
 sg13g2_nand3_1 _18348_ (.B(_11544_),
    .C(_11546_),
    .A(_11541_),
    .Y(\cpu.ex.c_mult[15] ));
 sg13g2_inv_1 _18349_ (.Y(_00000_),
    .A(net2));
 sg13g2_inv_1 _18350_ (.Y(_11547_),
    .A(\cpu.qspi.r_state[11] ));
 sg13g2_nor2_1 _18351_ (.A(_11547_),
    .B(net667),
    .Y(_00004_));
 sg13g2_nor2_1 _18352_ (.A(_09622_),
    .B(_09624_),
    .Y(_00007_));
 sg13g2_inv_1 _18353_ (.Y(_11548_),
    .A(_09598_));
 sg13g2_nor3_1 _18354_ (.A(_11548_),
    .B(net690),
    .C(net128),
    .Y(_00008_));
 sg13g2_buf_2 _18355_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11549_));
 sg13g2_buf_1 _18356_ (.A(net761),
    .X(_11550_));
 sg13g2_and2_1 _18357_ (.A(_11549_),
    .B(_11550_),
    .X(_00003_));
 sg13g2_buf_1 _18358_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11551_));
 sg13g2_and2_1 _18359_ (.A(_11551_),
    .B(net759),
    .X(_00002_));
 sg13g2_inv_1 _18360_ (.Y(_11552_),
    .A(_09593_));
 sg13g2_nor3_1 _18361_ (.A(_11552_),
    .B(_09097_),
    .C(net584),
    .Y(_00001_));
 sg13g2_inv_2 _18362_ (.Y(_11553_),
    .A(_08592_));
 sg13g2_nor2_1 _18363_ (.A(_10822_),
    .B(_10857_),
    .Y(_11554_));
 sg13g2_nor4_1 _18364_ (.A(_10742_),
    .B(_10646_),
    .C(_10942_),
    .D(_10960_),
    .Y(_11555_));
 sg13g2_inv_1 _18365_ (.Y(_11556_),
    .A(_10765_));
 sg13g2_and2_1 _18366_ (.A(_10541_),
    .B(_10611_),
    .X(_11557_));
 sg13g2_buf_1 _18367_ (.A(_11557_),
    .X(_11558_));
 sg13g2_nor4_1 _18368_ (.A(_11556_),
    .B(_11558_),
    .C(_10795_),
    .D(_10922_),
    .Y(_11559_));
 sg13g2_nand3_1 _18369_ (.B(_11555_),
    .C(_11559_),
    .A(_11554_),
    .Y(_11560_));
 sg13g2_or4_1 _18370_ (.A(_10711_),
    .B(_10979_),
    .C(_10997_),
    .D(_10874_),
    .X(_11561_));
 sg13g2_nor3_1 _18371_ (.A(_10676_),
    .B(_11560_),
    .C(_11561_),
    .Y(_11562_));
 sg13g2_o21ai_1 _18372_ (.B1(_10898_),
    .Y(_11563_),
    .A1(\cpu.cond[1] ),
    .A2(_11562_));
 sg13g2_xnor2_1 _18373_ (.Y(_11564_),
    .A(_11553_),
    .B(_11563_));
 sg13g2_inv_1 _18374_ (.Y(_11565_),
    .A(_10521_));
 sg13g2_a21o_1 _18375_ (.A2(_11564_),
    .A1(_10503_),
    .B1(_11565_),
    .X(_11566_));
 sg13g2_buf_1 _18376_ (.A(_11566_),
    .X(_11567_));
 sg13g2_nor2b_1 _18377_ (.A(\cpu.dec.jmp ),
    .B_N(_11567_),
    .Y(_11568_));
 sg13g2_nor2b_1 _18378_ (.A(_11568_),
    .B_N(net646),
    .Y(_00053_));
 sg13g2_buf_2 _18379_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11569_));
 sg13g2_and2_1 _18380_ (.A(_11569_),
    .B(net759),
    .X(_00009_));
 sg13g2_buf_2 _18381_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11570_));
 sg13g2_and2_1 _18382_ (.A(_11570_),
    .B(net759),
    .X(_00010_));
 sg13g2_and3_1 _18383_ (.X(_00005_),
    .A(net1082),
    .B(net759),
    .C(_09587_));
 sg13g2_buf_1 _18384_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11571_));
 sg13g2_and2_1 _18385_ (.A(_11571_),
    .B(net759),
    .X(_00006_));
 sg13g2_and2_1 _18386_ (.A(net112),
    .B(_09093_),
    .X(_00052_));
 sg13g2_nor3_1 _18387_ (.A(_09045_),
    .B(net1083),
    .C(_09088_),
    .Y(_11572_));
 sg13g2_nand2_1 _18388_ (.Y(_11573_),
    .A(_09032_),
    .B(_11572_));
 sg13g2_o21ai_1 _18389_ (.B1(net406),
    .Y(_11574_),
    .A1(net1017),
    .A2(net1083));
 sg13g2_nand3_1 _18390_ (.B(_11573_),
    .C(_11574_),
    .A(_09034_),
    .Y(_11575_));
 sg13g2_buf_1 _18391_ (.A(_11575_),
    .X(_11576_));
 sg13g2_inv_1 _18392_ (.Y(_11577_),
    .A(_00226_));
 sg13g2_nor3_2 _18393_ (.A(_09092_),
    .B(_09088_),
    .C(_11577_),
    .Y(_11578_));
 sg13g2_buf_1 _18394_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11579_));
 sg13g2_buf_1 _18395_ (.A(_11579_),
    .X(_11580_));
 sg13g2_inv_1 _18396_ (.Y(_11581_),
    .A(_00282_));
 sg13g2_buf_1 _18397_ (.A(\cpu.spi.r_src[2] ),
    .X(_11582_));
 sg13g2_buf_1 _18398_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11583_));
 sg13g2_inv_1 _18399_ (.Y(_11584_),
    .A(_11583_));
 sg13g2_mux2_1 _18400_ (.A0(_11581_),
    .A1(_11582_),
    .S(_11584_),
    .X(_11585_));
 sg13g2_buf_1 _18401_ (.A(_11583_),
    .X(_11586_));
 sg13g2_buf_1 _18402_ (.A(net987),
    .X(_11587_));
 sg13g2_nand2_1 _18403_ (.Y(_11588_),
    .A(net853),
    .B(_00283_));
 sg13g2_o21ai_1 _18404_ (.B1(_11588_),
    .Y(_11589_),
    .A1(net853),
    .A2(_11581_));
 sg13g2_nor2_1 _18405_ (.A(net988),
    .B(_11589_),
    .Y(_11590_));
 sg13g2_a21oi_2 _18406_ (.B1(_11590_),
    .Y(_11591_),
    .A2(_11585_),
    .A1(_11580_));
 sg13g2_nor2_1 _18407_ (.A(_11578_),
    .B(_11591_),
    .Y(_11592_));
 sg13g2_nor2_1 _18408_ (.A(net1017),
    .B(_09088_),
    .Y(_11593_));
 sg13g2_inv_1 _18409_ (.Y(_11594_),
    .A(_11579_));
 sg13g2_buf_1 _18410_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11595_));
 sg13g2_buf_1 _18411_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11596_));
 sg13g2_mux2_1 _18412_ (.A0(_11595_),
    .A1(_11596_),
    .S(net853),
    .X(_11597_));
 sg13g2_nor2_1 _18413_ (.A(_11594_),
    .B(_11583_),
    .Y(_11598_));
 sg13g2_buf_1 _18414_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11599_));
 sg13g2_a22oi_1 _18415_ (.Y(_11600_),
    .B1(_11598_),
    .B2(_11599_),
    .A2(_11597_),
    .A1(_11594_));
 sg13g2_xnor2_1 _18416_ (.Y(_11601_),
    .A(_11593_),
    .B(_11600_));
 sg13g2_buf_1 _18417_ (.A(_09733_),
    .X(_11602_));
 sg13g2_buf_1 _18418_ (.A(net875),
    .X(_11603_));
 sg13g2_buf_1 _18419_ (.A(net726),
    .X(_11604_));
 sg13g2_nand2_1 _18420_ (.Y(_11605_),
    .A(net644),
    .B(_00283_));
 sg13g2_o21ai_1 _18421_ (.B1(_11605_),
    .Y(_11606_),
    .A1(net644),
    .A2(_11581_));
 sg13g2_buf_1 _18422_ (.A(_09163_),
    .X(_11607_));
 sg13g2_nand3_1 _18423_ (.B(net851),
    .C(_11582_),
    .A(net852),
    .Y(_11608_));
 sg13g2_o21ai_1 _18424_ (.B1(_11608_),
    .Y(_11609_),
    .A1(net852),
    .A2(_11606_));
 sg13g2_and2_1 _18425_ (.A(_11578_),
    .B(_11609_),
    .X(_11610_));
 sg13g2_buf_1 _18426_ (.A(net852),
    .X(_11611_));
 sg13g2_buf_1 _18427_ (.A(net725),
    .X(_11612_));
 sg13g2_buf_2 _18428_ (.A(net644),
    .X(_11613_));
 sg13g2_buf_1 _18429_ (.A(net644),
    .X(_11614_));
 sg13g2_nand2b_1 _18430_ (.Y(_11615_),
    .B(net572),
    .A_N(_11595_));
 sg13g2_o21ai_1 _18431_ (.B1(_11615_),
    .Y(_11616_),
    .A1(net573),
    .A2(_11599_));
 sg13g2_buf_1 _18432_ (.A(net644),
    .X(_11617_));
 sg13g2_mux2_1 _18433_ (.A0(_11595_),
    .A1(_11596_),
    .S(_11617_),
    .X(_11618_));
 sg13g2_nor2_1 _18434_ (.A(net643),
    .B(_11618_),
    .Y(_11619_));
 sg13g2_a21oi_1 _18435_ (.A1(net643),
    .A2(_11616_),
    .Y(_11620_),
    .B1(_11619_));
 sg13g2_a22oi_1 _18436_ (.Y(_11621_),
    .B1(_11610_),
    .B2(_11620_),
    .A2(_11601_),
    .A1(_11592_));
 sg13g2_nor2_1 _18437_ (.A(_11592_),
    .B(_11610_),
    .Y(_11622_));
 sg13g2_buf_1 _18438_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11623_));
 sg13g2_o21ai_1 _18439_ (.B1(_11623_),
    .Y(_11624_),
    .A1(_11576_),
    .A2(_11622_));
 sg13g2_o21ai_1 _18440_ (.B1(_11624_),
    .Y(_00318_),
    .A1(_11576_),
    .A2(_11621_));
 sg13g2_nor2b_1 _18441_ (.A(_11576_),
    .B_N(_11622_),
    .Y(_11625_));
 sg13g2_or3_1 _18442_ (.A(_09092_),
    .B(_09088_),
    .C(_11577_),
    .X(_11626_));
 sg13g2_buf_1 _18443_ (.A(_11626_),
    .X(_11627_));
 sg13g2_and2_1 _18444_ (.A(_11578_),
    .B(_11620_),
    .X(_11628_));
 sg13g2_a21oi_1 _18445_ (.A1(net850),
    .A2(_11601_),
    .Y(_11629_),
    .B1(_11628_));
 sg13g2_buf_1 _18446_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11630_));
 sg13g2_nor2_1 _18447_ (.A(net1068),
    .B(_11625_),
    .Y(_11631_));
 sg13g2_a21oi_1 _18448_ (.A1(_11625_),
    .A2(_11629_),
    .Y(_00319_),
    .B1(_11631_));
 sg13g2_buf_1 _18449_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11632_));
 sg13g2_mux2_1 _18450_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_09856_),
    .S(net878),
    .X(_11633_));
 sg13g2_nor2_1 _18451_ (.A(_11584_),
    .B(\cpu.spi.r_mode[1][0] ),
    .Y(_11634_));
 sg13g2_a21oi_1 _18452_ (.A1(_11584_),
    .A2(_00224_),
    .Y(_11635_),
    .B1(_11634_));
 sg13g2_a22oi_1 _18453_ (.Y(_11636_),
    .B1(_11635_),
    .B2(_11594_),
    .A2(_11598_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18454_ (.A(_11636_),
    .X(_11637_));
 sg13g2_buf_1 _18455_ (.A(_11637_),
    .X(_11638_));
 sg13g2_nand3_1 _18456_ (.B(_09086_),
    .C(net520),
    .A(net1084),
    .Y(_11639_));
 sg13g2_o21ai_1 _18457_ (.B1(_11639_),
    .Y(_11640_),
    .A1(net1016),
    .A2(_11572_));
 sg13g2_nand2_1 _18458_ (.Y(_11641_),
    .A(net405),
    .B(_11637_));
 sg13g2_a21o_1 _18459_ (.A2(_09052_),
    .A1(_00221_),
    .B1(net1083),
    .X(_11642_));
 sg13g2_o21ai_1 _18460_ (.B1(net1083),
    .Y(_11643_),
    .A1(_08940_),
    .A2(_11637_));
 sg13g2_nand2_1 _18461_ (.Y(_11644_),
    .A(_09089_),
    .B(_11643_));
 sg13g2_o21ai_1 _18462_ (.B1(_11644_),
    .Y(_11645_),
    .A1(_11641_),
    .A2(_11642_));
 sg13g2_nand3_1 _18463_ (.B(_11640_),
    .C(_11645_),
    .A(net879),
    .Y(_11646_));
 sg13g2_nor2_1 _18464_ (.A(_11591_),
    .B(_11646_),
    .Y(_11647_));
 sg13g2_mux2_1 _18465_ (.A0(_11632_),
    .A1(_11633_),
    .S(_11647_),
    .X(_00320_));
 sg13g2_buf_1 _18466_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_11648_));
 sg13g2_inv_1 _18467_ (.Y(_11649_),
    .A(_11591_));
 sg13g2_nor2_1 _18468_ (.A(_11649_),
    .B(_11646_),
    .Y(_11650_));
 sg13g2_mux2_1 _18469_ (.A0(_11648_),
    .A1(_11633_),
    .S(_11650_),
    .X(_00321_));
 sg13g2_nand2_1 _18470_ (.Y(_11651_),
    .A(net760),
    .B(_09143_));
 sg13g2_buf_2 _18471_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_11652_));
 sg13g2_buf_1 _18472_ (.A(\cpu.d_wstrobe_d ),
    .X(_11653_));
 sg13g2_buf_1 _18473_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_11654_));
 sg13g2_buf_2 _18474_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_11655_));
 sg13g2_and2_1 _18475_ (.A(_11654_),
    .B(_11655_),
    .X(_11656_));
 sg13g2_buf_1 _18476_ (.A(_11656_),
    .X(_11657_));
 sg13g2_and3_1 _18477_ (.X(_11658_),
    .A(_11652_),
    .B(_11653_),
    .C(_11657_));
 sg13g2_buf_1 _18478_ (.A(_11658_),
    .X(_11659_));
 sg13g2_nor3_1 _18479_ (.A(_09131_),
    .B(_08536_),
    .C(_09572_),
    .Y(_11660_));
 sg13g2_o21ai_1 _18480_ (.B1(_11660_),
    .Y(_11661_),
    .A1(_09568_),
    .A2(_11659_));
 sg13g2_buf_1 _18481_ (.A(_11661_),
    .X(_11662_));
 sg13g2_or2_1 _18482_ (.X(_11663_),
    .B(_11662_),
    .A(_11651_));
 sg13g2_buf_1 _18483_ (.A(_11663_),
    .X(_11664_));
 sg13g2_buf_1 _18484_ (.A(_08534_),
    .X(_11665_));
 sg13g2_nand2b_1 _18485_ (.Y(_11666_),
    .B(\cpu.ex.r_wmask[1] ),
    .A_N(net986));
 sg13g2_buf_2 _18486_ (.A(_11666_),
    .X(_11667_));
 sg13g2_buf_2 _18487_ (.A(_00275_),
    .X(_11668_));
 sg13g2_o21ai_1 _18488_ (.B1(_11668_),
    .Y(_11669_),
    .A1(_08535_),
    .A2(_11667_));
 sg13g2_nor2_1 _18489_ (.A(_11664_),
    .B(_11669_),
    .Y(_11670_));
 sg13g2_buf_2 _18490_ (.A(_11670_),
    .X(_11671_));
 sg13g2_buf_1 _18491_ (.A(_11671_),
    .X(_11672_));
 sg13g2_buf_1 _18492_ (.A(uio_in[0]),
    .X(_11673_));
 sg13g2_buf_1 _18493_ (.A(_11673_),
    .X(_11674_));
 sg13g2_buf_1 _18494_ (.A(_11651_),
    .X(_11675_));
 sg13g2_buf_1 _18495_ (.A(_11653_),
    .X(_11676_));
 sg13g2_buf_1 _18496_ (.A(_00276_),
    .X(_11677_));
 sg13g2_buf_1 _18497_ (.A(_11677_),
    .X(_11678_));
 sg13g2_nor2b_1 _18498_ (.A(_11654_),
    .B_N(_11655_),
    .Y(_11679_));
 sg13g2_buf_1 _18499_ (.A(_11679_),
    .X(_11680_));
 sg13g2_nand3_1 _18500_ (.B(net984),
    .C(_11680_),
    .A(net985),
    .Y(_11681_));
 sg13g2_buf_2 _18501_ (.A(_11681_),
    .X(_11682_));
 sg13g2_nor2_1 _18502_ (.A(net570),
    .B(_11682_),
    .Y(_11683_));
 sg13g2_buf_2 _18503_ (.A(_11683_),
    .X(_11684_));
 sg13g2_mux2_1 _18504_ (.A0(\cpu.dcache.r_data[0][0] ),
    .A1(net1065),
    .S(_11684_),
    .X(_11685_));
 sg13g2_nor2_1 _18505_ (.A(_11671_),
    .B(_11685_),
    .Y(_11686_));
 sg13g2_a21oi_1 _18506_ (.A1(net745),
    .A2(net67),
    .Y(_00322_),
    .B1(_11686_));
 sg13g2_buf_1 _18507_ (.A(net744),
    .X(_11687_));
 sg13g2_inv_2 _18508_ (.Y(_11688_),
    .A(_11668_));
 sg13g2_mux2_1 _18509_ (.A0(net642),
    .A1(net983),
    .S(_08560_),
    .X(_11689_));
 sg13g2_or3_1 _18510_ (.A(_11664_),
    .B(_11667_),
    .C(_11689_),
    .X(_11690_));
 sg13g2_buf_2 _18511_ (.A(_11690_),
    .X(_11691_));
 sg13g2_buf_1 _18512_ (.A(_11691_),
    .X(_11692_));
 sg13g2_buf_1 _18513_ (.A(uio_in[2]),
    .X(_11693_));
 sg13g2_buf_1 _18514_ (.A(_11693_),
    .X(_11694_));
 sg13g2_buf_2 _18515_ (.A(net1064),
    .X(_11695_));
 sg13g2_nand3_1 _18516_ (.B(net984),
    .C(_11657_),
    .A(net985),
    .Y(_11696_));
 sg13g2_buf_2 _18517_ (.A(_11696_),
    .X(_11697_));
 sg13g2_nor2_1 _18518_ (.A(net570),
    .B(_11697_),
    .Y(_11698_));
 sg13g2_buf_2 _18519_ (.A(_11698_),
    .X(_11699_));
 sg13g2_nor2b_1 _18520_ (.A(_11699_),
    .B_N(\cpu.dcache.r_data[0][10] ),
    .Y(_11700_));
 sg13g2_a21oi_1 _18521_ (.A1(net982),
    .A2(_11699_),
    .Y(_11701_),
    .B1(_11700_));
 sg13g2_inv_2 _18522_ (.Y(_11702_),
    .A(\cpu.dcache.wdata[10] ));
 sg13g2_or2_1 _18523_ (.X(_11703_),
    .B(_11667_),
    .A(_08560_));
 sg13g2_buf_1 _18524_ (.A(_11703_),
    .X(_11704_));
 sg13g2_nand2_1 _18525_ (.Y(_11705_),
    .A(_09825_),
    .B(_11704_));
 sg13g2_o21ai_1 _18526_ (.B1(_11705_),
    .Y(_11706_),
    .A1(_11702_),
    .A2(_11704_));
 sg13g2_buf_2 _18527_ (.A(_11706_),
    .X(_11707_));
 sg13g2_buf_1 _18528_ (.A(_11707_),
    .X(_11708_));
 sg13g2_nor2_1 _18529_ (.A(net360),
    .B(_11691_),
    .Y(_11709_));
 sg13g2_a21oi_1 _18530_ (.A1(net66),
    .A2(_11701_),
    .Y(_00323_),
    .B1(_11709_));
 sg13g2_buf_1 _18531_ (.A(uio_in[3]),
    .X(_11710_));
 sg13g2_buf_1 _18532_ (.A(_11710_),
    .X(_11711_));
 sg13g2_buf_2 _18533_ (.A(net1063),
    .X(_11712_));
 sg13g2_nor2b_1 _18534_ (.A(_11699_),
    .B_N(\cpu.dcache.r_data[0][11] ),
    .Y(_11713_));
 sg13g2_a21oi_1 _18535_ (.A1(net981),
    .A2(_11699_),
    .Y(_11714_),
    .B1(_11713_));
 sg13g2_inv_1 _18536_ (.Y(_11715_),
    .A(net1078));
 sg13g2_buf_1 _18537_ (.A(_11715_),
    .X(_11716_));
 sg13g2_nor2_1 _18538_ (.A(_08560_),
    .B(_11667_),
    .Y(_11717_));
 sg13g2_buf_1 _18539_ (.A(_11717_),
    .X(_11718_));
 sg13g2_nand2_1 _18540_ (.Y(_11719_),
    .A(_09937_),
    .B(net569));
 sg13g2_o21ai_1 _18541_ (.B1(_11719_),
    .Y(_11720_),
    .A1(_11716_),
    .A2(net569));
 sg13g2_buf_2 _18542_ (.A(_11720_),
    .X(_11721_));
 sg13g2_buf_1 _18543_ (.A(_11721_),
    .X(_11722_));
 sg13g2_nor2_1 _18544_ (.A(_11691_),
    .B(net359),
    .Y(_11723_));
 sg13g2_a21oi_1 _18545_ (.A1(net66),
    .A2(_11714_),
    .Y(_00324_),
    .B1(_11723_));
 sg13g2_and2_1 _18546_ (.A(_09942_),
    .B(net569),
    .X(_11724_));
 sg13g2_a21oi_1 _18547_ (.A1(_09839_),
    .A2(_11704_),
    .Y(_11725_),
    .B1(_11724_));
 sg13g2_buf_2 _18548_ (.A(_11725_),
    .X(_11726_));
 sg13g2_buf_1 _18549_ (.A(_11726_),
    .X(_11727_));
 sg13g2_buf_1 _18550_ (.A(_11673_),
    .X(_11728_));
 sg13g2_buf_1 _18551_ (.A(_11655_),
    .X(_11729_));
 sg13g2_buf_1 _18552_ (.A(_11654_),
    .X(_11730_));
 sg13g2_nor2b_1 _18553_ (.A(net980),
    .B_N(_11730_),
    .Y(_11731_));
 sg13g2_nand3_1 _18554_ (.B(net984),
    .C(_11731_),
    .A(net985),
    .Y(_11732_));
 sg13g2_buf_4 _18555_ (.X(_11733_),
    .A(_11732_));
 sg13g2_nor2_2 _18556_ (.A(_11675_),
    .B(_11733_),
    .Y(_11734_));
 sg13g2_mux2_1 _18557_ (.A0(\cpu.dcache.r_data[0][12] ),
    .A1(_11728_),
    .S(_11734_),
    .X(_11735_));
 sg13g2_nand2_1 _18558_ (.Y(_11736_),
    .A(net66),
    .B(_11735_));
 sg13g2_o21ai_1 _18559_ (.B1(_11736_),
    .Y(_00325_),
    .A1(net66),
    .A2(net358));
 sg13g2_inv_2 _18560_ (.Y(_11737_),
    .A(\cpu.dcache.wdata[13] ));
 sg13g2_nor2_1 _18561_ (.A(_11737_),
    .B(_11704_),
    .Y(_11738_));
 sg13g2_a21oi_1 _18562_ (.A1(_09845_),
    .A2(_11704_),
    .Y(_11739_),
    .B1(_11738_));
 sg13g2_buf_2 _18563_ (.A(_11739_),
    .X(_11740_));
 sg13g2_buf_1 _18564_ (.A(_11740_),
    .X(_11741_));
 sg13g2_buf_1 _18565_ (.A(uio_in[1]),
    .X(_11742_));
 sg13g2_buf_1 _18566_ (.A(_11742_),
    .X(_11743_));
 sg13g2_mux2_1 _18567_ (.A0(\cpu.dcache.r_data[0][13] ),
    .A1(net1061),
    .S(_11734_),
    .X(_11744_));
 sg13g2_nand2_1 _18568_ (.Y(_11745_),
    .A(net66),
    .B(_11744_));
 sg13g2_o21ai_1 _18569_ (.B1(_11745_),
    .Y(_00326_),
    .A1(net66),
    .A2(net357));
 sg13g2_inv_1 _18570_ (.Y(_11746_),
    .A(_09851_));
 sg13g2_inv_2 _18571_ (.Y(_11747_),
    .A(\cpu.dcache.wdata[14] ));
 sg13g2_mux2_1 _18572_ (.A0(_11746_),
    .A1(_11747_),
    .S(net569),
    .X(_11748_));
 sg13g2_buf_2 _18573_ (.A(_11748_),
    .X(_11749_));
 sg13g2_buf_1 _18574_ (.A(_11749_),
    .X(_11750_));
 sg13g2_buf_1 _18575_ (.A(net1064),
    .X(_11751_));
 sg13g2_mux2_1 _18576_ (.A0(\cpu.dcache.r_data[0][14] ),
    .A1(net978),
    .S(_11734_),
    .X(_11752_));
 sg13g2_nand2_1 _18577_ (.Y(_11753_),
    .A(_11691_),
    .B(_11752_));
 sg13g2_o21ai_1 _18578_ (.B1(_11753_),
    .Y(_00327_),
    .A1(net66),
    .A2(net397));
 sg13g2_inv_1 _18579_ (.Y(_11754_),
    .A(_09856_));
 sg13g2_buf_1 _18580_ (.A(_11754_),
    .X(_11755_));
 sg13g2_nor2_1 _18581_ (.A(_11755_),
    .B(net569),
    .Y(_11756_));
 sg13g2_a21oi_1 _18582_ (.A1(_09958_),
    .A2(_11718_),
    .Y(_11757_),
    .B1(_11756_));
 sg13g2_buf_2 _18583_ (.A(_11757_),
    .X(_11758_));
 sg13g2_buf_1 _18584_ (.A(_11758_),
    .X(_11759_));
 sg13g2_buf_1 _18585_ (.A(net1063),
    .X(_11760_));
 sg13g2_mux2_1 _18586_ (.A0(\cpu.dcache.r_data[0][15] ),
    .A1(_11760_),
    .S(_11734_),
    .X(_11761_));
 sg13g2_nand2_1 _18587_ (.Y(_11762_),
    .A(_11691_),
    .B(_11761_));
 sg13g2_o21ai_1 _18588_ (.B1(_11762_),
    .Y(_00328_),
    .A1(net66),
    .A2(net356));
 sg13g2_o21ai_1 _18589_ (.B1(net642),
    .Y(_11763_),
    .A1(_08535_),
    .A2(_11667_));
 sg13g2_nor2_1 _18590_ (.A(_11664_),
    .B(_11763_),
    .Y(_11764_));
 sg13g2_buf_2 _18591_ (.A(_11764_),
    .X(_11765_));
 sg13g2_buf_1 _18592_ (.A(_11765_),
    .X(_11766_));
 sg13g2_buf_1 _18593_ (.A(_11652_),
    .X(_11767_));
 sg13g2_nand3_1 _18594_ (.B(net985),
    .C(_11680_),
    .A(net976),
    .Y(_11768_));
 sg13g2_buf_2 _18595_ (.A(_11768_),
    .X(_11769_));
 sg13g2_nor2_1 _18596_ (.A(net570),
    .B(_11769_),
    .Y(_11770_));
 sg13g2_buf_2 _18597_ (.A(_11770_),
    .X(_11771_));
 sg13g2_mux2_1 _18598_ (.A0(\cpu.dcache.r_data[0][16] ),
    .A1(net1065),
    .S(_11771_),
    .X(_11772_));
 sg13g2_nor2_1 _18599_ (.A(_11765_),
    .B(_11772_),
    .Y(_11773_));
 sg13g2_a21oi_1 _18600_ (.A1(net745),
    .A2(net65),
    .Y(_00329_),
    .B1(_11773_));
 sg13g2_buf_1 _18601_ (.A(_11742_),
    .X(_11774_));
 sg13g2_buf_1 _18602_ (.A(net1060),
    .X(_11775_));
 sg13g2_nor2b_1 _18603_ (.A(_11771_),
    .B_N(\cpu.dcache.r_data[0][17] ),
    .Y(_11776_));
 sg13g2_a21oi_1 _18604_ (.A1(net975),
    .A2(_11771_),
    .Y(_11777_),
    .B1(_11776_));
 sg13g2_buf_1 _18605_ (.A(net1009),
    .X(_11778_));
 sg13g2_nand2_1 _18606_ (.Y(_11779_),
    .A(net847),
    .B(net65));
 sg13g2_o21ai_1 _18607_ (.B1(_11779_),
    .Y(_00330_),
    .A1(net65),
    .A2(_11777_));
 sg13g2_buf_1 _18608_ (.A(net1064),
    .X(_11780_));
 sg13g2_nor2b_1 _18609_ (.A(_11771_),
    .B_N(\cpu.dcache.r_data[0][18] ),
    .Y(_11781_));
 sg13g2_a21oi_1 _18610_ (.A1(net974),
    .A2(_11771_),
    .Y(_11782_),
    .B1(_11781_));
 sg13g2_buf_1 _18611_ (.A(net1008),
    .X(_11783_));
 sg13g2_nand2_1 _18612_ (.Y(_11784_),
    .A(net846),
    .B(net65));
 sg13g2_o21ai_1 _18613_ (.B1(_11784_),
    .Y(_00331_),
    .A1(net65),
    .A2(_11782_));
 sg13g2_buf_1 _18614_ (.A(net849),
    .X(_11785_));
 sg13g2_buf_1 _18615_ (.A(net1063),
    .X(_11786_));
 sg13g2_mux2_1 _18616_ (.A0(\cpu.dcache.r_data[0][19] ),
    .A1(net973),
    .S(_11771_),
    .X(_11787_));
 sg13g2_nor2_1 _18617_ (.A(_11765_),
    .B(_11787_),
    .Y(_11788_));
 sg13g2_a21oi_1 _18618_ (.A1(net724),
    .A2(net65),
    .Y(_00332_),
    .B1(_11788_));
 sg13g2_nor2b_1 _18619_ (.A(_11684_),
    .B_N(\cpu.dcache.r_data[0][1] ),
    .Y(_11789_));
 sg13g2_a21oi_1 _18620_ (.A1(net975),
    .A2(_11684_),
    .Y(_11790_),
    .B1(_11789_));
 sg13g2_nand2_1 _18621_ (.Y(_11791_),
    .A(_11778_),
    .B(net67));
 sg13g2_o21ai_1 _18622_ (.B1(_11791_),
    .Y(_00333_),
    .A1(net67),
    .A2(_11790_));
 sg13g2_buf_1 _18623_ (.A(_11673_),
    .X(_11792_));
 sg13g2_buf_1 _18624_ (.A(net1059),
    .X(_11793_));
 sg13g2_nor2_1 _18625_ (.A(_11654_),
    .B(_11655_),
    .Y(_11794_));
 sg13g2_nand3_1 _18626_ (.B(net985),
    .C(_11794_),
    .A(net976),
    .Y(_11795_));
 sg13g2_buf_2 _18627_ (.A(_11795_),
    .X(_11796_));
 sg13g2_nor2_1 _18628_ (.A(net570),
    .B(_11796_),
    .Y(_11797_));
 sg13g2_buf_2 _18629_ (.A(_11797_),
    .X(_11798_));
 sg13g2_nor2b_1 _18630_ (.A(_11798_),
    .B_N(\cpu.dcache.r_data[0][20] ),
    .Y(_11799_));
 sg13g2_a21oi_1 _18631_ (.A1(net972),
    .A2(_11798_),
    .Y(_11800_),
    .B1(_11799_));
 sg13g2_buf_1 _18632_ (.A(_09839_),
    .X(_11801_));
 sg13g2_nand2_1 _18633_ (.Y(_11802_),
    .A(net971),
    .B(_11765_));
 sg13g2_o21ai_1 _18634_ (.B1(_11802_),
    .Y(_00334_),
    .A1(_11766_),
    .A2(_11800_));
 sg13g2_buf_1 _18635_ (.A(_11774_),
    .X(_11803_));
 sg13g2_nor2b_1 _18636_ (.A(_11798_),
    .B_N(\cpu.dcache.r_data[0][21] ),
    .Y(_11804_));
 sg13g2_a21oi_1 _18637_ (.A1(net970),
    .A2(_11798_),
    .Y(_11805_),
    .B1(_11804_));
 sg13g2_buf_1 _18638_ (.A(_09845_),
    .X(_11806_));
 sg13g2_nand2_1 _18639_ (.Y(_11807_),
    .A(net969),
    .B(_11765_));
 sg13g2_o21ai_1 _18640_ (.B1(_11807_),
    .Y(_00335_),
    .A1(net65),
    .A2(_11805_));
 sg13g2_buf_1 _18641_ (.A(_11746_),
    .X(_11808_));
 sg13g2_buf_1 _18642_ (.A(net845),
    .X(_11809_));
 sg13g2_buf_1 _18643_ (.A(_11693_),
    .X(_11810_));
 sg13g2_mux2_1 _18644_ (.A0(\cpu.dcache.r_data[0][22] ),
    .A1(net1058),
    .S(_11798_),
    .X(_11811_));
 sg13g2_nor2_1 _18645_ (.A(_11765_),
    .B(_11811_),
    .Y(_11812_));
 sg13g2_a21oi_1 _18646_ (.A1(net723),
    .A2(net65),
    .Y(_00336_),
    .B1(_11812_));
 sg13g2_buf_1 _18647_ (.A(net848),
    .X(_11813_));
 sg13g2_mux2_1 _18648_ (.A0(\cpu.dcache.r_data[0][23] ),
    .A1(net973),
    .S(_11798_),
    .X(_11814_));
 sg13g2_nor2_1 _18649_ (.A(_11765_),
    .B(_11814_),
    .Y(_11815_));
 sg13g2_a21oi_1 _18650_ (.A1(net722),
    .A2(_11766_),
    .Y(_00337_),
    .B1(_11815_));
 sg13g2_nand2_1 _18651_ (.Y(_11816_),
    .A(_09921_),
    .B(net569));
 sg13g2_o21ai_1 _18652_ (.B1(_11816_),
    .Y(_11817_),
    .A1(_09809_),
    .A2(net569));
 sg13g2_buf_2 _18653_ (.A(_11817_),
    .X(_11818_));
 sg13g2_buf_1 _18654_ (.A(_11818_),
    .X(_11819_));
 sg13g2_nand2b_1 _18655_ (.Y(_11820_),
    .B(_11659_),
    .A_N(net570));
 sg13g2_buf_1 _18656_ (.A(_11820_),
    .X(_11821_));
 sg13g2_mux2_1 _18657_ (.A0(_11674_),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net459),
    .X(_11822_));
 sg13g2_nor2_1 _18658_ (.A(_08535_),
    .B(net642),
    .Y(_11823_));
 sg13g2_nor2_1 _18659_ (.A(_08560_),
    .B(net983),
    .Y(_11824_));
 sg13g2_or4_1 _18660_ (.A(_11664_),
    .B(_11667_),
    .C(_11823_),
    .D(_11824_),
    .X(_11825_));
 sg13g2_buf_1 _18661_ (.A(_11825_),
    .X(_11826_));
 sg13g2_buf_1 _18662_ (.A(_11826_),
    .X(_11827_));
 sg13g2_mux2_1 _18663_ (.A0(net355),
    .A1(_11822_),
    .S(net64),
    .X(_00338_));
 sg13g2_mux2_1 _18664_ (.A0(_09818_),
    .A1(_09926_),
    .S(net569),
    .X(_11828_));
 sg13g2_buf_2 _18665_ (.A(_11828_),
    .X(_11829_));
 sg13g2_buf_1 _18666_ (.A(_11829_),
    .X(_11830_));
 sg13g2_mux2_1 _18667_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net459),
    .X(_11831_));
 sg13g2_mux2_1 _18668_ (.A0(net396),
    .A1(_11831_),
    .S(net64),
    .X(_00339_));
 sg13g2_mux2_1 _18669_ (.A0(net1058),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net459),
    .X(_11832_));
 sg13g2_mux2_1 _18670_ (.A0(net360),
    .A1(_11832_),
    .S(_11827_),
    .X(_00340_));
 sg13g2_buf_1 _18671_ (.A(_11710_),
    .X(_11833_));
 sg13g2_mux2_1 _18672_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(net459),
    .X(_11834_));
 sg13g2_mux2_1 _18673_ (.A0(net359),
    .A1(_11834_),
    .S(_11827_),
    .X(_00341_));
 sg13g2_nand3_1 _18674_ (.B(net985),
    .C(_11731_),
    .A(net976),
    .Y(_11835_));
 sg13g2_buf_4 _18675_ (.X(_11836_),
    .A(_11835_));
 sg13g2_nor2_2 _18676_ (.A(_11675_),
    .B(_11836_),
    .Y(_11837_));
 sg13g2_mux2_1 _18677_ (.A0(\cpu.dcache.r_data[0][28] ),
    .A1(net1062),
    .S(_11837_),
    .X(_11838_));
 sg13g2_nand2_1 _18678_ (.Y(_11839_),
    .A(net64),
    .B(_11838_));
 sg13g2_o21ai_1 _18679_ (.B1(_11839_),
    .Y(_00342_),
    .A1(_11727_),
    .A2(net64));
 sg13g2_mux2_1 _18680_ (.A0(\cpu.dcache.r_data[0][29] ),
    .A1(net1061),
    .S(_11837_),
    .X(_11840_));
 sg13g2_nand2_1 _18681_ (.Y(_11841_),
    .A(net64),
    .B(_11840_));
 sg13g2_o21ai_1 _18682_ (.B1(_11841_),
    .Y(_00343_),
    .A1(_11741_),
    .A2(net64));
 sg13g2_nor2b_1 _18683_ (.A(_11684_),
    .B_N(\cpu.dcache.r_data[0][2] ),
    .Y(_11842_));
 sg13g2_a21oi_1 _18684_ (.A1(net974),
    .A2(_11684_),
    .Y(_11843_),
    .B1(_11842_));
 sg13g2_nand2_1 _18685_ (.Y(_11844_),
    .A(net846),
    .B(net67));
 sg13g2_o21ai_1 _18686_ (.B1(_11844_),
    .Y(_00344_),
    .A1(net67),
    .A2(_11843_));
 sg13g2_buf_1 _18687_ (.A(_11693_),
    .X(_11845_));
 sg13g2_mux2_1 _18688_ (.A0(\cpu.dcache.r_data[0][30] ),
    .A1(net1056),
    .S(_11837_),
    .X(_11846_));
 sg13g2_nand2_1 _18689_ (.Y(_11847_),
    .A(_11826_),
    .B(_11846_));
 sg13g2_o21ai_1 _18690_ (.B1(_11847_),
    .Y(_00345_),
    .A1(_11750_),
    .A2(net64));
 sg13g2_mux2_1 _18691_ (.A0(\cpu.dcache.r_data[0][31] ),
    .A1(_11760_),
    .S(_11837_),
    .X(_11848_));
 sg13g2_nand2_1 _18692_ (.Y(_11849_),
    .A(_11826_),
    .B(_11848_));
 sg13g2_o21ai_1 _18693_ (.B1(_11849_),
    .Y(_00346_),
    .A1(_11759_),
    .A2(net64));
 sg13g2_mux2_1 _18694_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(_11786_),
    .S(_11684_),
    .X(_11850_));
 sg13g2_nor2_1 _18695_ (.A(_11671_),
    .B(_11850_),
    .Y(_11851_));
 sg13g2_a21oi_1 _18696_ (.A1(_11785_),
    .A2(net67),
    .Y(_00347_),
    .B1(_11851_));
 sg13g2_nand3_1 _18697_ (.B(net984),
    .C(_11794_),
    .A(net985),
    .Y(_11852_));
 sg13g2_buf_2 _18698_ (.A(_11852_),
    .X(_11853_));
 sg13g2_nor2_1 _18699_ (.A(net570),
    .B(_11853_),
    .Y(_11854_));
 sg13g2_buf_2 _18700_ (.A(_11854_),
    .X(_11855_));
 sg13g2_nor2b_1 _18701_ (.A(_11855_),
    .B_N(\cpu.dcache.r_data[0][4] ),
    .Y(_11856_));
 sg13g2_a21oi_1 _18702_ (.A1(net972),
    .A2(_11855_),
    .Y(_11857_),
    .B1(_11856_));
 sg13g2_nand2_1 _18703_ (.Y(_11858_),
    .A(net971),
    .B(_11671_));
 sg13g2_o21ai_1 _18704_ (.B1(_11858_),
    .Y(_00348_),
    .A1(_11672_),
    .A2(_11857_));
 sg13g2_nor2b_1 _18705_ (.A(_11855_),
    .B_N(\cpu.dcache.r_data[0][5] ),
    .Y(_11859_));
 sg13g2_a21oi_1 _18706_ (.A1(net970),
    .A2(_11855_),
    .Y(_11860_),
    .B1(_11859_));
 sg13g2_nand2_1 _18707_ (.Y(_11861_),
    .A(net969),
    .B(_11671_));
 sg13g2_o21ai_1 _18708_ (.B1(_11861_),
    .Y(_00349_),
    .A1(_11672_),
    .A2(_11860_));
 sg13g2_mux2_1 _18709_ (.A0(\cpu.dcache.r_data[0][6] ),
    .A1(net1058),
    .S(_11855_),
    .X(_11862_));
 sg13g2_nor2_1 _18710_ (.A(_11671_),
    .B(_11862_),
    .Y(_11863_));
 sg13g2_a21oi_1 _18711_ (.A1(_11809_),
    .A2(net67),
    .Y(_00350_),
    .B1(_11863_));
 sg13g2_mux2_1 _18712_ (.A0(\cpu.dcache.r_data[0][7] ),
    .A1(_11786_),
    .S(_11855_),
    .X(_11864_));
 sg13g2_nor2_1 _18713_ (.A(_11671_),
    .B(_11864_),
    .Y(_11865_));
 sg13g2_a21oi_1 _18714_ (.A1(net722),
    .A2(net67),
    .Y(_00351_),
    .B1(_11865_));
 sg13g2_buf_2 _18715_ (.A(net1059),
    .X(_11866_));
 sg13g2_nor2b_1 _18716_ (.A(_11699_),
    .B_N(\cpu.dcache.r_data[0][8] ),
    .Y(_11867_));
 sg13g2_a21oi_1 _18717_ (.A1(net968),
    .A2(_11699_),
    .Y(_11868_),
    .B1(_11867_));
 sg13g2_nor2_1 _18718_ (.A(_11691_),
    .B(net355),
    .Y(_11869_));
 sg13g2_a21oi_1 _18719_ (.A1(_11692_),
    .A2(_11868_),
    .Y(_00352_),
    .B1(_11869_));
 sg13g2_buf_2 _18720_ (.A(net1060),
    .X(_11870_));
 sg13g2_nor2b_1 _18721_ (.A(_11699_),
    .B_N(\cpu.dcache.r_data[0][9] ),
    .Y(_11871_));
 sg13g2_a21oi_1 _18722_ (.A1(net967),
    .A2(_11699_),
    .Y(_11872_),
    .B1(_11871_));
 sg13g2_nor2_1 _18723_ (.A(_11691_),
    .B(_11830_),
    .Y(_11873_));
 sg13g2_a21oi_1 _18724_ (.A1(_11692_),
    .A2(_11872_),
    .Y(_00353_),
    .B1(_11873_));
 sg13g2_buf_1 _18725_ (.A(_09430_),
    .X(_11874_));
 sg13g2_or2_1 _18726_ (.X(_11875_),
    .B(_11669_),
    .A(_11662_));
 sg13g2_buf_2 _18727_ (.A(_11875_),
    .X(_11876_));
 sg13g2_nor2_1 _18728_ (.A(net568),
    .B(_11876_),
    .Y(_11877_));
 sg13g2_buf_2 _18729_ (.A(_11877_),
    .X(_11878_));
 sg13g2_buf_1 _18730_ (.A(_11878_),
    .X(_11879_));
 sg13g2_nor2_1 _18731_ (.A(net568),
    .B(_11682_),
    .Y(_11880_));
 sg13g2_buf_2 _18732_ (.A(_11880_),
    .X(_11881_));
 sg13g2_mux2_1 _18733_ (.A0(\cpu.dcache.r_data[1][0] ),
    .A1(net1065),
    .S(_11881_),
    .X(_11882_));
 sg13g2_nor2_1 _18734_ (.A(_11878_),
    .B(_11882_),
    .Y(_11883_));
 sg13g2_a21oi_1 _18735_ (.A1(net745),
    .A2(net63),
    .Y(_00354_),
    .B1(_11883_));
 sg13g2_buf_1 _18736_ (.A(net534),
    .X(_11884_));
 sg13g2_buf_1 _18737_ (.A(net458),
    .X(_11885_));
 sg13g2_buf_1 _18738_ (.A(net395),
    .X(_11886_));
 sg13g2_nor3_1 _18739_ (.A(_11662_),
    .B(_11667_),
    .C(_11689_),
    .Y(_11887_));
 sg13g2_buf_2 _18740_ (.A(_11887_),
    .X(_11888_));
 sg13g2_nand2_1 _18741_ (.Y(_11889_),
    .A(net354),
    .B(_11888_));
 sg13g2_buf_1 _18742_ (.A(_11889_),
    .X(_11890_));
 sg13g2_buf_1 _18743_ (.A(_11890_),
    .X(_11891_));
 sg13g2_nor2_1 _18744_ (.A(net568),
    .B(_11697_),
    .Y(_11892_));
 sg13g2_buf_2 _18745_ (.A(_11892_),
    .X(_11893_));
 sg13g2_nor2b_1 _18746_ (.A(_11893_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_11894_));
 sg13g2_a21oi_1 _18747_ (.A1(net982),
    .A2(_11893_),
    .Y(_11895_),
    .B1(_11894_));
 sg13g2_nor2_1 _18748_ (.A(net360),
    .B(_11890_),
    .Y(_11896_));
 sg13g2_a21oi_1 _18749_ (.A1(net62),
    .A2(_11895_),
    .Y(_00355_),
    .B1(_11896_));
 sg13g2_nor2b_1 _18750_ (.A(_11893_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_11897_));
 sg13g2_a21oi_1 _18751_ (.A1(net981),
    .A2(_11893_),
    .Y(_11898_),
    .B1(_11897_));
 sg13g2_nor2_1 _18752_ (.A(net359),
    .B(_11890_),
    .Y(_11899_));
 sg13g2_a21oi_1 _18753_ (.A1(net62),
    .A2(_11898_),
    .Y(_00356_),
    .B1(_11899_));
 sg13g2_nor2_2 _18754_ (.A(_11874_),
    .B(_11733_),
    .Y(_11900_));
 sg13g2_mux2_1 _18755_ (.A0(\cpu.dcache.r_data[1][12] ),
    .A1(net1062),
    .S(_11900_),
    .X(_11901_));
 sg13g2_nand2_1 _18756_ (.Y(_11902_),
    .A(net62),
    .B(_11901_));
 sg13g2_o21ai_1 _18757_ (.B1(_11902_),
    .Y(_00357_),
    .A1(net358),
    .A2(net62));
 sg13g2_buf_1 _18758_ (.A(_11742_),
    .X(_11903_));
 sg13g2_mux2_1 _18759_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(net1055),
    .S(_11900_),
    .X(_11904_));
 sg13g2_nand2_1 _18760_ (.Y(_11905_),
    .A(net62),
    .B(_11904_));
 sg13g2_o21ai_1 _18761_ (.B1(_11905_),
    .Y(_00358_),
    .A1(net357),
    .A2(net62));
 sg13g2_mux2_1 _18762_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(net1056),
    .S(_11900_),
    .X(_11906_));
 sg13g2_nand2_1 _18763_ (.Y(_11907_),
    .A(_11890_),
    .B(_11906_));
 sg13g2_o21ai_1 _18764_ (.B1(_11907_),
    .Y(_00359_),
    .A1(net397),
    .A2(_11891_));
 sg13g2_buf_1 _18765_ (.A(_11710_),
    .X(_11908_));
 sg13g2_mux2_1 _18766_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(net1054),
    .S(_11900_),
    .X(_11909_));
 sg13g2_nand2_1 _18767_ (.Y(_11910_),
    .A(_11890_),
    .B(_11909_));
 sg13g2_o21ai_1 _18768_ (.B1(_11910_),
    .Y(_00360_),
    .A1(net356),
    .A2(net62));
 sg13g2_or2_1 _18769_ (.X(_11911_),
    .B(_11763_),
    .A(_11662_));
 sg13g2_buf_2 _18770_ (.A(_11911_),
    .X(_11912_));
 sg13g2_nor2_1 _18771_ (.A(net568),
    .B(_11912_),
    .Y(_11913_));
 sg13g2_buf_2 _18772_ (.A(_11913_),
    .X(_11914_));
 sg13g2_buf_1 _18773_ (.A(_11914_),
    .X(_11915_));
 sg13g2_nor2_1 _18774_ (.A(net568),
    .B(_11769_),
    .Y(_11916_));
 sg13g2_buf_2 _18775_ (.A(_11916_),
    .X(_11917_));
 sg13g2_mux2_1 _18776_ (.A0(\cpu.dcache.r_data[1][16] ),
    .A1(net1065),
    .S(_11917_),
    .X(_11918_));
 sg13g2_nor2_1 _18777_ (.A(_11914_),
    .B(_11918_),
    .Y(_11919_));
 sg13g2_a21oi_1 _18778_ (.A1(net745),
    .A2(net61),
    .Y(_00361_),
    .B1(_11919_));
 sg13g2_nor2b_1 _18779_ (.A(_11917_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_11920_));
 sg13g2_a21oi_1 _18780_ (.A1(net970),
    .A2(_11917_),
    .Y(_11921_),
    .B1(_11920_));
 sg13g2_nand2_1 _18781_ (.Y(_11922_),
    .A(net847),
    .B(net61));
 sg13g2_o21ai_1 _18782_ (.B1(_11922_),
    .Y(_00362_),
    .A1(net61),
    .A2(_11921_));
 sg13g2_buf_1 _18783_ (.A(net1064),
    .X(_11923_));
 sg13g2_nor2b_1 _18784_ (.A(_11917_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_11924_));
 sg13g2_a21oi_1 _18785_ (.A1(net966),
    .A2(_11917_),
    .Y(_11925_),
    .B1(_11924_));
 sg13g2_nand2_1 _18786_ (.Y(_11926_),
    .A(net846),
    .B(net61));
 sg13g2_o21ai_1 _18787_ (.B1(_11926_),
    .Y(_00363_),
    .A1(net61),
    .A2(_11925_));
 sg13g2_mux2_1 _18788_ (.A0(\cpu.dcache.r_data[1][19] ),
    .A1(net973),
    .S(_11917_),
    .X(_11927_));
 sg13g2_nor2_1 _18789_ (.A(_11914_),
    .B(_11927_),
    .Y(_11928_));
 sg13g2_a21oi_1 _18790_ (.A1(net724),
    .A2(net61),
    .Y(_00364_),
    .B1(_11928_));
 sg13g2_nor2b_1 _18791_ (.A(_11881_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_11929_));
 sg13g2_a21oi_1 _18792_ (.A1(net970),
    .A2(_11881_),
    .Y(_11930_),
    .B1(_11929_));
 sg13g2_nand2_1 _18793_ (.Y(_11931_),
    .A(net847),
    .B(net63));
 sg13g2_o21ai_1 _18794_ (.B1(_11931_),
    .Y(_00365_),
    .A1(net63),
    .A2(_11930_));
 sg13g2_buf_1 _18795_ (.A(net1059),
    .X(_11932_));
 sg13g2_nor2_1 _18796_ (.A(net568),
    .B(_11796_),
    .Y(_11933_));
 sg13g2_buf_2 _18797_ (.A(_11933_),
    .X(_11934_));
 sg13g2_nor2b_1 _18798_ (.A(_11934_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_11935_));
 sg13g2_a21oi_1 _18799_ (.A1(net965),
    .A2(_11934_),
    .Y(_11936_),
    .B1(_11935_));
 sg13g2_nand2_1 _18800_ (.Y(_11937_),
    .A(net971),
    .B(_11914_));
 sg13g2_o21ai_1 _18801_ (.B1(_11937_),
    .Y(_00366_),
    .A1(_11915_),
    .A2(_11936_));
 sg13g2_nor2b_1 _18802_ (.A(_11934_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_11938_));
 sg13g2_a21oi_1 _18803_ (.A1(net970),
    .A2(_11934_),
    .Y(_11939_),
    .B1(_11938_));
 sg13g2_nand2_1 _18804_ (.Y(_11940_),
    .A(net969),
    .B(_11914_));
 sg13g2_o21ai_1 _18805_ (.B1(_11940_),
    .Y(_00367_),
    .A1(_11915_),
    .A2(_11939_));
 sg13g2_mux2_1 _18806_ (.A0(\cpu.dcache.r_data[1][22] ),
    .A1(net1058),
    .S(_11934_),
    .X(_11941_));
 sg13g2_nor2_1 _18807_ (.A(_11914_),
    .B(_11941_),
    .Y(_11942_));
 sg13g2_a21oi_1 _18808_ (.A1(net723),
    .A2(net61),
    .Y(_00368_),
    .B1(_11942_));
 sg13g2_mux2_1 _18809_ (.A0(\cpu.dcache.r_data[1][23] ),
    .A1(net973),
    .S(_11934_),
    .X(_11943_));
 sg13g2_nor2_1 _18810_ (.A(_11914_),
    .B(_11943_),
    .Y(_11944_));
 sg13g2_a21oi_1 _18811_ (.A1(net722),
    .A2(net61),
    .Y(_00369_),
    .B1(_11944_));
 sg13g2_nor4_1 _18812_ (.A(_11662_),
    .B(_11667_),
    .C(_11823_),
    .D(_11824_),
    .Y(_11945_));
 sg13g2_buf_2 _18813_ (.A(_11945_),
    .X(_11946_));
 sg13g2_nand2_1 _18814_ (.Y(_11947_),
    .A(net354),
    .B(_11946_));
 sg13g2_buf_2 _18815_ (.A(_11947_),
    .X(_11948_));
 sg13g2_buf_1 _18816_ (.A(_11948_),
    .X(_11949_));
 sg13g2_nand3_1 _18817_ (.B(_11653_),
    .C(_11657_),
    .A(_11652_),
    .Y(_11950_));
 sg13g2_buf_1 _18818_ (.A(_11950_),
    .X(_11951_));
 sg13g2_nor2_1 _18819_ (.A(net668),
    .B(_11951_),
    .Y(_11952_));
 sg13g2_buf_1 _18820_ (.A(_11952_),
    .X(_11953_));
 sg13g2_nor2b_1 _18821_ (.A(_11953_),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_11954_));
 sg13g2_a21oi_1 _18822_ (.A1(net968),
    .A2(_11953_),
    .Y(_11955_),
    .B1(_11954_));
 sg13g2_nor2_1 _18823_ (.A(net355),
    .B(_11948_),
    .Y(_11956_));
 sg13g2_a21oi_1 _18824_ (.A1(net60),
    .A2(_11955_),
    .Y(_00370_),
    .B1(_11956_));
 sg13g2_nor2b_1 _18825_ (.A(net519),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_11957_));
 sg13g2_a21oi_1 _18826_ (.A1(net967),
    .A2(net519),
    .Y(_11958_),
    .B1(_11957_));
 sg13g2_nor2_1 _18827_ (.A(net396),
    .B(_11948_),
    .Y(_11959_));
 sg13g2_a21oi_1 _18828_ (.A1(net60),
    .A2(_11958_),
    .Y(_00371_),
    .B1(_11959_));
 sg13g2_nor2b_1 _18829_ (.A(net519),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_11960_));
 sg13g2_a21oi_1 _18830_ (.A1(net982),
    .A2(net519),
    .Y(_11961_),
    .B1(_11960_));
 sg13g2_nor2_1 _18831_ (.A(_11708_),
    .B(_11948_),
    .Y(_11962_));
 sg13g2_a21oi_1 _18832_ (.A1(_11949_),
    .A2(_11961_),
    .Y(_00372_),
    .B1(_11962_));
 sg13g2_nor2b_1 _18833_ (.A(net519),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_11963_));
 sg13g2_a21oi_1 _18834_ (.A1(net981),
    .A2(net519),
    .Y(_11964_),
    .B1(_11963_));
 sg13g2_nor2_1 _18835_ (.A(_11722_),
    .B(_11948_),
    .Y(_11965_));
 sg13g2_a21oi_1 _18836_ (.A1(_11949_),
    .A2(_11964_),
    .Y(_00373_),
    .B1(_11965_));
 sg13g2_nor2_2 _18837_ (.A(_11874_),
    .B(_11836_),
    .Y(_11966_));
 sg13g2_mux2_1 _18838_ (.A0(\cpu.dcache.r_data[1][28] ),
    .A1(net1062),
    .S(_11966_),
    .X(_11967_));
 sg13g2_nand2_1 _18839_ (.Y(_11968_),
    .A(net60),
    .B(_11967_));
 sg13g2_o21ai_1 _18840_ (.B1(_11968_),
    .Y(_00374_),
    .A1(net358),
    .A2(net60));
 sg13g2_mux2_1 _18841_ (.A0(\cpu.dcache.r_data[1][29] ),
    .A1(net1055),
    .S(_11966_),
    .X(_11969_));
 sg13g2_nand2_1 _18842_ (.Y(_11970_),
    .A(net60),
    .B(_11969_));
 sg13g2_o21ai_1 _18843_ (.B1(_11970_),
    .Y(_00375_),
    .A1(net357),
    .A2(net60));
 sg13g2_nor2b_1 _18844_ (.A(_11881_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_11971_));
 sg13g2_a21oi_1 _18845_ (.A1(net966),
    .A2(_11881_),
    .Y(_11972_),
    .B1(_11971_));
 sg13g2_nand2_1 _18846_ (.Y(_11973_),
    .A(net846),
    .B(net63));
 sg13g2_o21ai_1 _18847_ (.B1(_11973_),
    .Y(_00376_),
    .A1(net63),
    .A2(_11972_));
 sg13g2_mux2_1 _18848_ (.A0(\cpu.dcache.r_data[1][30] ),
    .A1(net1056),
    .S(_11966_),
    .X(_11974_));
 sg13g2_nand2_1 _18849_ (.Y(_11975_),
    .A(_11948_),
    .B(_11974_));
 sg13g2_o21ai_1 _18850_ (.B1(_11975_),
    .Y(_00377_),
    .A1(net397),
    .A2(net60));
 sg13g2_mux2_1 _18851_ (.A0(\cpu.dcache.r_data[1][31] ),
    .A1(net1054),
    .S(_11966_),
    .X(_11976_));
 sg13g2_nand2_1 _18852_ (.Y(_11977_),
    .A(_11948_),
    .B(_11976_));
 sg13g2_o21ai_1 _18853_ (.B1(_11977_),
    .Y(_00378_),
    .A1(net356),
    .A2(net60));
 sg13g2_mux2_1 _18854_ (.A0(\cpu.dcache.r_data[1][3] ),
    .A1(net973),
    .S(_11881_),
    .X(_11978_));
 sg13g2_nor2_1 _18855_ (.A(_11878_),
    .B(_11978_),
    .Y(_11979_));
 sg13g2_a21oi_1 _18856_ (.A1(net724),
    .A2(net63),
    .Y(_00379_),
    .B1(_11979_));
 sg13g2_nor2_1 _18857_ (.A(net668),
    .B(_11853_),
    .Y(_11980_));
 sg13g2_buf_2 _18858_ (.A(_11980_),
    .X(_11981_));
 sg13g2_nor2b_1 _18859_ (.A(_11981_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_11982_));
 sg13g2_a21oi_1 _18860_ (.A1(net965),
    .A2(_11981_),
    .Y(_11983_),
    .B1(_11982_));
 sg13g2_buf_1 _18861_ (.A(_09839_),
    .X(_11984_));
 sg13g2_nand2_1 _18862_ (.Y(_11985_),
    .A(net964),
    .B(_11878_));
 sg13g2_o21ai_1 _18863_ (.B1(_11985_),
    .Y(_00380_),
    .A1(_11879_),
    .A2(_11983_));
 sg13g2_nor2b_1 _18864_ (.A(_11981_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_11986_));
 sg13g2_a21oi_1 _18865_ (.A1(net970),
    .A2(_11981_),
    .Y(_11987_),
    .B1(_11986_));
 sg13g2_buf_1 _18866_ (.A(_09845_),
    .X(_11988_));
 sg13g2_nand2_1 _18867_ (.Y(_11989_),
    .A(net963),
    .B(_11878_));
 sg13g2_o21ai_1 _18868_ (.B1(_11989_),
    .Y(_00381_),
    .A1(net63),
    .A2(_11987_));
 sg13g2_mux2_1 _18869_ (.A0(\cpu.dcache.r_data[1][6] ),
    .A1(net978),
    .S(_11981_),
    .X(_11990_));
 sg13g2_nor2_1 _18870_ (.A(_11878_),
    .B(_11990_),
    .Y(_11991_));
 sg13g2_a21oi_1 _18871_ (.A1(net723),
    .A2(net63),
    .Y(_00382_),
    .B1(_11991_));
 sg13g2_mux2_1 _18872_ (.A0(\cpu.dcache.r_data[1][7] ),
    .A1(net973),
    .S(_11981_),
    .X(_11992_));
 sg13g2_nor2_1 _18873_ (.A(_11878_),
    .B(_11992_),
    .Y(_11993_));
 sg13g2_a21oi_1 _18874_ (.A1(net722),
    .A2(_11879_),
    .Y(_00383_),
    .B1(_11993_));
 sg13g2_nor2b_1 _18875_ (.A(_11893_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_11994_));
 sg13g2_a21oi_1 _18876_ (.A1(net968),
    .A2(_11893_),
    .Y(_11995_),
    .B1(_11994_));
 sg13g2_nor2_1 _18877_ (.A(net355),
    .B(_11890_),
    .Y(_11996_));
 sg13g2_a21oi_1 _18878_ (.A1(net62),
    .A2(_11995_),
    .Y(_00384_),
    .B1(_11996_));
 sg13g2_nor2b_1 _18879_ (.A(_11893_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_11997_));
 sg13g2_a21oi_1 _18880_ (.A1(net967),
    .A2(_11893_),
    .Y(_11998_),
    .B1(_11997_));
 sg13g2_nor2_1 _18881_ (.A(net396),
    .B(_11890_),
    .Y(_11999_));
 sg13g2_a21oi_1 _18882_ (.A1(_11891_),
    .A2(_11998_),
    .Y(_00385_),
    .B1(_11999_));
 sg13g2_buf_1 _18883_ (.A(_09440_),
    .X(_12000_));
 sg13g2_nor2_1 _18884_ (.A(net641),
    .B(_11876_),
    .Y(_12001_));
 sg13g2_buf_2 _18885_ (.A(_12001_),
    .X(_12002_));
 sg13g2_buf_1 _18886_ (.A(_12002_),
    .X(_12003_));
 sg13g2_nor2_1 _18887_ (.A(net641),
    .B(_11682_),
    .Y(_12004_));
 sg13g2_buf_2 _18888_ (.A(_12004_),
    .X(_12005_));
 sg13g2_mux2_1 _18889_ (.A0(\cpu.dcache.r_data[2][0] ),
    .A1(net1065),
    .S(_12005_),
    .X(_12006_));
 sg13g2_nor2_1 _18890_ (.A(_12002_),
    .B(_12006_),
    .Y(_12007_));
 sg13g2_a21oi_1 _18891_ (.A1(_09811_),
    .A2(net59),
    .Y(_00386_),
    .B1(_12007_));
 sg13g2_buf_1 _18892_ (.A(net592),
    .X(_12008_));
 sg13g2_buf_1 _18893_ (.A(net518),
    .X(_12009_));
 sg13g2_buf_1 _18894_ (.A(net457),
    .X(_12010_));
 sg13g2_nand2_1 _18895_ (.Y(_12011_),
    .A(net394),
    .B(_11888_));
 sg13g2_buf_2 _18896_ (.A(_12011_),
    .X(_12012_));
 sg13g2_buf_1 _18897_ (.A(_12012_),
    .X(_12013_));
 sg13g2_nor2_1 _18898_ (.A(net641),
    .B(_11697_),
    .Y(_12014_));
 sg13g2_buf_2 _18899_ (.A(_12014_),
    .X(_12015_));
 sg13g2_nor2b_1 _18900_ (.A(_12015_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12016_));
 sg13g2_a21oi_1 _18901_ (.A1(net982),
    .A2(_12015_),
    .Y(_12017_),
    .B1(_12016_));
 sg13g2_nor2_1 _18902_ (.A(net360),
    .B(_12012_),
    .Y(_12018_));
 sg13g2_a21oi_1 _18903_ (.A1(net58),
    .A2(_12017_),
    .Y(_00387_),
    .B1(_12018_));
 sg13g2_nor2b_1 _18904_ (.A(_12015_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12019_));
 sg13g2_a21oi_1 _18905_ (.A1(net981),
    .A2(_12015_),
    .Y(_12020_),
    .B1(_12019_));
 sg13g2_nor2_1 _18906_ (.A(net359),
    .B(_12012_),
    .Y(_12021_));
 sg13g2_a21oi_1 _18907_ (.A1(_12013_),
    .A2(_12020_),
    .Y(_00388_),
    .B1(_12021_));
 sg13g2_nor2_2 _18908_ (.A(_12000_),
    .B(_11733_),
    .Y(_12022_));
 sg13g2_mux2_1 _18909_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(net1062),
    .S(_12022_),
    .X(_12023_));
 sg13g2_nand2_1 _18910_ (.Y(_12024_),
    .A(net58),
    .B(_12023_));
 sg13g2_o21ai_1 _18911_ (.B1(_12024_),
    .Y(_00389_),
    .A1(net358),
    .A2(net58));
 sg13g2_mux2_1 _18912_ (.A0(\cpu.dcache.r_data[2][13] ),
    .A1(net1055),
    .S(_12022_),
    .X(_12025_));
 sg13g2_nand2_1 _18913_ (.Y(_12026_),
    .A(net58),
    .B(_12025_));
 sg13g2_o21ai_1 _18914_ (.B1(_12026_),
    .Y(_00390_),
    .A1(net357),
    .A2(net58));
 sg13g2_mux2_1 _18915_ (.A0(\cpu.dcache.r_data[2][14] ),
    .A1(net1056),
    .S(_12022_),
    .X(_12027_));
 sg13g2_nand2_1 _18916_ (.Y(_12028_),
    .A(_12012_),
    .B(_12027_));
 sg13g2_o21ai_1 _18917_ (.B1(_12028_),
    .Y(_00391_),
    .A1(net397),
    .A2(net58));
 sg13g2_mux2_1 _18918_ (.A0(\cpu.dcache.r_data[2][15] ),
    .A1(net1054),
    .S(_12022_),
    .X(_12029_));
 sg13g2_nand2_1 _18919_ (.Y(_12030_),
    .A(_12012_),
    .B(_12029_));
 sg13g2_o21ai_1 _18920_ (.B1(_12030_),
    .Y(_00392_),
    .A1(net356),
    .A2(net58));
 sg13g2_nor2_1 _18921_ (.A(net641),
    .B(_11912_),
    .Y(_12031_));
 sg13g2_buf_1 _18922_ (.A(_12031_),
    .X(_12032_));
 sg13g2_buf_1 _18923_ (.A(_12032_),
    .X(_12033_));
 sg13g2_nor2_1 _18924_ (.A(net641),
    .B(_11769_),
    .Y(_12034_));
 sg13g2_buf_2 _18925_ (.A(_12034_),
    .X(_12035_));
 sg13g2_mux2_1 _18926_ (.A0(\cpu.dcache.r_data[2][16] ),
    .A1(net1065),
    .S(_12035_),
    .X(_12036_));
 sg13g2_nor2_1 _18927_ (.A(_12032_),
    .B(_12036_),
    .Y(_12037_));
 sg13g2_a21oi_1 _18928_ (.A1(net745),
    .A2(_12033_),
    .Y(_00393_),
    .B1(_12037_));
 sg13g2_nor2b_1 _18929_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12038_));
 sg13g2_a21oi_1 _18930_ (.A1(net970),
    .A2(_12035_),
    .Y(_12039_),
    .B1(_12038_));
 sg13g2_nand2_1 _18931_ (.Y(_12040_),
    .A(net847),
    .B(net57));
 sg13g2_o21ai_1 _18932_ (.B1(_12040_),
    .Y(_00394_),
    .A1(net57),
    .A2(_12039_));
 sg13g2_nor2b_1 _18933_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12041_));
 sg13g2_a21oi_1 _18934_ (.A1(net966),
    .A2(_12035_),
    .Y(_12042_),
    .B1(_12041_));
 sg13g2_nand2_1 _18935_ (.Y(_12043_),
    .A(net846),
    .B(net57));
 sg13g2_o21ai_1 _18936_ (.B1(_12043_),
    .Y(_00395_),
    .A1(net57),
    .A2(_12042_));
 sg13g2_mux2_1 _18937_ (.A0(\cpu.dcache.r_data[2][19] ),
    .A1(net973),
    .S(_12035_),
    .X(_12044_));
 sg13g2_nor2_1 _18938_ (.A(_12032_),
    .B(_12044_),
    .Y(_12045_));
 sg13g2_a21oi_1 _18939_ (.A1(net724),
    .A2(_12033_),
    .Y(_00396_),
    .B1(_12045_));
 sg13g2_nor2b_1 _18940_ (.A(_12005_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12046_));
 sg13g2_a21oi_1 _18941_ (.A1(_11803_),
    .A2(_12005_),
    .Y(_12047_),
    .B1(_12046_));
 sg13g2_nand2_1 _18942_ (.Y(_12048_),
    .A(_11778_),
    .B(net59));
 sg13g2_o21ai_1 _18943_ (.B1(_12048_),
    .Y(_00397_),
    .A1(net59),
    .A2(_12047_));
 sg13g2_nor2_1 _18944_ (.A(_09440_),
    .B(_11796_),
    .Y(_12049_));
 sg13g2_buf_2 _18945_ (.A(_12049_),
    .X(_12050_));
 sg13g2_nor2b_1 _18946_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12051_));
 sg13g2_a21oi_1 _18947_ (.A1(net965),
    .A2(_12050_),
    .Y(_12052_),
    .B1(_12051_));
 sg13g2_nand2_1 _18948_ (.Y(_12053_),
    .A(net964),
    .B(_12032_));
 sg13g2_o21ai_1 _18949_ (.B1(_12053_),
    .Y(_00398_),
    .A1(net57),
    .A2(_12052_));
 sg13g2_nor2b_1 _18950_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12054_));
 sg13g2_a21oi_1 _18951_ (.A1(net970),
    .A2(_12050_),
    .Y(_12055_),
    .B1(_12054_));
 sg13g2_nand2_1 _18952_ (.Y(_12056_),
    .A(net963),
    .B(_12032_));
 sg13g2_o21ai_1 _18953_ (.B1(_12056_),
    .Y(_00399_),
    .A1(net57),
    .A2(_12055_));
 sg13g2_mux2_1 _18954_ (.A0(\cpu.dcache.r_data[2][22] ),
    .A1(net978),
    .S(_12050_),
    .X(_12057_));
 sg13g2_nor2_1 _18955_ (.A(_12032_),
    .B(_12057_),
    .Y(_12058_));
 sg13g2_a21oi_1 _18956_ (.A1(net723),
    .A2(net57),
    .Y(_00400_),
    .B1(_12058_));
 sg13g2_mux2_1 _18957_ (.A0(\cpu.dcache.r_data[2][23] ),
    .A1(net973),
    .S(_12050_),
    .X(_12059_));
 sg13g2_nor2_1 _18958_ (.A(_12032_),
    .B(_12059_),
    .Y(_12060_));
 sg13g2_a21oi_1 _18959_ (.A1(net722),
    .A2(net57),
    .Y(_00401_),
    .B1(_12060_));
 sg13g2_nand2_1 _18960_ (.Y(_12061_),
    .A(net394),
    .B(_11946_));
 sg13g2_buf_1 _18961_ (.A(_12061_),
    .X(_12062_));
 sg13g2_buf_1 _18962_ (.A(_12062_),
    .X(_12063_));
 sg13g2_nor2_1 _18963_ (.A(net641),
    .B(_11951_),
    .Y(_12064_));
 sg13g2_buf_1 _18964_ (.A(_12064_),
    .X(_12065_));
 sg13g2_nor2b_1 _18965_ (.A(net517),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12066_));
 sg13g2_a21oi_1 _18966_ (.A1(net968),
    .A2(net517),
    .Y(_12067_),
    .B1(_12066_));
 sg13g2_nor2_1 _18967_ (.A(_11819_),
    .B(_12062_),
    .Y(_12068_));
 sg13g2_a21oi_1 _18968_ (.A1(net56),
    .A2(_12067_),
    .Y(_00402_),
    .B1(_12068_));
 sg13g2_nor2b_1 _18969_ (.A(net517),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12069_));
 sg13g2_a21oi_1 _18970_ (.A1(net967),
    .A2(net517),
    .Y(_12070_),
    .B1(_12069_));
 sg13g2_nor2_1 _18971_ (.A(_11830_),
    .B(_12062_),
    .Y(_12071_));
 sg13g2_a21oi_1 _18972_ (.A1(net56),
    .A2(_12070_),
    .Y(_00403_),
    .B1(_12071_));
 sg13g2_nor2b_1 _18973_ (.A(net517),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12072_));
 sg13g2_a21oi_1 _18974_ (.A1(net982),
    .A2(net517),
    .Y(_12073_),
    .B1(_12072_));
 sg13g2_nor2_1 _18975_ (.A(net360),
    .B(_12062_),
    .Y(_12074_));
 sg13g2_a21oi_1 _18976_ (.A1(_12063_),
    .A2(_12073_),
    .Y(_00404_),
    .B1(_12074_));
 sg13g2_nor2b_1 _18977_ (.A(net517),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12075_));
 sg13g2_a21oi_1 _18978_ (.A1(net981),
    .A2(net517),
    .Y(_12076_),
    .B1(_12075_));
 sg13g2_nor2_1 _18979_ (.A(net359),
    .B(_12062_),
    .Y(_12077_));
 sg13g2_a21oi_1 _18980_ (.A1(_12063_),
    .A2(_12076_),
    .Y(_00405_),
    .B1(_12077_));
 sg13g2_nor2_2 _18981_ (.A(_12000_),
    .B(_11836_),
    .Y(_12078_));
 sg13g2_mux2_1 _18982_ (.A0(\cpu.dcache.r_data[2][28] ),
    .A1(net1062),
    .S(_12078_),
    .X(_12079_));
 sg13g2_nand2_1 _18983_ (.Y(_12080_),
    .A(net56),
    .B(_12079_));
 sg13g2_o21ai_1 _18984_ (.B1(_12080_),
    .Y(_00406_),
    .A1(net358),
    .A2(net56));
 sg13g2_mux2_1 _18985_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(net1055),
    .S(_12078_),
    .X(_12081_));
 sg13g2_nand2_1 _18986_ (.Y(_12082_),
    .A(net56),
    .B(_12081_));
 sg13g2_o21ai_1 _18987_ (.B1(_12082_),
    .Y(_00407_),
    .A1(net357),
    .A2(net56));
 sg13g2_nor2b_1 _18988_ (.A(_12005_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12083_));
 sg13g2_a21oi_1 _18989_ (.A1(net966),
    .A2(_12005_),
    .Y(_12084_),
    .B1(_12083_));
 sg13g2_nand2_1 _18990_ (.Y(_12085_),
    .A(_11783_),
    .B(net59));
 sg13g2_o21ai_1 _18991_ (.B1(_12085_),
    .Y(_00408_),
    .A1(net59),
    .A2(_12084_));
 sg13g2_mux2_1 _18992_ (.A0(\cpu.dcache.r_data[2][30] ),
    .A1(net1056),
    .S(_12078_),
    .X(_12086_));
 sg13g2_nand2_1 _18993_ (.Y(_12087_),
    .A(_12062_),
    .B(_12086_));
 sg13g2_o21ai_1 _18994_ (.B1(_12087_),
    .Y(_00409_),
    .A1(net397),
    .A2(net56));
 sg13g2_mux2_1 _18995_ (.A0(\cpu.dcache.r_data[2][31] ),
    .A1(_11908_),
    .S(_12078_),
    .X(_12088_));
 sg13g2_nand2_1 _18996_ (.Y(_12089_),
    .A(_12062_),
    .B(_12088_));
 sg13g2_o21ai_1 _18997_ (.B1(_12089_),
    .Y(_00410_),
    .A1(net356),
    .A2(net56));
 sg13g2_buf_1 _18998_ (.A(net1063),
    .X(_12090_));
 sg13g2_mux2_1 _18999_ (.A0(\cpu.dcache.r_data[2][3] ),
    .A1(_12090_),
    .S(_12005_),
    .X(_12091_));
 sg13g2_nor2_1 _19000_ (.A(_12002_),
    .B(_12091_),
    .Y(_12092_));
 sg13g2_a21oi_1 _19001_ (.A1(net724),
    .A2(net59),
    .Y(_00411_),
    .B1(_12092_));
 sg13g2_nor2_1 _19002_ (.A(_09440_),
    .B(_11853_),
    .Y(_12093_));
 sg13g2_buf_2 _19003_ (.A(_12093_),
    .X(_12094_));
 sg13g2_nor2b_1 _19004_ (.A(_12094_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12095_));
 sg13g2_a21oi_1 _19005_ (.A1(net965),
    .A2(_12094_),
    .Y(_12096_),
    .B1(_12095_));
 sg13g2_nand2_1 _19006_ (.Y(_12097_),
    .A(_11984_),
    .B(_12002_));
 sg13g2_o21ai_1 _19007_ (.B1(_12097_),
    .Y(_00412_),
    .A1(_12003_),
    .A2(_12096_));
 sg13g2_nor2b_1 _19008_ (.A(_12094_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12098_));
 sg13g2_a21oi_1 _19009_ (.A1(_11803_),
    .A2(_12094_),
    .Y(_12099_),
    .B1(_12098_));
 sg13g2_nand2_1 _19010_ (.Y(_12100_),
    .A(net963),
    .B(_12002_));
 sg13g2_o21ai_1 _19011_ (.B1(_12100_),
    .Y(_00413_),
    .A1(net59),
    .A2(_12099_));
 sg13g2_mux2_1 _19012_ (.A0(\cpu.dcache.r_data[2][6] ),
    .A1(net978),
    .S(_12094_),
    .X(_12101_));
 sg13g2_nor2_1 _19013_ (.A(_12002_),
    .B(_12101_),
    .Y(_12102_));
 sg13g2_a21oi_1 _19014_ (.A1(net723),
    .A2(net59),
    .Y(_00414_),
    .B1(_12102_));
 sg13g2_mux2_1 _19015_ (.A0(\cpu.dcache.r_data[2][7] ),
    .A1(net962),
    .S(_12094_),
    .X(_12103_));
 sg13g2_nor2_1 _19016_ (.A(_12002_),
    .B(_12103_),
    .Y(_12104_));
 sg13g2_a21oi_1 _19017_ (.A1(_11813_),
    .A2(_12003_),
    .Y(_00415_),
    .B1(_12104_));
 sg13g2_nor2b_1 _19018_ (.A(_12015_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12105_));
 sg13g2_a21oi_1 _19019_ (.A1(net968),
    .A2(_12015_),
    .Y(_12106_),
    .B1(_12105_));
 sg13g2_nor2_1 _19020_ (.A(net355),
    .B(_12012_),
    .Y(_12107_));
 sg13g2_a21oi_1 _19021_ (.A1(_12013_),
    .A2(_12106_),
    .Y(_00416_),
    .B1(_12107_));
 sg13g2_nor2b_1 _19022_ (.A(_12015_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12108_));
 sg13g2_a21oi_1 _19023_ (.A1(net967),
    .A2(_12015_),
    .Y(_12109_),
    .B1(_12108_));
 sg13g2_nor2_1 _19024_ (.A(net396),
    .B(_12012_),
    .Y(_12110_));
 sg13g2_a21oi_1 _19025_ (.A1(net58),
    .A2(_12109_),
    .Y(_00417_),
    .B1(_12110_));
 sg13g2_nand2_1 _19026_ (.Y(_12111_),
    .A(net1013),
    .B(_09157_));
 sg13g2_buf_1 _19027_ (.A(_12111_),
    .X(_12112_));
 sg13g2_nor2_1 _19028_ (.A(net640),
    .B(_11876_),
    .Y(_12113_));
 sg13g2_buf_1 _19029_ (.A(_12113_),
    .X(_12114_));
 sg13g2_buf_1 _19030_ (.A(_12114_),
    .X(_12115_));
 sg13g2_buf_1 _19031_ (.A(_11673_),
    .X(_12116_));
 sg13g2_nor2_1 _19032_ (.A(net640),
    .B(_11682_),
    .Y(_12117_));
 sg13g2_buf_2 _19033_ (.A(_12117_),
    .X(_12118_));
 sg13g2_mux2_1 _19034_ (.A0(\cpu.dcache.r_data[3][0] ),
    .A1(net1053),
    .S(_12118_),
    .X(_12119_));
 sg13g2_nor2_1 _19035_ (.A(_12114_),
    .B(_12119_),
    .Y(_12120_));
 sg13g2_a21oi_1 _19036_ (.A1(net745),
    .A2(net55),
    .Y(_00418_),
    .B1(_12120_));
 sg13g2_buf_1 _19037_ (.A(_09161_),
    .X(_12121_));
 sg13g2_buf_1 _19038_ (.A(net456),
    .X(_12122_));
 sg13g2_nand2_1 _19039_ (.Y(_12123_),
    .A(net393),
    .B(_11888_));
 sg13g2_buf_1 _19040_ (.A(_12123_),
    .X(_12124_));
 sg13g2_buf_1 _19041_ (.A(_12124_),
    .X(_12125_));
 sg13g2_nor2_1 _19042_ (.A(net640),
    .B(_11697_),
    .Y(_12126_));
 sg13g2_buf_2 _19043_ (.A(_12126_),
    .X(_12127_));
 sg13g2_nor2b_1 _19044_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12128_));
 sg13g2_a21oi_1 _19045_ (.A1(net982),
    .A2(_12127_),
    .Y(_12129_),
    .B1(_12128_));
 sg13g2_nor2_1 _19046_ (.A(net360),
    .B(_12124_),
    .Y(_12130_));
 sg13g2_a21oi_1 _19047_ (.A1(_12125_),
    .A2(_12129_),
    .Y(_00419_),
    .B1(_12130_));
 sg13g2_nor2b_1 _19048_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12131_));
 sg13g2_a21oi_1 _19049_ (.A1(net981),
    .A2(_12127_),
    .Y(_12132_),
    .B1(_12131_));
 sg13g2_nor2_1 _19050_ (.A(net359),
    .B(_12124_),
    .Y(_12133_));
 sg13g2_a21oi_1 _19051_ (.A1(_12125_),
    .A2(_12132_),
    .Y(_00420_),
    .B1(_12133_));
 sg13g2_nor2_2 _19052_ (.A(_12112_),
    .B(_11733_),
    .Y(_12134_));
 sg13g2_mux2_1 _19053_ (.A0(\cpu.dcache.r_data[3][12] ),
    .A1(net1062),
    .S(_12134_),
    .X(_12135_));
 sg13g2_nand2_1 _19054_ (.Y(_12136_),
    .A(net54),
    .B(_12135_));
 sg13g2_o21ai_1 _19055_ (.B1(_12136_),
    .Y(_00421_),
    .A1(net358),
    .A2(net54));
 sg13g2_mux2_1 _19056_ (.A0(\cpu.dcache.r_data[3][13] ),
    .A1(net1055),
    .S(_12134_),
    .X(_12137_));
 sg13g2_nand2_1 _19057_ (.Y(_12138_),
    .A(net54),
    .B(_12137_));
 sg13g2_o21ai_1 _19058_ (.B1(_12138_),
    .Y(_00422_),
    .A1(net357),
    .A2(net54));
 sg13g2_mux2_1 _19059_ (.A0(\cpu.dcache.r_data[3][14] ),
    .A1(net1056),
    .S(_12134_),
    .X(_12139_));
 sg13g2_nand2_1 _19060_ (.Y(_12140_),
    .A(_12124_),
    .B(_12139_));
 sg13g2_o21ai_1 _19061_ (.B1(_12140_),
    .Y(_00423_),
    .A1(net397),
    .A2(net54));
 sg13g2_mux2_1 _19062_ (.A0(\cpu.dcache.r_data[3][15] ),
    .A1(net1054),
    .S(_12134_),
    .X(_12141_));
 sg13g2_nand2_1 _19063_ (.Y(_12142_),
    .A(_12124_),
    .B(_12141_));
 sg13g2_o21ai_1 _19064_ (.B1(_12142_),
    .Y(_00424_),
    .A1(net356),
    .A2(net54));
 sg13g2_nor2_1 _19065_ (.A(net640),
    .B(_11912_),
    .Y(_12143_));
 sg13g2_buf_1 _19066_ (.A(_12143_),
    .X(_12144_));
 sg13g2_buf_1 _19067_ (.A(_12144_),
    .X(_12145_));
 sg13g2_nor2_1 _19068_ (.A(net640),
    .B(_11769_),
    .Y(_12146_));
 sg13g2_buf_2 _19069_ (.A(_12146_),
    .X(_12147_));
 sg13g2_mux2_1 _19070_ (.A0(\cpu.dcache.r_data[3][16] ),
    .A1(net1053),
    .S(_12147_),
    .X(_12148_));
 sg13g2_nor2_1 _19071_ (.A(_12144_),
    .B(_12148_),
    .Y(_12149_));
 sg13g2_a21oi_1 _19072_ (.A1(net745),
    .A2(net53),
    .Y(_00425_),
    .B1(_12149_));
 sg13g2_buf_1 _19073_ (.A(net1060),
    .X(_12150_));
 sg13g2_nor2b_1 _19074_ (.A(_12147_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12151_));
 sg13g2_a21oi_1 _19075_ (.A1(net961),
    .A2(_12147_),
    .Y(_12152_),
    .B1(_12151_));
 sg13g2_nand2_1 _19076_ (.Y(_12153_),
    .A(net847),
    .B(net53));
 sg13g2_o21ai_1 _19077_ (.B1(_12153_),
    .Y(_00426_),
    .A1(net53),
    .A2(_12152_));
 sg13g2_nor2b_1 _19078_ (.A(_12147_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12154_));
 sg13g2_a21oi_1 _19079_ (.A1(net966),
    .A2(_12147_),
    .Y(_12155_),
    .B1(_12154_));
 sg13g2_nand2_1 _19080_ (.Y(_12156_),
    .A(net846),
    .B(net53));
 sg13g2_o21ai_1 _19081_ (.B1(_12156_),
    .Y(_00427_),
    .A1(net53),
    .A2(_12155_));
 sg13g2_mux2_1 _19082_ (.A0(\cpu.dcache.r_data[3][19] ),
    .A1(net962),
    .S(_12147_),
    .X(_12157_));
 sg13g2_nor2_1 _19083_ (.A(_12144_),
    .B(_12157_),
    .Y(_12158_));
 sg13g2_a21oi_1 _19084_ (.A1(net724),
    .A2(net53),
    .Y(_00428_),
    .B1(_12158_));
 sg13g2_nor2b_1 _19085_ (.A(_12118_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12159_));
 sg13g2_a21oi_1 _19086_ (.A1(net961),
    .A2(_12118_),
    .Y(_12160_),
    .B1(_12159_));
 sg13g2_nand2_1 _19087_ (.Y(_12161_),
    .A(net847),
    .B(net55));
 sg13g2_o21ai_1 _19088_ (.B1(_12161_),
    .Y(_00429_),
    .A1(net55),
    .A2(_12160_));
 sg13g2_buf_2 _19089_ (.A(net1059),
    .X(_12162_));
 sg13g2_or2_1 _19090_ (.X(_12163_),
    .B(_11796_),
    .A(_12111_));
 sg13g2_buf_1 _19091_ (.A(_12163_),
    .X(_12164_));
 sg13g2_mux2_1 _19092_ (.A0(_12162_),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12164_),
    .X(_12165_));
 sg13g2_mux2_1 _19093_ (.A0(_12165_),
    .A1(net971),
    .S(net53),
    .X(_00430_));
 sg13g2_mux2_1 _19094_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12164_),
    .X(_12166_));
 sg13g2_mux2_1 _19095_ (.A0(_12166_),
    .A1(net969),
    .S(_12145_),
    .X(_00431_));
 sg13g2_mux2_1 _19096_ (.A0(net1058),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12164_),
    .X(_12167_));
 sg13g2_nor2_1 _19097_ (.A(_12144_),
    .B(_12167_),
    .Y(_12168_));
 sg13g2_a21oi_1 _19098_ (.A1(net723),
    .A2(net53),
    .Y(_00432_),
    .B1(_12168_));
 sg13g2_mux2_1 _19099_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12164_),
    .X(_12169_));
 sg13g2_nor2_1 _19100_ (.A(_12144_),
    .B(_12169_),
    .Y(_12170_));
 sg13g2_a21oi_1 _19101_ (.A1(net722),
    .A2(_12145_),
    .Y(_00433_),
    .B1(_12170_));
 sg13g2_nand2_1 _19102_ (.Y(_12171_),
    .A(net393),
    .B(_11946_));
 sg13g2_buf_2 _19103_ (.A(_12171_),
    .X(_12172_));
 sg13g2_buf_1 _19104_ (.A(_12172_),
    .X(_12173_));
 sg13g2_nor2_1 _19105_ (.A(net640),
    .B(_11951_),
    .Y(_12174_));
 sg13g2_buf_1 _19106_ (.A(_12174_),
    .X(_12175_));
 sg13g2_nor2b_1 _19107_ (.A(net516),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12176_));
 sg13g2_a21oi_1 _19108_ (.A1(net968),
    .A2(net516),
    .Y(_12177_),
    .B1(_12176_));
 sg13g2_nor2_1 _19109_ (.A(_11819_),
    .B(_12172_),
    .Y(_12178_));
 sg13g2_a21oi_1 _19110_ (.A1(net52),
    .A2(_12177_),
    .Y(_00434_),
    .B1(_12178_));
 sg13g2_nor2b_1 _19111_ (.A(net516),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12179_));
 sg13g2_a21oi_1 _19112_ (.A1(net967),
    .A2(net516),
    .Y(_12180_),
    .B1(_12179_));
 sg13g2_nor2_1 _19113_ (.A(net396),
    .B(_12172_),
    .Y(_12181_));
 sg13g2_a21oi_1 _19114_ (.A1(net52),
    .A2(_12180_),
    .Y(_00435_),
    .B1(_12181_));
 sg13g2_nor2b_1 _19115_ (.A(net516),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12182_));
 sg13g2_a21oi_1 _19116_ (.A1(net974),
    .A2(net516),
    .Y(_12183_),
    .B1(_12182_));
 sg13g2_nor2_1 _19117_ (.A(_11708_),
    .B(_12172_),
    .Y(_12184_));
 sg13g2_a21oi_1 _19118_ (.A1(_12173_),
    .A2(_12183_),
    .Y(_00436_),
    .B1(_12184_));
 sg13g2_buf_1 _19119_ (.A(net1063),
    .X(_12185_));
 sg13g2_nor2b_1 _19120_ (.A(_12175_),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12186_));
 sg13g2_a21oi_1 _19121_ (.A1(net960),
    .A2(_12175_),
    .Y(_12187_),
    .B1(_12186_));
 sg13g2_nor2_1 _19122_ (.A(net359),
    .B(_12172_),
    .Y(_12188_));
 sg13g2_a21oi_1 _19123_ (.A1(_12173_),
    .A2(_12187_),
    .Y(_00437_),
    .B1(_12188_));
 sg13g2_nor2_2 _19124_ (.A(_12112_),
    .B(_11836_),
    .Y(_12189_));
 sg13g2_mux2_1 _19125_ (.A0(\cpu.dcache.r_data[3][28] ),
    .A1(net1062),
    .S(_12189_),
    .X(_12190_));
 sg13g2_nand2_1 _19126_ (.Y(_12191_),
    .A(net52),
    .B(_12190_));
 sg13g2_o21ai_1 _19127_ (.B1(_12191_),
    .Y(_00438_),
    .A1(net358),
    .A2(net52));
 sg13g2_mux2_1 _19128_ (.A0(\cpu.dcache.r_data[3][29] ),
    .A1(_11903_),
    .S(_12189_),
    .X(_12192_));
 sg13g2_nand2_1 _19129_ (.Y(_12193_),
    .A(net52),
    .B(_12192_));
 sg13g2_o21ai_1 _19130_ (.B1(_12193_),
    .Y(_00439_),
    .A1(net357),
    .A2(net52));
 sg13g2_nor2b_1 _19131_ (.A(_12118_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12194_));
 sg13g2_a21oi_1 _19132_ (.A1(_11923_),
    .A2(_12118_),
    .Y(_12195_),
    .B1(_12194_));
 sg13g2_nand2_1 _19133_ (.Y(_12196_),
    .A(_11783_),
    .B(net55));
 sg13g2_o21ai_1 _19134_ (.B1(_12196_),
    .Y(_00440_),
    .A1(net55),
    .A2(_12195_));
 sg13g2_mux2_1 _19135_ (.A0(\cpu.dcache.r_data[3][30] ),
    .A1(_11845_),
    .S(_12189_),
    .X(_12197_));
 sg13g2_nand2_1 _19136_ (.Y(_12198_),
    .A(_12172_),
    .B(_12197_));
 sg13g2_o21ai_1 _19137_ (.B1(_12198_),
    .Y(_00441_),
    .A1(_11750_),
    .A2(net52));
 sg13g2_mux2_1 _19138_ (.A0(\cpu.dcache.r_data[3][31] ),
    .A1(_11908_),
    .S(_12189_),
    .X(_12199_));
 sg13g2_nand2_1 _19139_ (.Y(_12200_),
    .A(_12172_),
    .B(_12199_));
 sg13g2_o21ai_1 _19140_ (.B1(_12200_),
    .Y(_00442_),
    .A1(net356),
    .A2(net52));
 sg13g2_mux2_1 _19141_ (.A0(\cpu.dcache.r_data[3][3] ),
    .A1(_12090_),
    .S(_12118_),
    .X(_12201_));
 sg13g2_nor2_1 _19142_ (.A(_12114_),
    .B(_12201_),
    .Y(_12202_));
 sg13g2_a21oi_1 _19143_ (.A1(_11785_),
    .A2(net55),
    .Y(_00443_),
    .B1(_12202_));
 sg13g2_or2_1 _19144_ (.X(_12203_),
    .B(_11853_),
    .A(_12111_));
 sg13g2_buf_1 _19145_ (.A(_12203_),
    .X(_12204_));
 sg13g2_mux2_1 _19146_ (.A0(_12162_),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12204_),
    .X(_12205_));
 sg13g2_mux2_1 _19147_ (.A0(_12205_),
    .A1(net971),
    .S(net55),
    .X(_00444_));
 sg13g2_mux2_1 _19148_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12204_),
    .X(_12206_));
 sg13g2_mux2_1 _19149_ (.A0(_12206_),
    .A1(net969),
    .S(_12115_),
    .X(_00445_));
 sg13g2_mux2_1 _19150_ (.A0(net1058),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12204_),
    .X(_12207_));
 sg13g2_nor2_1 _19151_ (.A(_12114_),
    .B(_12207_),
    .Y(_12208_));
 sg13g2_a21oi_1 _19152_ (.A1(_11809_),
    .A2(_12115_),
    .Y(_00446_),
    .B1(_12208_));
 sg13g2_mux2_1 _19153_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12204_),
    .X(_12209_));
 sg13g2_nor2_1 _19154_ (.A(_12114_),
    .B(_12209_),
    .Y(_12210_));
 sg13g2_a21oi_1 _19155_ (.A1(net722),
    .A2(net55),
    .Y(_00447_),
    .B1(_12210_));
 sg13g2_nor2b_1 _19156_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12211_));
 sg13g2_a21oi_1 _19157_ (.A1(net972),
    .A2(_12127_),
    .Y(_12212_),
    .B1(_12211_));
 sg13g2_nor2_1 _19158_ (.A(net355),
    .B(_12124_),
    .Y(_12213_));
 sg13g2_a21oi_1 _19159_ (.A1(net54),
    .A2(_12212_),
    .Y(_00448_),
    .B1(_12213_));
 sg13g2_nor2b_1 _19160_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12214_));
 sg13g2_a21oi_1 _19161_ (.A1(net975),
    .A2(_12127_),
    .Y(_12215_),
    .B1(_12214_));
 sg13g2_nor2_1 _19162_ (.A(net396),
    .B(_12124_),
    .Y(_12216_));
 sg13g2_a21oi_1 _19163_ (.A1(net54),
    .A2(_12215_),
    .Y(_00449_),
    .B1(_12216_));
 sg13g2_buf_1 _19164_ (.A(_09871_),
    .X(_12217_));
 sg13g2_nor2_1 _19165_ (.A(net639),
    .B(_11876_),
    .Y(_12218_));
 sg13g2_buf_1 _19166_ (.A(_12218_),
    .X(_12219_));
 sg13g2_buf_1 _19167_ (.A(_12219_),
    .X(_12220_));
 sg13g2_nor2_1 _19168_ (.A(net639),
    .B(_11682_),
    .Y(_12221_));
 sg13g2_buf_2 _19169_ (.A(_12221_),
    .X(_12222_));
 sg13g2_mux2_1 _19170_ (.A0(\cpu.dcache.r_data[4][0] ),
    .A1(net1053),
    .S(_12222_),
    .X(_12223_));
 sg13g2_nor2_1 _19171_ (.A(_12219_),
    .B(_12223_),
    .Y(_12224_));
 sg13g2_a21oi_1 _19172_ (.A1(_09811_),
    .A2(net51),
    .Y(_00450_),
    .B1(_12224_));
 sg13g2_nand2_1 _19173_ (.Y(_12225_),
    .A(net400),
    .B(_11888_));
 sg13g2_buf_1 _19174_ (.A(_12225_),
    .X(_12226_));
 sg13g2_buf_1 _19175_ (.A(_12226_),
    .X(_12227_));
 sg13g2_nor2_1 _19176_ (.A(net639),
    .B(_11697_),
    .Y(_12228_));
 sg13g2_buf_2 _19177_ (.A(_12228_),
    .X(_12229_));
 sg13g2_nor2b_1 _19178_ (.A(_12229_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12230_));
 sg13g2_a21oi_1 _19179_ (.A1(net974),
    .A2(_12229_),
    .Y(_12231_),
    .B1(_12230_));
 sg13g2_nor2_1 _19180_ (.A(net360),
    .B(_12226_),
    .Y(_12232_));
 sg13g2_a21oi_1 _19181_ (.A1(net50),
    .A2(_12231_),
    .Y(_00451_),
    .B1(_12232_));
 sg13g2_nor2b_1 _19182_ (.A(_12229_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12233_));
 sg13g2_a21oi_1 _19183_ (.A1(net960),
    .A2(_12229_),
    .Y(_12234_),
    .B1(_12233_));
 sg13g2_nor2_1 _19184_ (.A(net359),
    .B(_12226_),
    .Y(_12235_));
 sg13g2_a21oi_1 _19185_ (.A1(net50),
    .A2(_12234_),
    .Y(_00452_),
    .B1(_12235_));
 sg13g2_nor2_2 _19186_ (.A(net639),
    .B(_11733_),
    .Y(_12236_));
 sg13g2_mux2_1 _19187_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(net1062),
    .S(_12236_),
    .X(_12237_));
 sg13g2_nand2_1 _19188_ (.Y(_12238_),
    .A(net50),
    .B(_12237_));
 sg13g2_o21ai_1 _19189_ (.B1(_12238_),
    .Y(_00453_),
    .A1(net358),
    .A2(net50));
 sg13g2_mux2_1 _19190_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(net1055),
    .S(_12236_),
    .X(_12239_));
 sg13g2_nand2_1 _19191_ (.Y(_12240_),
    .A(net50),
    .B(_12239_));
 sg13g2_o21ai_1 _19192_ (.B1(_12240_),
    .Y(_00454_),
    .A1(net357),
    .A2(net50));
 sg13g2_mux2_1 _19193_ (.A0(\cpu.dcache.r_data[4][14] ),
    .A1(net1056),
    .S(_12236_),
    .X(_12241_));
 sg13g2_nand2_1 _19194_ (.Y(_12242_),
    .A(_12226_),
    .B(_12241_));
 sg13g2_o21ai_1 _19195_ (.B1(_12242_),
    .Y(_00455_),
    .A1(net397),
    .A2(net50));
 sg13g2_mux2_1 _19196_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(net1054),
    .S(_12236_),
    .X(_12243_));
 sg13g2_nand2_1 _19197_ (.Y(_12244_),
    .A(_12226_),
    .B(_12243_));
 sg13g2_o21ai_1 _19198_ (.B1(_12244_),
    .Y(_00456_),
    .A1(net356),
    .A2(_12227_));
 sg13g2_buf_1 _19199_ (.A(_09810_),
    .X(_12245_));
 sg13g2_nor2_1 _19200_ (.A(net639),
    .B(_11912_),
    .Y(_12246_));
 sg13g2_buf_2 _19201_ (.A(_12246_),
    .X(_12247_));
 sg13g2_buf_1 _19202_ (.A(_12247_),
    .X(_12248_));
 sg13g2_nor2_1 _19203_ (.A(net639),
    .B(_11769_),
    .Y(_12249_));
 sg13g2_buf_2 _19204_ (.A(_12249_),
    .X(_12250_));
 sg13g2_mux2_1 _19205_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(net1053),
    .S(_12250_),
    .X(_12251_));
 sg13g2_nor2_1 _19206_ (.A(_12247_),
    .B(_12251_),
    .Y(_12252_));
 sg13g2_a21oi_1 _19207_ (.A1(net721),
    .A2(net49),
    .Y(_00457_),
    .B1(_12252_));
 sg13g2_nor2b_1 _19208_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12253_));
 sg13g2_a21oi_1 _19209_ (.A1(net961),
    .A2(_12250_),
    .Y(_12254_),
    .B1(_12253_));
 sg13g2_nand2_1 _19210_ (.Y(_12255_),
    .A(net847),
    .B(net49));
 sg13g2_o21ai_1 _19211_ (.B1(_12255_),
    .Y(_00458_),
    .A1(net49),
    .A2(_12254_));
 sg13g2_nor2b_1 _19212_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12256_));
 sg13g2_a21oi_1 _19213_ (.A1(net966),
    .A2(_12250_),
    .Y(_12257_),
    .B1(_12256_));
 sg13g2_nand2_1 _19214_ (.Y(_12258_),
    .A(net846),
    .B(net49));
 sg13g2_o21ai_1 _19215_ (.B1(_12258_),
    .Y(_00459_),
    .A1(net49),
    .A2(_12257_));
 sg13g2_mux2_1 _19216_ (.A0(\cpu.dcache.r_data[4][19] ),
    .A1(net962),
    .S(_12250_),
    .X(_12259_));
 sg13g2_nor2_1 _19217_ (.A(_12247_),
    .B(_12259_),
    .Y(_12260_));
 sg13g2_a21oi_1 _19218_ (.A1(net724),
    .A2(net49),
    .Y(_00460_),
    .B1(_12260_));
 sg13g2_nor2b_1 _19219_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12261_));
 sg13g2_a21oi_1 _19220_ (.A1(_12150_),
    .A2(_12222_),
    .Y(_12262_),
    .B1(_12261_));
 sg13g2_buf_1 _19221_ (.A(_09818_),
    .X(_12263_));
 sg13g2_nand2_1 _19222_ (.Y(_12264_),
    .A(net959),
    .B(net51));
 sg13g2_o21ai_1 _19223_ (.B1(_12264_),
    .Y(_00461_),
    .A1(net51),
    .A2(_12262_));
 sg13g2_nor2_1 _19224_ (.A(net639),
    .B(_11796_),
    .Y(_12265_));
 sg13g2_buf_2 _19225_ (.A(_12265_),
    .X(_12266_));
 sg13g2_nor2b_1 _19226_ (.A(_12266_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12267_));
 sg13g2_a21oi_1 _19227_ (.A1(net965),
    .A2(_12266_),
    .Y(_12268_),
    .B1(_12267_));
 sg13g2_nand2_1 _19228_ (.Y(_12269_),
    .A(net964),
    .B(_12247_));
 sg13g2_o21ai_1 _19229_ (.B1(_12269_),
    .Y(_00462_),
    .A1(_12248_),
    .A2(_12268_));
 sg13g2_nor2b_1 _19230_ (.A(_12266_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12270_));
 sg13g2_a21oi_1 _19231_ (.A1(net961),
    .A2(_12266_),
    .Y(_12271_),
    .B1(_12270_));
 sg13g2_nand2_1 _19232_ (.Y(_12272_),
    .A(net963),
    .B(_12247_));
 sg13g2_o21ai_1 _19233_ (.B1(_12272_),
    .Y(_00463_),
    .A1(net49),
    .A2(_12271_));
 sg13g2_mux2_1 _19234_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(net978),
    .S(_12266_),
    .X(_12273_));
 sg13g2_nor2_1 _19235_ (.A(_12247_),
    .B(_12273_),
    .Y(_12274_));
 sg13g2_a21oi_1 _19236_ (.A1(net723),
    .A2(net49),
    .Y(_00464_),
    .B1(_12274_));
 sg13g2_mux2_1 _19237_ (.A0(\cpu.dcache.r_data[4][23] ),
    .A1(net962),
    .S(_12266_),
    .X(_12275_));
 sg13g2_nor2_1 _19238_ (.A(_12247_),
    .B(_12275_),
    .Y(_12276_));
 sg13g2_a21oi_1 _19239_ (.A1(net722),
    .A2(_12248_),
    .Y(_00465_),
    .B1(_12276_));
 sg13g2_nand2_1 _19240_ (.Y(_12277_),
    .A(net400),
    .B(_11659_));
 sg13g2_buf_1 _19241_ (.A(_12277_),
    .X(_12278_));
 sg13g2_mux2_1 _19242_ (.A0(_11674_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net331),
    .X(_12279_));
 sg13g2_nand2_1 _19243_ (.Y(_12280_),
    .A(net400),
    .B(_11946_));
 sg13g2_buf_1 _19244_ (.A(_12280_),
    .X(_12281_));
 sg13g2_mux2_1 _19245_ (.A0(net355),
    .A1(_12279_),
    .S(net76),
    .X(_00466_));
 sg13g2_mux2_1 _19246_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net331),
    .X(_12282_));
 sg13g2_mux2_1 _19247_ (.A0(net396),
    .A1(_12282_),
    .S(net76),
    .X(_00467_));
 sg13g2_mux2_1 _19248_ (.A0(_11810_),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net331),
    .X(_12283_));
 sg13g2_mux2_1 _19249_ (.A0(net360),
    .A1(_12283_),
    .S(_12281_),
    .X(_00468_));
 sg13g2_mux2_1 _19250_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(net331),
    .X(_12284_));
 sg13g2_mux2_1 _19251_ (.A0(_11722_),
    .A1(_12284_),
    .S(_12281_),
    .X(_00469_));
 sg13g2_nor2_2 _19252_ (.A(_12217_),
    .B(_11836_),
    .Y(_12285_));
 sg13g2_mux2_1 _19253_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(_11728_),
    .S(_12285_),
    .X(_12286_));
 sg13g2_nand2_1 _19254_ (.Y(_12287_),
    .A(net76),
    .B(_12286_));
 sg13g2_o21ai_1 _19255_ (.B1(_12287_),
    .Y(_00470_),
    .A1(_11727_),
    .A2(net76));
 sg13g2_mux2_1 _19256_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(_11903_),
    .S(_12285_),
    .X(_12288_));
 sg13g2_nand2_1 _19257_ (.Y(_12289_),
    .A(net76),
    .B(_12288_));
 sg13g2_o21ai_1 _19258_ (.B1(_12289_),
    .Y(_00471_),
    .A1(_11741_),
    .A2(net76));
 sg13g2_nor2b_1 _19259_ (.A(_12222_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12290_));
 sg13g2_a21oi_1 _19260_ (.A1(_11923_),
    .A2(_12222_),
    .Y(_12291_),
    .B1(_12290_));
 sg13g2_buf_1 _19261_ (.A(_09826_),
    .X(_12292_));
 sg13g2_nand2_1 _19262_ (.Y(_12293_),
    .A(net844),
    .B(net51));
 sg13g2_o21ai_1 _19263_ (.B1(_12293_),
    .Y(_00472_),
    .A1(net51),
    .A2(_12291_));
 sg13g2_mux2_1 _19264_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(_11845_),
    .S(_12285_),
    .X(_12294_));
 sg13g2_nand2_1 _19265_ (.Y(_12295_),
    .A(_12280_),
    .B(_12294_));
 sg13g2_o21ai_1 _19266_ (.B1(_12295_),
    .Y(_00473_),
    .A1(net397),
    .A2(net76));
 sg13g2_mux2_1 _19267_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(net1054),
    .S(_12285_),
    .X(_12296_));
 sg13g2_nand2_1 _19268_ (.Y(_12297_),
    .A(_12280_),
    .B(_12296_));
 sg13g2_o21ai_1 _19269_ (.B1(_12297_),
    .Y(_00474_),
    .A1(_11759_),
    .A2(net76));
 sg13g2_mux2_1 _19270_ (.A0(\cpu.dcache.r_data[4][3] ),
    .A1(net962),
    .S(_12222_),
    .X(_12298_));
 sg13g2_nor2_1 _19271_ (.A(_12219_),
    .B(_12298_),
    .Y(_12299_));
 sg13g2_a21oi_1 _19272_ (.A1(net724),
    .A2(net51),
    .Y(_00475_),
    .B1(_12299_));
 sg13g2_nor2_1 _19273_ (.A(net639),
    .B(_11853_),
    .Y(_12300_));
 sg13g2_buf_2 _19274_ (.A(_12300_),
    .X(_12301_));
 sg13g2_nor2b_1 _19275_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12302_));
 sg13g2_a21oi_1 _19276_ (.A1(net965),
    .A2(_12301_),
    .Y(_12303_),
    .B1(_12302_));
 sg13g2_nand2_1 _19277_ (.Y(_12304_),
    .A(net964),
    .B(_12219_));
 sg13g2_o21ai_1 _19278_ (.B1(_12304_),
    .Y(_00476_),
    .A1(net51),
    .A2(_12303_));
 sg13g2_nor2b_1 _19279_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12305_));
 sg13g2_a21oi_1 _19280_ (.A1(_12150_),
    .A2(_12301_),
    .Y(_12306_),
    .B1(_12305_));
 sg13g2_nand2_1 _19281_ (.Y(_12307_),
    .A(_11988_),
    .B(_12219_));
 sg13g2_o21ai_1 _19282_ (.B1(_12307_),
    .Y(_00477_),
    .A1(net51),
    .A2(_12306_));
 sg13g2_mux2_1 _19283_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(net978),
    .S(_12301_),
    .X(_12308_));
 sg13g2_nor2_1 _19284_ (.A(_12219_),
    .B(_12308_),
    .Y(_12309_));
 sg13g2_a21oi_1 _19285_ (.A1(net723),
    .A2(_12220_),
    .Y(_00478_),
    .B1(_12309_));
 sg13g2_mux2_1 _19286_ (.A0(\cpu.dcache.r_data[4][7] ),
    .A1(net962),
    .S(_12301_),
    .X(_12310_));
 sg13g2_nor2_1 _19287_ (.A(_12219_),
    .B(_12310_),
    .Y(_12311_));
 sg13g2_a21oi_1 _19288_ (.A1(_11813_),
    .A2(_12220_),
    .Y(_00479_),
    .B1(_12311_));
 sg13g2_nor2b_1 _19289_ (.A(_12229_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12312_));
 sg13g2_a21oi_1 _19290_ (.A1(net972),
    .A2(_12229_),
    .Y(_12313_),
    .B1(_12312_));
 sg13g2_nor2_1 _19291_ (.A(net355),
    .B(_12226_),
    .Y(_12314_));
 sg13g2_a21oi_1 _19292_ (.A1(_12227_),
    .A2(_12313_),
    .Y(_00480_),
    .B1(_12314_));
 sg13g2_nor2b_1 _19293_ (.A(_12229_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12315_));
 sg13g2_a21oi_1 _19294_ (.A1(net975),
    .A2(_12229_),
    .Y(_12316_),
    .B1(_12315_));
 sg13g2_nor2_1 _19295_ (.A(net396),
    .B(_12226_),
    .Y(_12317_));
 sg13g2_a21oi_1 _19296_ (.A1(net50),
    .A2(_12316_),
    .Y(_00481_),
    .B1(_12317_));
 sg13g2_buf_1 _19297_ (.A(_09444_),
    .X(_12318_));
 sg13g2_nor2_1 _19298_ (.A(net638),
    .B(_11876_),
    .Y(_12319_));
 sg13g2_buf_2 _19299_ (.A(_12319_),
    .X(_12320_));
 sg13g2_buf_1 _19300_ (.A(_12320_),
    .X(_12321_));
 sg13g2_nor2_1 _19301_ (.A(net638),
    .B(_11682_),
    .Y(_12322_));
 sg13g2_buf_2 _19302_ (.A(_12322_),
    .X(_12323_));
 sg13g2_mux2_1 _19303_ (.A0(\cpu.dcache.r_data[5][0] ),
    .A1(net1053),
    .S(_12323_),
    .X(_12324_));
 sg13g2_nor2_1 _19304_ (.A(_12320_),
    .B(_12324_),
    .Y(_12325_));
 sg13g2_a21oi_1 _19305_ (.A1(net721),
    .A2(_12321_),
    .Y(_00482_),
    .B1(_12325_));
 sg13g2_buf_1 _19306_ (.A(net591),
    .X(_12326_));
 sg13g2_buf_1 _19307_ (.A(net515),
    .X(_12327_));
 sg13g2_buf_1 _19308_ (.A(net455),
    .X(_12328_));
 sg13g2_nand2_1 _19309_ (.Y(_12329_),
    .A(_12328_),
    .B(_11888_));
 sg13g2_buf_2 _19310_ (.A(_12329_),
    .X(_12330_));
 sg13g2_buf_1 _19311_ (.A(_12330_),
    .X(_12331_));
 sg13g2_nor2_1 _19312_ (.A(_12318_),
    .B(_11697_),
    .Y(_12332_));
 sg13g2_buf_2 _19313_ (.A(_12332_),
    .X(_12333_));
 sg13g2_nor2b_1 _19314_ (.A(_12333_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12334_));
 sg13g2_a21oi_1 _19315_ (.A1(net974),
    .A2(_12333_),
    .Y(_12335_),
    .B1(_12334_));
 sg13g2_nor2_1 _19316_ (.A(_11707_),
    .B(_12330_),
    .Y(_12336_));
 sg13g2_a21oi_1 _19317_ (.A1(net47),
    .A2(_12335_),
    .Y(_00483_),
    .B1(_12336_));
 sg13g2_nor2b_1 _19318_ (.A(_12333_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12337_));
 sg13g2_a21oi_1 _19319_ (.A1(net960),
    .A2(_12333_),
    .Y(_12338_),
    .B1(_12337_));
 sg13g2_nor2_1 _19320_ (.A(_11721_),
    .B(_12330_),
    .Y(_12339_));
 sg13g2_a21oi_1 _19321_ (.A1(net47),
    .A2(_12338_),
    .Y(_00484_),
    .B1(_12339_));
 sg13g2_nor2_2 _19322_ (.A(net638),
    .B(_11733_),
    .Y(_12340_));
 sg13g2_mux2_1 _19323_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(net1059),
    .S(_12340_),
    .X(_12341_));
 sg13g2_nand2_1 _19324_ (.Y(_12342_),
    .A(net47),
    .B(_12341_));
 sg13g2_o21ai_1 _19325_ (.B1(_12342_),
    .Y(_00485_),
    .A1(_11726_),
    .A2(net47));
 sg13g2_mux2_1 _19326_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(net1055),
    .S(_12340_),
    .X(_12343_));
 sg13g2_nand2_1 _19327_ (.Y(_12344_),
    .A(net47),
    .B(_12343_));
 sg13g2_o21ai_1 _19328_ (.B1(_12344_),
    .Y(_00486_),
    .A1(_11740_),
    .A2(net47));
 sg13g2_mux2_1 _19329_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(net1056),
    .S(_12340_),
    .X(_12345_));
 sg13g2_nand2_1 _19330_ (.Y(_12346_),
    .A(_12330_),
    .B(_12345_));
 sg13g2_o21ai_1 _19331_ (.B1(_12346_),
    .Y(_00487_),
    .A1(_11749_),
    .A2(net47));
 sg13g2_mux2_1 _19332_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(net1054),
    .S(_12340_),
    .X(_12347_));
 sg13g2_nand2_1 _19333_ (.Y(_12348_),
    .A(_12330_),
    .B(_12347_));
 sg13g2_o21ai_1 _19334_ (.B1(_12348_),
    .Y(_00488_),
    .A1(_11758_),
    .A2(net47));
 sg13g2_nor2_1 _19335_ (.A(net638),
    .B(_11912_),
    .Y(_12349_));
 sg13g2_buf_1 _19336_ (.A(_12349_),
    .X(_12350_));
 sg13g2_buf_1 _19337_ (.A(_12350_),
    .X(_12351_));
 sg13g2_nor2_1 _19338_ (.A(net638),
    .B(_11769_),
    .Y(_12352_));
 sg13g2_buf_2 _19339_ (.A(_12352_),
    .X(_12353_));
 sg13g2_mux2_1 _19340_ (.A0(\cpu.dcache.r_data[5][16] ),
    .A1(net1053),
    .S(_12353_),
    .X(_12354_));
 sg13g2_nor2_1 _19341_ (.A(_12350_),
    .B(_12354_),
    .Y(_12355_));
 sg13g2_a21oi_1 _19342_ (.A1(net721),
    .A2(net46),
    .Y(_00489_),
    .B1(_12355_));
 sg13g2_nor2b_1 _19343_ (.A(_12353_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12356_));
 sg13g2_a21oi_1 _19344_ (.A1(net961),
    .A2(_12353_),
    .Y(_12357_),
    .B1(_12356_));
 sg13g2_nand2_1 _19345_ (.Y(_12358_),
    .A(net959),
    .B(net46));
 sg13g2_o21ai_1 _19346_ (.B1(_12358_),
    .Y(_00490_),
    .A1(net46),
    .A2(_12357_));
 sg13g2_nor2b_1 _19347_ (.A(_12353_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12359_));
 sg13g2_a21oi_1 _19348_ (.A1(net966),
    .A2(_12353_),
    .Y(_12360_),
    .B1(_12359_));
 sg13g2_nand2_1 _19349_ (.Y(_12361_),
    .A(net844),
    .B(net46));
 sg13g2_o21ai_1 _19350_ (.B1(_12361_),
    .Y(_00491_),
    .A1(net46),
    .A2(_12360_));
 sg13g2_buf_1 _19351_ (.A(net849),
    .X(_12362_));
 sg13g2_mux2_1 _19352_ (.A0(\cpu.dcache.r_data[5][19] ),
    .A1(net962),
    .S(_12353_),
    .X(_12363_));
 sg13g2_nor2_1 _19353_ (.A(_12350_),
    .B(_12363_),
    .Y(_12364_));
 sg13g2_a21oi_1 _19354_ (.A1(net720),
    .A2(_12351_),
    .Y(_00492_),
    .B1(_12364_));
 sg13g2_nor2b_1 _19355_ (.A(_12323_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12365_));
 sg13g2_a21oi_1 _19356_ (.A1(net961),
    .A2(_12323_),
    .Y(_12366_),
    .B1(_12365_));
 sg13g2_nand2_1 _19357_ (.Y(_12367_),
    .A(net959),
    .B(net48));
 sg13g2_o21ai_1 _19358_ (.B1(_12367_),
    .Y(_00493_),
    .A1(net48),
    .A2(_12366_));
 sg13g2_nor2_1 _19359_ (.A(net748),
    .B(_11796_),
    .Y(_12368_));
 sg13g2_buf_2 _19360_ (.A(_12368_),
    .X(_12369_));
 sg13g2_nor2b_1 _19361_ (.A(_12369_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_12370_));
 sg13g2_a21oi_1 _19362_ (.A1(net965),
    .A2(_12369_),
    .Y(_12371_),
    .B1(_12370_));
 sg13g2_nand2_1 _19363_ (.Y(_12372_),
    .A(net964),
    .B(_12350_));
 sg13g2_o21ai_1 _19364_ (.B1(_12372_),
    .Y(_00494_),
    .A1(_12351_),
    .A2(_12371_));
 sg13g2_nor2b_1 _19365_ (.A(_12369_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_12373_));
 sg13g2_a21oi_1 _19366_ (.A1(net961),
    .A2(_12369_),
    .Y(_12374_),
    .B1(_12373_));
 sg13g2_nand2_1 _19367_ (.Y(_12375_),
    .A(net963),
    .B(_12350_));
 sg13g2_o21ai_1 _19368_ (.B1(_12375_),
    .Y(_00495_),
    .A1(net46),
    .A2(_12374_));
 sg13g2_buf_1 _19369_ (.A(net845),
    .X(_12376_));
 sg13g2_mux2_1 _19370_ (.A0(\cpu.dcache.r_data[5][22] ),
    .A1(net978),
    .S(_12369_),
    .X(_12377_));
 sg13g2_nor2_1 _19371_ (.A(_12350_),
    .B(_12377_),
    .Y(_12378_));
 sg13g2_a21oi_1 _19372_ (.A1(net719),
    .A2(net46),
    .Y(_00496_),
    .B1(_12378_));
 sg13g2_buf_1 _19373_ (.A(net848),
    .X(_12379_));
 sg13g2_mux2_1 _19374_ (.A0(\cpu.dcache.r_data[5][23] ),
    .A1(net962),
    .S(_12369_),
    .X(_12380_));
 sg13g2_nor2_1 _19375_ (.A(_12350_),
    .B(_12380_),
    .Y(_12381_));
 sg13g2_a21oi_1 _19376_ (.A1(net718),
    .A2(net46),
    .Y(_00497_),
    .B1(_12381_));
 sg13g2_nand2_1 _19377_ (.Y(_12382_),
    .A(_12328_),
    .B(_11946_));
 sg13g2_buf_2 _19378_ (.A(_12382_),
    .X(_12383_));
 sg13g2_buf_1 _19379_ (.A(_12383_),
    .X(_12384_));
 sg13g2_nor2_1 _19380_ (.A(net638),
    .B(_11951_),
    .Y(_12385_));
 sg13g2_buf_1 _19381_ (.A(_12385_),
    .X(_12386_));
 sg13g2_nor2b_1 _19382_ (.A(net514),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_12387_));
 sg13g2_a21oi_1 _19383_ (.A1(net972),
    .A2(net514),
    .Y(_12388_),
    .B1(_12387_));
 sg13g2_nor2_1 _19384_ (.A(_11818_),
    .B(_12383_),
    .Y(_12389_));
 sg13g2_a21oi_1 _19385_ (.A1(net45),
    .A2(_12388_),
    .Y(_00498_),
    .B1(_12389_));
 sg13g2_nor2b_1 _19386_ (.A(net514),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_12390_));
 sg13g2_a21oi_1 _19387_ (.A1(net975),
    .A2(net514),
    .Y(_12391_),
    .B1(_12390_));
 sg13g2_nor2_1 _19388_ (.A(_11829_),
    .B(_12383_),
    .Y(_12392_));
 sg13g2_a21oi_1 _19389_ (.A1(net45),
    .A2(_12391_),
    .Y(_00499_),
    .B1(_12392_));
 sg13g2_nor2b_1 _19390_ (.A(net514),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_12393_));
 sg13g2_a21oi_1 _19391_ (.A1(net974),
    .A2(net514),
    .Y(_12394_),
    .B1(_12393_));
 sg13g2_nor2_1 _19392_ (.A(_11707_),
    .B(_12383_),
    .Y(_12395_));
 sg13g2_a21oi_1 _19393_ (.A1(net45),
    .A2(_12394_),
    .Y(_00500_),
    .B1(_12395_));
 sg13g2_nor2b_1 _19394_ (.A(net514),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_12396_));
 sg13g2_a21oi_1 _19395_ (.A1(net960),
    .A2(net514),
    .Y(_12397_),
    .B1(_12396_));
 sg13g2_nor2_1 _19396_ (.A(_11721_),
    .B(_12383_),
    .Y(_12398_));
 sg13g2_a21oi_1 _19397_ (.A1(net45),
    .A2(_12397_),
    .Y(_00501_),
    .B1(_12398_));
 sg13g2_nor2_2 _19398_ (.A(_12318_),
    .B(_11836_),
    .Y(_12399_));
 sg13g2_mux2_1 _19399_ (.A0(\cpu.dcache.r_data[5][28] ),
    .A1(net1059),
    .S(_12399_),
    .X(_12400_));
 sg13g2_nand2_1 _19400_ (.Y(_12401_),
    .A(net45),
    .B(_12400_));
 sg13g2_o21ai_1 _19401_ (.B1(_12401_),
    .Y(_00502_),
    .A1(_11726_),
    .A2(net45));
 sg13g2_mux2_1 _19402_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(net1055),
    .S(_12399_),
    .X(_12402_));
 sg13g2_nand2_1 _19403_ (.Y(_12403_),
    .A(net45),
    .B(_12402_));
 sg13g2_o21ai_1 _19404_ (.B1(_12403_),
    .Y(_00503_),
    .A1(_11740_),
    .A2(net45));
 sg13g2_nor2b_1 _19405_ (.A(_12323_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_12404_));
 sg13g2_a21oi_1 _19406_ (.A1(net966),
    .A2(_12323_),
    .Y(_12405_),
    .B1(_12404_));
 sg13g2_nand2_1 _19407_ (.Y(_12406_),
    .A(net844),
    .B(net48));
 sg13g2_o21ai_1 _19408_ (.B1(_12406_),
    .Y(_00504_),
    .A1(net48),
    .A2(_12405_));
 sg13g2_mux2_1 _19409_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(_11694_),
    .S(_12399_),
    .X(_12407_));
 sg13g2_nand2_1 _19410_ (.Y(_12408_),
    .A(_12383_),
    .B(_12407_));
 sg13g2_o21ai_1 _19411_ (.B1(_12408_),
    .Y(_00505_),
    .A1(_11749_),
    .A2(_12384_));
 sg13g2_mux2_1 _19412_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(net1054),
    .S(_12399_),
    .X(_12409_));
 sg13g2_nand2_1 _19413_ (.Y(_12410_),
    .A(_12383_),
    .B(_12409_));
 sg13g2_o21ai_1 _19414_ (.B1(_12410_),
    .Y(_00506_),
    .A1(_11758_),
    .A2(_12384_));
 sg13g2_mux2_1 _19415_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(net977),
    .S(_12323_),
    .X(_12411_));
 sg13g2_nor2_1 _19416_ (.A(_12320_),
    .B(_12411_),
    .Y(_12412_));
 sg13g2_a21oi_1 _19417_ (.A1(_12362_),
    .A2(net48),
    .Y(_00507_),
    .B1(_12412_));
 sg13g2_nor2_1 _19418_ (.A(net748),
    .B(_11853_),
    .Y(_12413_));
 sg13g2_buf_2 _19419_ (.A(_12413_),
    .X(_12414_));
 sg13g2_nor2b_1 _19420_ (.A(_12414_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_12415_));
 sg13g2_a21oi_1 _19421_ (.A1(_11932_),
    .A2(_12414_),
    .Y(_12416_),
    .B1(_12415_));
 sg13g2_nand2_1 _19422_ (.Y(_12417_),
    .A(net964),
    .B(_12320_));
 sg13g2_o21ai_1 _19423_ (.B1(_12417_),
    .Y(_00508_),
    .A1(_12321_),
    .A2(_12416_));
 sg13g2_nor2b_1 _19424_ (.A(_12414_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_12418_));
 sg13g2_a21oi_1 _19425_ (.A1(net961),
    .A2(_12414_),
    .Y(_12419_),
    .B1(_12418_));
 sg13g2_nand2_1 _19426_ (.Y(_12420_),
    .A(net963),
    .B(_12320_));
 sg13g2_o21ai_1 _19427_ (.B1(_12420_),
    .Y(_00509_),
    .A1(net48),
    .A2(_12419_));
 sg13g2_mux2_1 _19428_ (.A0(\cpu.dcache.r_data[5][6] ),
    .A1(_11751_),
    .S(_12414_),
    .X(_12421_));
 sg13g2_nor2_1 _19429_ (.A(_12320_),
    .B(_12421_),
    .Y(_12422_));
 sg13g2_a21oi_1 _19430_ (.A1(net719),
    .A2(net48),
    .Y(_00510_),
    .B1(_12422_));
 sg13g2_mux2_1 _19431_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(net977),
    .S(_12414_),
    .X(_12423_));
 sg13g2_nor2_1 _19432_ (.A(_12320_),
    .B(_12423_),
    .Y(_12424_));
 sg13g2_a21oi_1 _19433_ (.A1(net718),
    .A2(net48),
    .Y(_00511_),
    .B1(_12424_));
 sg13g2_nor2b_1 _19434_ (.A(_12333_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_12425_));
 sg13g2_a21oi_1 _19435_ (.A1(net972),
    .A2(_12333_),
    .Y(_12426_),
    .B1(_12425_));
 sg13g2_nor2_1 _19436_ (.A(_11818_),
    .B(_12330_),
    .Y(_12427_));
 sg13g2_a21oi_1 _19437_ (.A1(_12331_),
    .A2(_12426_),
    .Y(_00512_),
    .B1(_12427_));
 sg13g2_nor2b_1 _19438_ (.A(_12333_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_12428_));
 sg13g2_a21oi_1 _19439_ (.A1(net975),
    .A2(_12333_),
    .Y(_12429_),
    .B1(_12428_));
 sg13g2_nor2_1 _19440_ (.A(_11829_),
    .B(_12330_),
    .Y(_12430_));
 sg13g2_a21oi_1 _19441_ (.A1(_12331_),
    .A2(_12429_),
    .Y(_00513_),
    .B1(_12430_));
 sg13g2_buf_1 _19442_ (.A(_09433_),
    .X(_12431_));
 sg13g2_nor2_1 _19443_ (.A(net717),
    .B(_11876_),
    .Y(_12432_));
 sg13g2_buf_1 _19444_ (.A(_12432_),
    .X(_12433_));
 sg13g2_buf_1 _19445_ (.A(_12433_),
    .X(_12434_));
 sg13g2_nor2_1 _19446_ (.A(net717),
    .B(_11682_),
    .Y(_12435_));
 sg13g2_buf_2 _19447_ (.A(_12435_),
    .X(_12436_));
 sg13g2_mux2_1 _19448_ (.A0(\cpu.dcache.r_data[6][0] ),
    .A1(net1053),
    .S(_12436_),
    .X(_12437_));
 sg13g2_nor2_1 _19449_ (.A(_12433_),
    .B(_12437_),
    .Y(_12438_));
 sg13g2_a21oi_1 _19450_ (.A1(net721),
    .A2(net44),
    .Y(_00514_),
    .B1(_12438_));
 sg13g2_buf_1 _19451_ (.A(net533),
    .X(_12439_));
 sg13g2_buf_1 _19452_ (.A(net454),
    .X(_12440_));
 sg13g2_buf_1 _19453_ (.A(net391),
    .X(_12441_));
 sg13g2_nand2_1 _19454_ (.Y(_12442_),
    .A(net353),
    .B(_11888_));
 sg13g2_buf_2 _19455_ (.A(_12442_),
    .X(_12443_));
 sg13g2_buf_1 _19456_ (.A(_12443_),
    .X(_12444_));
 sg13g2_nor2_1 _19457_ (.A(net717),
    .B(_11697_),
    .Y(_12445_));
 sg13g2_buf_2 _19458_ (.A(_12445_),
    .X(_12446_));
 sg13g2_nor2b_1 _19459_ (.A(_12446_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_12447_));
 sg13g2_a21oi_1 _19460_ (.A1(net974),
    .A2(_12446_),
    .Y(_12448_),
    .B1(_12447_));
 sg13g2_nor2_1 _19461_ (.A(_11707_),
    .B(_12443_),
    .Y(_12449_));
 sg13g2_a21oi_1 _19462_ (.A1(_12444_),
    .A2(_12448_),
    .Y(_00515_),
    .B1(_12449_));
 sg13g2_nor2b_1 _19463_ (.A(_12446_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_12450_));
 sg13g2_a21oi_1 _19464_ (.A1(net960),
    .A2(_12446_),
    .Y(_12451_),
    .B1(_12450_));
 sg13g2_nor2_1 _19465_ (.A(_11721_),
    .B(_12443_),
    .Y(_12452_));
 sg13g2_a21oi_1 _19466_ (.A1(net43),
    .A2(_12451_),
    .Y(_00516_),
    .B1(_12452_));
 sg13g2_nor2_2 _19467_ (.A(net717),
    .B(_11733_),
    .Y(_12453_));
 sg13g2_mux2_1 _19468_ (.A0(\cpu.dcache.r_data[6][12] ),
    .A1(net1059),
    .S(_12453_),
    .X(_12454_));
 sg13g2_nand2_1 _19469_ (.Y(_12455_),
    .A(net43),
    .B(_12454_));
 sg13g2_o21ai_1 _19470_ (.B1(_12455_),
    .Y(_00517_),
    .A1(_11726_),
    .A2(net43));
 sg13g2_mux2_1 _19471_ (.A0(\cpu.dcache.r_data[6][13] ),
    .A1(net1060),
    .S(_12453_),
    .X(_12456_));
 sg13g2_nand2_1 _19472_ (.Y(_12457_),
    .A(net43),
    .B(_12456_));
 sg13g2_o21ai_1 _19473_ (.B1(_12457_),
    .Y(_00518_),
    .A1(_11740_),
    .A2(net43));
 sg13g2_mux2_1 _19474_ (.A0(\cpu.dcache.r_data[6][14] ),
    .A1(net1064),
    .S(_12453_),
    .X(_12458_));
 sg13g2_nand2_1 _19475_ (.Y(_12459_),
    .A(_12443_),
    .B(_12458_));
 sg13g2_o21ai_1 _19476_ (.B1(_12459_),
    .Y(_00519_),
    .A1(_11749_),
    .A2(net43));
 sg13g2_mux2_1 _19477_ (.A0(\cpu.dcache.r_data[6][15] ),
    .A1(_11711_),
    .S(_12453_),
    .X(_12460_));
 sg13g2_nand2_1 _19478_ (.Y(_12461_),
    .A(_12443_),
    .B(_12460_));
 sg13g2_o21ai_1 _19479_ (.B1(_12461_),
    .Y(_00520_),
    .A1(_11758_),
    .A2(net43));
 sg13g2_nor2_1 _19480_ (.A(net717),
    .B(_11912_),
    .Y(_12462_));
 sg13g2_buf_2 _19481_ (.A(_12462_),
    .X(_12463_));
 sg13g2_buf_1 _19482_ (.A(_12463_),
    .X(_12464_));
 sg13g2_nor2_1 _19483_ (.A(net717),
    .B(_11769_),
    .Y(_12465_));
 sg13g2_buf_2 _19484_ (.A(_12465_),
    .X(_12466_));
 sg13g2_mux2_1 _19485_ (.A0(\cpu.dcache.r_data[6][16] ),
    .A1(net1053),
    .S(_12466_),
    .X(_12467_));
 sg13g2_nor2_1 _19486_ (.A(_12463_),
    .B(_12467_),
    .Y(_12468_));
 sg13g2_a21oi_1 _19487_ (.A1(net721),
    .A2(net42),
    .Y(_00521_),
    .B1(_12468_));
 sg13g2_buf_1 _19488_ (.A(net1060),
    .X(_12469_));
 sg13g2_nor2b_1 _19489_ (.A(_12466_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_12470_));
 sg13g2_a21oi_1 _19490_ (.A1(net958),
    .A2(_12466_),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_nand2_1 _19491_ (.Y(_12472_),
    .A(net959),
    .B(net42));
 sg13g2_o21ai_1 _19492_ (.B1(_12472_),
    .Y(_00522_),
    .A1(net42),
    .A2(_12471_));
 sg13g2_buf_1 _19493_ (.A(net1064),
    .X(_12473_));
 sg13g2_nor2b_1 _19494_ (.A(_12466_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_12474_));
 sg13g2_a21oi_1 _19495_ (.A1(net957),
    .A2(_12466_),
    .Y(_12475_),
    .B1(_12474_));
 sg13g2_nand2_1 _19496_ (.Y(_12476_),
    .A(net844),
    .B(net42));
 sg13g2_o21ai_1 _19497_ (.B1(_12476_),
    .Y(_00523_),
    .A1(net42),
    .A2(_12475_));
 sg13g2_mux2_1 _19498_ (.A0(\cpu.dcache.r_data[6][19] ),
    .A1(net977),
    .S(_12466_),
    .X(_12477_));
 sg13g2_nor2_1 _19499_ (.A(_12463_),
    .B(_12477_),
    .Y(_12478_));
 sg13g2_a21oi_1 _19500_ (.A1(net720),
    .A2(net42),
    .Y(_00524_),
    .B1(_12478_));
 sg13g2_nor2b_1 _19501_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_12479_));
 sg13g2_a21oi_1 _19502_ (.A1(net958),
    .A2(_12436_),
    .Y(_12480_),
    .B1(_12479_));
 sg13g2_nand2_1 _19503_ (.Y(_12481_),
    .A(net959),
    .B(net44));
 sg13g2_o21ai_1 _19504_ (.B1(_12481_),
    .Y(_00525_),
    .A1(net44),
    .A2(_12480_));
 sg13g2_nor2_1 _19505_ (.A(_09433_),
    .B(_11796_),
    .Y(_12482_));
 sg13g2_buf_2 _19506_ (.A(_12482_),
    .X(_12483_));
 sg13g2_nor2b_1 _19507_ (.A(_12483_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_12484_));
 sg13g2_a21oi_1 _19508_ (.A1(net965),
    .A2(_12483_),
    .Y(_12485_),
    .B1(_12484_));
 sg13g2_nand2_1 _19509_ (.Y(_12486_),
    .A(net964),
    .B(_12463_));
 sg13g2_o21ai_1 _19510_ (.B1(_12486_),
    .Y(_00526_),
    .A1(_12464_),
    .A2(_12485_));
 sg13g2_nor2b_1 _19511_ (.A(_12483_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_12487_));
 sg13g2_a21oi_1 _19512_ (.A1(net958),
    .A2(_12483_),
    .Y(_12488_),
    .B1(_12487_));
 sg13g2_nand2_1 _19513_ (.Y(_12489_),
    .A(net963),
    .B(_12463_));
 sg13g2_o21ai_1 _19514_ (.B1(_12489_),
    .Y(_00527_),
    .A1(_12464_),
    .A2(_12488_));
 sg13g2_mux2_1 _19515_ (.A0(\cpu.dcache.r_data[6][22] ),
    .A1(net978),
    .S(_12483_),
    .X(_12490_));
 sg13g2_nor2_1 _19516_ (.A(_12463_),
    .B(_12490_),
    .Y(_12491_));
 sg13g2_a21oi_1 _19517_ (.A1(net719),
    .A2(net42),
    .Y(_00528_),
    .B1(_12491_));
 sg13g2_mux2_1 _19518_ (.A0(\cpu.dcache.r_data[6][23] ),
    .A1(net977),
    .S(_12483_),
    .X(_12492_));
 sg13g2_nor2_1 _19519_ (.A(_12463_),
    .B(_12492_),
    .Y(_02684_));
 sg13g2_a21oi_1 _19520_ (.A1(net718),
    .A2(net42),
    .Y(_00529_),
    .B1(_02684_));
 sg13g2_nand2_1 _19521_ (.Y(_02685_),
    .A(net353),
    .B(_11946_));
 sg13g2_buf_2 _19522_ (.A(_02685_),
    .X(_02686_));
 sg13g2_buf_1 _19523_ (.A(_02686_),
    .X(_02687_));
 sg13g2_nor2_1 _19524_ (.A(_09433_),
    .B(_11951_),
    .Y(_02688_));
 sg13g2_buf_1 _19525_ (.A(_02688_),
    .X(_02689_));
 sg13g2_buf_1 _19526_ (.A(_02689_),
    .X(_02690_));
 sg13g2_nor2b_1 _19527_ (.A(net453),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02691_));
 sg13g2_a21oi_1 _19528_ (.A1(net972),
    .A2(net453),
    .Y(_02692_),
    .B1(_02691_));
 sg13g2_nor2_1 _19529_ (.A(_11818_),
    .B(_02686_),
    .Y(_02693_));
 sg13g2_a21oi_1 _19530_ (.A1(net41),
    .A2(_02692_),
    .Y(_00530_),
    .B1(_02693_));
 sg13g2_nor2b_1 _19531_ (.A(net453),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02694_));
 sg13g2_a21oi_1 _19532_ (.A1(net975),
    .A2(net453),
    .Y(_02695_),
    .B1(_02694_));
 sg13g2_nor2_1 _19533_ (.A(_11829_),
    .B(_02686_),
    .Y(_02696_));
 sg13g2_a21oi_1 _19534_ (.A1(net41),
    .A2(_02695_),
    .Y(_00531_),
    .B1(_02696_));
 sg13g2_nor2b_1 _19535_ (.A(net453),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02697_));
 sg13g2_a21oi_1 _19536_ (.A1(_11780_),
    .A2(net453),
    .Y(_02698_),
    .B1(_02697_));
 sg13g2_nor2_1 _19537_ (.A(_11707_),
    .B(_02686_),
    .Y(_02699_));
 sg13g2_a21oi_1 _19538_ (.A1(_02687_),
    .A2(_02698_),
    .Y(_00532_),
    .B1(_02699_));
 sg13g2_nor2b_1 _19539_ (.A(_02689_),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02700_));
 sg13g2_a21oi_1 _19540_ (.A1(net960),
    .A2(net453),
    .Y(_02701_),
    .B1(_02700_));
 sg13g2_nor2_1 _19541_ (.A(_11721_),
    .B(_02686_),
    .Y(_02702_));
 sg13g2_a21oi_1 _19542_ (.A1(_02687_),
    .A2(_02701_),
    .Y(_00533_),
    .B1(_02702_));
 sg13g2_nor2_2 _19543_ (.A(net717),
    .B(_11836_),
    .Y(_02703_));
 sg13g2_mux2_1 _19544_ (.A0(\cpu.dcache.r_data[6][28] ),
    .A1(_11792_),
    .S(_02703_),
    .X(_02704_));
 sg13g2_nand2_1 _19545_ (.Y(_02705_),
    .A(net41),
    .B(_02704_));
 sg13g2_o21ai_1 _19546_ (.B1(_02705_),
    .Y(_00534_),
    .A1(_11726_),
    .A2(net41));
 sg13g2_mux2_1 _19547_ (.A0(\cpu.dcache.r_data[6][29] ),
    .A1(net1060),
    .S(_02703_),
    .X(_02706_));
 sg13g2_nand2_1 _19548_ (.Y(_02707_),
    .A(net41),
    .B(_02706_));
 sg13g2_o21ai_1 _19549_ (.B1(_02707_),
    .Y(_00535_),
    .A1(_11740_),
    .A2(net41));
 sg13g2_nor2b_1 _19550_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02708_));
 sg13g2_a21oi_1 _19551_ (.A1(net957),
    .A2(_12436_),
    .Y(_02709_),
    .B1(_02708_));
 sg13g2_nand2_1 _19552_ (.Y(_02710_),
    .A(net844),
    .B(net44));
 sg13g2_o21ai_1 _19553_ (.B1(_02710_),
    .Y(_00536_),
    .A1(net44),
    .A2(_02709_));
 sg13g2_mux2_1 _19554_ (.A0(\cpu.dcache.r_data[6][30] ),
    .A1(net1064),
    .S(_02703_),
    .X(_02711_));
 sg13g2_nand2_1 _19555_ (.Y(_02712_),
    .A(_02686_),
    .B(_02711_));
 sg13g2_o21ai_1 _19556_ (.B1(_02712_),
    .Y(_00537_),
    .A1(_11749_),
    .A2(net41));
 sg13g2_mux2_1 _19557_ (.A0(\cpu.dcache.r_data[6][31] ),
    .A1(net1063),
    .S(_02703_),
    .X(_02713_));
 sg13g2_nand2_1 _19558_ (.Y(_02714_),
    .A(_02686_),
    .B(_02713_));
 sg13g2_o21ai_1 _19559_ (.B1(_02714_),
    .Y(_00538_),
    .A1(_11758_),
    .A2(net41));
 sg13g2_mux2_1 _19560_ (.A0(\cpu.dcache.r_data[6][3] ),
    .A1(net977),
    .S(_12436_),
    .X(_02715_));
 sg13g2_nor2_1 _19561_ (.A(_12433_),
    .B(_02715_),
    .Y(_02716_));
 sg13g2_a21oi_1 _19562_ (.A1(net720),
    .A2(_12434_),
    .Y(_00539_),
    .B1(_02716_));
 sg13g2_nor2_1 _19563_ (.A(_09433_),
    .B(_11853_),
    .Y(_02717_));
 sg13g2_buf_2 _19564_ (.A(_02717_),
    .X(_02718_));
 sg13g2_nor2b_1 _19565_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02719_));
 sg13g2_a21oi_1 _19566_ (.A1(_11932_),
    .A2(_02718_),
    .Y(_02720_),
    .B1(_02719_));
 sg13g2_nand2_1 _19567_ (.Y(_02721_),
    .A(_11984_),
    .B(_12433_));
 sg13g2_o21ai_1 _19568_ (.B1(_02721_),
    .Y(_00540_),
    .A1(net44),
    .A2(_02720_));
 sg13g2_nor2b_1 _19569_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02722_));
 sg13g2_a21oi_1 _19570_ (.A1(net958),
    .A2(_02718_),
    .Y(_02723_),
    .B1(_02722_));
 sg13g2_nand2_1 _19571_ (.Y(_02724_),
    .A(net963),
    .B(_12433_));
 sg13g2_o21ai_1 _19572_ (.B1(_02724_),
    .Y(_00541_),
    .A1(net44),
    .A2(_02723_));
 sg13g2_mux2_1 _19573_ (.A0(\cpu.dcache.r_data[6][6] ),
    .A1(_11751_),
    .S(_02718_),
    .X(_02725_));
 sg13g2_nor2_1 _19574_ (.A(_12433_),
    .B(_02725_),
    .Y(_02726_));
 sg13g2_a21oi_1 _19575_ (.A1(net719),
    .A2(net44),
    .Y(_00542_),
    .B1(_02726_));
 sg13g2_mux2_1 _19576_ (.A0(\cpu.dcache.r_data[6][7] ),
    .A1(net977),
    .S(_02718_),
    .X(_02727_));
 sg13g2_nor2_1 _19577_ (.A(_12433_),
    .B(_02727_),
    .Y(_02728_));
 sg13g2_a21oi_1 _19578_ (.A1(_12379_),
    .A2(_12434_),
    .Y(_00543_),
    .B1(_02728_));
 sg13g2_nor2b_1 _19579_ (.A(_12446_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02729_));
 sg13g2_a21oi_1 _19580_ (.A1(net972),
    .A2(_12446_),
    .Y(_02730_),
    .B1(_02729_));
 sg13g2_nor2_1 _19581_ (.A(_11818_),
    .B(_12443_),
    .Y(_02731_));
 sg13g2_a21oi_1 _19582_ (.A1(_12444_),
    .A2(_02730_),
    .Y(_00544_),
    .B1(_02731_));
 sg13g2_nor2b_1 _19583_ (.A(_12446_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02732_));
 sg13g2_a21oi_1 _19584_ (.A1(net975),
    .A2(_12446_),
    .Y(_02733_),
    .B1(_02732_));
 sg13g2_nor2_1 _19585_ (.A(_11829_),
    .B(_12443_),
    .Y(_02734_));
 sg13g2_a21oi_1 _19586_ (.A1(net43),
    .A2(_02733_),
    .Y(_00545_),
    .B1(_02734_));
 sg13g2_buf_1 _19587_ (.A(_09731_),
    .X(_02735_));
 sg13g2_nor2_1 _19588_ (.A(net567),
    .B(_11876_),
    .Y(_02736_));
 sg13g2_buf_1 _19589_ (.A(_02736_),
    .X(_02737_));
 sg13g2_buf_1 _19590_ (.A(_02737_),
    .X(_02738_));
 sg13g2_nor2_1 _19591_ (.A(net567),
    .B(_11682_),
    .Y(_02739_));
 sg13g2_buf_2 _19592_ (.A(_02739_),
    .X(_02740_));
 sg13g2_mux2_1 _19593_ (.A0(\cpu.dcache.r_data[7][0] ),
    .A1(_12116_),
    .S(_02740_),
    .X(_02741_));
 sg13g2_nor2_1 _19594_ (.A(_02737_),
    .B(_02741_),
    .Y(_02742_));
 sg13g2_a21oi_1 _19595_ (.A1(net721),
    .A2(net40),
    .Y(_00546_),
    .B1(_02742_));
 sg13g2_buf_1 _19596_ (.A(_09212_),
    .X(_02743_));
 sg13g2_buf_1 _19597_ (.A(net513),
    .X(_02744_));
 sg13g2_buf_1 _19598_ (.A(net452),
    .X(_02745_));
 sg13g2_nand2_1 _19599_ (.Y(_02746_),
    .A(net390),
    .B(_11888_));
 sg13g2_buf_1 _19600_ (.A(_02746_),
    .X(_02747_));
 sg13g2_buf_1 _19601_ (.A(_02747_),
    .X(_02748_));
 sg13g2_nor2_1 _19602_ (.A(net567),
    .B(_11697_),
    .Y(_02749_));
 sg13g2_buf_2 _19603_ (.A(_02749_),
    .X(_02750_));
 sg13g2_nor2b_1 _19604_ (.A(_02750_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02751_));
 sg13g2_a21oi_1 _19605_ (.A1(net974),
    .A2(_02750_),
    .Y(_02752_),
    .B1(_02751_));
 sg13g2_nor2_1 _19606_ (.A(_11707_),
    .B(_02747_),
    .Y(_02753_));
 sg13g2_a21oi_1 _19607_ (.A1(net39),
    .A2(_02752_),
    .Y(_00547_),
    .B1(_02753_));
 sg13g2_nor2b_1 _19608_ (.A(_02750_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02754_));
 sg13g2_a21oi_1 _19609_ (.A1(net960),
    .A2(_02750_),
    .Y(_02755_),
    .B1(_02754_));
 sg13g2_nor2_1 _19610_ (.A(_11721_),
    .B(_02747_),
    .Y(_02756_));
 sg13g2_a21oi_1 _19611_ (.A1(net39),
    .A2(_02755_),
    .Y(_00548_),
    .B1(_02756_));
 sg13g2_nor2_2 _19612_ (.A(_02735_),
    .B(_11733_),
    .Y(_02757_));
 sg13g2_mux2_1 _19613_ (.A0(\cpu.dcache.r_data[7][12] ),
    .A1(net1059),
    .S(_02757_),
    .X(_02758_));
 sg13g2_nand2_1 _19614_ (.Y(_02759_),
    .A(net39),
    .B(_02758_));
 sg13g2_o21ai_1 _19615_ (.B1(_02759_),
    .Y(_00549_),
    .A1(_11726_),
    .A2(net39));
 sg13g2_mux2_1 _19616_ (.A0(\cpu.dcache.r_data[7][13] ),
    .A1(net1060),
    .S(_02757_),
    .X(_02760_));
 sg13g2_nand2_1 _19617_ (.Y(_02761_),
    .A(net39),
    .B(_02760_));
 sg13g2_o21ai_1 _19618_ (.B1(_02761_),
    .Y(_00550_),
    .A1(_11740_),
    .A2(net39));
 sg13g2_mux2_1 _19619_ (.A0(\cpu.dcache.r_data[7][14] ),
    .A1(net1064),
    .S(_02757_),
    .X(_02762_));
 sg13g2_nand2_1 _19620_ (.Y(_02763_),
    .A(_02747_),
    .B(_02762_));
 sg13g2_o21ai_1 _19621_ (.B1(_02763_),
    .Y(_00551_),
    .A1(_11749_),
    .A2(net39));
 sg13g2_mux2_1 _19622_ (.A0(\cpu.dcache.r_data[7][15] ),
    .A1(net1063),
    .S(_02757_),
    .X(_02764_));
 sg13g2_nand2_1 _19623_ (.Y(_02765_),
    .A(_02747_),
    .B(_02764_));
 sg13g2_o21ai_1 _19624_ (.B1(_02765_),
    .Y(_00552_),
    .A1(_11758_),
    .A2(net39));
 sg13g2_nor2_1 _19625_ (.A(net567),
    .B(_11912_),
    .Y(_02766_));
 sg13g2_buf_1 _19626_ (.A(_02766_),
    .X(_02767_));
 sg13g2_buf_1 _19627_ (.A(_02767_),
    .X(_02768_));
 sg13g2_nor2_1 _19628_ (.A(net567),
    .B(_11769_),
    .Y(_02769_));
 sg13g2_buf_2 _19629_ (.A(_02769_),
    .X(_02770_));
 sg13g2_mux2_1 _19630_ (.A0(\cpu.dcache.r_data[7][16] ),
    .A1(_12116_),
    .S(_02770_),
    .X(_02771_));
 sg13g2_nor2_1 _19631_ (.A(_02767_),
    .B(_02771_),
    .Y(_02772_));
 sg13g2_a21oi_1 _19632_ (.A1(net721),
    .A2(net38),
    .Y(_00553_),
    .B1(_02772_));
 sg13g2_nor2b_1 _19633_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02773_));
 sg13g2_a21oi_1 _19634_ (.A1(net958),
    .A2(_02770_),
    .Y(_02774_),
    .B1(_02773_));
 sg13g2_nand2_1 _19635_ (.Y(_02775_),
    .A(net959),
    .B(net38));
 sg13g2_o21ai_1 _19636_ (.B1(_02775_),
    .Y(_00554_),
    .A1(net38),
    .A2(_02774_));
 sg13g2_nor2b_1 _19637_ (.A(_02770_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02776_));
 sg13g2_a21oi_1 _19638_ (.A1(net957),
    .A2(_02770_),
    .Y(_02777_),
    .B1(_02776_));
 sg13g2_nand2_1 _19639_ (.Y(_02778_),
    .A(net844),
    .B(net38));
 sg13g2_o21ai_1 _19640_ (.B1(_02778_),
    .Y(_00555_),
    .A1(net38),
    .A2(_02777_));
 sg13g2_mux2_1 _19641_ (.A0(\cpu.dcache.r_data[7][19] ),
    .A1(net977),
    .S(_02770_),
    .X(_02779_));
 sg13g2_nor2_1 _19642_ (.A(_02767_),
    .B(_02779_),
    .Y(_02780_));
 sg13g2_a21oi_1 _19643_ (.A1(net720),
    .A2(net38),
    .Y(_00556_),
    .B1(_02780_));
 sg13g2_nor2b_1 _19644_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02781_));
 sg13g2_a21oi_1 _19645_ (.A1(net958),
    .A2(_02740_),
    .Y(_02782_),
    .B1(_02781_));
 sg13g2_nand2_1 _19646_ (.Y(_02783_),
    .A(net959),
    .B(net40));
 sg13g2_o21ai_1 _19647_ (.B1(_02783_),
    .Y(_00557_),
    .A1(net40),
    .A2(_02782_));
 sg13g2_or2_1 _19648_ (.X(_02784_),
    .B(_11796_),
    .A(_09731_));
 sg13g2_buf_1 _19649_ (.A(_02784_),
    .X(_02785_));
 sg13g2_mux2_1 _19650_ (.A0(net1065),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02785_),
    .X(_02786_));
 sg13g2_mux2_1 _19651_ (.A0(_02786_),
    .A1(_11801_),
    .S(_02768_),
    .X(_00558_));
 sg13g2_mux2_1 _19652_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02785_),
    .X(_02787_));
 sg13g2_mux2_1 _19653_ (.A0(_02787_),
    .A1(net969),
    .S(net38),
    .X(_00559_));
 sg13g2_mux2_1 _19654_ (.A0(net1058),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02785_),
    .X(_02788_));
 sg13g2_nor2_1 _19655_ (.A(_02767_),
    .B(_02788_),
    .Y(_02789_));
 sg13g2_a21oi_1 _19656_ (.A1(net719),
    .A2(net38),
    .Y(_00560_),
    .B1(_02789_));
 sg13g2_mux2_1 _19657_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02785_),
    .X(_02790_));
 sg13g2_nor2_1 _19658_ (.A(_02767_),
    .B(_02790_),
    .Y(_02791_));
 sg13g2_a21oi_1 _19659_ (.A1(net718),
    .A2(_02768_),
    .Y(_00561_),
    .B1(_02791_));
 sg13g2_nand2_1 _19660_ (.Y(_02792_),
    .A(net390),
    .B(_11946_));
 sg13g2_buf_1 _19661_ (.A(_02792_),
    .X(_02793_));
 sg13g2_buf_1 _19662_ (.A(_02793_),
    .X(_02794_));
 sg13g2_nor2_1 _19663_ (.A(net567),
    .B(_11951_),
    .Y(_02795_));
 sg13g2_buf_1 _19664_ (.A(_02795_),
    .X(_02796_));
 sg13g2_nor2b_1 _19665_ (.A(net451),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02797_));
 sg13g2_a21oi_1 _19666_ (.A1(_11793_),
    .A2(net451),
    .Y(_02798_),
    .B1(_02797_));
 sg13g2_nor2_1 _19667_ (.A(_11818_),
    .B(_02793_),
    .Y(_02799_));
 sg13g2_a21oi_1 _19668_ (.A1(net37),
    .A2(_02798_),
    .Y(_00562_),
    .B1(_02799_));
 sg13g2_nor2b_1 _19669_ (.A(net451),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02800_));
 sg13g2_a21oi_1 _19670_ (.A1(_11775_),
    .A2(net451),
    .Y(_02801_),
    .B1(_02800_));
 sg13g2_nor2_1 _19671_ (.A(_11829_),
    .B(_02793_),
    .Y(_02802_));
 sg13g2_a21oi_1 _19672_ (.A1(net37),
    .A2(_02801_),
    .Y(_00563_),
    .B1(_02802_));
 sg13g2_nor2b_1 _19673_ (.A(net451),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02803_));
 sg13g2_a21oi_1 _19674_ (.A1(_11780_),
    .A2(net451),
    .Y(_02804_),
    .B1(_02803_));
 sg13g2_nor2_1 _19675_ (.A(_11707_),
    .B(_02793_),
    .Y(_02805_));
 sg13g2_a21oi_1 _19676_ (.A1(net37),
    .A2(_02804_),
    .Y(_00564_),
    .B1(_02805_));
 sg13g2_nor2b_1 _19677_ (.A(net451),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02806_));
 sg13g2_a21oi_1 _19678_ (.A1(net960),
    .A2(net451),
    .Y(_02807_),
    .B1(_02806_));
 sg13g2_nor2_1 _19679_ (.A(_11721_),
    .B(_02793_),
    .Y(_02808_));
 sg13g2_a21oi_1 _19680_ (.A1(_02794_),
    .A2(_02807_),
    .Y(_00565_),
    .B1(_02808_));
 sg13g2_nor2_2 _19681_ (.A(net567),
    .B(_11836_),
    .Y(_02809_));
 sg13g2_mux2_1 _19682_ (.A0(\cpu.dcache.r_data[7][28] ),
    .A1(_11792_),
    .S(_02809_),
    .X(_02810_));
 sg13g2_nand2_1 _19683_ (.Y(_02811_),
    .A(net37),
    .B(_02810_));
 sg13g2_o21ai_1 _19684_ (.B1(_02811_),
    .Y(_00566_),
    .A1(_11726_),
    .A2(net37));
 sg13g2_mux2_1 _19685_ (.A0(\cpu.dcache.r_data[7][29] ),
    .A1(net1060),
    .S(_02809_),
    .X(_02812_));
 sg13g2_nand2_1 _19686_ (.Y(_02813_),
    .A(net37),
    .B(_02812_));
 sg13g2_o21ai_1 _19687_ (.B1(_02813_),
    .Y(_00567_),
    .A1(_11740_),
    .A2(net37));
 sg13g2_nor2b_1 _19688_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02814_));
 sg13g2_a21oi_1 _19689_ (.A1(net957),
    .A2(_02740_),
    .Y(_02815_),
    .B1(_02814_));
 sg13g2_nand2_1 _19690_ (.Y(_02816_),
    .A(net844),
    .B(net40));
 sg13g2_o21ai_1 _19691_ (.B1(_02816_),
    .Y(_00568_),
    .A1(net40),
    .A2(_02815_));
 sg13g2_mux2_1 _19692_ (.A0(\cpu.dcache.r_data[7][30] ),
    .A1(_11694_),
    .S(_02809_),
    .X(_02817_));
 sg13g2_nand2_1 _19693_ (.Y(_02818_),
    .A(_02793_),
    .B(_02817_));
 sg13g2_o21ai_1 _19694_ (.B1(_02818_),
    .Y(_00569_),
    .A1(_11749_),
    .A2(net37));
 sg13g2_mux2_1 _19695_ (.A0(\cpu.dcache.r_data[7][31] ),
    .A1(net1063),
    .S(_02809_),
    .X(_02819_));
 sg13g2_nand2_1 _19696_ (.Y(_02820_),
    .A(_02793_),
    .B(_02819_));
 sg13g2_o21ai_1 _19697_ (.B1(_02820_),
    .Y(_00570_),
    .A1(_11758_),
    .A2(_02794_));
 sg13g2_mux2_1 _19698_ (.A0(\cpu.dcache.r_data[7][3] ),
    .A1(net977),
    .S(_02740_),
    .X(_02821_));
 sg13g2_nor2_1 _19699_ (.A(_02737_),
    .B(_02821_),
    .Y(_02822_));
 sg13g2_a21oi_1 _19700_ (.A1(net720),
    .A2(net40),
    .Y(_00571_),
    .B1(_02822_));
 sg13g2_or2_1 _19701_ (.X(_02823_),
    .B(_11853_),
    .A(_09731_));
 sg13g2_buf_1 _19702_ (.A(_02823_),
    .X(_02824_));
 sg13g2_mux2_1 _19703_ (.A0(net1065),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02824_),
    .X(_02825_));
 sg13g2_mux2_1 _19704_ (.A0(_02825_),
    .A1(net971),
    .S(net40),
    .X(_00572_));
 sg13g2_mux2_1 _19705_ (.A0(net1061),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02824_),
    .X(_02826_));
 sg13g2_mux2_1 _19706_ (.A0(_02826_),
    .A1(net969),
    .S(net40),
    .X(_00573_));
 sg13g2_mux2_1 _19707_ (.A0(net1058),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02824_),
    .X(_02827_));
 sg13g2_nor2_1 _19708_ (.A(_02737_),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_a21oi_1 _19709_ (.A1(_12376_),
    .A2(_02738_),
    .Y(_00574_),
    .B1(_02828_));
 sg13g2_mux2_1 _19710_ (.A0(net1057),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02824_),
    .X(_02829_));
 sg13g2_nor2_1 _19711_ (.A(_02737_),
    .B(_02829_),
    .Y(_02830_));
 sg13g2_a21oi_1 _19712_ (.A1(_12379_),
    .A2(_02738_),
    .Y(_00575_),
    .B1(_02830_));
 sg13g2_nor2b_1 _19713_ (.A(_02750_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02831_));
 sg13g2_a21oi_1 _19714_ (.A1(_11793_),
    .A2(_02750_),
    .Y(_02832_),
    .B1(_02831_));
 sg13g2_nor2_1 _19715_ (.A(_11818_),
    .B(_02747_),
    .Y(_02833_));
 sg13g2_a21oi_1 _19716_ (.A1(_02748_),
    .A2(_02832_),
    .Y(_00576_),
    .B1(_02833_));
 sg13g2_nor2b_1 _19717_ (.A(_02750_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02834_));
 sg13g2_a21oi_1 _19718_ (.A1(_11775_),
    .A2(_02750_),
    .Y(_02835_),
    .B1(_02834_));
 sg13g2_nor2_1 _19719_ (.A(_11829_),
    .B(_02747_),
    .Y(_02836_));
 sg13g2_a21oi_1 _19720_ (.A1(_02748_),
    .A2(_02835_),
    .Y(_00577_),
    .B1(_02836_));
 sg13g2_nand2_1 _19721_ (.Y(_02837_),
    .A(_09568_),
    .B(_11660_));
 sg13g2_buf_1 _19722_ (.A(\cpu.d_rstrobe_d ),
    .X(_02838_));
 sg13g2_nor2_1 _19723_ (.A(net986),
    .B(_02838_),
    .Y(_02839_));
 sg13g2_nand4_1 _19724_ (.B(_11676_),
    .C(_08561_),
    .A(_09132_),
    .Y(_02840_),
    .D(_02839_));
 sg13g2_nand2_1 _19725_ (.Y(_02841_),
    .A(_02837_),
    .B(_02840_));
 sg13g2_buf_2 _19726_ (.A(_02841_),
    .X(_02842_));
 sg13g2_xor2_1 _19727_ (.B(_11676_),
    .A(_02838_),
    .X(_02843_));
 sg13g2_nand3_1 _19728_ (.B(_11657_),
    .C(_02843_),
    .A(net976),
    .Y(_02844_));
 sg13g2_and2_1 _19729_ (.A(_02844_),
    .B(_02837_),
    .X(_02845_));
 sg13g2_buf_2 _19730_ (.A(_02845_),
    .X(_02846_));
 sg13g2_nor2_1 _19731_ (.A(net570),
    .B(_02846_),
    .Y(_02847_));
 sg13g2_mux2_1 _19732_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02842_),
    .S(_02847_),
    .X(_00578_));
 sg13g2_nor2_1 _19733_ (.A(net568),
    .B(_02846_),
    .Y(_02848_));
 sg13g2_mux2_1 _19734_ (.A0(\cpu.dcache.r_dirty[1] ),
    .A1(_02842_),
    .S(_02848_),
    .X(_00579_));
 sg13g2_nor2_1 _19735_ (.A(net641),
    .B(_02846_),
    .Y(_02849_));
 sg13g2_mux2_1 _19736_ (.A0(\cpu.dcache.r_dirty[2] ),
    .A1(_02842_),
    .S(_02849_),
    .X(_00580_));
 sg13g2_nor2_1 _19737_ (.A(net640),
    .B(_02846_),
    .Y(_02850_));
 sg13g2_mux2_1 _19738_ (.A0(\cpu.dcache.r_dirty[3] ),
    .A1(_02842_),
    .S(_02850_),
    .X(_00581_));
 sg13g2_nor2_1 _19739_ (.A(_12217_),
    .B(_02846_),
    .Y(_02851_));
 sg13g2_mux2_1 _19740_ (.A0(\cpu.dcache.r_dirty[4] ),
    .A1(_02842_),
    .S(_02851_),
    .X(_00582_));
 sg13g2_nor2_1 _19741_ (.A(net638),
    .B(_02846_),
    .Y(_02852_));
 sg13g2_mux2_1 _19742_ (.A0(\cpu.dcache.r_dirty[5] ),
    .A1(_02842_),
    .S(_02852_),
    .X(_00583_));
 sg13g2_nor2_1 _19743_ (.A(_12431_),
    .B(_02846_),
    .Y(_02853_));
 sg13g2_mux2_1 _19744_ (.A0(\cpu.dcache.r_dirty[6] ),
    .A1(_02842_),
    .S(_02853_),
    .X(_00584_));
 sg13g2_nor2_1 _19745_ (.A(_02735_),
    .B(_02846_),
    .Y(_02854_));
 sg13g2_mux2_1 _19746_ (.A0(\cpu.dcache.r_dirty[7] ),
    .A1(_02842_),
    .S(_02854_),
    .X(_00585_));
 sg13g2_inv_2 _19747_ (.Y(_02855_),
    .A(net1010));
 sg13g2_buf_2 _19748_ (.A(_02855_),
    .X(_02856_));
 sg13g2_buf_1 _19749_ (.A(_02856_),
    .X(_02857_));
 sg13g2_buf_1 _19750_ (.A(net459),
    .X(_02858_));
 sg13g2_buf_1 _19751_ (.A(net459),
    .X(_02859_));
 sg13g2_nand2_1 _19752_ (.Y(_02860_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net388));
 sg13g2_o21ai_1 _19753_ (.B1(_02860_),
    .Y(_00589_),
    .A1(net637),
    .A2(net389));
 sg13g2_mux2_1 _19754_ (.A0(net364),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net389),
    .X(_00590_));
 sg13g2_mux2_1 _19755_ (.A0(net368),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net389),
    .X(_00591_));
 sg13g2_mux2_1 _19756_ (.A0(net403),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net389),
    .X(_00592_));
 sg13g2_mux2_1 _19757_ (.A0(net365),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net389),
    .X(_00593_));
 sg13g2_mux2_1 _19758_ (.A0(net367),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net389),
    .X(_00594_));
 sg13g2_mux2_1 _19759_ (.A0(net401),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(_02858_),
    .X(_00595_));
 sg13g2_mux2_1 _19760_ (.A0(net369),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net389),
    .X(_00596_));
 sg13g2_mux2_1 _19761_ (.A0(net402),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(_02859_),
    .X(_00597_));
 sg13g2_inv_1 _19762_ (.Y(_02861_),
    .A(net404));
 sg13g2_nand2_1 _19763_ (.Y(_02862_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(net459));
 sg13g2_o21ai_1 _19764_ (.B1(_02862_),
    .Y(_00598_),
    .A1(_02861_),
    .A2(net389));
 sg13g2_buf_1 _19765_ (.A(_08950_),
    .X(_02863_));
 sg13g2_buf_1 _19766_ (.A(net715),
    .X(_02864_));
 sg13g2_nand2_1 _19767_ (.Y(_02865_),
    .A(\cpu.dcache.r_tag[0][6] ),
    .B(_11821_));
 sg13g2_o21ai_1 _19768_ (.B1(_02865_),
    .Y(_00599_),
    .A1(net636),
    .A2(_02858_));
 sg13g2_buf_2 _19769_ (.A(_08952_),
    .X(_02866_));
 sg13g2_buf_1 _19770_ (.A(net956),
    .X(_02867_));
 sg13g2_buf_1 _19771_ (.A(net843),
    .X(_02868_));
 sg13g2_mux2_1 _19772_ (.A0(net714),
    .A1(\cpu.dcache.r_tag[0][7] ),
    .S(net388),
    .X(_00600_));
 sg13g2_buf_1 _19773_ (.A(net1085),
    .X(_02869_));
 sg13g2_buf_1 _19774_ (.A(net955),
    .X(_02870_));
 sg13g2_mux2_1 _19775_ (.A0(net842),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(net388),
    .X(_00601_));
 sg13g2_buf_1 _19776_ (.A(_09985_),
    .X(_02871_));
 sg13g2_buf_1 _19777_ (.A(net954),
    .X(_02872_));
 sg13g2_mux2_1 _19778_ (.A0(net841),
    .A1(\cpu.dcache.r_tag[0][9] ),
    .S(net388),
    .X(_00602_));
 sg13g2_buf_1 _19779_ (.A(net1075),
    .X(_02873_));
 sg13g2_buf_1 _19780_ (.A(net953),
    .X(_02874_));
 sg13g2_mux2_1 _19781_ (.A0(net840),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(_02859_),
    .X(_00603_));
 sg13g2_buf_1 _19782_ (.A(_10147_),
    .X(_02875_));
 sg13g2_buf_1 _19783_ (.A(net952),
    .X(_02876_));
 sg13g2_mux2_1 _19784_ (.A0(net839),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net388),
    .X(_00604_));
 sg13g2_mux2_1 _19785_ (.A0(_09235_),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net388),
    .X(_00605_));
 sg13g2_mux2_1 _19786_ (.A0(net370),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net388),
    .X(_00606_));
 sg13g2_mux2_1 _19787_ (.A0(net366),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net388),
    .X(_00607_));
 sg13g2_buf_2 _19788_ (.A(net725),
    .X(_02877_));
 sg13g2_buf_1 _19789_ (.A(net635),
    .X(_02878_));
 sg13g2_buf_1 _19790_ (.A(_02878_),
    .X(_02879_));
 sg13g2_buf_1 _19791_ (.A(net519),
    .X(_02880_));
 sg13g2_mux2_1 _19792_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net512),
    .S(net450),
    .X(_00608_));
 sg13g2_mux2_1 _19793_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net364),
    .S(net450),
    .X(_00609_));
 sg13g2_mux2_1 _19794_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net368),
    .S(net450),
    .X(_00610_));
 sg13g2_mux2_1 _19795_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net403),
    .S(net450),
    .X(_00611_));
 sg13g2_mux2_1 _19796_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net365),
    .S(net450),
    .X(_00612_));
 sg13g2_mux2_1 _19797_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net367),
    .S(net450),
    .X(_00613_));
 sg13g2_mux2_1 _19798_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net401),
    .S(_02880_),
    .X(_00614_));
 sg13g2_mux2_1 _19799_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net369),
    .S(net450),
    .X(_00615_));
 sg13g2_mux2_1 _19800_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net402),
    .S(_02880_),
    .X(_00616_));
 sg13g2_mux2_1 _19801_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net404),
    .S(net450),
    .X(_00617_));
 sg13g2_buf_1 _19802_ (.A(net1022),
    .X(_02881_));
 sg13g2_buf_1 _19803_ (.A(net838),
    .X(_02882_));
 sg13g2_buf_1 _19804_ (.A(net519),
    .X(_02883_));
 sg13g2_mux2_1 _19805_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net713),
    .S(net449),
    .X(_00618_));
 sg13g2_buf_1 _19806_ (.A(net843),
    .X(_02884_));
 sg13g2_mux2_1 _19807_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net712),
    .S(net449),
    .X(_00619_));
 sg13g2_buf_1 _19808_ (.A(net955),
    .X(_02885_));
 sg13g2_mux2_1 _19809_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net837),
    .S(net449),
    .X(_00620_));
 sg13g2_buf_1 _19810_ (.A(net954),
    .X(_02886_));
 sg13g2_mux2_1 _19811_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net836),
    .S(_02883_),
    .X(_00621_));
 sg13g2_buf_1 _19812_ (.A(net953),
    .X(_02887_));
 sg13g2_mux2_1 _19813_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net835),
    .S(net449),
    .X(_00622_));
 sg13g2_buf_1 _19814_ (.A(net952),
    .X(_02888_));
 sg13g2_mux2_1 _19815_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net834),
    .S(net449),
    .X(_00623_));
 sg13g2_mux2_1 _19816_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net338),
    .S(net449),
    .X(_00624_));
 sg13g2_mux2_1 _19817_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net370),
    .S(net449),
    .X(_00625_));
 sg13g2_mux2_1 _19818_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net366),
    .S(net449),
    .X(_00626_));
 sg13g2_buf_1 _19819_ (.A(_12065_),
    .X(_02889_));
 sg13g2_mux2_1 _19820_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net512),
    .S(net448),
    .X(_00627_));
 sg13g2_mux2_1 _19821_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net364),
    .S(net448),
    .X(_00628_));
 sg13g2_mux2_1 _19822_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net368),
    .S(net448),
    .X(_00629_));
 sg13g2_mux2_1 _19823_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net403),
    .S(net448),
    .X(_00630_));
 sg13g2_mux2_1 _19824_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net365),
    .S(net448),
    .X(_00631_));
 sg13g2_mux2_1 _19825_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net367),
    .S(_02889_),
    .X(_00632_));
 sg13g2_mux2_1 _19826_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net401),
    .S(net448),
    .X(_00633_));
 sg13g2_mux2_1 _19827_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net369),
    .S(net448),
    .X(_00634_));
 sg13g2_mux2_1 _19828_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net402),
    .S(_02889_),
    .X(_00635_));
 sg13g2_buf_1 _19829_ (.A(_12064_),
    .X(_02890_));
 sg13g2_mux2_1 _19830_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net404),
    .S(net511),
    .X(_00636_));
 sg13g2_mux2_1 _19831_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net713),
    .S(net511),
    .X(_00637_));
 sg13g2_mux2_1 _19832_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net712),
    .S(net511),
    .X(_00638_));
 sg13g2_mux2_1 _19833_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net837),
    .S(_02890_),
    .X(_00639_));
 sg13g2_nand2_1 _19834_ (.Y(_02891_),
    .A(net954),
    .B(net511));
 sg13g2_o21ai_1 _19835_ (.B1(_02891_),
    .Y(_00640_),
    .A1(_09438_),
    .A2(net448));
 sg13g2_mux2_1 _19836_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net835),
    .S(net511),
    .X(_00641_));
 sg13g2_mux2_1 _19837_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net834),
    .S(_02890_),
    .X(_00642_));
 sg13g2_mux2_1 _19838_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net338),
    .S(net511),
    .X(_00643_));
 sg13g2_mux2_1 _19839_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net370),
    .S(net511),
    .X(_00644_));
 sg13g2_mux2_1 _19840_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net366),
    .S(net511),
    .X(_00645_));
 sg13g2_buf_1 _19841_ (.A(net516),
    .X(_02892_));
 sg13g2_mux2_1 _19842_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net512),
    .S(net447),
    .X(_00646_));
 sg13g2_mux2_1 _19843_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net364),
    .S(_02892_),
    .X(_00647_));
 sg13g2_mux2_1 _19844_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net368),
    .S(net447),
    .X(_00648_));
 sg13g2_mux2_1 _19845_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net403),
    .S(net447),
    .X(_00649_));
 sg13g2_mux2_1 _19846_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net365),
    .S(net447),
    .X(_00650_));
 sg13g2_mux2_1 _19847_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net367),
    .S(net447),
    .X(_00651_));
 sg13g2_mux2_1 _19848_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net401),
    .S(_02892_),
    .X(_00652_));
 sg13g2_mux2_1 _19849_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net369),
    .S(net447),
    .X(_00653_));
 sg13g2_mux2_1 _19850_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net402),
    .S(net447),
    .X(_00654_));
 sg13g2_mux2_1 _19851_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(net404),
    .S(net447),
    .X(_00655_));
 sg13g2_buf_1 _19852_ (.A(net516),
    .X(_02893_));
 sg13g2_mux2_1 _19853_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net713),
    .S(net446),
    .X(_00656_));
 sg13g2_mux2_1 _19854_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net712),
    .S(net446),
    .X(_00657_));
 sg13g2_mux2_1 _19855_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net837),
    .S(net446),
    .X(_00658_));
 sg13g2_mux2_1 _19856_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net836),
    .S(net446),
    .X(_00659_));
 sg13g2_mux2_1 _19857_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net835),
    .S(_02893_),
    .X(_00660_));
 sg13g2_mux2_1 _19858_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net834),
    .S(net446),
    .X(_00661_));
 sg13g2_mux2_1 _19859_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net338),
    .S(net446),
    .X(_00662_));
 sg13g2_mux2_1 _19860_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net370),
    .S(net446),
    .X(_00663_));
 sg13g2_mux2_1 _19861_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net366),
    .S(net446),
    .X(_00664_));
 sg13g2_buf_1 _19862_ (.A(net331),
    .X(_02894_));
 sg13g2_nand2_1 _19863_ (.Y(_02895_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net331));
 sg13g2_o21ai_1 _19864_ (.B1(_02895_),
    .Y(_00665_),
    .A1(net637),
    .A2(net288));
 sg13g2_mux2_1 _19865_ (.A0(net364),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net288),
    .X(_00666_));
 sg13g2_mux2_1 _19866_ (.A0(net368),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net288),
    .X(_00667_));
 sg13g2_mux2_1 _19867_ (.A0(net403),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(net288),
    .X(_00668_));
 sg13g2_mux2_1 _19868_ (.A0(net365),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net288),
    .X(_00669_));
 sg13g2_mux2_1 _19869_ (.A0(net367),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net288),
    .X(_00670_));
 sg13g2_mux2_1 _19870_ (.A0(net401),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(net288),
    .X(_00671_));
 sg13g2_buf_1 _19871_ (.A(net331),
    .X(_02896_));
 sg13g2_mux2_1 _19872_ (.A0(net369),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net287),
    .X(_00672_));
 sg13g2_mux2_1 _19873_ (.A0(_09371_),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(_02896_),
    .X(_00673_));
 sg13g2_nand2_1 _19874_ (.Y(_02897_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(net331));
 sg13g2_o21ai_1 _19875_ (.B1(_02897_),
    .Y(_00674_),
    .A1(_02861_),
    .A2(net288));
 sg13g2_nand2_1 _19876_ (.Y(_02898_),
    .A(\cpu.dcache.r_tag[4][6] ),
    .B(_12278_));
 sg13g2_o21ai_1 _19877_ (.B1(_02898_),
    .Y(_00675_),
    .A1(net636),
    .A2(_02894_));
 sg13g2_mux2_1 _19878_ (.A0(net714),
    .A1(\cpu.dcache.r_tag[4][7] ),
    .S(net287),
    .X(_00676_));
 sg13g2_mux2_1 _19879_ (.A0(net842),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(net287),
    .X(_00677_));
 sg13g2_mux2_1 _19880_ (.A0(net841),
    .A1(\cpu.dcache.r_tag[4][9] ),
    .S(net287),
    .X(_00678_));
 sg13g2_mux2_1 _19881_ (.A0(net840),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(_02896_),
    .X(_00679_));
 sg13g2_mux2_1 _19882_ (.A0(net839),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net287),
    .X(_00680_));
 sg13g2_mux2_1 _19883_ (.A0(net338),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net287),
    .X(_00681_));
 sg13g2_mux2_1 _19884_ (.A0(net370),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net287),
    .X(_00682_));
 sg13g2_mux2_1 _19885_ (.A0(net366),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net287),
    .X(_00683_));
 sg13g2_buf_1 _19886_ (.A(_12386_),
    .X(_02899_));
 sg13g2_mux2_1 _19887_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net512),
    .S(net445),
    .X(_00684_));
 sg13g2_mux2_1 _19888_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net364),
    .S(_02899_),
    .X(_00685_));
 sg13g2_mux2_1 _19889_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net368),
    .S(net445),
    .X(_00686_));
 sg13g2_mux2_1 _19890_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(net403),
    .S(net445),
    .X(_00687_));
 sg13g2_mux2_1 _19891_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net365),
    .S(net445),
    .X(_00688_));
 sg13g2_mux2_1 _19892_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net367),
    .S(_02899_),
    .X(_00689_));
 sg13g2_mux2_1 _19893_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net401),
    .S(net445),
    .X(_00690_));
 sg13g2_mux2_1 _19894_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net369),
    .S(net445),
    .X(_00691_));
 sg13g2_mux2_1 _19895_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net402),
    .S(net445),
    .X(_00692_));
 sg13g2_buf_1 _19896_ (.A(_12385_),
    .X(_02900_));
 sg13g2_mux2_1 _19897_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net404),
    .S(net510),
    .X(_00693_));
 sg13g2_mux2_1 _19898_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(net713),
    .S(net510),
    .X(_00694_));
 sg13g2_mux2_1 _19899_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(net712),
    .S(net510),
    .X(_00695_));
 sg13g2_mux2_1 _19900_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net837),
    .S(net510),
    .X(_00696_));
 sg13g2_nand2_1 _19901_ (.Y(_02901_),
    .A(net954),
    .B(net510));
 sg13g2_o21ai_1 _19902_ (.B1(_02901_),
    .Y(_00697_),
    .A1(_09442_),
    .A2(net445));
 sg13g2_mux2_1 _19903_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(net835),
    .S(_02900_),
    .X(_00698_));
 sg13g2_mux2_1 _19904_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net834),
    .S(_02900_),
    .X(_00699_));
 sg13g2_mux2_1 _19905_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net338),
    .S(net510),
    .X(_00700_));
 sg13g2_mux2_1 _19906_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net370),
    .S(net510),
    .X(_00701_));
 sg13g2_mux2_1 _19907_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(_09427_),
    .S(net510),
    .X(_00702_));
 sg13g2_buf_1 _19908_ (.A(_02690_),
    .X(_02902_));
 sg13g2_mux2_1 _19909_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net512),
    .S(net387),
    .X(_00703_));
 sg13g2_mux2_1 _19910_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net364),
    .S(net387),
    .X(_00704_));
 sg13g2_mux2_1 _19911_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(net368),
    .S(net387),
    .X(_00705_));
 sg13g2_mux2_1 _19912_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(net403),
    .S(net387),
    .X(_00706_));
 sg13g2_mux2_1 _19913_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net365),
    .S(net387),
    .X(_00707_));
 sg13g2_mux2_1 _19914_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(net367),
    .S(net387),
    .X(_00708_));
 sg13g2_mux2_1 _19915_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(_09395_),
    .S(net387),
    .X(_00709_));
 sg13g2_mux2_1 _19916_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net369),
    .S(_02902_),
    .X(_00710_));
 sg13g2_buf_1 _19917_ (.A(_02689_),
    .X(_02903_));
 sg13g2_mux2_1 _19918_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(net402),
    .S(_02903_),
    .X(_00711_));
 sg13g2_mux2_1 _19919_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(net404),
    .S(net444),
    .X(_00712_));
 sg13g2_mux2_1 _19920_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net713),
    .S(net444),
    .X(_00713_));
 sg13g2_mux2_1 _19921_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net712),
    .S(net444),
    .X(_00714_));
 sg13g2_mux2_1 _19922_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net837),
    .S(net444),
    .X(_00715_));
 sg13g2_nand2_1 _19923_ (.Y(_02904_),
    .A(net954),
    .B(net444));
 sg13g2_o21ai_1 _19924_ (.B1(_02904_),
    .Y(_00716_),
    .A1(_09431_),
    .A2(_02902_));
 sg13g2_inv_1 _19925_ (.Y(_02905_),
    .A(\cpu.dcache.r_tag[6][10] ));
 sg13g2_nand2_1 _19926_ (.Y(_02906_),
    .A(net953),
    .B(_02690_));
 sg13g2_o21ai_1 _19927_ (.B1(_02906_),
    .Y(_00717_),
    .A1(_02905_),
    .A2(net387));
 sg13g2_mux2_1 _19928_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net834),
    .S(_02903_),
    .X(_00718_));
 sg13g2_mux2_1 _19929_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net338),
    .S(net444),
    .X(_00719_));
 sg13g2_mux2_1 _19930_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(net370),
    .S(net444),
    .X(_00720_));
 sg13g2_mux2_1 _19931_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net366),
    .S(net444),
    .X(_00721_));
 sg13g2_buf_1 _19932_ (.A(_02796_),
    .X(_02907_));
 sg13g2_mux2_1 _19933_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net512),
    .S(net386),
    .X(_00722_));
 sg13g2_mux2_1 _19934_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net364),
    .S(net386),
    .X(_00723_));
 sg13g2_mux2_1 _19935_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net368),
    .S(net386),
    .X(_00724_));
 sg13g2_mux2_1 _19936_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net403),
    .S(net386),
    .X(_00725_));
 sg13g2_mux2_1 _19937_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(net365),
    .S(net386),
    .X(_00726_));
 sg13g2_mux2_1 _19938_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net367),
    .S(_02907_),
    .X(_00727_));
 sg13g2_mux2_1 _19939_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net401),
    .S(_02907_),
    .X(_00728_));
 sg13g2_mux2_1 _19940_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(_09254_),
    .S(net386),
    .X(_00729_));
 sg13g2_mux2_1 _19941_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net402),
    .S(net386),
    .X(_00730_));
 sg13g2_mux2_1 _19942_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(net404),
    .S(net386),
    .X(_00731_));
 sg13g2_buf_1 _19943_ (.A(_02796_),
    .X(_02908_));
 sg13g2_mux2_1 _19944_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net713),
    .S(net385),
    .X(_00732_));
 sg13g2_buf_1 _19945_ (.A(net843),
    .X(_02909_));
 sg13g2_mux2_1 _19946_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net711),
    .S(net385),
    .X(_00733_));
 sg13g2_buf_1 _19947_ (.A(net955),
    .X(_02910_));
 sg13g2_mux2_1 _19948_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net833),
    .S(net385),
    .X(_00734_));
 sg13g2_mux2_1 _19949_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net836),
    .S(net385),
    .X(_00735_));
 sg13g2_mux2_1 _19950_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net835),
    .S(_02908_),
    .X(_00736_));
 sg13g2_buf_1 _19951_ (.A(net952),
    .X(_02911_));
 sg13g2_mux2_1 _19952_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(_02911_),
    .S(_02908_),
    .X(_00737_));
 sg13g2_mux2_1 _19953_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net338),
    .S(net385),
    .X(_00738_));
 sg13g2_mux2_1 _19954_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net370),
    .S(net385),
    .X(_00739_));
 sg13g2_mux2_1 _19955_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(_09427_),
    .S(net385),
    .X(_00740_));
 sg13g2_buf_1 _19956_ (.A(_08622_),
    .X(_02912_));
 sg13g2_buf_1 _19957_ (.A(_08833_),
    .X(_02913_));
 sg13g2_buf_1 _19958_ (.A(_08663_),
    .X(_02914_));
 sg13g2_nor2_2 _19959_ (.A(net177),
    .B(net176),
    .Y(_02915_));
 sg13g2_nand2_1 _19960_ (.Y(_02916_),
    .A(_08832_),
    .B(_02915_));
 sg13g2_buf_1 _19961_ (.A(_08662_),
    .X(_02917_));
 sg13g2_nand2_1 _19962_ (.Y(_02918_),
    .A(_08642_),
    .B(net198));
 sg13g2_buf_2 _19963_ (.A(_02918_),
    .X(_02919_));
 sg13g2_buf_1 _19964_ (.A(_08642_),
    .X(_02920_));
 sg13g2_nor2_1 _19965_ (.A(_08681_),
    .B(net339),
    .Y(_02921_));
 sg13g2_buf_1 _19966_ (.A(_02921_),
    .X(_02922_));
 sg13g2_a21o_1 _19967_ (.A2(_08672_),
    .A1(net1025),
    .B1(_08679_),
    .X(_02923_));
 sg13g2_buf_1 _19968_ (.A(_02923_),
    .X(_02924_));
 sg13g2_buf_1 _19969_ (.A(_02924_),
    .X(_02925_));
 sg13g2_nor2_1 _19970_ (.A(net212),
    .B(net286),
    .Y(_02926_));
 sg13g2_buf_1 _19971_ (.A(_02926_),
    .X(_02927_));
 sg13g2_a21oi_1 _19972_ (.A1(net198),
    .A2(_02922_),
    .Y(_02928_),
    .B1(net150));
 sg13g2_or2_1 _19973_ (.X(_02929_),
    .B(_02928_),
    .A(net197));
 sg13g2_buf_1 _19974_ (.A(_02929_),
    .X(_02930_));
 sg13g2_nand2_1 _19975_ (.Y(_02931_),
    .A(_02919_),
    .B(_02930_));
 sg13g2_nand3b_1 _19976_ (.B(_02916_),
    .C(_02931_),
    .Y(_02932_),
    .A_N(_02912_));
 sg13g2_o21ai_1 _19977_ (.B1(_02932_),
    .Y(_00749_),
    .A1(_11565_),
    .A2(_08852_));
 sg13g2_buf_1 _19978_ (.A(_08681_),
    .X(_02933_));
 sg13g2_buf_1 _19979_ (.A(net198),
    .X(_02934_));
 sg13g2_nand2_1 _19980_ (.Y(_02935_),
    .A(net176),
    .B(net214));
 sg13g2_buf_1 _19981_ (.A(net197),
    .X(_02936_));
 sg13g2_a22oi_1 _19982_ (.Y(_02937_),
    .B1(_02935_),
    .B2(net174),
    .A2(net339),
    .A1(net175));
 sg13g2_buf_1 _19983_ (.A(net252),
    .X(_02938_));
 sg13g2_nor2_1 _19984_ (.A(net176),
    .B(net196),
    .Y(_02939_));
 sg13g2_nand2_1 _19985_ (.Y(_02940_),
    .A(net177),
    .B(net212));
 sg13g2_nor2_1 _19986_ (.A(_02924_),
    .B(net339),
    .Y(_02941_));
 sg13g2_buf_1 _19987_ (.A(_02941_),
    .X(_02942_));
 sg13g2_a22oi_1 _19988_ (.Y(_02943_),
    .B1(_02940_),
    .B2(_02942_),
    .A2(_02939_),
    .A1(net177));
 sg13g2_o21ai_1 _19989_ (.B1(_02943_),
    .Y(_02944_),
    .A1(net285),
    .A2(_02937_));
 sg13g2_nand2_1 _19990_ (.Y(_02945_),
    .A(net111),
    .B(_02944_));
 sg13g2_o21ai_1 _19991_ (.B1(_02945_),
    .Y(_00750_),
    .A1(_11553_),
    .A2(net112));
 sg13g2_nand2_1 _19992_ (.Y(_02946_),
    .A(_08699_),
    .B(_08681_));
 sg13g2_buf_1 _19993_ (.A(_02946_),
    .X(_02947_));
 sg13g2_nor3_1 _19994_ (.A(net108),
    .B(net126),
    .C(_02947_),
    .Y(_02948_));
 sg13g2_a21o_1 _19995_ (.A2(net89),
    .A1(\cpu.cond[1] ),
    .B1(_02948_),
    .X(_00751_));
 sg13g2_a21oi_1 _19996_ (.A1(net285),
    .A2(_02940_),
    .Y(_02949_),
    .B1(net176));
 sg13g2_buf_1 _19997_ (.A(_08622_),
    .X(_02950_));
 sg13g2_mux2_1 _19998_ (.A0(_02949_),
    .A1(\cpu.cond[2] ),
    .S(net103),
    .X(_00752_));
 sg13g2_nor3_1 _19999_ (.A(net108),
    .B(_08837_),
    .C(_08858_),
    .Y(_02951_));
 sg13g2_a21o_1 _20000_ (.A2(net89),
    .A1(_09113_),
    .B1(_02951_),
    .X(_00753_));
 sg13g2_nor2_1 _20001_ (.A(_08642_),
    .B(_02917_),
    .Y(_02952_));
 sg13g2_nor3_2 _20002_ (.A(_08699_),
    .B(_08681_),
    .C(_08828_),
    .Y(_02953_));
 sg13g2_nand2_1 _20003_ (.Y(_02954_),
    .A(_02952_),
    .B(_02953_));
 sg13g2_buf_1 _20004_ (.A(_02954_),
    .X(_02955_));
 sg13g2_nor2_1 _20005_ (.A(_00175_),
    .B(net539),
    .Y(_02956_));
 sg13g2_mux2_1 _20006_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_08163_),
    .X(_02957_));
 sg13g2_a22oi_1 _20007_ (.Y(_02958_),
    .B1(_02957_),
    .B2(net771),
    .A2(_08650_),
    .A1(\cpu.icache.r_data[5][24] ));
 sg13g2_nor2_1 _20008_ (.A(_08162_),
    .B(_02958_),
    .Y(_02959_));
 sg13g2_and2_1 _20009_ (.A(net775),
    .B(\cpu.icache.r_data[3][24] ),
    .X(_02960_));
 sg13g2_a21oi_1 _20010_ (.A1(net777),
    .A2(\cpu.icache.r_data[7][24] ),
    .Y(_02961_),
    .B1(_02960_));
 sg13g2_a22oi_1 _20011_ (.Y(_02962_),
    .B1(_08208_),
    .B2(\cpu.icache.r_data[1][24] ),
    .A2(net472),
    .A1(\cpu.icache.r_data[2][24] ));
 sg13g2_o21ai_1 _20012_ (.B1(_02962_),
    .Y(_02963_),
    .A1(net765),
    .A2(_02961_));
 sg13g2_nor3_1 _20013_ (.A(_02956_),
    .B(_02959_),
    .C(_02963_),
    .Y(_02964_));
 sg13g2_nand2_1 _20014_ (.Y(_02965_),
    .A(_00174_),
    .B(net541));
 sg13g2_a22oi_1 _20015_ (.Y(_02966_),
    .B1(net700),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(net546),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_a22oi_1 _20016_ (.Y(_02967_),
    .B1(net598),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net702),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_mux2_1 _20017_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_08110_),
    .X(_02968_));
 sg13g2_a22oi_1 _20018_ (.Y(_02969_),
    .B1(_02968_),
    .B2(_08385_),
    .A2(_08235_),
    .A1(\cpu.icache.r_data[7][8] ));
 sg13g2_or2_1 _20019_ (.X(_02970_),
    .B(_02969_),
    .A(net775));
 sg13g2_nand4_1 _20020_ (.B(_02966_),
    .C(_02967_),
    .A(net476),
    .Y(_02971_),
    .D(_02970_));
 sg13g2_a21oi_1 _20021_ (.A1(_02965_),
    .A2(_02971_),
    .Y(_02972_),
    .B1(net1025));
 sg13g2_a21oi_1 _20022_ (.A1(net1025),
    .A2(_02964_),
    .Y(_02973_),
    .B1(_02972_));
 sg13g2_buf_2 _20023_ (.A(_02973_),
    .X(_02974_));
 sg13g2_inv_1 _20024_ (.Y(_02975_),
    .A(_00176_));
 sg13g2_mux4_1 _20025_ (.S0(_08109_),
    .A0(\cpu.icache.r_data[4][9] ),
    .A1(\cpu.icache.r_data[5][9] ),
    .A2(\cpu.icache.r_data[6][9] ),
    .A3(\cpu.icache.r_data[7][9] ),
    .S1(_08112_),
    .X(_02976_));
 sg13g2_nand2_1 _20026_ (.Y(_02977_),
    .A(net777),
    .B(_02976_));
 sg13g2_nand2_1 _20027_ (.Y(_02978_),
    .A(\cpu.icache.r_data[2][9] ),
    .B(net475));
 sg13g2_a22oi_1 _20028_ (.Y(_02979_),
    .B1(net545),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(net596),
    .A1(\cpu.icache.r_data[1][9] ));
 sg13g2_nand4_1 _20029_ (.B(_02977_),
    .C(_02978_),
    .A(net410),
    .Y(_02980_),
    .D(_02979_));
 sg13g2_o21ai_1 _20030_ (.B1(_02980_),
    .Y(_02981_),
    .A1(_02975_),
    .A2(_08101_));
 sg13g2_nor2_1 _20031_ (.A(_00177_),
    .B(net410),
    .Y(_02982_));
 sg13g2_mux2_1 _20032_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(net776),
    .X(_02983_));
 sg13g2_a22oi_1 _20033_ (.Y(_02984_),
    .B1(_02983_),
    .B2(_08258_),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][25] ));
 sg13g2_nand2_1 _20034_ (.Y(_02985_),
    .A(net775),
    .B(\cpu.icache.r_data[3][25] ));
 sg13g2_nand2_1 _20035_ (.Y(_02986_),
    .A(net906),
    .B(\cpu.icache.r_data[7][25] ));
 sg13g2_a21oi_1 _20036_ (.A1(_02985_),
    .A2(_02986_),
    .Y(_02987_),
    .B1(net765));
 sg13g2_a221oi_1 _20037_ (.B2(\cpu.icache.r_data[1][25] ),
    .C1(_02987_),
    .B1(net599),
    .A1(\cpu.icache.r_data[2][25] ),
    .Y(_02988_),
    .A2(net472));
 sg13g2_o21ai_1 _20038_ (.B1(_02988_),
    .Y(_02989_),
    .A1(net701),
    .A2(_02984_));
 sg13g2_nor3_1 _20039_ (.A(net764),
    .B(_02982_),
    .C(_02989_),
    .Y(_02990_));
 sg13g2_a21oi_1 _20040_ (.A1(net764),
    .A2(_02981_),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_inv_1 _20041_ (.Y(_02992_),
    .A(_00172_));
 sg13g2_mux4_1 _20042_ (.S0(net905),
    .A0(\cpu.icache.r_data[4][7] ),
    .A1(\cpu.icache.r_data[5][7] ),
    .A2(\cpu.icache.r_data[6][7] ),
    .A3(\cpu.icache.r_data[7][7] ),
    .S1(_08113_),
    .X(_02993_));
 sg13g2_nand2_1 _20043_ (.Y(_02994_),
    .A(net777),
    .B(_02993_));
 sg13g2_nand2_1 _20044_ (.Y(_02995_),
    .A(\cpu.icache.r_data[2][7] ),
    .B(_08121_));
 sg13g2_a22oi_1 _20045_ (.Y(_02996_),
    .B1(net473),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(net599),
    .A1(\cpu.icache.r_data[1][7] ));
 sg13g2_nand4_1 _20046_ (.B(_02994_),
    .C(_02995_),
    .A(net410),
    .Y(_02997_),
    .D(_02996_));
 sg13g2_o21ai_1 _20047_ (.B1(_02997_),
    .Y(_02998_),
    .A1(_02992_),
    .A2(net411));
 sg13g2_nor2_1 _20048_ (.A(_00173_),
    .B(_08104_),
    .Y(_02999_));
 sg13g2_mux2_1 _20049_ (.A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_08113_),
    .X(_03000_));
 sg13g2_a22oi_1 _20050_ (.Y(_03001_),
    .B1(_03000_),
    .B2(_08258_),
    .A2(net694),
    .A1(\cpu.icache.r_data[5][23] ));
 sg13g2_nand2_1 _20051_ (.Y(_03002_),
    .A(_08306_),
    .B(\cpu.icache.r_data[3][23] ));
 sg13g2_nand2_1 _20052_ (.Y(_03003_),
    .A(_08107_),
    .B(\cpu.icache.r_data[7][23] ));
 sg13g2_a21oi_1 _20053_ (.A1(_03002_),
    .A2(_03003_),
    .Y(_03004_),
    .B1(_08654_));
 sg13g2_a221oi_1 _20054_ (.B2(\cpu.icache.r_data[1][23] ),
    .C1(_03004_),
    .B1(net599),
    .A1(\cpu.icache.r_data[2][23] ),
    .Y(_03005_),
    .A2(_08121_));
 sg13g2_o21ai_1 _20055_ (.B1(_03005_),
    .Y(_03006_),
    .A1(_08162_),
    .A2(_03001_));
 sg13g2_nor3_1 _20056_ (.A(_08821_),
    .B(_02999_),
    .C(_03006_),
    .Y(_03007_));
 sg13g2_a21oi_2 _20057_ (.B1(_03007_),
    .Y(_03008_),
    .A2(_02998_),
    .A1(_08821_));
 sg13g2_nor3_1 _20058_ (.A(_02974_),
    .B(_02991_),
    .C(_03008_),
    .Y(_03009_));
 sg13g2_nand2_1 _20059_ (.Y(_03010_),
    .A(_09633_),
    .B(_03009_));
 sg13g2_or3_1 _20060_ (.A(net247),
    .B(_08858_),
    .C(_03010_),
    .X(_03011_));
 sg13g2_nor2_1 _20061_ (.A(_02955_),
    .B(_03011_),
    .Y(_03012_));
 sg13g2_mux2_1 _20062_ (.A0(_03012_),
    .A1(\cpu.dec.do_flush_all ),
    .S(net103),
    .X(_00754_));
 sg13g2_nand2_1 _20063_ (.Y(_03013_),
    .A(net252),
    .B(_02922_));
 sg13g2_nor3_1 _20064_ (.A(net108),
    .B(_09645_),
    .C(_03013_),
    .Y(_03014_));
 sg13g2_a21o_1 _20065_ (.A2(net89),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03014_),
    .X(_00755_));
 sg13g2_nand2_1 _20066_ (.Y(_03015_),
    .A(net177),
    .B(_08662_));
 sg13g2_nor2_1 _20067_ (.A(_03015_),
    .B(net150),
    .Y(_03016_));
 sg13g2_a21o_1 _20068_ (.A2(_03016_),
    .A1(net339),
    .B1(_08836_),
    .X(_03017_));
 sg13g2_nor2_1 _20069_ (.A(net285),
    .B(net245),
    .Y(_03018_));
 sg13g2_a21oi_1 _20070_ (.A1(net211),
    .A2(_02942_),
    .Y(_03019_),
    .B1(_03018_));
 sg13g2_nand3_1 _20071_ (.B(net248),
    .C(_02942_),
    .A(net175),
    .Y(_03020_));
 sg13g2_o21ai_1 _20072_ (.B1(_03020_),
    .Y(_03021_),
    .A1(net175),
    .A2(_03019_));
 sg13g2_nor2_1 _20073_ (.A(net246),
    .B(_02955_),
    .Y(_03022_));
 sg13g2_a221oi_1 _20074_ (.B2(net174),
    .C1(_03022_),
    .B1(_03021_),
    .A1(net248),
    .Y(_03023_),
    .A2(_03017_));
 sg13g2_nand2_1 _20075_ (.Y(_03024_),
    .A(_11021_),
    .B(net109));
 sg13g2_o21ai_1 _20076_ (.B1(_03024_),
    .Y(_00756_),
    .A1(net90),
    .A2(_03023_));
 sg13g2_buf_1 _20077_ (.A(_08828_),
    .X(_03025_));
 sg13g2_nor2_2 _20078_ (.A(net252),
    .B(_03025_),
    .Y(_03026_));
 sg13g2_a21oi_1 _20079_ (.A1(_08881_),
    .A2(_03026_),
    .Y(_03027_),
    .B1(_03015_));
 sg13g2_buf_2 _20080_ (.A(_03027_),
    .X(_03028_));
 sg13g2_buf_1 _20081_ (.A(_02922_),
    .X(_03029_));
 sg13g2_nand2_1 _20082_ (.Y(_03030_),
    .A(net195),
    .B(_02974_));
 sg13g2_a21oi_1 _20083_ (.A1(_09647_),
    .A2(net150),
    .Y(_03031_),
    .B1(_03026_));
 sg13g2_nor2_1 _20084_ (.A(_08698_),
    .B(_02924_),
    .Y(_03032_));
 sg13g2_buf_2 _20085_ (.A(_03032_),
    .X(_03033_));
 sg13g2_inv_1 _20086_ (.Y(_03034_),
    .A(_03033_));
 sg13g2_nor2_2 _20087_ (.A(net339),
    .B(_03034_),
    .Y(_03035_));
 sg13g2_nand2_1 _20088_ (.Y(_03036_),
    .A(net211),
    .B(_03035_));
 sg13g2_nand3_1 _20089_ (.B(_03031_),
    .C(_03036_),
    .A(_03030_),
    .Y(_03037_));
 sg13g2_nand2_1 _20090_ (.Y(_03038_),
    .A(_03028_),
    .B(_03037_));
 sg13g2_nand2_1 _20091_ (.Y(_03039_),
    .A(net212),
    .B(_02922_));
 sg13g2_buf_2 _20092_ (.A(_03039_),
    .X(_03040_));
 sg13g2_nor2_1 _20093_ (.A(_08662_),
    .B(_03040_),
    .Y(_03041_));
 sg13g2_a21o_1 _20094_ (.A2(net155),
    .A1(net198),
    .B1(_03041_),
    .X(_03042_));
 sg13g2_nand3_1 _20095_ (.B(net247),
    .C(_03042_),
    .A(net197),
    .Y(_03043_));
 sg13g2_buf_1 _20096_ (.A(_03043_),
    .X(_03044_));
 sg13g2_nor2_1 _20097_ (.A(_08835_),
    .B(_02953_),
    .Y(_03045_));
 sg13g2_buf_2 _20098_ (.A(_03045_),
    .X(_03046_));
 sg13g2_nand2_1 _20099_ (.Y(_03047_),
    .A(_09647_),
    .B(net150));
 sg13g2_buf_2 _20100_ (.A(_03047_),
    .X(_03048_));
 sg13g2_nand2_1 _20101_ (.Y(_03049_),
    .A(_03048_),
    .B(_03036_));
 sg13g2_nand2_1 _20102_ (.Y(_03050_),
    .A(_03046_),
    .B(_03049_));
 sg13g2_nand3_1 _20103_ (.B(_03044_),
    .C(_03050_),
    .A(_03038_),
    .Y(_03051_));
 sg13g2_mux2_1 _20104_ (.A0(_03051_),
    .A1(\cpu.dec.imm[10] ),
    .S(_02950_),
    .X(_00757_));
 sg13g2_nand2_1 _20105_ (.Y(_03052_),
    .A(_08828_),
    .B(_03033_));
 sg13g2_buf_2 _20106_ (.A(_03052_),
    .X(_03053_));
 sg13g2_o21ai_1 _20107_ (.B1(_03048_),
    .Y(_03054_),
    .A1(net245),
    .A2(_03053_));
 sg13g2_nand2_1 _20108_ (.Y(_03055_),
    .A(_03046_),
    .B(_03054_));
 sg13g2_o21ai_1 _20109_ (.B1(net284),
    .Y(_03056_),
    .A1(net250),
    .A2(_03033_));
 sg13g2_o21ai_1 _20110_ (.B1(net252),
    .Y(_03057_),
    .A1(net249),
    .A2(net250));
 sg13g2_and2_1 _20111_ (.A(_03056_),
    .B(_03057_),
    .X(_03058_));
 sg13g2_buf_1 _20112_ (.A(_03058_),
    .X(_03059_));
 sg13g2_inv_1 _20113_ (.Y(_03060_),
    .A(_02974_));
 sg13g2_buf_1 _20114_ (.A(_02991_),
    .X(_03061_));
 sg13g2_or4_1 _20115_ (.A(net213),
    .B(_03060_),
    .C(net233),
    .D(_03008_),
    .X(_03062_));
 sg13g2_buf_1 _20116_ (.A(_03062_),
    .X(_03063_));
 sg13g2_buf_1 _20117_ (.A(_03063_),
    .X(_03064_));
 sg13g2_o21ai_1 _20118_ (.B1(_03035_),
    .Y(_03065_),
    .A1(net247),
    .A2(net121));
 sg13g2_buf_1 _20119_ (.A(_03065_),
    .X(_03066_));
 sg13g2_a21oi_1 _20120_ (.A1(net245),
    .A2(net121),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_o21ai_1 _20121_ (.B1(_03028_),
    .Y(_03068_),
    .A1(_03059_),
    .A2(_03067_));
 sg13g2_nand3_1 _20122_ (.B(_03055_),
    .C(_03068_),
    .A(_03044_),
    .Y(_03069_));
 sg13g2_mux2_1 _20123_ (.A0(_03069_),
    .A1(\cpu.dec.imm[11] ),
    .S(net103),
    .X(_00758_));
 sg13g2_o21ai_1 _20124_ (.B1(_03048_),
    .Y(_03070_),
    .A1(_08803_),
    .A2(_03053_));
 sg13g2_nand2_1 _20125_ (.Y(_03071_),
    .A(_03046_),
    .B(_03070_));
 sg13g2_a21oi_1 _20126_ (.A1(_08803_),
    .A2(net121),
    .Y(_03072_),
    .B1(_03066_));
 sg13g2_o21ai_1 _20127_ (.B1(_03028_),
    .Y(_03073_),
    .A1(_03059_),
    .A2(_03072_));
 sg13g2_nand3_1 _20128_ (.B(_03071_),
    .C(_03073_),
    .A(_03044_),
    .Y(_03074_));
 sg13g2_mux2_1 _20129_ (.A0(_03074_),
    .A1(\cpu.dec.imm[12] ),
    .S(net103),
    .X(_00759_));
 sg13g2_or4_1 _20130_ (.A(net286),
    .B(net214),
    .C(_08835_),
    .D(_03026_),
    .X(_03075_));
 sg13g2_a21oi_1 _20131_ (.A1(net214),
    .A2(net121),
    .Y(_03076_),
    .B1(_03066_));
 sg13g2_o21ai_1 _20132_ (.B1(_03028_),
    .Y(_03077_),
    .A1(_03059_),
    .A2(_03076_));
 sg13g2_nand3_1 _20133_ (.B(_03075_),
    .C(_03077_),
    .A(_03044_),
    .Y(_03078_));
 sg13g2_mux2_1 _20134_ (.A0(_03078_),
    .A1(\cpu.dec.imm[13] ),
    .S(net103),
    .X(_00760_));
 sg13g2_o21ai_1 _20135_ (.B1(_03048_),
    .Y(_03079_),
    .A1(net244),
    .A2(_03053_));
 sg13g2_nand2_1 _20136_ (.Y(_03080_),
    .A(_03046_),
    .B(_03079_));
 sg13g2_a21oi_1 _20137_ (.A1(net244),
    .A2(net121),
    .Y(_03081_),
    .B1(_03066_));
 sg13g2_o21ai_1 _20138_ (.B1(_03028_),
    .Y(_03082_),
    .A1(_03059_),
    .A2(_03081_));
 sg13g2_nand2_1 _20139_ (.Y(_03083_),
    .A(_03044_),
    .B(_03082_));
 sg13g2_nor2_1 _20140_ (.A(net104),
    .B(_03083_),
    .Y(_03084_));
 sg13g2_a22oi_1 _20141_ (.Y(_00761_),
    .B1(_03080_),
    .B2(_03084_),
    .A2(_09630_),
    .A1(_10265_));
 sg13g2_o21ai_1 _20142_ (.B1(_03048_),
    .Y(_03085_),
    .A1(_08741_),
    .A2(_03053_));
 sg13g2_a21oi_1 _20143_ (.A1(_03046_),
    .A2(_03085_),
    .Y(_03086_),
    .B1(_03083_));
 sg13g2_nand2_1 _20144_ (.Y(_03087_),
    .A(\cpu.dec.imm[15] ),
    .B(net109));
 sg13g2_o21ai_1 _20145_ (.B1(_03087_),
    .Y(_00762_),
    .A1(_09630_),
    .A2(_03086_));
 sg13g2_o21ai_1 _20146_ (.B1(net284),
    .Y(_03088_),
    .A1(net286),
    .A2(_03064_));
 sg13g2_nand2_1 _20147_ (.Y(_03089_),
    .A(net285),
    .B(net339));
 sg13g2_nand2_1 _20148_ (.Y(_03090_),
    .A(net176),
    .B(_02922_));
 sg13g2_nand2_1 _20149_ (.Y(_03091_),
    .A(_03089_),
    .B(_03090_));
 sg13g2_a21oi_1 _20150_ (.A1(net198),
    .A2(_03088_),
    .Y(_03092_),
    .B1(_03091_));
 sg13g2_nor2_1 _20151_ (.A(net197),
    .B(_08719_),
    .Y(_03093_));
 sg13g2_o21ai_1 _20152_ (.B1(_03093_),
    .Y(_03094_),
    .A1(net196),
    .A2(_03092_));
 sg13g2_nand2_1 _20153_ (.Y(_03095_),
    .A(_02930_),
    .B(_02955_));
 sg13g2_nor2_1 _20154_ (.A(_09680_),
    .B(_02915_),
    .Y(_03096_));
 sg13g2_a22oi_1 _20155_ (.Y(_03097_),
    .B1(_03095_),
    .B2(_03096_),
    .A2(_03094_),
    .A1(_08802_));
 sg13g2_nand2_1 _20156_ (.Y(_03098_),
    .A(_11048_),
    .B(net109));
 sg13g2_o21ai_1 _20157_ (.B1(_03098_),
    .Y(_00763_),
    .A1(net90),
    .A2(_03097_));
 sg13g2_nor2_1 _20158_ (.A(net177),
    .B(net198),
    .Y(_03099_));
 sg13g2_and2_1 _20159_ (.A(_03099_),
    .B(_03040_),
    .X(_03100_));
 sg13g2_nand2_1 _20160_ (.Y(_03101_),
    .A(net285),
    .B(net248));
 sg13g2_o21ai_1 _20161_ (.B1(_03101_),
    .Y(_03102_),
    .A1(net285),
    .A2(_09680_));
 sg13g2_or2_1 _20162_ (.X(_03103_),
    .B(_03026_),
    .A(net197));
 sg13g2_o21ai_1 _20163_ (.B1(_03090_),
    .Y(_03104_),
    .A1(net197),
    .A2(_03089_));
 sg13g2_a22oi_1 _20164_ (.Y(_03105_),
    .B1(_03104_),
    .B2(net212),
    .A2(_03103_),
    .A1(_02934_));
 sg13g2_nor2_1 _20165_ (.A(_03015_),
    .B(_03026_),
    .Y(_03106_));
 sg13g2_or2_1 _20166_ (.X(_03107_),
    .B(_03063_),
    .A(_03053_));
 sg13g2_buf_1 _20167_ (.A(_03107_),
    .X(_03108_));
 sg13g2_inv_1 _20168_ (.Y(_03109_),
    .A(_03108_));
 sg13g2_nand3_1 _20169_ (.B(_03109_),
    .C(_03106_),
    .A(net248),
    .Y(_03110_));
 sg13g2_o21ai_1 _20170_ (.B1(_03110_),
    .Y(_03111_),
    .A1(_08832_),
    .A2(net243));
 sg13g2_o21ai_1 _20171_ (.B1(_03111_),
    .Y(_03112_),
    .A1(_03046_),
    .A2(_03106_));
 sg13g2_o21ai_1 _20172_ (.B1(_03112_),
    .Y(_03113_),
    .A1(net251),
    .A2(_03105_));
 sg13g2_a221oi_1 _20173_ (.B2(_03102_),
    .C1(_03113_),
    .B1(_03100_),
    .A1(net211),
    .Y(_03114_),
    .A2(_03095_));
 sg13g2_nand2_1 _20174_ (.Y(_03115_),
    .A(_11078_),
    .B(_09636_));
 sg13g2_o21ai_1 _20175_ (.B1(_03115_),
    .Y(_00764_),
    .A1(net90),
    .A2(_03114_));
 sg13g2_a22oi_1 _20176_ (.Y(_03116_),
    .B1(net150),
    .B2(net213),
    .A2(net211),
    .A1(net155));
 sg13g2_nor3_1 _20177_ (.A(net244),
    .B(_03053_),
    .C(_03064_),
    .Y(_03117_));
 sg13g2_a21oi_1 _20178_ (.A1(_08856_),
    .A2(net195),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_nand2_1 _20179_ (.Y(_03119_),
    .A(_03116_),
    .B(_03118_));
 sg13g2_o21ai_1 _20180_ (.B1(_03116_),
    .Y(_03120_),
    .A1(net245),
    .A2(_09664_));
 sg13g2_nand2_1 _20181_ (.Y(_03121_),
    .A(net176),
    .B(net286));
 sg13g2_a21oi_1 _20182_ (.A1(_03121_),
    .A2(_03103_),
    .Y(_03122_),
    .B1(_03041_));
 sg13g2_nand3_1 _20183_ (.B(_09679_),
    .C(_03100_),
    .A(net286),
    .Y(_03123_));
 sg13g2_o21ai_1 _20184_ (.B1(_03123_),
    .Y(_03124_),
    .A1(net244),
    .A2(_03122_));
 sg13g2_a221oi_1 _20185_ (.B2(_02952_),
    .C1(_03124_),
    .B1(_03120_),
    .A1(_03106_),
    .Y(_03125_),
    .A2(_03119_));
 sg13g2_nand2_1 _20186_ (.Y(_03126_),
    .A(_11112_),
    .B(net104));
 sg13g2_o21ai_1 _20187_ (.B1(_03126_),
    .Y(_00765_),
    .A1(_08624_),
    .A2(_03125_));
 sg13g2_nand2_1 _20188_ (.Y(_03127_),
    .A(_02939_),
    .B(_03088_));
 sg13g2_a21o_1 _20189_ (.A2(_03127_),
    .A1(_03093_),
    .B1(net214),
    .X(_03128_));
 sg13g2_o21ai_1 _20190_ (.B1(_03128_),
    .Y(_03129_),
    .A1(net244),
    .A2(_02930_));
 sg13g2_mux2_1 _20191_ (.A0(_03129_),
    .A1(\cpu.dec.imm[4] ),
    .S(net103),
    .X(_00766_));
 sg13g2_a21oi_1 _20192_ (.A1(_02947_),
    .A2(_03093_),
    .Y(_03130_),
    .B1(net246));
 sg13g2_nor2_1 _20193_ (.A(net175),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_nand2_1 _20194_ (.Y(_03132_),
    .A(_02938_),
    .B(net286));
 sg13g2_o21ai_1 _20195_ (.B1(_03101_),
    .Y(_03133_),
    .A1(net246),
    .A2(_03132_));
 sg13g2_a221oi_1 _20196_ (.B2(net339),
    .C1(_02919_),
    .B1(_03133_),
    .A1(_08717_),
    .Y(_03134_),
    .A2(_03018_));
 sg13g2_nand3_1 _20197_ (.B(_03035_),
    .C(net121),
    .A(net175),
    .Y(_03135_));
 sg13g2_a21oi_1 _20198_ (.A1(_09678_),
    .A2(_03135_),
    .Y(_03136_),
    .B1(net174));
 sg13g2_nor4_1 _20199_ (.A(_08623_),
    .B(_03131_),
    .C(_03134_),
    .D(_03136_),
    .Y(_03137_));
 sg13g2_a21o_1 _20200_ (.A2(_09677_),
    .A1(\cpu.dec.imm[5] ),
    .B1(_03137_),
    .X(_00767_));
 sg13g2_buf_1 _20201_ (.A(_03008_),
    .X(_03138_));
 sg13g2_nand2_1 _20202_ (.Y(_03139_),
    .A(_03029_),
    .B(_03138_));
 sg13g2_o21ai_1 _20203_ (.B1(_03139_),
    .Y(_03140_),
    .A1(net243),
    .A2(_03108_));
 sg13g2_a21o_1 _20204_ (.A2(_03040_),
    .A1(net286),
    .B1(net243),
    .X(_03141_));
 sg13g2_nand3_1 _20205_ (.B(net176),
    .C(_03141_),
    .A(net174),
    .Y(_03142_));
 sg13g2_o21ai_1 _20206_ (.B1(_02913_),
    .Y(_03143_),
    .A1(net245),
    .A2(_02947_));
 sg13g2_nor4_1 _20207_ (.A(_02914_),
    .B(_02938_),
    .C(_03025_),
    .D(net243),
    .Y(_03144_));
 sg13g2_a221oi_1 _20208_ (.B2(_03143_),
    .C1(_03144_),
    .B1(_03142_),
    .A1(_03106_),
    .Y(_03145_),
    .A2(_03140_));
 sg13g2_nor2_1 _20209_ (.A(_08681_),
    .B(_08718_),
    .Y(_03146_));
 sg13g2_a221oi_1 _20210_ (.B2(_03146_),
    .C1(_02919_),
    .B1(net232),
    .A1(net127),
    .Y(_03147_),
    .A2(_09639_));
 sg13g2_nor3_1 _20211_ (.A(net108),
    .B(_03145_),
    .C(_03147_),
    .Y(_03148_));
 sg13g2_a21o_1 _20212_ (.A2(net89),
    .A1(\cpu.dec.imm[6] ),
    .B1(_03148_),
    .X(_00768_));
 sg13g2_inv_1 _20213_ (.Y(_03149_),
    .A(_02930_));
 sg13g2_a22oi_1 _20214_ (.Y(_03150_),
    .B1(_03088_),
    .B2(_08664_),
    .A2(_03029_),
    .A1(_03099_));
 sg13g2_or2_1 _20215_ (.X(_03151_),
    .B(_03089_),
    .A(_09666_));
 sg13g2_o21ai_1 _20216_ (.B1(_03151_),
    .Y(_03152_),
    .A1(net196),
    .A2(_03150_));
 sg13g2_a221oi_1 _20217_ (.B2(net211),
    .C1(_02915_),
    .B1(_03152_),
    .A1(_08802_),
    .Y(_03153_),
    .A2(_03149_));
 sg13g2_a221oi_1 _20218_ (.B2(_03146_),
    .C1(_02919_),
    .B1(_02974_),
    .A1(net127),
    .Y(_03154_),
    .A2(net211));
 sg13g2_nor3_1 _20219_ (.A(net108),
    .B(_03153_),
    .C(_03154_),
    .Y(_03155_));
 sg13g2_a21o_1 _20220_ (.A2(_09677_),
    .A1(\cpu.dec.imm[7] ),
    .B1(_03155_),
    .X(_00769_));
 sg13g2_o21ai_1 _20221_ (.B1(_03048_),
    .Y(_03156_),
    .A1(net246),
    .A2(_03053_));
 sg13g2_a21o_1 _20222_ (.A2(net121),
    .A1(net246),
    .B1(_03066_),
    .X(_03157_));
 sg13g2_nand2_1 _20223_ (.Y(_03158_),
    .A(net195),
    .B(net233));
 sg13g2_nand3_1 _20224_ (.B(_03157_),
    .C(_03158_),
    .A(_03031_),
    .Y(_03159_));
 sg13g2_nand3_1 _20225_ (.B(net233),
    .C(_03146_),
    .A(_02915_),
    .Y(_03160_));
 sg13g2_nand2_1 _20226_ (.Y(_03161_),
    .A(_03044_),
    .B(_03160_));
 sg13g2_a221oi_1 _20227_ (.B2(_03028_),
    .C1(_03161_),
    .B1(_03159_),
    .A1(_03046_),
    .Y(_03162_),
    .A2(_03156_));
 sg13g2_nand2_1 _20228_ (.Y(_03163_),
    .A(\cpu.dec.imm[8] ),
    .B(_02912_));
 sg13g2_o21ai_1 _20229_ (.B1(_03163_),
    .Y(_00770_),
    .A1(net91),
    .A2(_03162_));
 sg13g2_o21ai_1 _20230_ (.B1(_03048_),
    .Y(_03164_),
    .A1(net243),
    .A2(_03053_));
 sg13g2_nand2_1 _20231_ (.Y(_03165_),
    .A(_03046_),
    .B(_03164_));
 sg13g2_a21oi_1 _20232_ (.A1(net243),
    .A2(net121),
    .Y(_03166_),
    .B1(_03066_));
 sg13g2_inv_1 _20233_ (.Y(_03167_),
    .A(net195));
 sg13g2_o21ai_1 _20234_ (.B1(_03031_),
    .Y(_03168_),
    .A1(net251),
    .A2(_03167_));
 sg13g2_o21ai_1 _20235_ (.B1(_03028_),
    .Y(_03169_),
    .A1(_03166_),
    .A2(_03168_));
 sg13g2_nand3_1 _20236_ (.B(_03165_),
    .C(_03169_),
    .A(_03044_),
    .Y(_03170_));
 sg13g2_mux2_1 _20237_ (.A0(_03170_),
    .A1(\cpu.dec.imm[9] ),
    .S(_02950_),
    .X(_00771_));
 sg13g2_buf_2 _20238_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03171_));
 sg13g2_inv_1 _20239_ (.Y(_03172_),
    .A(_03171_));
 sg13g2_nand2_1 _20240_ (.Y(_03173_),
    .A(net896),
    .B(_02953_));
 sg13g2_nor4_1 _20241_ (.A(_09647_),
    .B(_08803_),
    .C(_03010_),
    .D(_03173_),
    .Y(_03174_));
 sg13g2_nand3_1 _20242_ (.B(_02952_),
    .C(_03174_),
    .A(net132),
    .Y(_03175_));
 sg13g2_o21ai_1 _20243_ (.B1(_03175_),
    .Y(_00772_),
    .A1(_03172_),
    .A2(net112));
 sg13g2_nor4_1 _20244_ (.A(net196),
    .B(net249),
    .C(net126),
    .D(_02942_),
    .Y(_03176_));
 sg13g2_mux2_1 _20245_ (.A0(_03176_),
    .A1(\cpu.dec.io ),
    .S(net103),
    .X(_00773_));
 sg13g2_or3_1 _20246_ (.A(_08825_),
    .B(net247),
    .C(_08924_),
    .X(_03177_));
 sg13g2_buf_2 _20247_ (.A(_03177_),
    .X(_03178_));
 sg13g2_nor3_1 _20248_ (.A(_08832_),
    .B(_09666_),
    .C(_03178_),
    .Y(_03179_));
 sg13g2_mux2_1 _20249_ (.A0(_03179_),
    .A1(\cpu.dec.jmp ),
    .S(_09636_),
    .X(_00774_));
 sg13g2_inv_1 _20250_ (.Y(_03180_),
    .A(_11205_));
 sg13g2_o21ai_1 _20251_ (.B1(net177),
    .Y(_03181_),
    .A1(net175),
    .A2(net284));
 sg13g2_nand3_1 _20252_ (.B(_03033_),
    .C(_03181_),
    .A(net132),
    .Y(_03182_));
 sg13g2_o21ai_1 _20253_ (.B1(_03182_),
    .Y(_00775_),
    .A1(_03180_),
    .A2(net112));
 sg13g2_nor4_1 _20254_ (.A(net113),
    .B(_09647_),
    .C(_08825_),
    .D(_08837_),
    .Y(_03183_));
 sg13g2_a21o_1 _20255_ (.A2(net89),
    .A1(_09106_),
    .B1(_03183_),
    .X(_00776_));
 sg13g2_a21oi_1 _20256_ (.A1(net244),
    .A2(_09647_),
    .Y(_03184_),
    .B1(_08826_));
 sg13g2_nand3_1 _20257_ (.B(net212),
    .C(net214),
    .A(net197),
    .Y(_03185_));
 sg13g2_nand3_1 _20258_ (.B(net196),
    .C(_09644_),
    .A(net177),
    .Y(_03186_));
 sg13g2_nand4_1 _20259_ (.B(net249),
    .C(_03185_),
    .A(net176),
    .Y(_03187_),
    .D(_03186_));
 sg13g2_o21ai_1 _20260_ (.B1(_03187_),
    .Y(_03188_),
    .A1(_08720_),
    .A2(_03184_));
 sg13g2_nand2_1 _20261_ (.Y(_03189_),
    .A(_08853_),
    .B(_03188_));
 sg13g2_o21ai_1 _20262_ (.B1(_03189_),
    .Y(_00777_),
    .A1(net858),
    .A2(_08852_));
 sg13g2_o21ai_1 _20263_ (.B1(net198),
    .Y(_03190_),
    .A1(_08642_),
    .A2(net232));
 sg13g2_nor3_1 _20264_ (.A(net150),
    .B(net195),
    .C(_03190_),
    .Y(_03191_));
 sg13g2_a21oi_1 _20265_ (.A1(net195),
    .A2(_02939_),
    .Y(_03192_),
    .B1(_03191_));
 sg13g2_nand2_1 _20266_ (.Y(_03193_),
    .A(_09647_),
    .B(_03179_));
 sg13g2_o21ai_1 _20267_ (.B1(_03193_),
    .Y(_03194_),
    .A1(net174),
    .A2(_03192_));
 sg13g2_nand2_1 _20268_ (.Y(_03195_),
    .A(net284),
    .B(net232));
 sg13g2_o21ai_1 _20269_ (.B1(_03195_),
    .Y(_03196_),
    .A1(net284),
    .A2(_08900_));
 sg13g2_a22oi_1 _20270_ (.Y(_03197_),
    .B1(_03033_),
    .B2(_03196_),
    .A2(net232),
    .A1(net127));
 sg13g2_o21ai_1 _20271_ (.B1(_03191_),
    .Y(_03198_),
    .A1(net196),
    .A2(_09678_));
 sg13g2_o21ai_1 _20272_ (.B1(_03198_),
    .Y(_03199_),
    .A1(net126),
    .A2(_03197_));
 sg13g2_a21oi_1 _20273_ (.A1(net249),
    .A2(_03178_),
    .Y(_03200_),
    .B1(net212));
 sg13g2_nor2_1 _20274_ (.A(_09666_),
    .B(_03200_),
    .Y(_03201_));
 sg13g2_and2_1 _20275_ (.A(net232),
    .B(_03201_),
    .X(_03202_));
 sg13g2_nor3_1 _20276_ (.A(_03194_),
    .B(_03199_),
    .C(_03202_),
    .Y(_03203_));
 sg13g2_nand2_1 _20277_ (.Y(_03204_),
    .A(\cpu.dec.r_rd[0] ),
    .B(net104));
 sg13g2_o21ai_1 _20278_ (.B1(_03204_),
    .Y(_00778_),
    .A1(net91),
    .A2(_03203_));
 sg13g2_nor3_1 _20279_ (.A(net196),
    .B(_02919_),
    .C(net195),
    .Y(_03205_));
 sg13g2_a21o_1 _20280_ (.A2(_03016_),
    .A1(_03167_),
    .B1(_03201_),
    .X(_03206_));
 sg13g2_nor2_1 _20281_ (.A(_02933_),
    .B(_03060_),
    .Y(_03207_));
 sg13g2_a21oi_1 _20282_ (.A1(_02933_),
    .A2(_08916_),
    .Y(_03208_),
    .B1(net196));
 sg13g2_o21ai_1 _20283_ (.B1(_08716_),
    .Y(_03209_),
    .A1(_03207_),
    .A2(_03208_));
 sg13g2_nand2_1 _20284_ (.Y(_03210_),
    .A(_02974_),
    .B(_03035_));
 sg13g2_nand4_1 _20285_ (.B(_08803_),
    .C(_08823_),
    .A(_08782_),
    .Y(_03211_),
    .D(_08880_));
 sg13g2_nor2_1 _20286_ (.A(_03010_),
    .B(_03211_),
    .Y(_03212_));
 sg13g2_nand3_1 _20287_ (.B(_09639_),
    .C(_03212_),
    .A(_08900_),
    .Y(_03213_));
 sg13g2_buf_1 _20288_ (.A(_03213_),
    .X(_03214_));
 sg13g2_a221oi_1 _20289_ (.B2(_02953_),
    .C1(net126),
    .B1(_03214_),
    .A1(_03209_),
    .Y(_03215_),
    .A2(_03210_));
 sg13g2_a221oi_1 _20290_ (.B2(_02974_),
    .C1(_03215_),
    .B1(_03206_),
    .A1(_09639_),
    .Y(_03216_),
    .A2(_03205_));
 sg13g2_nand2_1 _20291_ (.Y(_03217_),
    .A(\cpu.dec.r_rd[1] ),
    .B(net104));
 sg13g2_o21ai_1 _20292_ (.B1(_03217_),
    .Y(_00779_),
    .A1(net91),
    .A2(_03216_));
 sg13g2_nand2_1 _20293_ (.Y(_03218_),
    .A(net284),
    .B(net233));
 sg13g2_o21ai_1 _20294_ (.B1(_03218_),
    .Y(_03219_),
    .A1(net284),
    .A2(_08881_));
 sg13g2_a22oi_1 _20295_ (.Y(_03220_),
    .B1(_03033_),
    .B2(_03219_),
    .A2(net233),
    .A1(net127));
 sg13g2_nor2_1 _20296_ (.A(net126),
    .B(_03220_),
    .Y(_03221_));
 sg13g2_a221oi_1 _20297_ (.B2(net233),
    .C1(_03221_),
    .B1(_03206_),
    .A1(net211),
    .Y(_03222_),
    .A2(_03205_));
 sg13g2_nand2_1 _20298_ (.Y(_03223_),
    .A(\cpu.dec.r_rd[2] ),
    .B(net104));
 sg13g2_o21ai_1 _20299_ (.B1(_03223_),
    .Y(_00780_),
    .A1(_08624_),
    .A2(_03222_));
 sg13g2_inv_1 _20300_ (.Y(_03224_),
    .A(\cpu.dec.r_rd[3] ));
 sg13g2_o21ai_1 _20301_ (.B1(net213),
    .Y(_03225_),
    .A1(_09663_),
    .A2(net249));
 sg13g2_nand3_1 _20302_ (.B(_08719_),
    .C(_03178_),
    .A(_02920_),
    .Y(_03226_));
 sg13g2_a221oi_1 _20303_ (.B2(_03034_),
    .C1(net198),
    .B1(_03226_),
    .A1(_02920_),
    .Y(_03227_),
    .A2(_03225_));
 sg13g2_o21ai_1 _20304_ (.B1(net213),
    .Y(_03228_),
    .A1(net285),
    .A2(_03227_));
 sg13g2_nand2_1 _20305_ (.Y(_03229_),
    .A(net284),
    .B(_03228_));
 sg13g2_o21ai_1 _20306_ (.B1(_03229_),
    .Y(_03230_),
    .A1(_03016_),
    .A2(_03227_));
 sg13g2_nor4_1 _20307_ (.A(_08623_),
    .B(_08836_),
    .C(_09667_),
    .D(_03205_),
    .Y(_03231_));
 sg13g2_a22oi_1 _20308_ (.Y(_00781_),
    .B1(_03230_),
    .B2(_03231_),
    .A2(net90),
    .A1(_03224_));
 sg13g2_nand4_1 _20309_ (.B(_08826_),
    .C(_08861_),
    .A(net248),
    .Y(_03232_),
    .D(_08879_));
 sg13g2_o21ai_1 _20310_ (.B1(_08663_),
    .Y(_03233_),
    .A1(_08924_),
    .A2(_03232_));
 sg13g2_nand2_1 _20311_ (.Y(_03234_),
    .A(_02924_),
    .B(_03233_));
 sg13g2_nor3_1 _20312_ (.A(_08662_),
    .B(_08830_),
    .C(_02942_),
    .Y(_03235_));
 sg13g2_a221oi_1 _20313_ (.B2(net252),
    .C1(_03235_),
    .B1(_03234_),
    .A1(_08662_),
    .Y(_03236_),
    .A2(net249));
 sg13g2_a21oi_2 _20314_ (.B1(_08832_),
    .Y(_03237_),
    .A2(_03178_),
    .A1(net250));
 sg13g2_o21ai_1 _20315_ (.B1(_03099_),
    .Y(_03238_),
    .A1(_03146_),
    .A2(_03237_));
 sg13g2_o21ai_1 _20316_ (.B1(_03238_),
    .Y(_03239_),
    .A1(net197),
    .A2(_03236_));
 sg13g2_a21oi_1 _20317_ (.A1(net232),
    .A2(_03239_),
    .Y(_03240_),
    .B1(_02915_));
 sg13g2_a21oi_1 _20318_ (.A1(net285),
    .A2(net232),
    .Y(_03241_),
    .B1(_02916_));
 sg13g2_nor3_1 _20319_ (.A(net108),
    .B(_03240_),
    .C(_03241_),
    .Y(_03242_));
 sg13g2_a21o_1 _20320_ (.A2(net89),
    .A1(_10662_),
    .B1(_03242_),
    .X(_00782_));
 sg13g2_nor2_1 _20321_ (.A(_08642_),
    .B(_03236_),
    .Y(_03243_));
 sg13g2_nor3_1 _20322_ (.A(_08717_),
    .B(_03243_),
    .C(_03237_),
    .Y(_03244_));
 sg13g2_o21ai_1 _20323_ (.B1(_02925_),
    .Y(_03245_),
    .A1(_03060_),
    .A2(_03244_));
 sg13g2_o21ai_1 _20324_ (.B1(_03245_),
    .Y(_03246_),
    .A1(_03099_),
    .A2(_03243_));
 sg13g2_nor2_1 _20325_ (.A(_02925_),
    .B(_02974_),
    .Y(_03247_));
 sg13g2_a22oi_1 _20326_ (.Y(_03248_),
    .B1(_03247_),
    .B2(_09666_),
    .A2(_03246_),
    .A1(_02916_));
 sg13g2_o21ai_1 _20327_ (.B1(_02955_),
    .Y(_03249_),
    .A1(_03015_),
    .A2(_03108_));
 sg13g2_o21ai_1 _20328_ (.B1(net132),
    .Y(_03250_),
    .A1(_03248_),
    .A2(_03249_));
 sg13g2_o21ai_1 _20329_ (.B1(_03250_),
    .Y(_00783_),
    .A1(_10746_),
    .A2(net112));
 sg13g2_nor2_1 _20330_ (.A(net286),
    .B(_02919_),
    .Y(_03251_));
 sg13g2_o21ai_1 _20331_ (.B1(net233),
    .Y(_03252_),
    .A1(_03239_),
    .A2(_03251_));
 sg13g2_nor2b_1 _20332_ (.A(net104),
    .B_N(_02955_),
    .Y(_03253_));
 sg13g2_a22oi_1 _20333_ (.Y(_00784_),
    .B1(_03252_),
    .B2(_03253_),
    .A2(net90),
    .A1(_10733_));
 sg13g2_inv_1 _20334_ (.Y(_03254_),
    .A(_03013_));
 sg13g2_nor2_1 _20335_ (.A(_02953_),
    .B(_03254_),
    .Y(_03255_));
 sg13g2_nand2_1 _20336_ (.Y(_03256_),
    .A(_09632_),
    .B(_03237_));
 sg13g2_a21oi_1 _20337_ (.A1(_03255_),
    .A2(_03256_),
    .Y(_03257_),
    .B1(_09666_));
 sg13g2_nor4_1 _20338_ (.A(_09656_),
    .B(_03243_),
    .C(_03251_),
    .D(_03257_),
    .Y(_03258_));
 sg13g2_a21oi_1 _20339_ (.A1(_10575_),
    .A2(net90),
    .Y(_00785_),
    .B1(_03258_));
 sg13g2_nand2_1 _20340_ (.Y(_03259_),
    .A(_08916_),
    .B(net232));
 sg13g2_nand2_1 _20341_ (.Y(_03260_),
    .A(_09678_),
    .B(_09642_));
 sg13g2_o21ai_1 _20342_ (.B1(_03260_),
    .Y(_03261_),
    .A1(_03232_),
    .A2(_03259_));
 sg13g2_nor2_1 _20343_ (.A(_09638_),
    .B(_03040_),
    .Y(_03262_));
 sg13g2_a21oi_1 _20344_ (.A1(net127),
    .A2(_03261_),
    .Y(_03263_),
    .B1(_03262_));
 sg13g2_nor2_1 _20345_ (.A(_02917_),
    .B(_02947_),
    .Y(_03264_));
 sg13g2_nand2_1 _20346_ (.Y(_03265_),
    .A(_03138_),
    .B(_03264_));
 sg13g2_o21ai_1 _20347_ (.B1(_03265_),
    .Y(_03266_),
    .A1(_09638_),
    .A2(net150));
 sg13g2_a22oi_1 _20348_ (.Y(_03267_),
    .B1(_03266_),
    .B2(net174),
    .A2(_09678_),
    .A1(net175));
 sg13g2_o21ai_1 _20349_ (.B1(_03267_),
    .Y(_03268_),
    .A1(_09645_),
    .A2(_03263_));
 sg13g2_nand2_1 _20350_ (.Y(_03269_),
    .A(net111),
    .B(_03268_));
 sg13g2_o21ai_1 _20351_ (.B1(_03269_),
    .Y(_00786_),
    .A1(_10028_),
    .A2(net111));
 sg13g2_a22oi_1 _20352_ (.Y(_03270_),
    .B1(_02927_),
    .B2(_02936_),
    .A2(_08925_),
    .A1(net246));
 sg13g2_nor3_1 _20353_ (.A(_02934_),
    .B(_03060_),
    .C(_03270_),
    .Y(_03271_));
 sg13g2_nand2_1 _20354_ (.Y(_03272_),
    .A(_02952_),
    .B(_03040_));
 sg13g2_o21ai_1 _20355_ (.B1(_03272_),
    .Y(_03273_),
    .A1(_09666_),
    .A2(_02947_));
 sg13g2_o21ai_1 _20356_ (.B1(_09631_),
    .Y(_03274_),
    .A1(_09642_),
    .A2(_03272_));
 sg13g2_a21oi_1 _20357_ (.A1(_03273_),
    .A2(_03274_),
    .Y(_03275_),
    .B1(net243));
 sg13g2_o21ai_1 _20358_ (.B1(net132),
    .Y(_03276_),
    .A1(_03271_),
    .A2(_03275_));
 sg13g2_o21ai_1 _20359_ (.B1(_03276_),
    .Y(_00787_),
    .A1(net664),
    .A2(net111));
 sg13g2_a22oi_1 _20360_ (.Y(_03277_),
    .B1(_03061_),
    .B2(_03264_),
    .A2(_02947_),
    .A1(_09679_));
 sg13g2_nor2_1 _20361_ (.A(_02913_),
    .B(_03277_),
    .Y(_03278_));
 sg13g2_nor3_1 _20362_ (.A(_08924_),
    .B(_09640_),
    .C(_03061_),
    .Y(_03279_));
 sg13g2_o21ai_1 _20363_ (.B1(_03040_),
    .Y(_03280_),
    .A1(_08832_),
    .A2(_03279_));
 sg13g2_a21oi_1 _20364_ (.A1(net177),
    .A2(_03280_),
    .Y(_03281_),
    .B1(net175));
 sg13g2_nor2_1 _20365_ (.A(_08881_),
    .B(_03281_),
    .Y(_03282_));
 sg13g2_o21ai_1 _20366_ (.B1(net132),
    .Y(_03283_),
    .A1(_03278_),
    .A2(_03282_));
 sg13g2_o21ai_1 _20367_ (.B1(_03283_),
    .Y(_00788_),
    .A1(net738),
    .A2(net111));
 sg13g2_nand2b_1 _20368_ (.Y(_03284_),
    .B(_08924_),
    .A_N(_09642_));
 sg13g2_a21oi_1 _20369_ (.A1(_09631_),
    .A2(_03284_),
    .Y(_03285_),
    .B1(_03272_));
 sg13g2_a22oi_1 _20370_ (.Y(_03286_),
    .B1(_02927_),
    .B2(_08760_),
    .A2(_09646_),
    .A1(net127));
 sg13g2_nor2_1 _20371_ (.A(_09666_),
    .B(_03286_),
    .Y(_03287_));
 sg13g2_nor3_1 _20372_ (.A(_09656_),
    .B(_03285_),
    .C(_03287_),
    .Y(_03288_));
 sg13g2_a21o_1 _20373_ (.A2(net89),
    .A1(net656),
    .B1(_03288_),
    .X(_00789_));
 sg13g2_nand2_1 _20374_ (.Y(_03289_),
    .A(_09979_),
    .B(net104));
 sg13g2_o21ai_1 _20375_ (.B1(_03289_),
    .Y(_00790_),
    .A1(net91),
    .A2(_08918_));
 sg13g2_nor4_1 _20376_ (.A(_08832_),
    .B(net126),
    .C(_08924_),
    .D(_09642_),
    .Y(_03290_));
 sg13g2_mux2_1 _20377_ (.A0(_03290_),
    .A1(_09978_),
    .S(net109),
    .X(_00791_));
 sg13g2_nor3_1 _20378_ (.A(_08784_),
    .B(_08802_),
    .C(_08860_),
    .Y(_03291_));
 sg13g2_mux2_1 _20379_ (.A0(_03291_),
    .A1(\cpu.dec.r_set_cc ),
    .S(net109),
    .X(_00792_));
 sg13g2_nand2_1 _20380_ (.Y(_03292_),
    .A(net174),
    .B(net150));
 sg13g2_o21ai_1 _20381_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net174),
    .A2(_03090_));
 sg13g2_buf_1 _20382_ (.A(\cpu.dec.r_store ),
    .X(_03294_));
 sg13g2_mux2_1 _20383_ (.A0(_03293_),
    .A1(_03294_),
    .S(net109),
    .X(_00793_));
 sg13g2_nor3_1 _20384_ (.A(net108),
    .B(_02955_),
    .C(_03214_),
    .Y(_03295_));
 sg13g2_a21o_1 _20385_ (.A2(net103),
    .A1(\cpu.dec.r_swapsp ),
    .B1(_03295_),
    .X(_00794_));
 sg13g2_inv_1 _20386_ (.Y(_03296_),
    .A(\cpu.dec.r_sys_call ));
 sg13g2_nor4_1 _20387_ (.A(net126),
    .B(net246),
    .C(_09639_),
    .D(_09664_),
    .Y(_03297_));
 sg13g2_nand3_1 _20388_ (.B(_03212_),
    .C(_03297_),
    .A(_08851_),
    .Y(_03298_));
 sg13g2_o21ai_1 _20389_ (.B1(_03298_),
    .Y(_00795_),
    .A1(_03296_),
    .A2(_08853_));
 sg13g2_a21oi_1 _20390_ (.A1(_03011_),
    .A2(_03214_),
    .Y(_03299_),
    .B1(_03173_));
 sg13g2_nor3_1 _20391_ (.A(_08835_),
    .B(_03174_),
    .C(_03299_),
    .Y(_03300_));
 sg13g2_nand3_1 _20392_ (.B(net247),
    .C(_08924_),
    .A(net248),
    .Y(_03301_));
 sg13g2_nand2_1 _20393_ (.Y(_03302_),
    .A(net213),
    .B(_09647_));
 sg13g2_a21oi_1 _20394_ (.A1(_08803_),
    .A2(_03301_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_o21ai_1 _20395_ (.B1(net155),
    .Y(_03304_),
    .A1(_09657_),
    .A2(_03303_));
 sg13g2_buf_1 _20396_ (.A(net896),
    .X(_03305_));
 sg13g2_nand3_1 _20397_ (.B(net250),
    .C(_09633_),
    .A(_03305_),
    .Y(_03306_));
 sg13g2_o21ai_1 _20398_ (.B1(_03254_),
    .Y(_03307_),
    .A1(_03178_),
    .A2(_03306_));
 sg13g2_nor3_1 _20399_ (.A(_03305_),
    .B(_10388_),
    .C(_02942_),
    .Y(_03308_));
 sg13g2_o21ai_1 _20400_ (.B1(net212),
    .Y(_03309_),
    .A1(net249),
    .A2(_03308_));
 sg13g2_nand2_1 _20401_ (.Y(_03310_),
    .A(_02974_),
    .B(_03008_));
 sg13g2_xor2_1 _20402_ (.B(_03310_),
    .A(net233),
    .X(_03311_));
 sg13g2_nor2_1 _20403_ (.A(net896),
    .B(_03311_),
    .Y(_03312_));
 sg13g2_nand3_1 _20404_ (.B(_03035_),
    .C(_03312_),
    .A(_08760_),
    .Y(_03313_));
 sg13g2_nand4_1 _20405_ (.B(_03307_),
    .C(_03309_),
    .A(_03304_),
    .Y(_03314_),
    .D(_03313_));
 sg13g2_a22oi_1 _20406_ (.Y(_03315_),
    .B1(_08825_),
    .B2(_08740_),
    .A2(_08802_),
    .A1(net213));
 sg13g2_nand3_1 _20407_ (.B(net250),
    .C(_09678_),
    .A(_09657_),
    .Y(_03316_));
 sg13g2_o21ai_1 _20408_ (.B1(_03316_),
    .Y(_03317_),
    .A1(net214),
    .A2(_03315_));
 sg13g2_nand2_1 _20409_ (.Y(_03318_),
    .A(net155),
    .B(_03317_));
 sg13g2_nand2_1 _20410_ (.Y(_03319_),
    .A(_03313_),
    .B(_03318_));
 sg13g2_a22oi_1 _20411_ (.Y(_03320_),
    .B1(_03319_),
    .B2(_08664_),
    .A2(_03314_),
    .A1(_03300_));
 sg13g2_o21ai_1 _20412_ (.B1(net251),
    .Y(_03321_),
    .A1(_08681_),
    .A2(_03237_));
 sg13g2_nand2_1 _20413_ (.Y(_03322_),
    .A(_03040_),
    .B(_03321_));
 sg13g2_and2_1 _20414_ (.A(_03312_),
    .B(_03322_),
    .X(_03323_));
 sg13g2_xor2_1 _20415_ (.B(_08917_),
    .A(net247),
    .X(_03324_));
 sg13g2_nand2_1 _20416_ (.Y(_03325_),
    .A(_08514_),
    .B(_08783_));
 sg13g2_o21ai_1 _20417_ (.B1(_03325_),
    .Y(_03326_),
    .A1(net710),
    .A2(_08783_));
 sg13g2_nand4_1 _20418_ (.B(_09646_),
    .C(_03324_),
    .A(net155),
    .Y(_03327_),
    .D(_03326_));
 sg13g2_a21oi_1 _20419_ (.A1(net214),
    .A2(_08900_),
    .Y(_03328_),
    .B1(_09664_));
 sg13g2_o21ai_1 _20420_ (.B1(_03328_),
    .Y(_03329_),
    .A1(net214),
    .A2(_08825_));
 sg13g2_nand4_1 _20421_ (.B(_03013_),
    .C(_03327_),
    .A(_02914_),
    .Y(_03330_),
    .D(_03329_));
 sg13g2_o21ai_1 _20422_ (.B1(_02936_),
    .Y(_03331_),
    .A1(_03323_),
    .A2(_03330_));
 sg13g2_a21oi_1 _20423_ (.A1(net245),
    .A2(_03009_),
    .Y(_03332_),
    .B1(_08832_));
 sg13g2_nor3_1 _20424_ (.A(_09664_),
    .B(_03010_),
    .C(_03178_),
    .Y(_03333_));
 sg13g2_nor4_1 _20425_ (.A(_02919_),
    .B(net195),
    .C(_03332_),
    .D(_03333_),
    .Y(_03334_));
 sg13g2_a21oi_1 _20426_ (.A1(_03320_),
    .A2(_03331_),
    .Y(_03335_),
    .B1(_03334_));
 sg13g2_nand2_1 _20427_ (.Y(_03336_),
    .A(net132),
    .B(_03335_));
 sg13g2_o21ai_1 _20428_ (.B1(_03336_),
    .Y(_00796_),
    .A1(_10515_),
    .A2(net111));
 sg13g2_buf_1 _20429_ (.A(_08588_),
    .X(_03337_));
 sg13g2_buf_1 _20430_ (.A(net951),
    .X(_03338_));
 sg13g2_buf_1 _20431_ (.A(net831),
    .X(_03339_));
 sg13g2_nand2b_1 _20432_ (.Y(_03340_),
    .B(net1077),
    .A_N(net1003));
 sg13g2_buf_1 _20433_ (.A(_03340_),
    .X(_03341_));
 sg13g2_nand3_1 _20434_ (.B(_09968_),
    .C(_09960_),
    .A(net1076),
    .Y(_03342_));
 sg13g2_buf_1 _20435_ (.A(_03342_),
    .X(_03343_));
 sg13g2_nor2_1 _20436_ (.A(_03341_),
    .B(_03343_),
    .Y(_03344_));
 sg13g2_buf_4 _20437_ (.X(_03345_),
    .A(_03344_));
 sg13g2_buf_1 _20438_ (.A(_03345_),
    .X(_03346_));
 sg13g2_mux2_1 _20439_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net709),
    .S(net509),
    .X(_00801_));
 sg13g2_buf_1 _20440_ (.A(net953),
    .X(_03347_));
 sg13g2_mux2_1 _20441_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net830),
    .S(net509),
    .X(_00802_));
 sg13g2_mux2_1 _20442_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net832),
    .S(net509),
    .X(_00803_));
 sg13g2_buf_1 _20443_ (.A(net576),
    .X(_03348_));
 sg13g2_nand2_1 _20444_ (.Y(_03349_),
    .A(net508),
    .B(_03345_));
 sg13g2_o21ai_1 _20445_ (.B1(_03349_),
    .Y(_00804_),
    .A1(_10333_),
    .A2(_03346_));
 sg13g2_buf_1 _20446_ (.A(net577),
    .X(_03350_));
 sg13g2_buf_1 _20447_ (.A(net507),
    .X(_03351_));
 sg13g2_mux2_1 _20448_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net443),
    .S(net509),
    .X(_00805_));
 sg13g2_buf_1 _20449_ (.A(net578),
    .X(_03352_));
 sg13g2_buf_1 _20450_ (.A(net506),
    .X(_03353_));
 sg13g2_mux2_1 _20451_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net442),
    .S(net509),
    .X(_00806_));
 sg13g2_buf_1 _20452_ (.A(net994),
    .X(_03354_));
 sg13g2_mux2_1 _20453_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net829),
    .S(_03346_),
    .X(_00807_));
 sg13g2_buf_1 _20454_ (.A(net530),
    .X(_03355_));
 sg13g2_mux2_1 _20455_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net441),
    .S(net509),
    .X(_00808_));
 sg13g2_buf_2 _20456_ (.A(net692),
    .X(_03356_));
 sg13g2_buf_1 _20457_ (.A(_03356_),
    .X(_03357_));
 sg13g2_mux2_1 _20458_ (.A0(\cpu.ex.r_10[2] ),
    .A1(_03357_),
    .S(net509),
    .X(_00809_));
 sg13g2_buf_1 _20459_ (.A(net538),
    .X(_03358_));
 sg13g2_mux2_1 _20460_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net440),
    .S(net509),
    .X(_00810_));
 sg13g2_buf_1 _20461_ (.A(net573),
    .X(_03359_));
 sg13g2_mux2_1 _20462_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net504),
    .S(_03345_),
    .X(_00811_));
 sg13g2_mux2_1 _20463_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net512),
    .S(_03345_),
    .X(_00812_));
 sg13g2_mux2_1 _20464_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net713),
    .S(_03345_),
    .X(_00813_));
 sg13g2_mux2_1 _20465_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net711),
    .S(_03345_),
    .X(_00814_));
 sg13g2_mux2_1 _20466_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net833),
    .S(_03345_),
    .X(_00815_));
 sg13g2_mux2_1 _20467_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net836),
    .S(_03345_),
    .X(_00816_));
 sg13g2_nor2_1 _20468_ (.A(_09965_),
    .B(_03343_),
    .Y(_03360_));
 sg13g2_buf_2 _20469_ (.A(_03360_),
    .X(_03361_));
 sg13g2_buf_1 _20470_ (.A(_03361_),
    .X(_03362_));
 sg13g2_mux2_1 _20471_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net709),
    .S(net503),
    .X(_00817_));
 sg13g2_mux2_1 _20472_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net830),
    .S(net503),
    .X(_00818_));
 sg13g2_mux2_1 _20473_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net832),
    .S(net503),
    .X(_00819_));
 sg13g2_buf_1 _20474_ (.A(net508),
    .X(_03363_));
 sg13g2_mux2_1 _20475_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net439),
    .S(net503),
    .X(_00820_));
 sg13g2_mux2_1 _20476_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net443),
    .S(net503),
    .X(_00821_));
 sg13g2_mux2_1 _20477_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net442),
    .S(_03362_),
    .X(_00822_));
 sg13g2_mux2_1 _20478_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net829),
    .S(net503),
    .X(_00823_));
 sg13g2_mux2_1 _20479_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net441),
    .S(net503),
    .X(_00824_));
 sg13g2_mux2_1 _20480_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net505),
    .S(net503),
    .X(_00825_));
 sg13g2_mux2_1 _20481_ (.A0(\cpu.ex.r_11[3] ),
    .A1(net440),
    .S(_03362_),
    .X(_00826_));
 sg13g2_mux2_1 _20482_ (.A0(\cpu.ex.r_11[4] ),
    .A1(_03359_),
    .S(_03361_),
    .X(_00827_));
 sg13g2_mux2_1 _20483_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net512),
    .S(_03361_),
    .X(_00828_));
 sg13g2_mux2_1 _20484_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net713),
    .S(_03361_),
    .X(_00829_));
 sg13g2_mux2_1 _20485_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net711),
    .S(_03361_),
    .X(_00830_));
 sg13g2_mux2_1 _20486_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net833),
    .S(_03361_),
    .X(_00831_));
 sg13g2_mux2_1 _20487_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net836),
    .S(_03361_),
    .X(_00832_));
 sg13g2_nand3_1 _20488_ (.B(_09967_),
    .C(_09960_),
    .A(net1076),
    .Y(_03364_));
 sg13g2_buf_1 _20489_ (.A(_03364_),
    .X(_03365_));
 sg13g2_nor3_1 _20490_ (.A(net1077),
    .B(net1003),
    .C(_03365_),
    .Y(_03366_));
 sg13g2_buf_2 _20491_ (.A(_03366_),
    .X(_03367_));
 sg13g2_buf_1 _20492_ (.A(_03367_),
    .X(_03368_));
 sg13g2_mux2_1 _20493_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net709),
    .S(net564),
    .X(_00833_));
 sg13g2_mux2_1 _20494_ (.A0(\cpu.ex.r_12[10] ),
    .A1(_03347_),
    .S(net564),
    .X(_00834_));
 sg13g2_mux2_1 _20495_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net832),
    .S(net564),
    .X(_00835_));
 sg13g2_mux2_1 _20496_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net439),
    .S(net564),
    .X(_00836_));
 sg13g2_mux2_1 _20497_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net443),
    .S(net564),
    .X(_00837_));
 sg13g2_mux2_1 _20498_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net442),
    .S(_03368_),
    .X(_00838_));
 sg13g2_mux2_1 _20499_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net829),
    .S(_03368_),
    .X(_00839_));
 sg13g2_mux2_1 _20500_ (.A0(\cpu.ex.r_12[1] ),
    .A1(_03355_),
    .S(net564),
    .X(_00840_));
 sg13g2_mux2_1 _20501_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net505),
    .S(net564),
    .X(_00841_));
 sg13g2_mux2_1 _20502_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net440),
    .S(net564),
    .X(_00842_));
 sg13g2_mux2_1 _20503_ (.A0(\cpu.ex.r_12[4] ),
    .A1(net504),
    .S(_03367_),
    .X(_00843_));
 sg13g2_mux2_1 _20504_ (.A0(\cpu.ex.r_12[5] ),
    .A1(_02879_),
    .S(_03367_),
    .X(_00844_));
 sg13g2_mux2_1 _20505_ (.A0(\cpu.ex.r_12[6] ),
    .A1(_02882_),
    .S(_03367_),
    .X(_00845_));
 sg13g2_mux2_1 _20506_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net711),
    .S(_03367_),
    .X(_00846_));
 sg13g2_mux2_1 _20507_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net833),
    .S(_03367_),
    .X(_00847_));
 sg13g2_buf_1 _20508_ (.A(net954),
    .X(_03369_));
 sg13g2_mux2_1 _20509_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net828),
    .S(_03367_),
    .X(_00848_));
 sg13g2_inv_1 _20510_ (.Y(_03370_),
    .A(net1077));
 sg13g2_nand2_1 _20511_ (.Y(_03371_),
    .A(_03370_),
    .B(net1003));
 sg13g2_nor2_1 _20512_ (.A(_03365_),
    .B(_03371_),
    .Y(_03372_));
 sg13g2_buf_2 _20513_ (.A(_03372_),
    .X(_03373_));
 sg13g2_buf_1 _20514_ (.A(_03373_),
    .X(_03374_));
 sg13g2_mux2_1 _20515_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net709),
    .S(net563),
    .X(_00849_));
 sg13g2_mux2_1 _20516_ (.A0(\cpu.ex.r_13[10] ),
    .A1(_03347_),
    .S(_03374_),
    .X(_00850_));
 sg13g2_mux2_1 _20517_ (.A0(\cpu.ex.r_13[11] ),
    .A1(net832),
    .S(net563),
    .X(_00851_));
 sg13g2_mux2_1 _20518_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net439),
    .S(net563),
    .X(_00852_));
 sg13g2_mux2_1 _20519_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net443),
    .S(net563),
    .X(_00853_));
 sg13g2_mux2_1 _20520_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net442),
    .S(net563),
    .X(_00854_));
 sg13g2_mux2_1 _20521_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net829),
    .S(_03374_),
    .X(_00855_));
 sg13g2_mux2_1 _20522_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net441),
    .S(net563),
    .X(_00856_));
 sg13g2_mux2_1 _20523_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net505),
    .S(net563),
    .X(_00857_));
 sg13g2_mux2_1 _20524_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net440),
    .S(net563),
    .X(_00858_));
 sg13g2_mux2_1 _20525_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net504),
    .S(_03373_),
    .X(_00859_));
 sg13g2_mux2_1 _20526_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_02879_),
    .S(_03373_),
    .X(_00860_));
 sg13g2_mux2_1 _20527_ (.A0(\cpu.ex.r_13[6] ),
    .A1(_02882_),
    .S(_03373_),
    .X(_00861_));
 sg13g2_mux2_1 _20528_ (.A0(\cpu.ex.r_13[7] ),
    .A1(net711),
    .S(_03373_),
    .X(_00862_));
 sg13g2_mux2_1 _20529_ (.A0(\cpu.ex.r_13[8] ),
    .A1(net833),
    .S(_03373_),
    .X(_00863_));
 sg13g2_mux2_1 _20530_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net828),
    .S(_03373_),
    .X(_00864_));
 sg13g2_nor2_1 _20531_ (.A(_03341_),
    .B(_03365_),
    .Y(_03375_));
 sg13g2_buf_2 _20532_ (.A(_03375_),
    .X(_03376_));
 sg13g2_buf_1 _20533_ (.A(_03376_),
    .X(_03377_));
 sg13g2_mux2_1 _20534_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net709),
    .S(net502),
    .X(_00865_));
 sg13g2_mux2_1 _20535_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net830),
    .S(net502),
    .X(_00866_));
 sg13g2_mux2_1 _20536_ (.A0(\cpu.ex.r_14[11] ),
    .A1(_02911_),
    .S(_03377_),
    .X(_00867_));
 sg13g2_mux2_1 _20537_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net439),
    .S(net502),
    .X(_00868_));
 sg13g2_mux2_1 _20538_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net443),
    .S(net502),
    .X(_00869_));
 sg13g2_mux2_1 _20539_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net442),
    .S(net502),
    .X(_00870_));
 sg13g2_mux2_1 _20540_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net829),
    .S(_03377_),
    .X(_00871_));
 sg13g2_mux2_1 _20541_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net441),
    .S(net502),
    .X(_00872_));
 sg13g2_mux2_1 _20542_ (.A0(\cpu.ex.r_14[2] ),
    .A1(net505),
    .S(net502),
    .X(_00873_));
 sg13g2_mux2_1 _20543_ (.A0(\cpu.ex.r_14[3] ),
    .A1(_03358_),
    .S(net502),
    .X(_00874_));
 sg13g2_mux2_1 _20544_ (.A0(\cpu.ex.r_14[4] ),
    .A1(_03359_),
    .S(_03376_),
    .X(_00875_));
 sg13g2_buf_1 _20545_ (.A(net566),
    .X(_03378_));
 sg13g2_mux2_1 _20546_ (.A0(\cpu.ex.r_14[5] ),
    .A1(net501),
    .S(_03376_),
    .X(_00876_));
 sg13g2_buf_1 _20547_ (.A(net1022),
    .X(_03379_));
 sg13g2_mux2_1 _20548_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net827),
    .S(_03376_),
    .X(_00877_));
 sg13g2_mux2_1 _20549_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net711),
    .S(_03376_),
    .X(_00878_));
 sg13g2_mux2_1 _20550_ (.A0(\cpu.ex.r_14[8] ),
    .A1(_02910_),
    .S(_03376_),
    .X(_00879_));
 sg13g2_mux2_1 _20551_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net828),
    .S(_03376_),
    .X(_00880_));
 sg13g2_nor2_1 _20552_ (.A(_09965_),
    .B(_03365_),
    .Y(_03380_));
 sg13g2_buf_2 _20553_ (.A(_03380_),
    .X(_03381_));
 sg13g2_buf_1 _20554_ (.A(_03381_),
    .X(_03382_));
 sg13g2_mux2_1 _20555_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net709),
    .S(net562),
    .X(_00881_));
 sg13g2_mux2_1 _20556_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net830),
    .S(net562),
    .X(_00882_));
 sg13g2_mux2_1 _20557_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net832),
    .S(net562),
    .X(_00883_));
 sg13g2_mux2_1 _20558_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net439),
    .S(net562),
    .X(_00884_));
 sg13g2_mux2_1 _20559_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net443),
    .S(net562),
    .X(_00885_));
 sg13g2_mux2_1 _20560_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net442),
    .S(net562),
    .X(_00886_));
 sg13g2_mux2_1 _20561_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net829),
    .S(_03382_),
    .X(_00887_));
 sg13g2_mux2_1 _20562_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net441),
    .S(net562),
    .X(_00888_));
 sg13g2_mux2_1 _20563_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net505),
    .S(_03382_),
    .X(_00889_));
 sg13g2_mux2_1 _20564_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net440),
    .S(net562),
    .X(_00890_));
 sg13g2_mux2_1 _20565_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net504),
    .S(_03381_),
    .X(_00891_));
 sg13g2_mux2_1 _20566_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net501),
    .S(_03381_),
    .X(_00892_));
 sg13g2_mux2_1 _20567_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net827),
    .S(_03381_),
    .X(_00893_));
 sg13g2_mux2_1 _20568_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net711),
    .S(_03381_),
    .X(_00894_));
 sg13g2_mux2_1 _20569_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net833),
    .S(_03381_),
    .X(_00895_));
 sg13g2_mux2_1 _20570_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net828),
    .S(_03381_),
    .X(_00896_));
 sg13g2_nor3_1 _20571_ (.A(net1077),
    .B(net1003),
    .C(_03343_),
    .Y(_03383_));
 sg13g2_buf_2 _20572_ (.A(_03383_),
    .X(_03384_));
 sg13g2_buf_1 _20573_ (.A(_03384_),
    .X(_03385_));
 sg13g2_mux2_1 _20574_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net709),
    .S(net500),
    .X(_00897_));
 sg13g2_mux2_1 _20575_ (.A0(\cpu.ex.r_8[10] ),
    .A1(net830),
    .S(_03385_),
    .X(_00898_));
 sg13g2_mux2_1 _20576_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net832),
    .S(net500),
    .X(_00899_));
 sg13g2_mux2_1 _20577_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net439),
    .S(net500),
    .X(_00900_));
 sg13g2_mux2_1 _20578_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net443),
    .S(net500),
    .X(_00901_));
 sg13g2_mux2_1 _20579_ (.A0(\cpu.ex.r_8[14] ),
    .A1(net442),
    .S(_03385_),
    .X(_00902_));
 sg13g2_mux2_1 _20580_ (.A0(\cpu.ex.r_8[15] ),
    .A1(_03354_),
    .S(net500),
    .X(_00903_));
 sg13g2_mux2_1 _20581_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net441),
    .S(net500),
    .X(_00904_));
 sg13g2_mux2_1 _20582_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net505),
    .S(net500),
    .X(_00905_));
 sg13g2_mux2_1 _20583_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net440),
    .S(net500),
    .X(_00906_));
 sg13g2_mux2_1 _20584_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net504),
    .S(_03384_),
    .X(_00907_));
 sg13g2_mux2_1 _20585_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net501),
    .S(_03384_),
    .X(_00908_));
 sg13g2_mux2_1 _20586_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net827),
    .S(_03384_),
    .X(_00909_));
 sg13g2_mux2_1 _20587_ (.A0(\cpu.ex.r_8[7] ),
    .A1(_02909_),
    .S(_03384_),
    .X(_00910_));
 sg13g2_mux2_1 _20588_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net833),
    .S(_03384_),
    .X(_00911_));
 sg13g2_mux2_1 _20589_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net828),
    .S(_03384_),
    .X(_00912_));
 sg13g2_nor2_1 _20590_ (.A(_03343_),
    .B(_03371_),
    .Y(_03386_));
 sg13g2_buf_2 _20591_ (.A(_03386_),
    .X(_03387_));
 sg13g2_buf_1 _20592_ (.A(_03387_),
    .X(_03388_));
 sg13g2_mux2_1 _20593_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net709),
    .S(net499),
    .X(_00913_));
 sg13g2_mux2_1 _20594_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net830),
    .S(net499),
    .X(_00914_));
 sg13g2_mux2_1 _20595_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net832),
    .S(net499),
    .X(_00915_));
 sg13g2_mux2_1 _20596_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net439),
    .S(net499),
    .X(_00916_));
 sg13g2_buf_1 _20597_ (.A(_10286_),
    .X(_03389_));
 sg13g2_mux2_1 _20598_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net498),
    .S(_03388_),
    .X(_00917_));
 sg13g2_buf_1 _20599_ (.A(net506),
    .X(_03390_));
 sg13g2_mux2_1 _20600_ (.A0(\cpu.ex.r_9[14] ),
    .A1(net438),
    .S(_03388_),
    .X(_00918_));
 sg13g2_mux2_1 _20601_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net829),
    .S(net499),
    .X(_00919_));
 sg13g2_mux2_1 _20602_ (.A0(\cpu.ex.r_9[1] ),
    .A1(_03355_),
    .S(net499),
    .X(_00920_));
 sg13g2_mux2_1 _20603_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net505),
    .S(net499),
    .X(_00921_));
 sg13g2_mux2_1 _20604_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net440),
    .S(net499),
    .X(_00922_));
 sg13g2_mux2_1 _20605_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net504),
    .S(_03387_),
    .X(_00923_));
 sg13g2_mux2_1 _20606_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net501),
    .S(_03387_),
    .X(_00924_));
 sg13g2_mux2_1 _20607_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net827),
    .S(_03387_),
    .X(_00925_));
 sg13g2_mux2_1 _20608_ (.A0(\cpu.ex.r_9[7] ),
    .A1(_02909_),
    .S(_03387_),
    .X(_00926_));
 sg13g2_mux2_1 _20609_ (.A0(\cpu.ex.r_9[8] ),
    .A1(_02910_),
    .S(_03387_),
    .X(_00927_));
 sg13g2_mux2_1 _20610_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net828),
    .S(_03387_),
    .X(_00928_));
 sg13g2_inv_1 _20611_ (.Y(_03391_),
    .A(\cpu.ex.r_cc ));
 sg13g2_inv_1 _20612_ (.Y(_03392_),
    .A(_11229_));
 sg13g2_nor2_1 _20613_ (.A(_10512_),
    .B(_03392_),
    .Y(_03393_));
 sg13g2_buf_1 _20614_ (.A(_03393_),
    .X(_03394_));
 sg13g2_nor2_1 _20615_ (.A(_11222_),
    .B(_03394_),
    .Y(_03395_));
 sg13g2_buf_1 _20616_ (.A(_03395_),
    .X(_03396_));
 sg13g2_nor2b_1 _20617_ (.A(_10899_),
    .B_N(_10901_),
    .Y(_03397_));
 sg13g2_buf_1 _20618_ (.A(_03397_),
    .X(_03398_));
 sg13g2_nand2_1 _20619_ (.Y(_03399_),
    .A(net241),
    .B(net231));
 sg13g2_buf_1 _20620_ (.A(_10859_),
    .X(_03400_));
 sg13g2_nor2_1 _20621_ (.A(_11514_),
    .B(net194),
    .Y(_03401_));
 sg13g2_buf_1 _20622_ (.A(_03400_),
    .X(_03402_));
 sg13g2_buf_1 _20623_ (.A(net294),
    .X(_03403_));
 sg13g2_a21oi_1 _20624_ (.A1(net230),
    .A2(_10874_),
    .Y(_03404_),
    .B1(_10875_));
 sg13g2_buf_1 _20625_ (.A(_03404_),
    .X(_03405_));
 sg13g2_mux2_1 _20626_ (.A0(_10770_),
    .A1(_10795_),
    .S(net336),
    .X(_03406_));
 sg13g2_buf_8 _20627_ (.A(_03406_),
    .X(_03407_));
 sg13g2_nor2_1 _20628_ (.A(_11271_),
    .B(net229),
    .Y(_03408_));
 sg13g2_or3_1 _20629_ (.A(net363),
    .B(_11558_),
    .C(_11082_),
    .X(_03409_));
 sg13g2_nand3_1 _20630_ (.B(net363),
    .C(_11179_),
    .A(_00297_),
    .Y(_03410_));
 sg13g2_a22oi_1 _20631_ (.Y(_03411_),
    .B1(_03409_),
    .B2(_03410_),
    .A2(_03407_),
    .A1(_11271_));
 sg13g2_nand2_1 _20632_ (.Y(_03412_),
    .A(_10981_),
    .B(_10487_));
 sg13g2_o21ai_1 _20633_ (.B1(_03412_),
    .Y(_03413_),
    .A1(_03408_),
    .A2(_03411_));
 sg13g2_nand2b_1 _20634_ (.Y(_03414_),
    .B(_11123_),
    .A_N(_10981_));
 sg13g2_nor2_1 _20635_ (.A(_11565_),
    .B(_10771_),
    .Y(_03415_));
 sg13g2_nand2_1 _20636_ (.Y(_03416_),
    .A(_10513_),
    .B(_03415_));
 sg13g2_o21ai_1 _20637_ (.B1(_03415_),
    .Y(_03417_),
    .A1(_08557_),
    .A2(_10520_));
 sg13g2_o21ai_1 _20638_ (.B1(_03417_),
    .Y(_03418_),
    .A1(_08615_),
    .A2(_03416_));
 sg13g2_a21o_1 _20639_ (.A2(_10822_),
    .A1(_10525_),
    .B1(_03418_),
    .X(_03419_));
 sg13g2_buf_2 _20640_ (.A(_03419_),
    .X(_03420_));
 sg13g2_nand4_1 _20641_ (.B(_10656_),
    .C(_10678_),
    .A(_10652_),
    .Y(_03421_),
    .D(_11171_));
 sg13g2_nand2_1 _20642_ (.Y(_03422_),
    .A(_03420_),
    .B(_03421_));
 sg13g2_o21ai_1 _20643_ (.B1(net334),
    .Y(_03423_),
    .A1(_03420_),
    .A2(_03421_));
 sg13g2_mux2_1 _20644_ (.A0(_10528_),
    .A1(_11558_),
    .S(net336),
    .X(_03424_));
 sg13g2_buf_2 _20645_ (.A(_03424_),
    .X(_03425_));
 sg13g2_a22oi_1 _20646_ (.Y(_03426_),
    .B1(_03425_),
    .B2(net333),
    .A2(net229),
    .A1(_11271_));
 sg13g2_nand4_1 _20647_ (.B(_03423_),
    .C(_03426_),
    .A(_03422_),
    .Y(_03427_),
    .D(_03412_));
 sg13g2_nand3_1 _20648_ (.B(_03414_),
    .C(_03427_),
    .A(_03413_),
    .Y(_03428_));
 sg13g2_buf_1 _20649_ (.A(_03428_),
    .X(_03429_));
 sg13g2_nor2_1 _20650_ (.A(_00296_),
    .B(net294),
    .Y(_03430_));
 sg13g2_a21oi_1 _20651_ (.A1(net294),
    .A2(_10942_),
    .Y(_03431_),
    .B1(_03430_));
 sg13g2_buf_2 _20652_ (.A(_03431_),
    .X(_03432_));
 sg13g2_nor2_1 _20653_ (.A(_03432_),
    .B(net295),
    .Y(_03433_));
 sg13g2_nor2_1 _20654_ (.A(_10999_),
    .B(_03433_),
    .Y(_03434_));
 sg13g2_buf_1 _20655_ (.A(_03434_),
    .X(_03435_));
 sg13g2_nor3_1 _20656_ (.A(_10944_),
    .B(_10999_),
    .C(_11127_),
    .Y(_03436_));
 sg13g2_o21ai_1 _20657_ (.B1(_10999_),
    .Y(_03437_),
    .A1(_10944_),
    .A2(_11127_));
 sg13g2_o21ai_1 _20658_ (.B1(_03437_),
    .Y(_03438_),
    .A1(_10435_),
    .A2(_03436_));
 sg13g2_nand4_1 _20659_ (.B(_03414_),
    .C(_03427_),
    .A(_03413_),
    .Y(_03439_),
    .D(_03438_));
 sg13g2_buf_2 _20660_ (.A(_03439_),
    .X(_03440_));
 sg13g2_nor2_1 _20661_ (.A(_10435_),
    .B(_03436_),
    .Y(_03441_));
 sg13g2_a21oi_1 _20662_ (.A1(_03433_),
    .A2(_03438_),
    .Y(_03442_),
    .B1(_03441_));
 sg13g2_buf_2 _20663_ (.A(_03442_),
    .X(_03443_));
 sg13g2_nand2_1 _20664_ (.Y(_03444_),
    .A(net182),
    .B(_11166_));
 sg13g2_a221oi_1 _20665_ (.B2(_03443_),
    .C1(_03444_),
    .B1(_03440_),
    .A1(net102),
    .Y(_03445_),
    .A2(_03435_));
 sg13g2_nand2_1 _20666_ (.Y(_03446_),
    .A(_11166_),
    .B(_10713_));
 sg13g2_a221oi_1 _20667_ (.B2(_03443_),
    .C1(_03446_),
    .B1(_03440_),
    .A1(net102),
    .Y(_03447_),
    .A2(_03435_));
 sg13g2_nand2_1 _20668_ (.Y(_03448_),
    .A(net182),
    .B(_10962_));
 sg13g2_a221oi_1 _20669_ (.B2(_03443_),
    .C1(_03448_),
    .B1(_03440_),
    .A1(net102),
    .Y(_03449_),
    .A2(_03435_));
 sg13g2_nand2_1 _20670_ (.Y(_03450_),
    .A(_10713_),
    .B(_10962_));
 sg13g2_a221oi_1 _20671_ (.B2(_03443_),
    .C1(_03450_),
    .B1(_03440_),
    .A1(_03429_),
    .Y(_03451_),
    .A2(_03435_));
 sg13g2_nor4_1 _20672_ (.A(_03445_),
    .B(_03447_),
    .C(_03449_),
    .D(_03451_),
    .Y(_03452_));
 sg13g2_buf_1 _20673_ (.A(_10713_),
    .X(_03453_));
 sg13g2_nor2_1 _20674_ (.A(_00294_),
    .B(net230),
    .Y(_03454_));
 sg13g2_a21oi_1 _20675_ (.A1(net230),
    .A2(_10960_),
    .Y(_03455_),
    .B1(_03454_));
 sg13g2_buf_1 _20676_ (.A(_03455_),
    .X(_03456_));
 sg13g2_nor2_1 _20677_ (.A(net240),
    .B(_03456_),
    .Y(_03457_));
 sg13g2_nand2_1 _20678_ (.Y(_03458_),
    .A(net182),
    .B(_03457_));
 sg13g2_o21ai_1 _20679_ (.B1(_03458_),
    .Y(_03459_),
    .A1(net240),
    .A2(_03450_));
 sg13g2_a21oi_1 _20680_ (.A1(_10116_),
    .A2(_03453_),
    .Y(_03460_),
    .B1(_03459_));
 sg13g2_nand2_1 _20681_ (.Y(_03461_),
    .A(_10526_),
    .B(_10646_));
 sg13g2_o21ai_1 _20682_ (.B1(_03461_),
    .Y(_03462_),
    .A1(_00291_),
    .A2(net230));
 sg13g2_buf_1 _20683_ (.A(_03462_),
    .X(_03463_));
 sg13g2_buf_1 _20684_ (.A(_03463_),
    .X(_03464_));
 sg13g2_inv_1 _20685_ (.Y(_03465_),
    .A(_00290_));
 sg13g2_nor2_1 _20686_ (.A(net363),
    .B(_10765_),
    .Y(_03466_));
 sg13g2_a21oi_1 _20687_ (.A1(_03465_),
    .A2(net363),
    .Y(_03467_),
    .B1(_03466_));
 sg13g2_buf_2 _20688_ (.A(_03467_),
    .X(_03468_));
 sg13g2_nand2_1 _20689_ (.Y(_03469_),
    .A(net209),
    .B(_03468_));
 sg13g2_buf_1 _20690_ (.A(_03469_),
    .X(_03470_));
 sg13g2_mux2_1 _20691_ (.A0(_10718_),
    .A1(_10742_),
    .S(net294),
    .X(_03471_));
 sg13g2_buf_1 _20692_ (.A(_03471_),
    .X(_03472_));
 sg13g2_buf_1 _20693_ (.A(_03472_),
    .X(_03473_));
 sg13g2_inv_1 _20694_ (.Y(_03474_),
    .A(net172));
 sg13g2_nand2_1 _20695_ (.Y(_03475_),
    .A(net234),
    .B(_03474_));
 sg13g2_nand3_1 _20696_ (.B(_03470_),
    .C(_03475_),
    .A(net149),
    .Y(_03476_));
 sg13g2_nand3_1 _20697_ (.B(_03470_),
    .C(_03475_),
    .A(net207),
    .Y(_03477_));
 sg13g2_a22oi_1 _20698_ (.Y(_03478_),
    .B1(_03476_),
    .B2(_03477_),
    .A2(_03460_),
    .A1(_03452_));
 sg13g2_buf_1 _20699_ (.A(_03478_),
    .X(_03479_));
 sg13g2_nand4_1 _20700_ (.B(net149),
    .C(_03470_),
    .A(net205),
    .Y(_03480_),
    .D(net172));
 sg13g2_nand4_1 _20701_ (.B(net205),
    .C(_03470_),
    .A(net207),
    .Y(_03481_),
    .D(net172));
 sg13g2_nand3_1 _20702_ (.B(net149),
    .C(_03470_),
    .A(net207),
    .Y(_03482_));
 sg13g2_nand3_1 _20703_ (.B(_03481_),
    .C(_03482_),
    .A(_03480_),
    .Y(_03483_));
 sg13g2_buf_1 _20704_ (.A(_03483_),
    .X(_03484_));
 sg13g2_nor2_2 _20705_ (.A(net209),
    .B(_03468_),
    .Y(_03485_));
 sg13g2_nor3_1 _20706_ (.A(_03479_),
    .B(_03484_),
    .C(_03485_),
    .Y(_03486_));
 sg13g2_nor2_1 _20707_ (.A(net179),
    .B(_03485_),
    .Y(_03487_));
 sg13g2_nor2_1 _20708_ (.A(_03479_),
    .B(_03484_),
    .Y(_03488_));
 sg13g2_buf_1 _20709_ (.A(_10877_),
    .X(_03489_));
 sg13g2_nor2_1 _20710_ (.A(net179),
    .B(net193),
    .Y(_03490_));
 sg13g2_a221oi_1 _20711_ (.B2(_03488_),
    .C1(_03490_),
    .B1(_03487_),
    .A1(_03405_),
    .Y(_03491_),
    .A2(_03486_));
 sg13g2_buf_1 _20712_ (.A(_03491_),
    .X(_03492_));
 sg13g2_a21oi_1 _20713_ (.A1(net230),
    .A2(_10922_),
    .Y(_03493_),
    .B1(_10923_));
 sg13g2_buf_1 _20714_ (.A(_03493_),
    .X(_03494_));
 sg13g2_nand2_1 _20715_ (.Y(_03495_),
    .A(net199),
    .B(net171));
 sg13g2_nor2_2 _20716_ (.A(net199),
    .B(net171),
    .Y(_03496_));
 sg13g2_a221oi_1 _20717_ (.B2(_03495_),
    .C1(_03496_),
    .B1(_03492_),
    .A1(net151),
    .Y(_03497_),
    .A2(net173));
 sg13g2_buf_1 _20718_ (.A(net239),
    .X(_03498_));
 sg13g2_nand2_1 _20719_ (.Y(_03499_),
    .A(_10275_),
    .B(net192));
 sg13g2_o21ai_1 _20720_ (.B1(_03499_),
    .Y(_03500_),
    .A1(_03401_),
    .A2(_03497_));
 sg13g2_a21o_1 _20721_ (.A2(_03500_),
    .A1(_03399_),
    .B1(_08922_),
    .X(_03501_));
 sg13g2_nand2_1 _20722_ (.Y(_03502_),
    .A(net241),
    .B(net192));
 sg13g2_nor2_1 _20723_ (.A(_00295_),
    .B(net230),
    .Y(_03503_));
 sg13g2_a21oi_1 _20724_ (.A1(net230),
    .A2(_10997_),
    .Y(_03504_),
    .B1(_03503_));
 sg13g2_buf_1 _20725_ (.A(_03504_),
    .X(_03505_));
 sg13g2_nor2_1 _20726_ (.A(_11150_),
    .B(net148),
    .Y(_03506_));
 sg13g2_buf_2 _20727_ (.A(_03506_),
    .X(_03507_));
 sg13g2_a22oi_1 _20728_ (.Y(_03508_),
    .B1(_11077_),
    .B2(_11081_),
    .A2(_10611_),
    .A1(_10541_));
 sg13g2_a21oi_1 _20729_ (.A1(_11077_),
    .A2(_11081_),
    .Y(_03509_),
    .B1(_10528_));
 sg13g2_mux2_1 _20730_ (.A0(_03508_),
    .A1(_03509_),
    .S(_10768_),
    .X(_03510_));
 sg13g2_a21o_1 _20731_ (.A2(_10793_),
    .A1(net525),
    .B1(_10794_),
    .X(_03511_));
 sg13g2_mux2_1 _20732_ (.A0(_00191_),
    .A1(_03511_),
    .S(net294),
    .X(_03512_));
 sg13g2_buf_2 _20733_ (.A(_03512_),
    .X(_03513_));
 sg13g2_o21ai_1 _20734_ (.B1(_03513_),
    .Y(_03514_),
    .A1(_11271_),
    .A2(_03510_));
 sg13g2_nand2_1 _20735_ (.Y(_03515_),
    .A(_11271_),
    .B(_03510_));
 sg13g2_a22oi_1 _20736_ (.Y(_03516_),
    .B1(_03514_),
    .B2(_03515_),
    .A2(_11123_),
    .A1(_10981_));
 sg13g2_nand2b_1 _20737_ (.Y(_03517_),
    .B(_10487_),
    .A_N(_10981_));
 sg13g2_nand2_1 _20738_ (.Y(_03518_),
    .A(_10981_),
    .B(_11123_));
 sg13g2_nand3_1 _20739_ (.B(_10656_),
    .C(_10678_),
    .A(_10652_),
    .Y(_03519_));
 sg13g2_buf_1 _20740_ (.A(_03519_),
    .X(_03520_));
 sg13g2_nand3_1 _20741_ (.B(_11171_),
    .C(_03420_),
    .A(_03520_),
    .Y(_03521_));
 sg13g2_nor2_1 _20742_ (.A(net335),
    .B(_11054_),
    .Y(_03522_));
 sg13g2_buf_1 _20743_ (.A(_03522_),
    .X(_03523_));
 sg13g2_a22oi_1 _20744_ (.Y(_03524_),
    .B1(_03523_),
    .B2(_03520_),
    .A2(_03420_),
    .A1(_11173_));
 sg13g2_a22oi_1 _20745_ (.Y(_03525_),
    .B1(_03425_),
    .B2(_11179_),
    .A2(net229),
    .A1(_11117_));
 sg13g2_nand4_1 _20746_ (.B(_03521_),
    .C(_03524_),
    .A(_03518_),
    .Y(_03526_),
    .D(_03525_));
 sg13g2_nand3b_1 _20747_ (.B(_03517_),
    .C(_03526_),
    .Y(_03527_),
    .A_N(_03516_));
 sg13g2_buf_1 _20748_ (.A(_03527_),
    .X(_03528_));
 sg13g2_buf_1 _20749_ (.A(_10944_),
    .X(_03529_));
 sg13g2_nand2_1 _20750_ (.Y(_03530_),
    .A(net191),
    .B(net295));
 sg13g2_nand2_1 _20751_ (.Y(_03531_),
    .A(_03432_),
    .B(net236));
 sg13g2_inv_1 _20752_ (.Y(_03532_),
    .A(_03531_));
 sg13g2_a221oi_1 _20753_ (.B2(_03530_),
    .C1(_03532_),
    .B1(_03528_),
    .A1(_11150_),
    .Y(_03533_),
    .A2(net148));
 sg13g2_buf_1 _20754_ (.A(_03533_),
    .X(_03534_));
 sg13g2_inv_1 _20755_ (.Y(_03535_),
    .A(_10711_));
 sg13g2_mux2_1 _20756_ (.A0(_00293_),
    .A1(_03535_),
    .S(net336),
    .X(_03536_));
 sg13g2_buf_2 _20757_ (.A(_03536_),
    .X(_03537_));
 sg13g2_nor3_1 _20758_ (.A(_10067_),
    .B(_10108_),
    .C(_03537_),
    .Y(_03538_));
 sg13g2_buf_2 _20759_ (.A(_03538_),
    .X(_03539_));
 sg13g2_nand2_1 _20760_ (.Y(_03540_),
    .A(_03472_),
    .B(_03539_));
 sg13g2_o21ai_1 _20761_ (.B1(net296),
    .Y(_03541_),
    .A1(_03472_),
    .A2(_03539_));
 sg13g2_or2_1 _20762_ (.X(_03542_),
    .B(_03472_),
    .A(net296));
 sg13g2_buf_1 _20763_ (.A(_03542_),
    .X(_03543_));
 sg13g2_o21ai_1 _20764_ (.B1(_03537_),
    .Y(_03544_),
    .A1(_10067_),
    .A2(_10108_));
 sg13g2_buf_2 _20765_ (.A(_03544_),
    .X(_03545_));
 sg13g2_a21oi_1 _20766_ (.A1(_03543_),
    .A2(_03545_),
    .Y(_03546_),
    .B1(_10183_));
 sg13g2_and3_1 _20767_ (.X(_03547_),
    .A(_03540_),
    .B(_03541_),
    .C(_03546_));
 sg13g2_buf_1 _20768_ (.A(_03547_),
    .X(_03548_));
 sg13g2_a21oi_1 _20769_ (.A1(_03543_),
    .A2(_03545_),
    .Y(_03549_),
    .B1(_03463_));
 sg13g2_and3_1 _20770_ (.X(_03550_),
    .A(_03540_),
    .B(_03541_),
    .C(_03549_));
 sg13g2_buf_1 _20771_ (.A(_03550_),
    .X(_03551_));
 sg13g2_nand2_1 _20772_ (.Y(_03552_),
    .A(_11166_),
    .B(_03456_));
 sg13g2_or2_1 _20773_ (.X(_03553_),
    .B(_03463_),
    .A(_10183_));
 sg13g2_buf_1 _20774_ (.A(_03553_),
    .X(_03554_));
 sg13g2_nand2_1 _20775_ (.Y(_03555_),
    .A(_03552_),
    .B(_03554_));
 sg13g2_nor4_1 _20776_ (.A(_03468_),
    .B(_03548_),
    .C(_03551_),
    .D(_03555_),
    .Y(_03556_));
 sg13g2_o21ai_1 _20777_ (.B1(_03556_),
    .Y(_03557_),
    .A1(_03507_),
    .A2(_03534_));
 sg13g2_nor4_1 _20778_ (.A(_10193_),
    .B(_03548_),
    .C(_03551_),
    .D(_03555_),
    .Y(_03558_));
 sg13g2_o21ai_1 _20779_ (.B1(_03558_),
    .Y(_03559_),
    .A1(_03507_),
    .A2(_03534_));
 sg13g2_a21o_1 _20780_ (.A2(net363),
    .A1(_03465_),
    .B1(_03466_),
    .X(_03560_));
 sg13g2_buf_2 _20781_ (.A(_03560_),
    .X(_03561_));
 sg13g2_nor2_1 _20782_ (.A(net172),
    .B(_03539_),
    .Y(_03562_));
 sg13g2_a21oi_1 _20783_ (.A1(_03472_),
    .A2(_03539_),
    .Y(_03563_),
    .B1(net234));
 sg13g2_o21ai_1 _20784_ (.B1(_03549_),
    .Y(_03564_),
    .A1(_03562_),
    .A2(_03563_));
 sg13g2_nand2_1 _20785_ (.Y(_03565_),
    .A(_03561_),
    .B(_03564_));
 sg13g2_nand2_1 _20786_ (.Y(_03566_),
    .A(_10154_),
    .B(_03564_));
 sg13g2_and2_1 _20787_ (.A(_10402_),
    .B(_10962_),
    .X(_03567_));
 sg13g2_buf_1 _20788_ (.A(_03567_),
    .X(_03568_));
 sg13g2_nand3_1 _20789_ (.B(_03545_),
    .C(_03568_),
    .A(_03543_),
    .Y(_03569_));
 sg13g2_o21ai_1 _20790_ (.B1(_10183_),
    .Y(_03570_),
    .A1(net149),
    .A2(_03568_));
 sg13g2_nand4_1 _20791_ (.B(_03541_),
    .C(_03569_),
    .A(_03540_),
    .Y(_03571_),
    .D(_03570_));
 sg13g2_nand2_1 _20792_ (.Y(_03572_),
    .A(_03571_),
    .B(_03554_));
 sg13g2_a21o_1 _20793_ (.A2(_03566_),
    .A1(_03565_),
    .B1(_03572_),
    .X(_03573_));
 sg13g2_nand2_1 _20794_ (.Y(_03574_),
    .A(net209),
    .B(_03561_));
 sg13g2_and4_1 _20795_ (.A(_03557_),
    .B(_03559_),
    .C(_03573_),
    .D(_03574_),
    .X(_03575_));
 sg13g2_buf_2 _20796_ (.A(_03575_),
    .X(_03576_));
 sg13g2_nor2_1 _20797_ (.A(_11476_),
    .B(_03405_),
    .Y(_03577_));
 sg13g2_buf_1 _20798_ (.A(_03577_),
    .X(_03578_));
 sg13g2_nor2_1 _20799_ (.A(_11184_),
    .B(net171),
    .Y(_03579_));
 sg13g2_nor2_1 _20800_ (.A(_03578_),
    .B(_03579_),
    .Y(_03580_));
 sg13g2_nor2_2 _20801_ (.A(net200),
    .B(_10877_),
    .Y(_03581_));
 sg13g2_o21ai_1 _20802_ (.B1(_11184_),
    .Y(_03582_),
    .A1(net171),
    .A2(_03581_));
 sg13g2_nand2_1 _20803_ (.Y(_03583_),
    .A(net171),
    .B(_03581_));
 sg13g2_nand2_1 _20804_ (.Y(_03584_),
    .A(_03582_),
    .B(_03583_));
 sg13g2_a21oi_1 _20805_ (.A1(_03576_),
    .A2(_03580_),
    .Y(_03585_),
    .B1(_03584_));
 sg13g2_nor3_1 _20806_ (.A(net173),
    .B(_03578_),
    .C(_03579_),
    .Y(_03586_));
 sg13g2_nand2_1 _20807_ (.Y(_03587_),
    .A(_03576_),
    .B(_03586_));
 sg13g2_a21oi_1 _20808_ (.A1(_03582_),
    .A2(_03583_),
    .Y(_03588_),
    .B1(net173));
 sg13g2_nor2_1 _20809_ (.A(_11514_),
    .B(_03588_),
    .Y(_03589_));
 sg13g2_a22oi_1 _20810_ (.Y(_03590_),
    .B1(_03587_),
    .B2(_03589_),
    .A2(_03585_),
    .A1(net173));
 sg13g2_nor2_1 _20811_ (.A(_10230_),
    .B(net239),
    .Y(_03591_));
 sg13g2_a21oi_1 _20812_ (.A1(_03502_),
    .A2(_03590_),
    .Y(_03592_),
    .B1(_03591_));
 sg13g2_a21oi_1 _20813_ (.A1(_08922_),
    .A2(_03592_),
    .Y(_03593_),
    .B1(net36));
 sg13g2_a22oi_1 _20814_ (.Y(_00929_),
    .B1(_03501_),
    .B2(_03593_),
    .A2(net36),
    .A1(_03391_));
 sg13g2_nand4_1 _20815_ (.B(net1003),
    .C(_09960_),
    .A(net1077),
    .Y(_03594_),
    .D(_09987_));
 sg13g2_nor2_1 _20816_ (.A(_08514_),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_buf_2 _20817_ (.A(_03595_),
    .X(_03596_));
 sg13g2_buf_1 _20818_ (.A(_03596_),
    .X(_03597_));
 sg13g2_mux2_1 _20819_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(net441),
    .S(net561),
    .X(_00931_));
 sg13g2_mux2_1 _20820_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(net832),
    .S(net561),
    .X(_00932_));
 sg13g2_buf_1 _20821_ (.A(net576),
    .X(_03598_));
 sg13g2_mux2_1 _20822_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(net497),
    .S(net561),
    .X(_00933_));
 sg13g2_mux2_1 _20823_ (.A0(\cpu.ex.r_epc[13] ),
    .A1(net498),
    .S(net561),
    .X(_00934_));
 sg13g2_mux2_1 _20824_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(net438),
    .S(_03597_),
    .X(_00935_));
 sg13g2_mux2_1 _20825_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(net829),
    .S(_03597_),
    .X(_00936_));
 sg13g2_mux2_1 _20826_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(_03357_),
    .S(net561),
    .X(_00937_));
 sg13g2_mux2_1 _20827_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(_03358_),
    .S(net561),
    .X(_00938_));
 sg13g2_mux2_1 _20828_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(net504),
    .S(net561),
    .X(_00939_));
 sg13g2_mux2_1 _20829_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(net501),
    .S(net561),
    .X(_00940_));
 sg13g2_mux2_1 _20830_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net827),
    .S(_03596_),
    .X(_00941_));
 sg13g2_mux2_1 _20831_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(net711),
    .S(_03596_),
    .X(_00942_));
 sg13g2_mux2_1 _20832_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net833),
    .S(_03596_),
    .X(_00943_));
 sg13g2_mux2_1 _20833_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(net828),
    .S(_03596_),
    .X(_00944_));
 sg13g2_mux2_1 _20834_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(net830),
    .S(_03596_),
    .X(_00945_));
 sg13g2_nand4_1 _20835_ (.B(net1003),
    .C(_09960_),
    .A(_03370_),
    .Y(_03599_),
    .D(_09987_));
 sg13g2_buf_1 _20836_ (.A(_03599_),
    .X(_03600_));
 sg13g2_buf_1 _20837_ (.A(_03600_),
    .X(_03601_));
 sg13g2_buf_1 _20838_ (.A(_03600_),
    .X(_03602_));
 sg13g2_nand2_1 _20839_ (.Y(_03603_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net633));
 sg13g2_o21ai_1 _20840_ (.B1(_03603_),
    .Y(_00951_),
    .A1(_09882_),
    .A2(net634));
 sg13g2_mux2_1 _20841_ (.A0(_02876_),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net634),
    .X(_00952_));
 sg13g2_buf_1 _20842_ (.A(_03348_),
    .X(_03604_));
 sg13g2_mux2_1 _20843_ (.A0(_03604_),
    .A1(\cpu.ex.r_lr[12] ),
    .S(net634),
    .X(_00953_));
 sg13g2_buf_1 _20844_ (.A(net507),
    .X(_03605_));
 sg13g2_mux2_1 _20845_ (.A0(net436),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net634),
    .X(_00954_));
 sg13g2_buf_1 _20846_ (.A(net506),
    .X(_03606_));
 sg13g2_mux2_1 _20847_ (.A0(net435),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net633),
    .X(_00955_));
 sg13g2_buf_1 _20848_ (.A(net679),
    .X(_03607_));
 sg13g2_nand2_1 _20849_ (.Y(_03608_),
    .A(\cpu.ex.r_lr[15] ),
    .B(net633));
 sg13g2_o21ai_1 _20850_ (.B1(_03608_),
    .Y(_00956_),
    .A1(net560),
    .A2(_03601_));
 sg13g2_buf_2 _20851_ (.A(_09470_),
    .X(_03609_));
 sg13g2_nand2_1 _20852_ (.Y(_03610_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net633));
 sg13g2_o21ai_1 _20853_ (.B1(_03610_),
    .Y(_00957_),
    .A1(_03609_),
    .A2(net634));
 sg13g2_nand2_1 _20854_ (.Y(_03611_),
    .A(\cpu.ex.r_lr[3] ),
    .B(net633));
 sg13g2_o21ai_1 _20855_ (.B1(_03611_),
    .Y(_00958_),
    .A1(net760),
    .A2(net634));
 sg13g2_buf_2 _20856_ (.A(_11607_),
    .X(_03612_));
 sg13g2_buf_1 _20857_ (.A(net708),
    .X(_03613_));
 sg13g2_nand2_1 _20858_ (.Y(_03614_),
    .A(\cpu.ex.r_lr[4] ),
    .B(_03602_));
 sg13g2_o21ai_1 _20859_ (.B1(_03614_),
    .Y(_00959_),
    .A1(net631),
    .A2(_03601_));
 sg13g2_nand2_1 _20860_ (.Y(_03615_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03600_));
 sg13g2_o21ai_1 _20861_ (.B1(_03615_),
    .Y(_00960_),
    .A1(net637),
    .A2(net634));
 sg13g2_nand2_1 _20862_ (.Y(_03616_),
    .A(\cpu.ex.r_lr[6] ),
    .B(_03600_));
 sg13g2_o21ai_1 _20863_ (.B1(_03616_),
    .Y(_00961_),
    .A1(net636),
    .A2(net634));
 sg13g2_mux2_1 _20864_ (.A0(net714),
    .A1(\cpu.ex.r_lr[7] ),
    .S(net633),
    .X(_00962_));
 sg13g2_mux2_1 _20865_ (.A0(net842),
    .A1(\cpu.ex.r_lr[8] ),
    .S(net633),
    .X(_00963_));
 sg13g2_mux2_1 _20866_ (.A0(net841),
    .A1(\cpu.ex.r_lr[9] ),
    .S(net633),
    .X(_00964_));
 sg13g2_mux2_1 _20867_ (.A0(_02874_),
    .A1(\cpu.ex.r_lr[10] ),
    .S(_03602_),
    .X(_00965_));
 sg13g2_buf_1 _20868_ (.A(net335),
    .X(_03617_));
 sg13g2_buf_1 _20869_ (.A(net33),
    .X(_03618_));
 sg13g2_nor2_1 _20870_ (.A(_03617_),
    .B(net31),
    .Y(_03619_));
 sg13g2_xnor2_1 _20871_ (.Y(_03620_),
    .A(net80),
    .B(_03619_));
 sg13g2_inv_1 _20872_ (.Y(_03621_),
    .A(net831));
 sg13g2_buf_1 _20873_ (.A(_09971_),
    .X(_03622_));
 sg13g2_mux2_1 _20874_ (.A0(_11539_),
    .A1(_11543_),
    .S(_10275_),
    .X(_03623_));
 sg13g2_a22oi_1 _20875_ (.Y(_03624_),
    .B1(_03623_),
    .B2(_11517_),
    .A2(_10229_),
    .A1(_11238_));
 sg13g2_nor2_1 _20876_ (.A(net151),
    .B(_03624_),
    .Y(_03625_));
 sg13g2_and4_1 _20877_ (.A(_11539_),
    .B(net241),
    .C(_10272_),
    .D(_11518_),
    .X(_03626_));
 sg13g2_o21ai_1 _20878_ (.B1(_11191_),
    .Y(_03627_),
    .A1(_03625_),
    .A2(_03626_));
 sg13g2_nor3_1 _20879_ (.A(_11517_),
    .B(_11539_),
    .C(net398),
    .Y(_03628_));
 sg13g2_o21ai_1 _20880_ (.B1(_03628_),
    .Y(_03629_),
    .A1(_10278_),
    .A2(_11003_));
 sg13g2_a221oi_1 _20881_ (.B2(_03629_),
    .C1(_11511_),
    .B1(_03627_),
    .A1(_11400_),
    .Y(_03630_),
    .A2(_11407_));
 sg13g2_buf_1 _20882_ (.A(_03630_),
    .X(_03631_));
 sg13g2_nand2_1 _20883_ (.Y(_03632_),
    .A(_03627_),
    .B(_03629_));
 sg13g2_nand2_1 _20884_ (.Y(_03633_),
    .A(_11505_),
    .B(_03632_));
 sg13g2_nand2_1 _20885_ (.Y(_03634_),
    .A(_11539_),
    .B(_10275_));
 sg13g2_nor2_1 _20886_ (.A(_11539_),
    .B(_10275_),
    .Y(_03635_));
 sg13g2_a21oi_1 _20887_ (.A1(_11534_),
    .A2(_03634_),
    .Y(_03636_),
    .B1(_03635_));
 sg13g2_or2_1 _20888_ (.X(_03637_),
    .B(_03636_),
    .A(net361));
 sg13g2_a21oi_1 _20889_ (.A1(_03633_),
    .A2(_03637_),
    .Y(_03638_),
    .B1(net80));
 sg13g2_or3_1 _20890_ (.A(_11545_),
    .B(_03631_),
    .C(_03638_),
    .X(_03639_));
 sg13g2_nand3b_1 _20891_ (.B(_03634_),
    .C(_11525_),
    .Y(_03640_),
    .A_N(_03635_));
 sg13g2_o21ai_1 _20892_ (.B1(_03640_),
    .Y(_03641_),
    .A1(net151),
    .A2(_03624_));
 sg13g2_o21ai_1 _20893_ (.B1(_03641_),
    .Y(_03642_),
    .A1(_11502_),
    .A2(_11503_));
 sg13g2_a21oi_1 _20894_ (.A1(_03636_),
    .A2(_03642_),
    .Y(_03643_),
    .B1(_11256_));
 sg13g2_or2_1 _20895_ (.X(_03644_),
    .B(_03643_),
    .A(_03631_));
 sg13g2_buf_1 _20896_ (.A(_03644_),
    .X(_03645_));
 sg13g2_o21ai_1 _20897_ (.B1(_11545_),
    .Y(_03646_),
    .A1(_11240_),
    .A2(_03645_));
 sg13g2_nand3_1 _20898_ (.B(_03639_),
    .C(_03646_),
    .A(_11196_),
    .Y(_03647_));
 sg13g2_a21oi_1 _20899_ (.A1(\cpu.ex.r_mult[16] ),
    .A2(_11199_),
    .Y(_03648_),
    .B1(net523));
 sg13g2_nor3_1 _20900_ (.A(\cpu.ex.r_cc ),
    .B(net559),
    .C(_09972_),
    .Y(_03649_));
 sg13g2_a221oi_1 _20901_ (.B2(_03648_),
    .C1(_03649_),
    .B1(_03647_),
    .A1(_03621_),
    .Y(_03650_),
    .A2(net559));
 sg13g2_a21o_1 _20902_ (.A2(_03620_),
    .A1(_11494_),
    .B1(_03650_),
    .X(_00966_));
 sg13g2_inv_1 _20903_ (.Y(_03651_),
    .A(\cpu.ex.r_mult[17] ));
 sg13g2_and2_1 _20904_ (.A(net463),
    .B(_11199_),
    .X(_03652_));
 sg13g2_buf_2 _20905_ (.A(_03652_),
    .X(_03653_));
 sg13g2_nor2_1 _20906_ (.A(_00309_),
    .B(_10197_),
    .Y(_03654_));
 sg13g2_nand2_1 _20907_ (.Y(_03655_),
    .A(_11256_),
    .B(net292));
 sg13g2_buf_1 _20908_ (.A(_11055_),
    .X(_03656_));
 sg13g2_xnor2_1 _20909_ (.Y(_03657_),
    .A(_03655_),
    .B(net282));
 sg13g2_nor2_1 _20910_ (.A(net33),
    .B(_03657_),
    .Y(_03658_));
 sg13g2_xor2_1 _20911_ (.B(_03658_),
    .A(_03654_),
    .X(_03659_));
 sg13g2_nor2b_1 _20912_ (.A(_00309_),
    .B_N(_11545_),
    .Y(_03660_));
 sg13g2_and2_1 _20913_ (.A(_03645_),
    .B(_03660_),
    .X(_03661_));
 sg13g2_buf_1 _20914_ (.A(_03661_),
    .X(_03662_));
 sg13g2_a21oi_1 _20915_ (.A1(_11545_),
    .A2(_03645_),
    .Y(_03663_),
    .B1(_11026_));
 sg13g2_nor3_1 _20916_ (.A(_11265_),
    .B(_03662_),
    .C(_03663_),
    .Y(_03664_));
 sg13g2_a21oi_1 _20917_ (.A1(net77),
    .A2(_03659_),
    .Y(_03665_),
    .B1(_03664_));
 sg13g2_nand2b_1 _20918_ (.Y(_03666_),
    .B(net463),
    .A_N(_03665_));
 sg13g2_buf_1 _20919_ (.A(net559),
    .X(_03667_));
 sg13g2_nand2_2 _20920_ (.Y(_03668_),
    .A(_09972_),
    .B(_11199_));
 sg13g2_nand4_1 _20921_ (.B(_09960_),
    .C(\cpu.ex.r_set_cc ),
    .A(net1086),
    .Y(_03669_),
    .D(\cpu.ex.r_cc ));
 sg13g2_a21oi_1 _20922_ (.A1(_03668_),
    .A2(_03669_),
    .Y(_03670_),
    .B1(_03622_));
 sg13g2_buf_2 _20923_ (.A(_03670_),
    .X(_03671_));
 sg13g2_buf_1 _20924_ (.A(_03671_),
    .X(_03672_));
 sg13g2_a21oi_1 _20925_ (.A1(net530),
    .A2(net496),
    .Y(_03673_),
    .B1(net227));
 sg13g2_a22oi_1 _20926_ (.Y(_00967_),
    .B1(_03666_),
    .B2(_03673_),
    .A2(_03653_),
    .A1(_03651_));
 sg13g2_inv_1 _20927_ (.Y(_03674_),
    .A(\cpu.ex.r_mult[18] ));
 sg13g2_nor2_1 _20928_ (.A(_09124_),
    .B(net361),
    .Y(_03675_));
 sg13g2_buf_2 _20929_ (.A(_03675_),
    .X(_03676_));
 sg13g2_nand2b_1 _20930_ (.Y(_03677_),
    .B(_03676_),
    .A_N(_03662_));
 sg13g2_a21o_1 _20931_ (.A2(net282),
    .A1(_03655_),
    .B1(_03654_),
    .X(_03678_));
 sg13g2_o21ai_1 _20932_ (.B1(_03678_),
    .Y(_03679_),
    .A1(_03655_),
    .A2(net282));
 sg13g2_xnor2_1 _20933_ (.Y(_03680_),
    .A(net289),
    .B(_03679_));
 sg13g2_nor2_1 _20934_ (.A(net33),
    .B(_03680_),
    .Y(_03681_));
 sg13g2_nand2_1 _20935_ (.Y(_03682_),
    .A(net526),
    .B(net77));
 sg13g2_or2_1 _20936_ (.X(_03683_),
    .B(_03682_),
    .A(_03681_));
 sg13g2_a21oi_1 _20937_ (.A1(_03677_),
    .A2(_03683_),
    .Y(_03684_),
    .B1(_00308_));
 sg13g2_a22oi_1 _20938_ (.Y(_03685_),
    .B1(_03681_),
    .B2(net77),
    .A2(_03662_),
    .A1(_03676_));
 sg13g2_nor2_1 _20939_ (.A(_11084_),
    .B(_03685_),
    .Y(_03686_));
 sg13g2_o21ai_1 _20940_ (.B1(net463),
    .Y(_03687_),
    .A1(_03684_),
    .A2(_03686_));
 sg13g2_a21oi_1 _20941_ (.A1(net565),
    .A2(net496),
    .Y(_03688_),
    .B1(net227));
 sg13g2_a22oi_1 _20942_ (.Y(_00968_),
    .B1(_03687_),
    .B2(_03688_),
    .A2(_03653_),
    .A1(_03674_));
 sg13g2_nand3b_1 _20943_ (.B(_11171_),
    .C(_11003_),
    .Y(_03689_),
    .A_N(_11086_));
 sg13g2_buf_1 _20944_ (.A(_03689_),
    .X(_03690_));
 sg13g2_and3_1 _20945_ (.X(_03691_),
    .A(net202),
    .B(_11136_),
    .C(_03690_));
 sg13g2_a21oi_1 _20946_ (.A1(_11136_),
    .A2(_03690_),
    .Y(_03692_),
    .B1(net235));
 sg13g2_nor3_1 _20947_ (.A(net31),
    .B(_03691_),
    .C(_03692_),
    .Y(_03693_));
 sg13g2_xnor2_1 _20948_ (.Y(_03694_),
    .A(_11119_),
    .B(_03693_));
 sg13g2_and3_1 _20949_ (.X(_03695_),
    .A(_11084_),
    .B(_03645_),
    .C(_03660_));
 sg13g2_xnor2_1 _20950_ (.Y(_03696_),
    .A(_11118_),
    .B(_03695_));
 sg13g2_a221oi_1 _20951_ (.B2(_03676_),
    .C1(net227),
    .B1(_03696_),
    .A1(_11372_),
    .Y(_03697_),
    .A2(_03694_));
 sg13g2_nor2_1 _20952_ (.A(_09972_),
    .B(_03671_),
    .Y(_03698_));
 sg13g2_nor2_1 _20953_ (.A(_03622_),
    .B(_03698_),
    .Y(_03699_));
 sg13g2_o21ai_1 _20954_ (.B1(_03699_),
    .Y(_03700_),
    .A1(\cpu.ex.r_mult[19] ),
    .A2(_03668_));
 sg13g2_nand2_1 _20955_ (.Y(_03701_),
    .A(_08947_),
    .B(net496));
 sg13g2_o21ai_1 _20956_ (.B1(_03701_),
    .Y(_00969_),
    .A1(_03697_),
    .A2(_03700_));
 sg13g2_nand3_1 _20957_ (.B(_11136_),
    .C(_03690_),
    .A(net202),
    .Y(_03702_));
 sg13g2_a21o_1 _20958_ (.A2(_03702_),
    .A1(_11119_),
    .B1(_03692_),
    .X(_03703_));
 sg13g2_buf_1 _20959_ (.A(_03703_),
    .X(_03704_));
 sg13g2_xnor2_1 _20960_ (.Y(_03705_),
    .A(net238),
    .B(_03704_));
 sg13g2_nor2_1 _20961_ (.A(_11164_),
    .B(_03705_),
    .Y(_03706_));
 sg13g2_xor2_1 _20962_ (.B(_03706_),
    .A(_11124_),
    .X(_03707_));
 sg13g2_nor2_1 _20963_ (.A(_11190_),
    .B(_03707_),
    .Y(_03708_));
 sg13g2_nand3b_1 _20964_ (.B(net460),
    .C(_03695_),
    .Y(_03709_),
    .A_N(_11118_));
 sg13g2_nand3b_1 _20965_ (.B(_11084_),
    .C(_03660_),
    .Y(_03710_),
    .A_N(_10461_));
 sg13g2_nor3_1 _20966_ (.A(_11118_),
    .B(_11239_),
    .C(_03710_),
    .Y(_03711_));
 sg13g2_o21ai_1 _20967_ (.B1(_03711_),
    .Y(_03712_),
    .A1(_03631_),
    .A2(_03643_));
 sg13g2_buf_2 _20968_ (.A(_03712_),
    .X(_03713_));
 sg13g2_nand2_1 _20969_ (.Y(_03714_),
    .A(_03676_),
    .B(_03713_));
 sg13g2_a21oi_1 _20970_ (.A1(_10461_),
    .A2(_03709_),
    .Y(_03715_),
    .B1(_03714_));
 sg13g2_nor3_1 _20971_ (.A(_03671_),
    .B(_03708_),
    .C(_03715_),
    .Y(_03716_));
 sg13g2_o21ai_1 _20972_ (.B1(_03699_),
    .Y(_03717_),
    .A1(\cpu.ex.r_mult[20] ),
    .A2(_03668_));
 sg13g2_nand2_1 _20973_ (.Y(_03718_),
    .A(net573),
    .B(_03667_));
 sg13g2_o21ai_1 _20974_ (.B1(_03718_),
    .Y(_00970_),
    .A1(_03716_),
    .A2(_03717_));
 sg13g2_nand2_1 _20975_ (.Y(_03719_),
    .A(net238),
    .B(_03704_));
 sg13g2_o21ai_1 _20976_ (.B1(_11124_),
    .Y(_03720_),
    .A1(_11167_),
    .A2(_03704_));
 sg13g2_and3_1 _20977_ (.X(_03721_),
    .A(net236),
    .B(_03719_),
    .C(_03720_));
 sg13g2_a21oi_1 _20978_ (.A1(_03719_),
    .A2(_03720_),
    .Y(_03722_),
    .B1(_11186_));
 sg13g2_nor3_1 _20979_ (.A(_03618_),
    .B(_03721_),
    .C(_03722_),
    .Y(_03723_));
 sg13g2_nor2_1 _20980_ (.A(_11265_),
    .B(_03713_),
    .Y(_03724_));
 sg13g2_a21oi_1 _20981_ (.A1(net77),
    .A2(_03723_),
    .Y(_03725_),
    .B1(_03724_));
 sg13g2_nand2_1 _20982_ (.Y(_03726_),
    .A(net463),
    .B(_11199_));
 sg13g2_nor2_1 _20983_ (.A(\cpu.ex.r_mult[21] ),
    .B(_03726_),
    .Y(_03727_));
 sg13g2_nand3b_1 _20984_ (.B(_09975_),
    .C(_10489_),
    .Y(_03728_),
    .A_N(_03727_));
 sg13g2_a21oi_1 _20985_ (.A1(net635),
    .A2(net559),
    .Y(_03729_),
    .B1(_03671_));
 sg13g2_or2_1 _20986_ (.X(_03730_),
    .B(_03729_),
    .A(_03727_));
 sg13g2_o21ai_1 _20987_ (.B1(_03730_),
    .Y(_03731_),
    .A1(_03725_),
    .A2(_03728_));
 sg13g2_o21ai_1 _20988_ (.B1(_03714_),
    .Y(_03732_),
    .A1(_03682_),
    .A2(_03723_));
 sg13g2_nor2_1 _20989_ (.A(net523),
    .B(_03727_),
    .Y(_03733_));
 sg13g2_nand3b_1 _20990_ (.B(_03732_),
    .C(_03733_),
    .Y(_03734_),
    .A_N(_10489_));
 sg13g2_nand2b_1 _20991_ (.Y(_00971_),
    .B(_03734_),
    .A_N(_03731_));
 sg13g2_inv_1 _20992_ (.Y(_03735_),
    .A(_10493_));
 sg13g2_nor2_1 _20993_ (.A(_11139_),
    .B(_03735_),
    .Y(_03736_));
 sg13g2_xnor2_1 _20994_ (.Y(_03737_),
    .A(_10435_),
    .B(_03736_));
 sg13g2_nor2_1 _20995_ (.A(_03618_),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_xnor2_1 _20996_ (.Y(_03739_),
    .A(_10496_),
    .B(_03738_));
 sg13g2_o21ai_1 _20997_ (.B1(_00304_),
    .Y(_03740_),
    .A1(_10489_),
    .A2(_03713_));
 sg13g2_or2_1 _20998_ (.X(_03741_),
    .B(_10489_),
    .A(_00304_));
 sg13g2_buf_1 _20999_ (.A(_03741_),
    .X(_03742_));
 sg13g2_nor2_1 _21000_ (.A(_03713_),
    .B(_03742_),
    .Y(_03743_));
 sg13g2_nor2_1 _21001_ (.A(_11265_),
    .B(_03743_),
    .Y(_03744_));
 sg13g2_a221oi_1 _21002_ (.B2(_03744_),
    .C1(_03672_),
    .B1(_03740_),
    .A1(net77),
    .Y(_03745_),
    .A2(_03739_));
 sg13g2_o21ai_1 _21003_ (.B1(_03699_),
    .Y(_03746_),
    .A1(_10415_),
    .A2(_03668_));
 sg13g2_nand2_1 _21004_ (.Y(_03747_),
    .A(net838),
    .B(net496));
 sg13g2_o21ai_1 _21005_ (.B1(_03747_),
    .Y(_00972_),
    .A1(_03745_),
    .A2(_03746_));
 sg13g2_o21ai_1 _21006_ (.B1(net204),
    .Y(_03748_),
    .A1(_11139_),
    .A2(_03735_));
 sg13g2_nor3_1 _21007_ (.A(net204),
    .B(_11139_),
    .C(_03735_),
    .Y(_03749_));
 sg13g2_a21oi_1 _21008_ (.A1(_10496_),
    .A2(_03748_),
    .Y(_03750_),
    .B1(_03749_));
 sg13g2_xnor2_1 _21009_ (.Y(_03751_),
    .A(_11166_),
    .B(_03750_));
 sg13g2_nor2_1 _21010_ (.A(net31),
    .B(_03751_),
    .Y(_03752_));
 sg13g2_xnor2_1 _21011_ (.Y(_03753_),
    .A(_11142_),
    .B(_03752_));
 sg13g2_nand2_1 _21012_ (.Y(_03754_),
    .A(_10415_),
    .B(net460));
 sg13g2_mux2_1 _21013_ (.A0(_03754_),
    .A1(_10415_),
    .S(_03743_),
    .X(_03755_));
 sg13g2_inv_1 _21014_ (.Y(_03756_),
    .A(_03755_));
 sg13g2_a221oi_1 _21015_ (.B2(net989),
    .C1(net227),
    .B1(_03756_),
    .A1(net77),
    .Y(_03757_),
    .A2(_03753_));
 sg13g2_o21ai_1 _21016_ (.B1(_03699_),
    .Y(_03758_),
    .A1(\cpu.ex.r_mult[23] ),
    .A2(_03668_));
 sg13g2_nand2_1 _21017_ (.Y(_03759_),
    .A(net843),
    .B(_03667_));
 sg13g2_o21ai_1 _21018_ (.B1(_03759_),
    .Y(_00973_),
    .A1(_03757_),
    .A2(_03758_));
 sg13g2_inv_1 _21019_ (.Y(_03760_),
    .A(\cpu.ex.r_mult[24] ));
 sg13g2_nor2_2 _21020_ (.A(_11240_),
    .B(_11418_),
    .Y(_03761_));
 sg13g2_nand2_1 _21021_ (.Y(_03762_),
    .A(_10415_),
    .B(_03743_));
 sg13g2_xnor2_1 _21022_ (.Y(_03763_),
    .A(_10110_),
    .B(_03762_));
 sg13g2_nand2_1 _21023_ (.Y(_03764_),
    .A(_03761_),
    .B(_03763_));
 sg13g2_nand3_1 _21024_ (.B(_11147_),
    .C(_11152_),
    .A(_11141_),
    .Y(_03765_));
 sg13g2_buf_2 _21025_ (.A(_03765_),
    .X(_03766_));
 sg13g2_nor2_1 _21026_ (.A(net181),
    .B(_03766_),
    .Y(_03767_));
 sg13g2_nor2_1 _21027_ (.A(net182),
    .B(_11153_),
    .Y(_03768_));
 sg13g2_nor3_1 _21028_ (.A(net31),
    .B(_03767_),
    .C(_03768_),
    .Y(_03769_));
 sg13g2_xor2_1 _21029_ (.B(_03769_),
    .A(_10366_),
    .X(_03770_));
 sg13g2_a221oi_1 _21030_ (.B2(_03770_),
    .C1(_03672_),
    .B1(_11494_),
    .A1(net1085),
    .Y(_03771_),
    .A2(net496));
 sg13g2_a22oi_1 _21031_ (.Y(_00974_),
    .B1(_03764_),
    .B2(_03771_),
    .A2(_03653_),
    .A1(_03760_));
 sg13g2_inv_1 _21032_ (.Y(_03772_),
    .A(\cpu.ex.r_mult[25] ));
 sg13g2_nand3b_1 _21033_ (.B(_10110_),
    .C(_10415_),
    .Y(_03773_),
    .A_N(_10112_));
 sg13g2_nor3_1 _21034_ (.A(_03713_),
    .B(_03742_),
    .C(_03773_),
    .Y(_03774_));
 sg13g2_o21ai_1 _21035_ (.B1(_10112_),
    .Y(_03775_),
    .A1(_10109_),
    .A2(_03762_));
 sg13g2_nand3b_1 _21036_ (.B(_03761_),
    .C(_03775_),
    .Y(_03776_),
    .A_N(_03774_));
 sg13g2_a221oi_1 _21037_ (.B2(_03766_),
    .C1(_10109_),
    .B1(net181),
    .A1(_09113_),
    .Y(_03777_),
    .A2(net646));
 sg13g2_o21ai_1 _21038_ (.B1(net234),
    .Y(_03778_),
    .A1(_03767_),
    .A2(_03777_));
 sg13g2_or3_1 _21039_ (.A(net234),
    .B(_03767_),
    .C(_03777_),
    .X(_03779_));
 sg13g2_a21oi_1 _21040_ (.A1(_03778_),
    .A2(_03779_),
    .Y(_03780_),
    .B1(net31));
 sg13g2_xor2_1 _21041_ (.B(_03780_),
    .A(_10372_),
    .X(_03781_));
 sg13g2_a221oi_1 _21042_ (.B2(_03781_),
    .C1(net227),
    .B1(_11494_),
    .A1(_09985_),
    .Y(_03782_),
    .A2(net496));
 sg13g2_a22oi_1 _21043_ (.Y(_00975_),
    .B1(_03776_),
    .B2(_03782_),
    .A2(_03653_),
    .A1(_03772_));
 sg13g2_and2_1 _21044_ (.A(_10361_),
    .B(_03774_),
    .X(_03783_));
 sg13g2_nand2b_1 _21045_ (.Y(_03784_),
    .B(_10190_),
    .A_N(_03774_));
 sg13g2_nand3b_1 _21046_ (.B(_03784_),
    .C(_03761_),
    .Y(_03785_),
    .A_N(_03783_));
 sg13g2_nand2_1 _21047_ (.Y(_03786_),
    .A(_10361_),
    .B(net526));
 sg13g2_buf_2 _21048_ (.A(_03786_),
    .X(_03787_));
 sg13g2_nand4_1 _21049_ (.B(_11141_),
    .C(_11147_),
    .A(_10375_),
    .Y(_03788_),
    .D(_11152_));
 sg13g2_nor2b_1 _21050_ (.A(_10119_),
    .B_N(_03788_),
    .Y(_03789_));
 sg13g2_buf_1 _21051_ (.A(_03789_),
    .X(_03790_));
 sg13g2_xnor2_1 _21052_ (.Y(_03791_),
    .A(net208),
    .B(_03790_));
 sg13g2_nor2_1 _21053_ (.A(net31),
    .B(_03791_),
    .Y(_03792_));
 sg13g2_xnor2_1 _21054_ (.Y(_03793_),
    .A(_03787_),
    .B(_03792_));
 sg13g2_a221oi_1 _21055_ (.B2(_03793_),
    .C1(net227),
    .B1(_11494_),
    .A1(net1075),
    .Y(_03794_),
    .A2(net496));
 sg13g2_a22oi_1 _21056_ (.Y(_00976_),
    .B1(_03785_),
    .B2(_03794_),
    .A2(_03653_),
    .A1(_10189_));
 sg13g2_nor2_1 _21057_ (.A(\cpu.ex.r_mult[27] ),
    .B(_03726_),
    .Y(_03795_));
 sg13g2_nor2_1 _21058_ (.A(net180),
    .B(net33),
    .Y(_03796_));
 sg13g2_nor2_1 _21059_ (.A(_10193_),
    .B(net33),
    .Y(_03797_));
 sg13g2_nor2_1 _21060_ (.A(_10190_),
    .B(net462),
    .Y(_03798_));
 sg13g2_nor2_1 _21061_ (.A(net207),
    .B(_03798_),
    .Y(_03799_));
 sg13g2_nand2_1 _21062_ (.Y(_03800_),
    .A(net207),
    .B(_03798_));
 sg13g2_o21ai_1 _21063_ (.B1(_03800_),
    .Y(_03801_),
    .A1(_03790_),
    .A2(_03799_));
 sg13g2_mux2_1 _21064_ (.A0(_03796_),
    .A1(_03797_),
    .S(_03801_),
    .X(_03802_));
 sg13g2_nand2_1 _21065_ (.Y(_03803_),
    .A(net995),
    .B(net526));
 sg13g2_xnor2_1 _21066_ (.Y(_03804_),
    .A(_03802_),
    .B(_03803_));
 sg13g2_a221oi_1 _21067_ (.B2(_03804_),
    .C1(net227),
    .B1(_11494_),
    .A1(_10147_),
    .Y(_03805_),
    .A2(net559));
 sg13g2_xnor2_1 _21068_ (.Y(_03806_),
    .A(_10189_),
    .B(_03783_));
 sg13g2_nand2_1 _21069_ (.Y(_03807_),
    .A(_03761_),
    .B(_03806_));
 sg13g2_o21ai_1 _21070_ (.B1(_03807_),
    .Y(_00977_),
    .A1(_03795_),
    .A2(_03805_));
 sg13g2_a21oi_1 _21071_ (.A1(net508),
    .A2(net496),
    .Y(_03808_),
    .B1(net227));
 sg13g2_nor2_1 _21072_ (.A(_10344_),
    .B(net462),
    .Y(_03809_));
 sg13g2_a21oi_1 _21073_ (.A1(_10119_),
    .A2(_10185_),
    .Y(_03810_),
    .B1(_10198_));
 sg13g2_nor2b_1 _21074_ (.A(_10363_),
    .B_N(_10375_),
    .Y(_03811_));
 sg13g2_nand4_1 _21075_ (.B(_11147_),
    .C(_11152_),
    .A(_11141_),
    .Y(_03812_),
    .D(_03811_));
 sg13g2_buf_1 _21076_ (.A(_03812_),
    .X(_03813_));
 sg13g2_a21o_1 _21077_ (.A2(_03813_),
    .A1(_03810_),
    .B1(net179),
    .X(_03814_));
 sg13g2_nand3_1 _21078_ (.B(_03810_),
    .C(_03813_),
    .A(net179),
    .Y(_03815_));
 sg13g2_a21oi_1 _21079_ (.A1(_03814_),
    .A2(_03815_),
    .Y(_03816_),
    .B1(net33));
 sg13g2_xor2_1 _21080_ (.B(_03816_),
    .A(_03809_),
    .X(_03817_));
 sg13g2_nand2_1 _21081_ (.Y(_03818_),
    .A(net995),
    .B(_10361_));
 sg13g2_nor4_2 _21082_ (.A(_03713_),
    .B(_03742_),
    .C(_03773_),
    .Y(_03819_),
    .D(_03818_));
 sg13g2_xnor2_1 _21083_ (.Y(_03820_),
    .A(_10344_),
    .B(_03819_));
 sg13g2_a22oi_1 _21084_ (.Y(_03821_),
    .B1(_03820_),
    .B2(_03676_),
    .A2(_03817_),
    .A1(net77));
 sg13g2_nand2b_1 _21085_ (.Y(_03822_),
    .B(_09975_),
    .A_N(_03821_));
 sg13g2_a22oi_1 _21086_ (.Y(_00978_),
    .B1(_03808_),
    .B2(_03822_),
    .A2(_03653_),
    .A1(_10343_));
 sg13g2_nor4_1 _21087_ (.A(net1071),
    .B(net462),
    .C(net203),
    .D(net31),
    .Y(_03823_));
 sg13g2_nor2_1 _21088_ (.A(_10343_),
    .B(net462),
    .Y(_03824_));
 sg13g2_and2_1 _21089_ (.A(net203),
    .B(_03824_),
    .X(_03825_));
 sg13g2_nand2_1 _21090_ (.Y(_03826_),
    .A(_10344_),
    .B(net200));
 sg13g2_nor2_1 _21091_ (.A(_10344_),
    .B(net180),
    .Y(_03827_));
 sg13g2_a21oi_1 _21092_ (.A1(net995),
    .A2(_03826_),
    .Y(_03828_),
    .B1(_03827_));
 sg13g2_nor2_1 _21093_ (.A(net208),
    .B(_03828_),
    .Y(_03829_));
 sg13g2_a221oi_1 _21094_ (.B2(_03829_),
    .C1(_10347_),
    .B1(_03798_),
    .A1(net995),
    .Y(_03830_),
    .A2(_10193_));
 sg13g2_a21oi_1 _21095_ (.A1(net995),
    .A2(_03798_),
    .Y(_03831_),
    .B1(_03829_));
 sg13g2_or2_1 _21096_ (.X(_03832_),
    .B(_03831_),
    .A(_03790_));
 sg13g2_nand3b_1 _21097_ (.B(_03788_),
    .C(_03787_),
    .Y(_03833_),
    .A_N(_10119_));
 sg13g2_nor2_1 _21098_ (.A(net180),
    .B(_03787_),
    .Y(_03834_));
 sg13g2_nand2_1 _21099_ (.Y(_03835_),
    .A(_10375_),
    .B(_03834_));
 sg13g2_a21oi_1 _21100_ (.A1(_10119_),
    .A2(_03834_),
    .Y(_03836_),
    .B1(net995));
 sg13g2_o21ai_1 _21101_ (.B1(_03836_),
    .Y(_03837_),
    .A1(_03766_),
    .A2(_03835_));
 sg13g2_nor2_1 _21102_ (.A(_10344_),
    .B(_03787_),
    .Y(_03838_));
 sg13g2_nand2_1 _21103_ (.Y(_03839_),
    .A(_10375_),
    .B(_03838_));
 sg13g2_a21oi_1 _21104_ (.A1(_10119_),
    .A2(_03838_),
    .Y(_03840_),
    .B1(_03827_));
 sg13g2_o21ai_1 _21105_ (.B1(_03840_),
    .Y(_03841_),
    .A1(_03766_),
    .A2(_03839_));
 sg13g2_a221oi_1 _21106_ (.B2(_03841_),
    .C1(net179),
    .B1(_03837_),
    .A1(_03833_),
    .Y(_03842_),
    .A2(_03829_));
 sg13g2_a21oi_1 _21107_ (.A1(_03830_),
    .A2(_03832_),
    .Y(_03843_),
    .B1(_03842_));
 sg13g2_o21ai_1 _21108_ (.B1(_03843_),
    .Y(_03844_),
    .A1(_03823_),
    .A2(_03825_));
 sg13g2_inv_1 _21109_ (.Y(_03845_),
    .A(net33));
 sg13g2_nand2_1 _21110_ (.Y(_03846_),
    .A(net179),
    .B(_10193_));
 sg13g2_nor2_1 _21111_ (.A(_03846_),
    .B(_03787_),
    .Y(_03847_));
 sg13g2_nand2_1 _21112_ (.Y(_03848_),
    .A(_10375_),
    .B(_03847_));
 sg13g2_nor2_1 _21113_ (.A(net208),
    .B(_03846_),
    .Y(_03849_));
 sg13g2_nand2_1 _21114_ (.Y(_03850_),
    .A(_10375_),
    .B(_03849_));
 sg13g2_a21oi_1 _21115_ (.A1(_03848_),
    .A2(_03850_),
    .Y(_03851_),
    .B1(_03766_));
 sg13g2_o21ai_1 _21116_ (.B1(_10119_),
    .Y(_03852_),
    .A1(_03847_),
    .A2(_03849_));
 sg13g2_o21ai_1 _21117_ (.B1(_03852_),
    .Y(_03853_),
    .A1(_03846_),
    .A2(_03800_));
 sg13g2_nor2_1 _21118_ (.A(_03851_),
    .B(_03853_),
    .Y(_03854_));
 sg13g2_nand4_1 _21119_ (.B(net203),
    .C(_03845_),
    .A(_10343_),
    .Y(_03855_),
    .D(_03854_));
 sg13g2_nand3_1 _21120_ (.B(_03854_),
    .C(_03824_),
    .A(net199),
    .Y(_03856_));
 sg13g2_a21o_1 _21121_ (.A2(_03856_),
    .A1(_03855_),
    .B1(_03843_),
    .X(_03857_));
 sg13g2_or2_1 _21122_ (.X(_03858_),
    .B(_03853_),
    .A(_03851_));
 sg13g2_nor2_1 _21123_ (.A(net1071),
    .B(net203),
    .Y(_03859_));
 sg13g2_nand3_1 _21124_ (.B(_03858_),
    .C(_03859_),
    .A(_03845_),
    .Y(_03860_));
 sg13g2_a22oi_1 _21125_ (.Y(_03861_),
    .B1(_03825_),
    .B2(_03858_),
    .A2(_03824_),
    .A1(net31));
 sg13g2_and4_1 _21126_ (.A(_03844_),
    .B(_03857_),
    .C(_03860_),
    .D(_03861_),
    .X(_03862_));
 sg13g2_nand2_1 _21127_ (.Y(_03863_),
    .A(_10347_),
    .B(_03819_));
 sg13g2_xnor2_1 _21128_ (.Y(_03864_),
    .A(net1071),
    .B(_03863_));
 sg13g2_a21oi_1 _21129_ (.A1(net577),
    .A2(net559),
    .Y(_03865_),
    .B1(_03671_));
 sg13g2_a21oi_1 _21130_ (.A1(_10271_),
    .A2(_03653_),
    .Y(_03866_),
    .B1(_03865_));
 sg13g2_a21oi_1 _21131_ (.A1(_03761_),
    .A2(_03864_),
    .Y(_03867_),
    .B1(_03866_));
 sg13g2_o21ai_1 _21132_ (.B1(_03867_),
    .Y(_00979_),
    .A1(_11413_),
    .A2(_03862_));
 sg13g2_a21oi_1 _21133_ (.A1(net578),
    .A2(net559),
    .Y(_03868_),
    .B1(_03671_));
 sg13g2_inv_1 _21134_ (.Y(_03869_),
    .A(_10355_));
 sg13g2_a21oi_1 _21135_ (.A1(_03810_),
    .A2(_03813_),
    .Y(_03870_),
    .B1(_03869_));
 sg13g2_nand2_1 _21136_ (.Y(_03871_),
    .A(net1074),
    .B(net526));
 sg13g2_a21oi_1 _21137_ (.A1(_10285_),
    .A2(_03870_),
    .Y(_03872_),
    .B1(_03871_));
 sg13g2_a21oi_1 _21138_ (.A1(_11155_),
    .A2(_11156_),
    .Y(_03873_),
    .B1(net462));
 sg13g2_nor2_1 _21139_ (.A(_03873_),
    .B(_03870_),
    .Y(_03874_));
 sg13g2_xor2_1 _21140_ (.B(_03871_),
    .A(net178),
    .X(_03875_));
 sg13g2_xnor2_1 _21141_ (.Y(_03876_),
    .A(_03874_),
    .B(_03875_));
 sg13g2_mux2_1 _21142_ (.A0(_03872_),
    .A1(_03876_),
    .S(_11162_),
    .X(_03877_));
 sg13g2_nand3_1 _21143_ (.B(_10347_),
    .C(_03819_),
    .A(net1071),
    .Y(_03878_));
 sg13g2_xnor2_1 _21144_ (.Y(_03879_),
    .A(_10231_),
    .B(_03878_));
 sg13g2_a22oi_1 _21145_ (.Y(_03880_),
    .B1(_03879_),
    .B2(_03676_),
    .A2(_03877_),
    .A1(net77));
 sg13g2_nand2_1 _21146_ (.Y(_03881_),
    .A(net523),
    .B(_03868_));
 sg13g2_o21ai_1 _21147_ (.B1(_03881_),
    .Y(_03882_),
    .A1(\cpu.ex.r_mult[30] ),
    .A2(_03726_));
 sg13g2_a21oi_1 _21148_ (.A1(_03868_),
    .A2(_03880_),
    .Y(_00980_),
    .B1(_03882_));
 sg13g2_a21oi_1 _21149_ (.A1(net994),
    .A2(net559),
    .Y(_03883_),
    .B1(_03671_));
 sg13g2_nand4_1 _21150_ (.B(net1074),
    .C(_10347_),
    .A(net1071),
    .Y(_03884_),
    .D(_03819_));
 sg13g2_xnor2_1 _21151_ (.Y(_03885_),
    .A(_10279_),
    .B(_03884_));
 sg13g2_nor2_1 _21152_ (.A(_10232_),
    .B(_03682_),
    .Y(_03886_));
 sg13g2_nor2_1 _21153_ (.A(_10189_),
    .B(net180),
    .Y(_03887_));
 sg13g2_o21ai_1 _21154_ (.B1(_03826_),
    .Y(_03888_),
    .A1(_11154_),
    .A2(_03887_));
 sg13g2_nand2_1 _21155_ (.Y(_03889_),
    .A(net1071),
    .B(net203));
 sg13g2_o21ai_1 _21156_ (.B1(_03889_),
    .Y(_03890_),
    .A1(_03859_),
    .A2(_03888_));
 sg13g2_a21oi_1 _21157_ (.A1(net1074),
    .A2(net151),
    .Y(_03891_),
    .B1(_03890_));
 sg13g2_a21oi_1 _21158_ (.A1(_10271_),
    .A2(net178),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_a21oi_1 _21159_ (.A1(_10189_),
    .A2(_10271_),
    .Y(_03893_),
    .B1(net462));
 sg13g2_nor3_1 _21160_ (.A(net178),
    .B(net180),
    .C(_03893_),
    .Y(_03894_));
 sg13g2_nand3_1 _21161_ (.B(_10273_),
    .C(_10193_),
    .A(_10189_),
    .Y(_03895_));
 sg13g2_xnor2_1 _21162_ (.Y(_03896_),
    .A(net1074),
    .B(net178));
 sg13g2_nand3_1 _21163_ (.B(net180),
    .C(_03896_),
    .A(net995),
    .Y(_03897_));
 sg13g2_a21oi_1 _21164_ (.A1(_03895_),
    .A2(_03897_),
    .Y(_03898_),
    .B1(net462));
 sg13g2_o21ai_1 _21165_ (.B1(_10355_),
    .Y(_03899_),
    .A1(_03894_),
    .A2(_03898_));
 sg13g2_nor2b_1 _21166_ (.A(_03899_),
    .B_N(_03833_),
    .Y(_03900_));
 sg13g2_o21ai_1 _21167_ (.B1(net208),
    .Y(_03901_),
    .A1(_03787_),
    .A2(_03790_));
 sg13g2_a22oi_1 _21168_ (.Y(_03902_),
    .B1(_03900_),
    .B2(_03901_),
    .A2(_03892_),
    .A1(net526));
 sg13g2_o21ai_1 _21169_ (.B1(_03845_),
    .Y(_03903_),
    .A1(net241),
    .A2(_03902_));
 sg13g2_a22oi_1 _21170_ (.Y(_03904_),
    .B1(_03886_),
    .B2(_03903_),
    .A2(_03885_),
    .A1(_03676_));
 sg13g2_nand2_1 _21171_ (.Y(_03905_),
    .A(_11233_),
    .B(_03883_));
 sg13g2_o21ai_1 _21172_ (.B1(_03905_),
    .Y(_03906_),
    .A1(\cpu.ex.r_mult[31] ),
    .A2(_03726_));
 sg13g2_a21oi_1 _21173_ (.A1(_03883_),
    .A2(_03904_),
    .Y(_00981_),
    .B1(_03906_));
 sg13g2_inv_1 _21174_ (.Y(_03907_),
    .A(_00258_));
 sg13g2_nand3_1 _21175_ (.B(_03907_),
    .C(_11567_),
    .A(_08589_),
    .Y(_03908_));
 sg13g2_o21ai_1 _21176_ (.B1(_03908_),
    .Y(_03909_),
    .A1(net1091),
    .A2(_11567_));
 sg13g2_and2_1 _21177_ (.A(_08619_),
    .B(_10654_),
    .X(_03910_));
 sg13g2_buf_1 _21178_ (.A(_03910_),
    .X(_03911_));
 sg13g2_nand3_1 _21179_ (.B(_03909_),
    .C(_03911_),
    .A(net646),
    .Y(_03912_));
 sg13g2_buf_1 _21180_ (.A(_03912_),
    .X(_03913_));
 sg13g2_buf_1 _21181_ (.A(_03913_),
    .X(_03914_));
 sg13g2_buf_1 _21182_ (.A(_11209_),
    .X(_03915_));
 sg13g2_nor2_2 _21183_ (.A(net290),
    .B(_11272_),
    .Y(_03916_));
 sg13g2_nor2b_1 _21184_ (.A(_03398_),
    .B_N(_08051_),
    .Y(_03917_));
 sg13g2_nand3_1 _21185_ (.B(_03916_),
    .C(_03917_),
    .A(net292),
    .Y(_03918_));
 sg13g2_buf_1 _21186_ (.A(_03407_),
    .X(_03919_));
 sg13g2_nand3_1 _21187_ (.B(_11182_),
    .C(net190),
    .A(net283),
    .Y(_03920_));
 sg13g2_a21oi_1 _21188_ (.A1(_03918_),
    .A2(_03920_),
    .Y(_03921_),
    .B1(net282));
 sg13g2_nor2_2 _21189_ (.A(net333),
    .B(net237),
    .Y(_03922_));
 sg13g2_and2_1 _21190_ (.A(_03523_),
    .B(_03922_),
    .X(_03923_));
 sg13g2_buf_1 _21191_ (.A(_03923_),
    .X(_03924_));
 sg13g2_nand2_1 _21192_ (.Y(_03925_),
    .A(net228),
    .B(_03924_));
 sg13g2_buf_1 _21193_ (.A(_10981_),
    .X(_03926_));
 sg13g2_nor4_1 _21194_ (.A(net335),
    .B(net334),
    .C(net332),
    .D(net237),
    .Y(_03927_));
 sg13g2_buf_1 _21195_ (.A(_03927_),
    .X(_03928_));
 sg13g2_nand2_1 _21196_ (.Y(_03929_),
    .A(net225),
    .B(net170));
 sg13g2_nand2_1 _21197_ (.Y(_03930_),
    .A(net335),
    .B(net334));
 sg13g2_nand2_1 _21198_ (.Y(_03931_),
    .A(net332),
    .B(net237));
 sg13g2_buf_1 _21199_ (.A(_03931_),
    .X(_03932_));
 sg13g2_nor2_1 _21200_ (.A(_03930_),
    .B(_03932_),
    .Y(_03933_));
 sg13g2_buf_1 _21201_ (.A(_03933_),
    .X(_03934_));
 sg13g2_nor2_1 _21202_ (.A(net332),
    .B(_11271_),
    .Y(_03935_));
 sg13g2_nor2_1 _21203_ (.A(net335),
    .B(net362),
    .Y(_03936_));
 sg13g2_buf_1 _21204_ (.A(_03936_),
    .X(_03937_));
 sg13g2_and2_1 _21205_ (.A(_03935_),
    .B(_03937_),
    .X(_03938_));
 sg13g2_buf_1 _21206_ (.A(_03938_),
    .X(_03939_));
 sg13g2_a22oi_1 _21207_ (.Y(_03940_),
    .B1(_03939_),
    .B2(net149),
    .A2(_03934_),
    .A1(_10925_));
 sg13g2_nand3_1 _21208_ (.B(_03929_),
    .C(_03940_),
    .A(_03925_),
    .Y(_03941_));
 sg13g2_nand2_1 _21209_ (.Y(_03942_),
    .A(net333),
    .B(_11271_));
 sg13g2_buf_1 _21210_ (.A(_03942_),
    .X(_03943_));
 sg13g2_nor2_1 _21211_ (.A(net292),
    .B(_03917_),
    .Y(_03944_));
 sg13g2_nor3_1 _21212_ (.A(net362),
    .B(_03943_),
    .C(_03944_),
    .Y(_03945_));
 sg13g2_nand2_1 _21213_ (.Y(_03946_),
    .A(_03922_),
    .B(net224));
 sg13g2_nor2_1 _21214_ (.A(_03505_),
    .B(_03946_),
    .Y(_03947_));
 sg13g2_nand2_1 _21215_ (.Y(_03948_),
    .A(_11175_),
    .B(_03922_));
 sg13g2_nor2_1 _21216_ (.A(_03432_),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_nor4_1 _21217_ (.A(_03941_),
    .B(_03945_),
    .C(_03947_),
    .D(_03949_),
    .Y(_03950_));
 sg13g2_and2_1 _21218_ (.A(_03523_),
    .B(_03935_),
    .X(_03951_));
 sg13g2_buf_1 _21219_ (.A(_03951_),
    .X(_03952_));
 sg13g2_nor2_1 _21220_ (.A(_11171_),
    .B(net334),
    .Y(_03953_));
 sg13g2_buf_1 _21221_ (.A(_03953_),
    .X(_03954_));
 sg13g2_nand3_1 _21222_ (.B(net235),
    .C(_03954_),
    .A(net332),
    .Y(_03955_));
 sg13g2_buf_1 _21223_ (.A(_03955_),
    .X(_03956_));
 sg13g2_nor2_1 _21224_ (.A(_03456_),
    .B(_03956_),
    .Y(_03957_));
 sg13g2_a21oi_1 _21225_ (.A1(net193),
    .A2(net169),
    .Y(_03958_),
    .B1(_03957_));
 sg13g2_a22oi_1 _21226_ (.Y(_03959_),
    .B1(_03954_),
    .B2(net192),
    .A2(net224),
    .A1(net194));
 sg13g2_nand2b_1 _21227_ (.Y(_03960_),
    .B(_03916_),
    .A_N(_03959_));
 sg13g2_buf_1 _21228_ (.A(_03561_),
    .X(_03961_));
 sg13g2_nand2_2 _21229_ (.Y(_03962_),
    .A(net335),
    .B(net362));
 sg13g2_nor3_1 _21230_ (.A(net332),
    .B(net235),
    .C(_03962_),
    .Y(_03963_));
 sg13g2_buf_1 _21231_ (.A(_03963_),
    .X(_03964_));
 sg13g2_nor3_1 _21232_ (.A(net332),
    .B(net235),
    .C(_03930_),
    .Y(_03965_));
 sg13g2_buf_1 _21233_ (.A(_03965_),
    .X(_03966_));
 sg13g2_buf_1 _21234_ (.A(_03966_),
    .X(_03967_));
 sg13g2_buf_1 _21235_ (.A(net172),
    .X(_03968_));
 sg13g2_a22oi_1 _21236_ (.Y(_03969_),
    .B1(net147),
    .B2(net146),
    .A2(net168),
    .A1(net189));
 sg13g2_nand4_1 _21237_ (.B(_03958_),
    .C(_03960_),
    .A(_03950_),
    .Y(_03970_),
    .D(_03969_));
 sg13g2_nor2_1 _21238_ (.A(_00297_),
    .B(net230),
    .Y(_03971_));
 sg13g2_a21oi_1 _21239_ (.A1(_03403_),
    .A2(_11558_),
    .Y(_03972_),
    .B1(_03971_));
 sg13g2_nor4_1 _21240_ (.A(net335),
    .B(net362),
    .C(net332),
    .D(net237),
    .Y(_03973_));
 sg13g2_buf_2 _21241_ (.A(_03973_),
    .X(_03974_));
 sg13g2_buf_1 _21242_ (.A(_03974_),
    .X(_03975_));
 sg13g2_buf_1 _21243_ (.A(net145),
    .X(_03976_));
 sg13g2_nor2_2 _21244_ (.A(_08051_),
    .B(_09635_),
    .Y(_03977_));
 sg13g2_a21oi_1 _21245_ (.A1(_03972_),
    .A2(net120),
    .Y(_03978_),
    .B1(_03977_));
 sg13g2_o21ai_1 _21246_ (.B1(_03978_),
    .Y(_03979_),
    .A1(_03921_),
    .A2(_03970_));
 sg13g2_nor2_1 _21247_ (.A(_09662_),
    .B(net293),
    .Y(_03980_));
 sg13g2_nor2b_1 _21248_ (.A(_11197_),
    .B_N(_11208_),
    .Y(_03981_));
 sg13g2_buf_1 _21249_ (.A(_03981_),
    .X(_03982_));
 sg13g2_a221oi_1 _21250_ (.B2(_03980_),
    .C1(_03982_),
    .B1(net120),
    .A1(_08763_),
    .Y(_03983_),
    .A2(net234));
 sg13g2_a21oi_2 _21251_ (.B1(_03418_),
    .Y(_03984_),
    .A2(_10822_),
    .A1(_03403_));
 sg13g2_nor2_1 _21252_ (.A(net282),
    .B(_03984_),
    .Y(_03985_));
 sg13g2_nand2_1 _21253_ (.Y(_03986_),
    .A(net282),
    .B(_03984_));
 sg13g2_nand2b_1 _21254_ (.Y(_03987_),
    .B(_03986_),
    .A_N(_03985_));
 sg13g2_nor4_1 _21255_ (.A(net1088),
    .B(_09654_),
    .C(_09661_),
    .D(_09672_),
    .Y(_03988_));
 sg13g2_nor4_1 _21256_ (.A(_08839_),
    .B(\cpu.dec.r_op[6] ),
    .C(_09652_),
    .D(_09676_),
    .Y(_03989_));
 sg13g2_and3_1 _21257_ (.X(_03990_),
    .A(_03977_),
    .B(_03988_),
    .C(_03989_));
 sg13g2_buf_1 _21258_ (.A(_03990_),
    .X(_03991_));
 sg13g2_nor3_2 _21259_ (.A(_09652_),
    .B(_09676_),
    .C(_03991_),
    .Y(_03992_));
 sg13g2_a21oi_1 _21260_ (.A1(net293),
    .A2(_03987_),
    .Y(_03993_),
    .B1(_03992_));
 sg13g2_or3_1 _21261_ (.A(_09652_),
    .B(_09676_),
    .C(_03991_),
    .X(_03994_));
 sg13g2_buf_2 _21262_ (.A(_03994_),
    .X(_03995_));
 sg13g2_o21ai_1 _21263_ (.B1(net292),
    .Y(_03996_),
    .A1(_10680_),
    .A2(_03995_));
 sg13g2_buf_1 _21264_ (.A(_03520_),
    .X(_03997_));
 sg13g2_nor2_1 _21265_ (.A(_03997_),
    .B(_03992_),
    .Y(_03998_));
 sg13g2_nor2_1 _21266_ (.A(_08922_),
    .B(_10680_),
    .Y(_03999_));
 sg13g2_nor3_1 _21267_ (.A(_03987_),
    .B(_03998_),
    .C(_03999_),
    .Y(_04000_));
 sg13g2_a22oi_1 _21268_ (.Y(_04001_),
    .B1(_04000_),
    .B2(net292),
    .A2(_03996_),
    .A1(_03987_));
 sg13g2_o21ai_1 _21269_ (.B1(_04001_),
    .Y(_04002_),
    .A1(net1086),
    .A2(_03993_));
 sg13g2_nand2_1 _21270_ (.Y(_04003_),
    .A(net1011),
    .B(_03985_));
 sg13g2_o21ai_1 _21271_ (.B1(_04003_),
    .Y(_04004_),
    .A1(net883),
    .A2(_03985_));
 sg13g2_o21ai_1 _21272_ (.B1(_03986_),
    .Y(_04005_),
    .A1(_09655_),
    .A2(_04004_));
 sg13g2_nand4_1 _21273_ (.B(_03983_),
    .C(_04002_),
    .A(_03979_),
    .Y(_04006_),
    .D(_04005_));
 sg13g2_o21ai_1 _21274_ (.B1(_04006_),
    .Y(_04007_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[1] ));
 sg13g2_nor3_1 _21275_ (.A(_09013_),
    .B(net1019),
    .C(_09108_),
    .Y(_04008_));
 sg13g2_and3_1 _21276_ (.X(_04009_),
    .A(_11568_),
    .B(_03911_),
    .C(_04008_));
 sg13g2_buf_1 _21277_ (.A(_04009_),
    .X(_04010_));
 sg13g2_nand2_1 _21278_ (.Y(_04011_),
    .A(\cpu.dec.iready ),
    .B(_00199_));
 sg13g2_nor2_1 _21279_ (.A(\cpu.ex.r_branch_stall ),
    .B(_04011_),
    .Y(_04012_));
 sg13g2_buf_1 _21280_ (.A(_04012_),
    .X(_04013_));
 sg13g2_nand3_1 _21281_ (.B(_08619_),
    .C(_04013_),
    .A(_08967_),
    .Y(_04014_));
 sg13g2_o21ai_1 _21282_ (.B1(_09108_),
    .Y(_04015_),
    .A1(_08557_),
    .A2(_08617_));
 sg13g2_a21oi_1 _21283_ (.A1(_04014_),
    .A2(_04015_),
    .Y(_04016_),
    .B1(_08558_));
 sg13g2_and4_1 _21284_ (.A(_10515_),
    .B(_08619_),
    .C(_09009_),
    .D(_04008_),
    .X(_04017_));
 sg13g2_nor4_1 _21285_ (.A(net1019),
    .B(net35),
    .C(_04016_),
    .D(_04017_),
    .Y(_04018_));
 sg13g2_and2_1 _21286_ (.A(_03913_),
    .B(_04018_),
    .X(_04019_));
 sg13g2_buf_1 _21287_ (.A(_04019_),
    .X(_04020_));
 sg13g2_buf_1 _21288_ (.A(_04020_),
    .X(_04021_));
 sg13g2_a22oi_1 _21289_ (.Y(_04022_),
    .B1(net28),
    .B2(net885),
    .A2(net35),
    .A1(_10771_));
 sg13g2_o21ai_1 _21290_ (.B1(_04022_),
    .Y(_00982_),
    .A1(_03914_),
    .A2(_04007_));
 sg13g2_nand2_1 _21291_ (.Y(_04023_),
    .A(_10193_),
    .B(_03468_));
 sg13g2_nand2_1 _21292_ (.Y(_04024_),
    .A(_03574_),
    .B(_04023_));
 sg13g2_buf_1 _21293_ (.A(_03464_),
    .X(_04025_));
 sg13g2_a221oi_1 _21294_ (.B2(_03443_),
    .C1(_03456_),
    .B1(_03440_),
    .A1(net102),
    .Y(_04026_),
    .A2(_03435_));
 sg13g2_buf_1 _21295_ (.A(_04026_),
    .X(_04027_));
 sg13g2_a221oi_1 _21296_ (.B2(_03443_),
    .C1(_10402_),
    .B1(_03440_),
    .A1(net102),
    .Y(_04028_),
    .A2(_03435_));
 sg13g2_buf_1 _21297_ (.A(_04028_),
    .X(_04029_));
 sg13g2_nand2_1 _21298_ (.Y(_04030_),
    .A(_10365_),
    .B(net172));
 sg13g2_nand2_1 _21299_ (.Y(_04031_),
    .A(net181),
    .B(_04030_));
 sg13g2_nor4_1 _21300_ (.A(_04027_),
    .B(_03457_),
    .C(_04029_),
    .D(_04031_),
    .Y(_04032_));
 sg13g2_nand2_1 _21301_ (.Y(_04033_),
    .A(_03537_),
    .B(_04030_));
 sg13g2_nor4_1 _21302_ (.A(_04027_),
    .B(_03457_),
    .C(_04029_),
    .D(_04033_),
    .Y(_04034_));
 sg13g2_nand3_1 _21303_ (.B(_03537_),
    .C(_04030_),
    .A(net181),
    .Y(_04035_));
 sg13g2_nand2_1 _21304_ (.Y(_04036_),
    .A(_03475_),
    .B(_04035_));
 sg13g2_nor3_2 _21305_ (.A(_04032_),
    .B(_04034_),
    .C(_04036_),
    .Y(_04037_));
 sg13g2_nor2_1 _21306_ (.A(net119),
    .B(_04037_),
    .Y(_04038_));
 sg13g2_a21oi_1 _21307_ (.A1(net119),
    .A2(_04037_),
    .Y(_04039_),
    .B1(_10188_));
 sg13g2_nor2_1 _21308_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_xnor2_1 _21309_ (.Y(_04041_),
    .A(_04024_),
    .B(_04040_));
 sg13g2_buf_1 _21310_ (.A(_03991_),
    .X(_04042_));
 sg13g2_nor2_1 _21311_ (.A(_03507_),
    .B(_03534_),
    .Y(_04043_));
 sg13g2_or3_1 _21312_ (.A(_04043_),
    .B(_03548_),
    .C(_03555_),
    .X(_04044_));
 sg13g2_a21o_1 _21313_ (.A2(_04044_),
    .A1(_03572_),
    .B1(_03551_),
    .X(_04045_));
 sg13g2_xor2_1 _21314_ (.B(_04024_),
    .A(_04045_),
    .X(_04046_));
 sg13g2_nand2b_1 _21315_ (.Y(_04047_),
    .B(_03552_),
    .A_N(_03568_));
 sg13g2_xor2_1 _21316_ (.B(_04047_),
    .A(_04043_),
    .X(_04048_));
 sg13g2_a21oi_1 _21317_ (.A1(_09652_),
    .A2(_04048_),
    .Y(_04049_),
    .B1(net223));
 sg13g2_buf_2 _21318_ (.A(_04049_),
    .X(_04050_));
 sg13g2_o21ai_1 _21319_ (.B1(net292),
    .Y(_04051_),
    .A1(_10859_),
    .A2(_11055_));
 sg13g2_o21ai_1 _21320_ (.B1(_04051_),
    .Y(_04052_),
    .A1(net171),
    .A2(_03962_));
 sg13g2_nand2_1 _21321_ (.Y(_04053_),
    .A(_11182_),
    .B(_04052_));
 sg13g2_o21ai_1 _21322_ (.B1(_04053_),
    .Y(_04054_),
    .A1(net231),
    .A2(_03948_));
 sg13g2_o21ai_1 _21323_ (.B1(_03498_),
    .Y(_04055_),
    .A1(_11175_),
    .A2(_03943_));
 sg13g2_nand2_1 _21324_ (.Y(_04056_),
    .A(_04053_),
    .B(_04055_));
 sg13g2_a22oi_1 _21325_ (.Y(_04057_),
    .B1(_04056_),
    .B2(net1043),
    .A2(_04054_),
    .A1(net1081));
 sg13g2_a21o_1 _21326_ (.A2(net120),
    .A1(_03405_),
    .B1(_04057_),
    .X(_04058_));
 sg13g2_mux2_1 _21327_ (.A0(net1011),
    .A1(net1087),
    .S(_03574_),
    .X(_04059_));
 sg13g2_inv_1 _21328_ (.Y(_04060_),
    .A(_09654_));
 sg13g2_nand2b_1 _21329_ (.Y(_04061_),
    .B(_04060_),
    .A_N(_04059_));
 sg13g2_a22oi_1 _21330_ (.Y(_04062_),
    .B1(_04023_),
    .B2(_04061_),
    .A2(net201),
    .A1(net1024));
 sg13g2_buf_1 _21331_ (.A(_03425_),
    .X(_04063_));
 sg13g2_buf_1 _21332_ (.A(_03939_),
    .X(_04064_));
 sg13g2_nor2_1 _21333_ (.A(_03943_),
    .B(_03962_),
    .Y(_04065_));
 sg13g2_buf_2 _21334_ (.A(_04065_),
    .X(_04066_));
 sg13g2_buf_1 _21335_ (.A(_04066_),
    .X(_04067_));
 sg13g2_nand3_1 _21336_ (.B(net235),
    .C(_03523_),
    .A(net290),
    .Y(_04068_));
 sg13g2_buf_1 _21337_ (.A(_04068_),
    .X(_04069_));
 sg13g2_nand3_1 _21338_ (.B(net235),
    .C(net224),
    .A(net290),
    .Y(_04070_));
 sg13g2_buf_1 _21339_ (.A(_04070_),
    .X(_04071_));
 sg13g2_buf_1 _21340_ (.A(_04071_),
    .X(_04072_));
 sg13g2_o21ai_1 _21341_ (.B1(net143),
    .Y(_04073_),
    .A1(_03537_),
    .A2(_04069_));
 sg13g2_a221oi_1 _21342_ (.B2(net146),
    .C1(_04073_),
    .B1(net118),
    .A1(net167),
    .Y(_04074_),
    .A2(net144));
 sg13g2_nor3_1 _21343_ (.A(net290),
    .B(net237),
    .C(_03962_),
    .Y(_04075_));
 sg13g2_buf_1 _21344_ (.A(_04075_),
    .X(_04076_));
 sg13g2_buf_1 _21345_ (.A(_04076_),
    .X(_04077_));
 sg13g2_a22oi_1 _21346_ (.Y(_04078_),
    .B1(net142),
    .B2(net191),
    .A2(net169),
    .A1(net222));
 sg13g2_buf_1 _21347_ (.A(_10962_),
    .X(_04079_));
 sg13g2_nor3_1 _21348_ (.A(net333),
    .B(net237),
    .C(_03930_),
    .Y(_04080_));
 sg13g2_buf_2 _21349_ (.A(_04080_),
    .X(_04081_));
 sg13g2_buf_1 _21350_ (.A(_04081_),
    .X(_04082_));
 sg13g2_a22oi_1 _21351_ (.Y(_04083_),
    .B1(net147),
    .B2(net190),
    .A2(net141),
    .A1(net221));
 sg13g2_and2_1 _21352_ (.A(_04078_),
    .B(_04083_),
    .X(_04084_));
 sg13g2_buf_1 _21353_ (.A(_03420_),
    .X(_04085_));
 sg13g2_nand2_1 _21354_ (.Y(_04086_),
    .A(net188),
    .B(net168));
 sg13g2_buf_1 _21355_ (.A(_03924_),
    .X(_04087_));
 sg13g2_a21oi_1 _21356_ (.A1(net225),
    .A2(net117),
    .Y(_04088_),
    .B1(_03947_));
 sg13g2_nand4_1 _21357_ (.B(_04084_),
    .C(_04086_),
    .A(_04074_),
    .Y(_04089_),
    .D(_04088_));
 sg13g2_nand2b_1 _21358_ (.Y(_04090_),
    .B(net120),
    .A_N(_04025_));
 sg13g2_nand3_1 _21359_ (.B(_04089_),
    .C(_04090_),
    .A(net1080),
    .Y(_04091_));
 sg13g2_nand4_1 _21360_ (.B(_04058_),
    .C(_04062_),
    .A(_04050_),
    .Y(_04092_),
    .D(_04091_));
 sg13g2_a21oi_1 _21361_ (.A1(net630),
    .A2(_04046_),
    .Y(_04093_),
    .B1(_04092_));
 sg13g2_o21ai_1 _21362_ (.B1(_04093_),
    .Y(_04094_),
    .A1(_08922_),
    .A2(_04041_));
 sg13g2_o21ai_1 _21363_ (.B1(_04094_),
    .Y(_04095_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[11] ));
 sg13g2_buf_1 _21364_ (.A(_08473_),
    .X(_04096_));
 sg13g2_nor2_2 _21365_ (.A(net884),
    .B(net765),
    .Y(_04097_));
 sg13g2_nand4_1 _21366_ (.B(_08482_),
    .C(_08435_),
    .A(net1038),
    .Y(_04098_),
    .D(_04097_));
 sg13g2_or2_1 _21367_ (.X(_04099_),
    .B(_04098_),
    .A(_08500_));
 sg13g2_buf_1 _21368_ (.A(_04099_),
    .X(_04100_));
 sg13g2_nor2_1 _21369_ (.A(net950),
    .B(_04100_),
    .Y(_04101_));
 sg13g2_nand3_1 _21370_ (.B(_08490_),
    .C(_04101_),
    .A(_08460_),
    .Y(_04102_));
 sg13g2_xnor2_1 _21371_ (.Y(_04103_),
    .A(_03465_),
    .B(_04102_));
 sg13g2_buf_1 _21372_ (.A(net35),
    .X(_04104_));
 sg13g2_a22oi_1 _21373_ (.Y(_04105_),
    .B1(_04103_),
    .B2(net32),
    .A2(net28),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_o21ai_1 _21374_ (.B1(_04105_),
    .Y(_00983_),
    .A1(net30),
    .A2(_04095_));
 sg13g2_nor2_1 _21375_ (.A(_03581_),
    .B(_03578_),
    .Y(_04106_));
 sg13g2_xnor2_1 _21376_ (.Y(_04107_),
    .A(_03486_),
    .B(_04106_));
 sg13g2_xnor2_1 _21377_ (.Y(_04108_),
    .A(_03576_),
    .B(_04106_));
 sg13g2_nand2_1 _21378_ (.Y(_04109_),
    .A(net1079),
    .B(_03578_));
 sg13g2_o21ai_1 _21379_ (.B1(_04109_),
    .Y(_04110_),
    .A1(net883),
    .A2(_03578_));
 sg13g2_nor2_1 _21380_ (.A(net1012),
    .B(_04110_),
    .Y(_04111_));
 sg13g2_or2_1 _21381_ (.X(_04112_),
    .B(_04111_),
    .A(_03581_));
 sg13g2_a21oi_1 _21382_ (.A1(_03402_),
    .A2(_03954_),
    .Y(_04113_),
    .B1(net224));
 sg13g2_o21ai_1 _21383_ (.B1(net1043),
    .Y(_04114_),
    .A1(net282),
    .A2(_03943_));
 sg13g2_o21ai_1 _21384_ (.B1(_04114_),
    .Y(_04115_),
    .A1(net283),
    .A2(_03943_));
 sg13g2_nand2_1 _21385_ (.Y(_04116_),
    .A(net192),
    .B(_04115_));
 sg13g2_o21ai_1 _21386_ (.B1(_04116_),
    .Y(_04117_),
    .A1(_03943_),
    .A2(_04113_));
 sg13g2_a21oi_1 _21387_ (.A1(_03494_),
    .A2(net120),
    .Y(_04118_),
    .B1(_03977_));
 sg13g2_a22oi_1 _21388_ (.Y(_04119_),
    .B1(_04117_),
    .B2(_04118_),
    .A2(_11167_),
    .A1(net1024));
 sg13g2_nand2_1 _21389_ (.Y(_04120_),
    .A(net225),
    .B(_03967_));
 sg13g2_nand2_1 _21390_ (.Y(_04121_),
    .A(net188),
    .B(net169));
 sg13g2_a22oi_1 _21391_ (.Y(_04122_),
    .B1(net141),
    .B2(net228),
    .A2(_03934_),
    .A1(net222));
 sg13g2_nor2_1 _21392_ (.A(net148),
    .B(_03956_),
    .Y(_04123_));
 sg13g2_a21oi_1 _21393_ (.A1(net191),
    .A2(net117),
    .Y(_04124_),
    .B1(_04123_));
 sg13g2_a22oi_1 _21394_ (.Y(_04125_),
    .B1(net144),
    .B2(net229),
    .A2(_03928_),
    .A1(net146));
 sg13g2_a21oi_1 _21395_ (.A1(_03464_),
    .A2(net118),
    .Y(_04126_),
    .B1(_03974_));
 sg13g2_nor4_1 _21396_ (.A(_11025_),
    .B(net362),
    .C(_11083_),
    .D(net237),
    .Y(_04127_));
 sg13g2_buf_2 _21397_ (.A(_04127_),
    .X(_04128_));
 sg13g2_a22oi_1 _21398_ (.Y(_04129_),
    .B1(net168),
    .B2(net167),
    .A2(_04128_),
    .A1(_04079_));
 sg13g2_and4_1 _21399_ (.A(_04124_),
    .B(_04125_),
    .C(_04126_),
    .D(_04129_),
    .X(_04130_));
 sg13g2_nand4_1 _21400_ (.B(_04121_),
    .C(_04122_),
    .A(_04120_),
    .Y(_04131_),
    .D(_04130_));
 sg13g2_nand2_1 _21401_ (.Y(_04132_),
    .A(_03468_),
    .B(net120));
 sg13g2_nand3_1 _21402_ (.B(_04131_),
    .C(_04132_),
    .A(net1080),
    .Y(_04133_));
 sg13g2_nand4_1 _21403_ (.B(_04112_),
    .C(_04119_),
    .A(_04050_),
    .Y(_04134_),
    .D(_04133_));
 sg13g2_a21oi_1 _21404_ (.A1(_04042_),
    .A2(_04108_),
    .Y(_04135_),
    .B1(_04134_));
 sg13g2_o21ai_1 _21405_ (.B1(_04135_),
    .Y(_04136_),
    .A1(_08922_),
    .A2(_04107_));
 sg13g2_o21ai_1 _21406_ (.B1(_04136_),
    .Y(_04137_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[12] ));
 sg13g2_nor2_1 _21407_ (.A(_08446_),
    .B(_04102_),
    .Y(_04138_));
 sg13g2_xnor2_1 _21408_ (.Y(_04139_),
    .A(_00289_),
    .B(_04138_));
 sg13g2_a22oi_1 _21409_ (.Y(_04140_),
    .B1(_04139_),
    .B2(net32),
    .A2(net28),
    .A1(net769));
 sg13g2_o21ai_1 _21410_ (.B1(_04140_),
    .Y(_00984_),
    .A1(net30),
    .A2(_04137_));
 sg13g2_buf_1 _21411_ (.A(net223),
    .X(_04141_));
 sg13g2_xnor2_1 _21412_ (.Y(_04142_),
    .A(net199),
    .B(net171));
 sg13g2_nor4_1 _21413_ (.A(_03468_),
    .B(_04038_),
    .C(_04039_),
    .D(_04142_),
    .Y(_04143_));
 sg13g2_nor4_1 _21414_ (.A(_11426_),
    .B(_04038_),
    .C(_04039_),
    .D(_04142_),
    .Y(_04144_));
 sg13g2_or3_1 _21415_ (.A(_03485_),
    .B(_04143_),
    .C(_04144_),
    .X(_04145_));
 sg13g2_nand2_1 _21416_ (.Y(_04146_),
    .A(net200),
    .B(_03405_));
 sg13g2_a21o_1 _21417_ (.A2(_03927_),
    .A1(net149),
    .B1(_03974_),
    .X(_04147_));
 sg13g2_nor2_1 _21418_ (.A(_10981_),
    .B(net289),
    .Y(_04148_));
 sg13g2_a21oi_1 _21419_ (.A1(net293),
    .A2(net289),
    .Y(_04149_),
    .B1(_04148_));
 sg13g2_nand3_1 _21420_ (.B(net224),
    .C(_04149_),
    .A(net201),
    .Y(_04150_));
 sg13g2_a21oi_1 _21421_ (.A1(net228),
    .A2(_04128_),
    .Y(_04151_),
    .B1(_03957_));
 sg13g2_nand2_1 _21422_ (.Y(_04152_),
    .A(_04150_),
    .B(_04151_));
 sg13g2_nand2_1 _21423_ (.Y(_04153_),
    .A(_03420_),
    .B(_03934_));
 sg13g2_a22oi_1 _21424_ (.Y(_04154_),
    .B1(_03964_),
    .B2(net229),
    .A2(_03924_),
    .A1(_10999_));
 sg13g2_a22oi_1 _21425_ (.Y(_04155_),
    .B1(_04066_),
    .B2(net189),
    .A2(_03966_),
    .A1(net191));
 sg13g2_a22oi_1 _21426_ (.Y(_04156_),
    .B1(net169),
    .B2(_03425_),
    .A2(_04081_),
    .A1(net172));
 sg13g2_nand4_1 _21427_ (.B(_04154_),
    .C(_04155_),
    .A(_04153_),
    .Y(_04157_),
    .D(_04156_));
 sg13g2_nor3_1 _21428_ (.A(_04147_),
    .B(_04152_),
    .C(_04157_),
    .Y(_04158_));
 sg13g2_o21ai_1 _21429_ (.B1(net1080),
    .Y(_04159_),
    .A1(_03489_),
    .A2(net143));
 sg13g2_nor2_1 _21430_ (.A(net200),
    .B(_03405_),
    .Y(_04160_));
 sg13g2_a21oi_1 _21431_ (.A1(_03485_),
    .A2(_04146_),
    .Y(_04161_),
    .B1(_04160_));
 sg13g2_o21ai_1 _21432_ (.B1(net883),
    .Y(_04162_),
    .A1(_08922_),
    .A2(_04161_));
 sg13g2_a22oi_1 _21433_ (.Y(_04163_),
    .B1(_04066_),
    .B2(net239),
    .A2(_03974_),
    .A1(_10859_));
 sg13g2_nand2b_1 _21434_ (.Y(_04164_),
    .B(net1081),
    .A_N(_04163_));
 sg13g2_a221oi_1 _21435_ (.B2(net1088),
    .C1(net630),
    .B1(net295),
    .A1(_09654_),
    .Y(_04165_),
    .A2(_11472_));
 sg13g2_nor2_1 _21436_ (.A(_10859_),
    .B(_04071_),
    .Y(_04166_));
 sg13g2_a21oi_1 _21437_ (.A1(net231),
    .A2(_04071_),
    .Y(_04167_),
    .B1(_04166_));
 sg13g2_a21o_1 _21438_ (.A2(_10315_),
    .A1(net1079),
    .B1(_09654_),
    .X(_04168_));
 sg13g2_buf_1 _21439_ (.A(_10925_),
    .X(_04169_));
 sg13g2_a22oi_1 _21440_ (.Y(_04170_),
    .B1(_04168_),
    .B2(net166),
    .A2(_04167_),
    .A1(net1043));
 sg13g2_nand3_1 _21441_ (.B(_04165_),
    .C(_04170_),
    .A(_04164_),
    .Y(_04171_));
 sg13g2_a21oi_1 _21442_ (.A1(_04142_),
    .A2(_04162_),
    .Y(_04172_),
    .B1(_04171_));
 sg13g2_o21ai_1 _21443_ (.B1(_04172_),
    .Y(_04173_),
    .A1(_04158_),
    .A2(_04159_));
 sg13g2_a21oi_1 _21444_ (.A1(_09652_),
    .A2(_04048_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_and2_1 _21445_ (.A(_04146_),
    .B(_04174_),
    .X(_04175_));
 sg13g2_nand2_1 _21446_ (.Y(_04176_),
    .A(_03470_),
    .B(_04146_));
 sg13g2_or3_1 _21447_ (.A(_04038_),
    .B(_04039_),
    .C(_04176_),
    .X(_04177_));
 sg13g2_buf_1 _21448_ (.A(net1086),
    .X(_04178_));
 sg13g2_o21ai_1 _21449_ (.B1(net949),
    .Y(_04179_),
    .A1(_11450_),
    .A2(_03405_));
 sg13g2_a21o_1 _21450_ (.A2(_04177_),
    .A1(_04142_),
    .B1(_04179_),
    .X(_04180_));
 sg13g2_inv_1 _21451_ (.Y(_04181_),
    .A(_03578_));
 sg13g2_o21ai_1 _21452_ (.B1(_04181_),
    .Y(_04182_),
    .A1(_03581_),
    .A2(_03576_));
 sg13g2_xnor2_1 _21453_ (.Y(_04183_),
    .A(_04182_),
    .B(_04142_));
 sg13g2_a21o_1 _21454_ (.A2(_04183_),
    .A1(_04042_),
    .B1(net187),
    .X(_04184_));
 sg13g2_a221oi_1 _21455_ (.B2(_04174_),
    .C1(_04184_),
    .B1(_04180_),
    .A1(_04145_),
    .Y(_04185_),
    .A2(_04175_));
 sg13g2_a21oi_1 _21456_ (.A1(net187),
    .A2(\cpu.ex.c_mult[13] ),
    .Y(_04186_),
    .B1(_04185_));
 sg13g2_nand2_1 _21457_ (.Y(_04187_),
    .A(net769),
    .B(_04138_));
 sg13g2_xor2_1 _21458_ (.B(_04187_),
    .A(_00196_),
    .X(_04188_));
 sg13g2_a22oi_1 _21459_ (.Y(_04189_),
    .B1(_04188_),
    .B2(net32),
    .A2(net28),
    .A1(net768));
 sg13g2_o21ai_1 _21460_ (.B1(_04189_),
    .Y(_00985_),
    .A1(net30),
    .A2(_04186_));
 sg13g2_xor2_1 _21461_ (.B(net194),
    .A(_10269_),
    .X(_04190_));
 sg13g2_buf_1 _21462_ (.A(_04190_),
    .X(_04191_));
 sg13g2_xor2_1 _21463_ (.B(_04191_),
    .A(_03585_),
    .X(_04192_));
 sg13g2_or2_1 _21464_ (.X(_04193_),
    .B(_03492_),
    .A(_03496_));
 sg13g2_nand3_1 _21465_ (.B(_03495_),
    .C(_04191_),
    .A(_03492_),
    .Y(_04194_));
 sg13g2_o21ai_1 _21466_ (.B1(_04194_),
    .Y(_04195_),
    .A1(_04191_),
    .A2(_04193_));
 sg13g2_nand2_2 _21467_ (.Y(_04196_),
    .A(_08051_),
    .B(_10903_));
 sg13g2_nand2_1 _21468_ (.Y(_04197_),
    .A(_03496_),
    .B(_04191_));
 sg13g2_o21ai_1 _21469_ (.B1(_04197_),
    .Y(_04198_),
    .A1(_03495_),
    .A2(_04191_));
 sg13g2_a22oi_1 _21470_ (.Y(_04199_),
    .B1(_04149_),
    .B2(net201),
    .A2(_03922_),
    .A1(_03453_));
 sg13g2_nor2_1 _21471_ (.A(net283),
    .B(_03984_),
    .Y(_04200_));
 sg13g2_a21oi_1 _21472_ (.A1(net283),
    .A2(_04063_),
    .Y(_04201_),
    .B1(_04200_));
 sg13g2_nor3_1 _21473_ (.A(net362),
    .B(_03932_),
    .C(_04201_),
    .Y(_04202_));
 sg13g2_nand2_1 _21474_ (.Y(_04203_),
    .A(_11175_),
    .B(_03935_));
 sg13g2_buf_1 _21475_ (.A(_04128_),
    .X(_04204_));
 sg13g2_a21oi_1 _21476_ (.A1(net146),
    .A2(net140),
    .Y(_04205_),
    .B1(_03975_));
 sg13g2_o21ai_1 _21477_ (.B1(_04205_),
    .Y(_04206_),
    .A1(_03505_),
    .A2(_04203_));
 sg13g2_nand2_1 _21478_ (.Y(_04207_),
    .A(_03523_),
    .B(_03922_));
 sg13g2_nor2_1 _21479_ (.A(_03456_),
    .B(_04207_),
    .Y(_04208_));
 sg13g2_a21o_1 _21480_ (.A2(net144),
    .A1(_03529_),
    .B1(_04208_),
    .X(_04209_));
 sg13g2_nand2_1 _21481_ (.Y(_04210_),
    .A(net193),
    .B(net118));
 sg13g2_nand2_1 _21482_ (.Y(_04211_),
    .A(net119),
    .B(net141));
 sg13g2_a22oi_1 _21483_ (.Y(_04212_),
    .B1(net169),
    .B2(net190),
    .A2(net170),
    .A1(net189));
 sg13g2_nand3_1 _21484_ (.B(_04211_),
    .C(_04212_),
    .A(_04210_),
    .Y(_04213_));
 sg13g2_nor4_1 _21485_ (.A(_04202_),
    .B(_04206_),
    .C(_04209_),
    .D(_04213_),
    .Y(_04214_));
 sg13g2_o21ai_1 _21486_ (.B1(_04214_),
    .Y(_04215_),
    .A1(_03962_),
    .A2(_04199_));
 sg13g2_a21oi_1 _21487_ (.A1(_03494_),
    .A2(_03976_),
    .Y(_04216_),
    .B1(_09662_));
 sg13g2_a21oi_1 _21488_ (.A1(net178),
    .A2(net173),
    .Y(_04217_),
    .B1(net883));
 sg13g2_and3_1 _21489_ (.X(_04218_),
    .A(_09673_),
    .B(net178),
    .C(net173));
 sg13g2_nor3_1 _21490_ (.A(_09655_),
    .B(_04217_),
    .C(_04218_),
    .Y(_04219_));
 sg13g2_nor2_1 _21491_ (.A(net178),
    .B(net173),
    .Y(_04220_));
 sg13g2_nor2b_1 _21492_ (.A(net231),
    .B_N(net1081),
    .Y(_04221_));
 sg13g2_a22oi_1 _21493_ (.Y(_04222_),
    .B1(_03976_),
    .B2(_04221_),
    .A2(_10435_),
    .A1(net1024));
 sg13g2_o21ai_1 _21494_ (.B1(_04222_),
    .Y(_04223_),
    .A1(_04219_),
    .A2(_04220_));
 sg13g2_a221oi_1 _21495_ (.B2(_04216_),
    .C1(_04223_),
    .B1(_04215_),
    .A1(net949),
    .Y(_04224_),
    .A2(_04198_));
 sg13g2_nand3_1 _21496_ (.B(_04050_),
    .C(_04224_),
    .A(_04196_),
    .Y(_04225_));
 sg13g2_a221oi_1 _21497_ (.B2(net949),
    .C1(_04225_),
    .B1(_04195_),
    .A1(net630),
    .Y(_04226_),
    .A2(_04192_));
 sg13g2_inv_1 _21498_ (.Y(_04227_),
    .A(_03913_));
 sg13g2_o21ai_1 _21499_ (.B1(_04227_),
    .Y(_04228_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_nand3_1 _21500_ (.B(net768),
    .C(_04138_),
    .A(net769),
    .Y(_04229_));
 sg13g2_xnor2_1 _21501_ (.Y(_04230_),
    .A(_10831_),
    .B(_04229_));
 sg13g2_a22oi_1 _21502_ (.Y(_04231_),
    .B1(_04230_),
    .B2(net32),
    .A2(_04021_),
    .A1(_08184_));
 sg13g2_o21ai_1 _21503_ (.B1(_04231_),
    .Y(_00986_),
    .A1(_04226_),
    .A2(_04228_));
 sg13g2_nor2_1 _21504_ (.A(_10275_),
    .B(net231),
    .Y(_04232_));
 sg13g2_nor2_2 _21505_ (.A(_04232_),
    .B(_03591_),
    .Y(_04233_));
 sg13g2_xnor2_1 _21506_ (.Y(_04234_),
    .A(_03590_),
    .B(_04233_));
 sg13g2_nor2b_1 _21507_ (.A(_11497_),
    .B_N(net173),
    .Y(_04235_));
 sg13g2_nor2_1 _21508_ (.A(_04235_),
    .B(_04233_),
    .Y(_04236_));
 sg13g2_nor2b_1 _21509_ (.A(_03401_),
    .B_N(_04233_),
    .Y(_04237_));
 sg13g2_nor2_1 _21510_ (.A(_03496_),
    .B(_03485_),
    .Y(_04238_));
 sg13g2_inv_1 _21511_ (.Y(_04239_),
    .A(_04238_));
 sg13g2_nor4_1 _21512_ (.A(_11476_),
    .B(_03479_),
    .C(_03484_),
    .D(_04239_),
    .Y(_04240_));
 sg13g2_nor4_1 _21513_ (.A(net193),
    .B(_03479_),
    .C(_03484_),
    .D(_04239_),
    .Y(_04241_));
 sg13g2_o21ai_1 _21514_ (.B1(_03495_),
    .Y(_04242_),
    .A1(_03496_),
    .A2(_04146_));
 sg13g2_nor3_1 _21515_ (.A(_04240_),
    .B(_04241_),
    .C(_04242_),
    .Y(_04243_));
 sg13g2_mux2_1 _21516_ (.A0(_04236_),
    .A1(_04237_),
    .S(_04243_),
    .X(_04244_));
 sg13g2_mux2_1 _21517_ (.A0(_03401_),
    .A1(_04235_),
    .S(_04233_),
    .X(_04245_));
 sg13g2_nand2_1 _21518_ (.Y(_04246_),
    .A(net883),
    .B(_03502_));
 sg13g2_o21ai_1 _21519_ (.B1(_04246_),
    .Y(_04247_),
    .A1(net1011),
    .A2(_03502_));
 sg13g2_a21oi_1 _21520_ (.A1(_04060_),
    .A2(_04247_),
    .Y(_04248_),
    .B1(_03591_));
 sg13g2_a221oi_1 _21521_ (.B2(net949),
    .C1(_04248_),
    .B1(_04245_),
    .A1(net1024),
    .Y(_04249_),
    .A2(net240));
 sg13g2_nor2_1 _21522_ (.A(net293),
    .B(_11025_),
    .Y(_04250_));
 sg13g2_nor2_1 _21523_ (.A(net292),
    .B(net289),
    .Y(_04251_));
 sg13g2_a22oi_1 _21524_ (.Y(_04252_),
    .B1(_04251_),
    .B2(net191),
    .A2(_04250_),
    .A1(net289));
 sg13g2_nor3_1 _21525_ (.A(net282),
    .B(net202),
    .C(_04252_),
    .Y(_04253_));
 sg13g2_a22oi_1 _21526_ (.Y(_04254_),
    .B1(net169),
    .B2(net225),
    .A2(_04082_),
    .A1(_03961_));
 sg13g2_nand2_1 _21527_ (.Y(_04255_),
    .A(_10877_),
    .B(_03928_));
 sg13g2_a22oi_1 _21528_ (.Y(_04256_),
    .B1(net142),
    .B2(net146),
    .A2(_03934_),
    .A1(net190));
 sg13g2_a22oi_1 _21529_ (.Y(_04257_),
    .B1(_04067_),
    .B2(net166),
    .A2(net147),
    .A1(net221));
 sg13g2_nand4_1 _21530_ (.B(_04255_),
    .C(_04256_),
    .A(_04254_),
    .Y(_04258_),
    .D(_04257_));
 sg13g2_nand2_1 _21531_ (.Y(_04259_),
    .A(net167),
    .B(net224));
 sg13g2_nand2_1 _21532_ (.Y(_04260_),
    .A(net188),
    .B(_03954_));
 sg13g2_a21oi_1 _21533_ (.A1(_04259_),
    .A2(_04260_),
    .Y(_04261_),
    .B1(_03932_));
 sg13g2_nand2_1 _21534_ (.Y(_04262_),
    .A(_10999_),
    .B(net144));
 sg13g2_a21oi_1 _21535_ (.A1(net119),
    .A2(net140),
    .Y(_04263_),
    .B1(_03975_));
 sg13g2_nand3_1 _21536_ (.B(_04262_),
    .C(_04263_),
    .A(_03925_),
    .Y(_04264_));
 sg13g2_nor4_1 _21537_ (.A(_04253_),
    .B(_04258_),
    .C(_04261_),
    .D(_04264_),
    .Y(_04265_));
 sg13g2_or3_1 _21538_ (.A(_09662_),
    .B(_04166_),
    .C(_04265_),
    .X(_04266_));
 sg13g2_nand4_1 _21539_ (.B(_04050_),
    .C(_04249_),
    .A(_04196_),
    .Y(_04267_),
    .D(_04266_));
 sg13g2_a221oi_1 _21540_ (.B2(net949),
    .C1(_04267_),
    .B1(_04244_),
    .A1(net630),
    .Y(_04268_),
    .A2(_04234_));
 sg13g2_nand4_1 _21541_ (.B(_11541_),
    .C(_11544_),
    .A(net187),
    .Y(_04269_),
    .D(_11546_));
 sg13g2_nand2b_1 _21542_ (.Y(_04270_),
    .B(_04269_),
    .A_N(_04268_));
 sg13g2_or2_1 _21543_ (.X(_04271_),
    .B(_04229_),
    .A(_08344_));
 sg13g2_xnor2_1 _21544_ (.Y(_04272_),
    .A(_10900_),
    .B(_04271_));
 sg13g2_a22oi_1 _21545_ (.Y(_04273_),
    .B1(_04272_),
    .B2(_04104_),
    .A2(_04021_),
    .A1(net1094));
 sg13g2_o21ai_1 _21546_ (.B1(_04273_),
    .Y(_00987_),
    .A1(net30),
    .A2(_04270_));
 sg13g2_and3_1 _21547_ (.X(_04274_),
    .A(_08967_),
    .B(net253),
    .C(_11212_));
 sg13g2_a21oi_1 _21548_ (.A1(net764),
    .A2(net35),
    .Y(_04275_),
    .B1(_04020_));
 sg13g2_a21oi_1 _21549_ (.A1(net885),
    .A2(net35),
    .Y(_04276_),
    .B1(_08282_));
 sg13g2_a21oi_1 _21550_ (.A1(net770),
    .A2(_04275_),
    .Y(_04277_),
    .B1(_04276_));
 sg13g2_nand2_1 _21551_ (.Y(_04278_),
    .A(_03916_),
    .B(_03917_));
 sg13g2_nand3_1 _21552_ (.B(net202),
    .C(_04251_),
    .A(_03926_),
    .Y(_04279_));
 sg13g2_a21oi_1 _21553_ (.A1(_04278_),
    .A2(_04279_),
    .Y(_04280_),
    .B1(_03656_));
 sg13g2_a22oi_1 _21554_ (.Y(_04281_),
    .B1(_03952_),
    .B2(net166),
    .A2(_04064_),
    .A1(net189));
 sg13g2_a22oi_1 _21555_ (.Y(_04282_),
    .B1(net142),
    .B2(net228),
    .A2(_03934_),
    .A1(net194));
 sg13g2_nand2_1 _21556_ (.Y(_04283_),
    .A(_04281_),
    .B(_04282_));
 sg13g2_nand2_1 _21557_ (.Y(_04284_),
    .A(net146),
    .B(net117));
 sg13g2_nand3_1 _21558_ (.B(_03916_),
    .C(net224),
    .A(net192),
    .Y(_04285_));
 sg13g2_nor2_1 _21559_ (.A(_03432_),
    .B(_04069_),
    .Y(_04286_));
 sg13g2_a21oi_1 _21560_ (.A1(net193),
    .A2(net168),
    .Y(_04287_),
    .B1(_04286_));
 sg13g2_nor2_1 _21561_ (.A(net148),
    .B(_03948_),
    .Y(_04288_));
 sg13g2_a221oi_1 _21562_ (.B2(net119),
    .C1(_04288_),
    .B1(net147),
    .A1(_04079_),
    .Y(_04289_),
    .A2(_04204_));
 sg13g2_nand4_1 _21563_ (.B(_04285_),
    .C(_04287_),
    .A(_04284_),
    .Y(_04290_),
    .D(_04289_));
 sg13g2_nor4_1 _21564_ (.A(_03945_),
    .B(_04280_),
    .C(_04283_),
    .D(_04290_),
    .Y(_04291_));
 sg13g2_or2_1 _21565_ (.X(_04292_),
    .B(net1081),
    .A(_08052_));
 sg13g2_buf_1 _21566_ (.A(_04292_),
    .X(_04293_));
 sg13g2_o21ai_1 _21567_ (.B1(_04293_),
    .Y(_04294_),
    .A1(net190),
    .A2(net143));
 sg13g2_and2_1 _21568_ (.A(_03422_),
    .B(_03423_),
    .X(_04295_));
 sg13g2_buf_1 _21569_ (.A(_04295_),
    .X(_04296_));
 sg13g2_nand2_1 _21570_ (.Y(_04297_),
    .A(_11254_),
    .B(_03972_));
 sg13g2_nand2_1 _21571_ (.Y(_04298_),
    .A(net289),
    .B(_03425_));
 sg13g2_nand2_1 _21572_ (.Y(_04299_),
    .A(_04297_),
    .B(_04298_));
 sg13g2_xnor2_1 _21573_ (.Y(_04300_),
    .A(_04296_),
    .B(_04299_));
 sg13g2_nand2_1 _21574_ (.Y(_04301_),
    .A(_03521_),
    .B(_03524_));
 sg13g2_xnor2_1 _21575_ (.Y(_04302_),
    .A(_04301_),
    .B(_04299_));
 sg13g2_nor2_1 _21576_ (.A(net1079),
    .B(_04298_),
    .Y(_04303_));
 sg13g2_a21oi_1 _21577_ (.A1(_08841_),
    .A2(_04298_),
    .Y(_04304_),
    .B1(_04303_));
 sg13g2_o21ai_1 _21578_ (.B1(_04297_),
    .Y(_04305_),
    .A1(net1012),
    .A2(_04304_));
 sg13g2_nand2_1 _21579_ (.Y(_04306_),
    .A(_03997_),
    .B(_04067_));
 sg13g2_o21ai_1 _21580_ (.B1(_04306_),
    .Y(_04307_),
    .A1(_03984_),
    .A2(net143));
 sg13g2_nand2_1 _21581_ (.Y(_04308_),
    .A(net1080),
    .B(_04307_));
 sg13g2_a21oi_1 _21582_ (.A1(net1088),
    .A2(_10184_),
    .Y(_04309_),
    .B1(net223));
 sg13g2_nand3_1 _21583_ (.B(_04308_),
    .C(_04309_),
    .A(_04305_),
    .Y(_04310_));
 sg13g2_a221oi_1 _21584_ (.B2(_03995_),
    .C1(_04310_),
    .B1(_04302_),
    .A1(_08921_),
    .Y(_04311_),
    .A2(_04300_));
 sg13g2_o21ai_1 _21585_ (.B1(_04311_),
    .Y(_04312_),
    .A1(_04291_),
    .A2(_04294_));
 sg13g2_o21ai_1 _21586_ (.B1(_04312_),
    .Y(_04313_),
    .A1(_03915_),
    .A2(\cpu.ex.c_mult[2] ));
 sg13g2_nor2_1 _21587_ (.A(_03913_),
    .B(_04313_),
    .Y(_04314_));
 sg13g2_or3_1 _21588_ (.A(_04274_),
    .B(_04277_),
    .C(_04314_),
    .X(_00988_));
 sg13g2_nor2_1 _21589_ (.A(net225),
    .B(net143),
    .Y(_04315_));
 sg13g2_o21ai_1 _21590_ (.B1(_11183_),
    .Y(_04316_),
    .A1(_11175_),
    .A2(_03932_));
 sg13g2_a22oi_1 _21591_ (.Y(_04317_),
    .B1(_04077_),
    .B2(_03968_),
    .A2(net140),
    .A1(net228));
 sg13g2_a22oi_1 _21592_ (.Y(_04318_),
    .B1(net168),
    .B2(_04169_),
    .A2(_03934_),
    .A1(net192));
 sg13g2_o21ai_1 _21593_ (.B1(_04071_),
    .Y(_04319_),
    .A1(net148),
    .A2(_04069_));
 sg13g2_a221oi_1 _21594_ (.B2(net194),
    .C1(_04319_),
    .B1(net169),
    .A1(net221),
    .Y(_04320_),
    .A2(_04081_));
 sg13g2_a22oi_1 _21595_ (.Y(_04321_),
    .B1(_03939_),
    .B2(_10877_),
    .A2(_03924_),
    .A1(net149));
 sg13g2_a22oi_1 _21596_ (.Y(_04322_),
    .B1(_04066_),
    .B2(_03529_),
    .A2(_03966_),
    .A1(_03561_));
 sg13g2_and2_1 _21597_ (.A(_04321_),
    .B(_04322_),
    .X(_04323_));
 sg13g2_nand4_1 _21598_ (.B(_04318_),
    .C(_04320_),
    .A(_04317_),
    .Y(_04324_),
    .D(_04323_));
 sg13g2_a21oi_1 _21599_ (.A1(net192),
    .A2(_04316_),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_a21oi_1 _21600_ (.A1(net1081),
    .A2(_04324_),
    .Y(_04326_),
    .B1(net1043));
 sg13g2_nor3_1 _21601_ (.A(_04315_),
    .B(_04325_),
    .C(_04326_),
    .Y(_04327_));
 sg13g2_o21ai_1 _21602_ (.B1(net1087),
    .Y(_04328_),
    .A1(net202),
    .A2(_03513_));
 sg13g2_nand3_1 _21603_ (.B(net201),
    .C(_03919_),
    .A(net1079),
    .Y(_04329_));
 sg13g2_nand3_1 _21604_ (.B(_04328_),
    .C(_04329_),
    .A(_04060_),
    .Y(_04330_));
 sg13g2_o21ai_1 _21605_ (.B1(_04330_),
    .Y(_04331_),
    .A1(net201),
    .A2(_03919_));
 sg13g2_a21oi_1 _21606_ (.A1(net1088),
    .A2(_11426_),
    .Y(_04332_),
    .B1(_03982_));
 sg13g2_a21oi_1 _21607_ (.A1(net283),
    .A2(_04085_),
    .Y(_04333_),
    .B1(_04250_));
 sg13g2_o21ai_1 _21608_ (.B1(_04259_),
    .Y(_04334_),
    .A1(_03656_),
    .A2(_04333_));
 sg13g2_nand3_1 _21609_ (.B(_11182_),
    .C(_04334_),
    .A(net1080),
    .Y(_04335_));
 sg13g2_nand3_1 _21610_ (.B(_04332_),
    .C(_04335_),
    .A(_04331_),
    .Y(_04336_));
 sg13g2_nor2_1 _21611_ (.A(_04327_),
    .B(_04336_),
    .Y(_04337_));
 sg13g2_o21ai_1 _21612_ (.B1(_04296_),
    .Y(_04338_),
    .A1(net289),
    .A2(_03972_));
 sg13g2_o21ai_1 _21613_ (.B1(_04338_),
    .Y(_04339_),
    .A1(net290),
    .A2(_04063_));
 sg13g2_xnor2_1 _21614_ (.Y(_04340_),
    .A(net201),
    .B(_03513_));
 sg13g2_xor2_1 _21615_ (.B(_04340_),
    .A(_04339_),
    .X(_04341_));
 sg13g2_inv_1 _21616_ (.Y(_04342_),
    .A(_04298_));
 sg13g2_a21oi_1 _21617_ (.A1(_04297_),
    .A2(_04301_),
    .Y(_04343_),
    .B1(_04342_));
 sg13g2_xnor2_1 _21618_ (.Y(_04344_),
    .A(_04340_),
    .B(_04343_));
 sg13g2_a22oi_1 _21619_ (.Y(_04345_),
    .B1(_04344_),
    .B2(_03995_),
    .A2(_04341_),
    .A1(_04178_));
 sg13g2_a22oi_1 _21620_ (.Y(_04346_),
    .B1(_04337_),
    .B2(_04345_),
    .A2(_11288_),
    .A1(net187));
 sg13g2_nand2_1 _21621_ (.Y(_04347_),
    .A(_08282_),
    .B(net885));
 sg13g2_a21oi_1 _21622_ (.A1(net35),
    .A2(_04347_),
    .Y(_04348_),
    .B1(_04020_));
 sg13g2_inv_1 _21623_ (.Y(_04349_),
    .A(_00274_));
 sg13g2_nor2_1 _21624_ (.A(net703),
    .B(_04347_),
    .Y(_04350_));
 sg13g2_a221oi_1 _21625_ (.B2(_04010_),
    .C1(_04017_),
    .B1(_04350_),
    .A1(_04349_),
    .Y(_04351_),
    .A2(_04274_));
 sg13g2_o21ai_1 _21626_ (.B1(_04351_),
    .Y(_04352_),
    .A1(_08090_),
    .A2(_04348_));
 sg13g2_a21o_1 _21627_ (.A2(_04346_),
    .A1(_04227_),
    .B1(_04352_),
    .X(_00989_));
 sg13g2_a221oi_1 _21628_ (.B2(_03426_),
    .C1(_03411_),
    .B1(_04296_),
    .A1(net201),
    .Y(_04353_),
    .A2(_03513_));
 sg13g2_nand2_1 _21629_ (.Y(_04354_),
    .A(_03518_),
    .B(_03517_));
 sg13g2_xor2_1 _21630_ (.B(_04354_),
    .A(_04353_),
    .X(_04355_));
 sg13g2_o21ai_1 _21631_ (.B1(_03513_),
    .Y(_04356_),
    .A1(net202),
    .A2(_04343_));
 sg13g2_nand2_1 _21632_ (.Y(_04357_),
    .A(_11273_),
    .B(_04343_));
 sg13g2_nand2_1 _21633_ (.Y(_04358_),
    .A(_04356_),
    .B(_04357_));
 sg13g2_xor2_1 _21634_ (.B(_04358_),
    .A(_04354_),
    .X(_04359_));
 sg13g2_and2_1 _21635_ (.A(_10999_),
    .B(_04066_),
    .X(_04360_));
 sg13g2_a221oi_1 _21636_ (.B2(net119),
    .C1(_04360_),
    .B1(_04077_),
    .A1(net166),
    .Y(_04361_),
    .A2(net144));
 sg13g2_a22oi_1 _21637_ (.Y(_04362_),
    .B1(_03966_),
    .B2(net193),
    .A2(net168),
    .A1(_10859_));
 sg13g2_a22oi_1 _21638_ (.Y(_04363_),
    .B1(net169),
    .B2(net239),
    .A2(net170),
    .A1(net221));
 sg13g2_and2_1 _21639_ (.A(_04362_),
    .B(_04363_),
    .X(_04364_));
 sg13g2_a21oi_1 _21640_ (.A1(_11183_),
    .A2(_03932_),
    .Y(_04365_),
    .B1(_04196_));
 sg13g2_a221oi_1 _21641_ (.B2(net228),
    .C1(_04365_),
    .B1(net141),
    .A1(_03961_),
    .Y(_04366_),
    .A2(_04087_));
 sg13g2_nand4_1 _21642_ (.B(_04361_),
    .C(_04364_),
    .A(_04205_),
    .Y(_04367_),
    .D(_04366_));
 sg13g2_nand2_1 _21643_ (.Y(_04368_),
    .A(_03432_),
    .B(net145));
 sg13g2_nand3_1 _21644_ (.B(_04367_),
    .C(_04368_),
    .A(_04293_),
    .Y(_04369_));
 sg13g2_nand2_1 _21645_ (.Y(_04370_),
    .A(_03425_),
    .B(_04066_));
 sg13g2_o21ai_1 _21646_ (.B1(_04370_),
    .Y(_04371_),
    .A1(_03984_),
    .A2(_04069_));
 sg13g2_o21ai_1 _21647_ (.B1(net143),
    .Y(_04372_),
    .A1(net293),
    .A2(_03948_));
 sg13g2_o21ai_1 _21648_ (.B1(net1080),
    .Y(_04373_),
    .A1(net190),
    .A2(_04072_));
 sg13g2_inv_1 _21649_ (.Y(_04374_),
    .A(_04373_));
 sg13g2_o21ai_1 _21650_ (.B1(_04374_),
    .Y(_04375_),
    .A1(_04371_),
    .A2(_04372_));
 sg13g2_nor2_1 _21651_ (.A(net1079),
    .B(_03518_),
    .Y(_04376_));
 sg13g2_a21oi_1 _21652_ (.A1(net883),
    .A2(_03518_),
    .Y(_04377_),
    .B1(_04376_));
 sg13g2_o21ai_1 _21653_ (.B1(_03517_),
    .Y(_04378_),
    .A1(net1012),
    .A2(_04377_));
 sg13g2_a21oi_1 _21654_ (.A1(_08762_),
    .A2(_11450_),
    .Y(_04379_),
    .B1(net223));
 sg13g2_nand4_1 _21655_ (.B(_04375_),
    .C(_04378_),
    .A(_04369_),
    .Y(_04380_),
    .D(_04379_));
 sg13g2_a221oi_1 _21656_ (.B2(_03995_),
    .C1(_04380_),
    .B1(_04359_),
    .A1(_04178_),
    .Y(_04381_),
    .A2(_04355_));
 sg13g2_a21o_1 _21657_ (.A2(_11306_),
    .A1(_04141_),
    .B1(_04381_),
    .X(_04382_));
 sg13g2_nand2_1 _21658_ (.Y(_04383_),
    .A(net885),
    .B(net696));
 sg13g2_a21o_1 _21659_ (.A2(_04383_),
    .A1(_04010_),
    .B1(_04020_),
    .X(_04384_));
 sg13g2_nor2_1 _21660_ (.A(net1038),
    .B(_04383_),
    .Y(_04385_));
 sg13g2_nor4_1 _21661_ (.A(net1091),
    .B(net253),
    .C(net877),
    .D(_04013_),
    .Y(_04386_));
 sg13g2_a221oi_1 _21662_ (.B2(net35),
    .C1(_04386_),
    .B1(_04385_),
    .A1(net1038),
    .Y(_04387_),
    .A2(_04384_));
 sg13g2_o21ai_1 _21663_ (.B1(_04387_),
    .Y(_00990_),
    .A1(_03914_),
    .A2(_04382_));
 sg13g2_nor2_1 _21664_ (.A(net1011),
    .B(_03530_),
    .Y(_04388_));
 sg13g2_a21oi_1 _21665_ (.A1(net883),
    .A2(_03530_),
    .Y(_04389_),
    .B1(_04388_));
 sg13g2_o21ai_1 _21666_ (.B1(_03531_),
    .Y(_04390_),
    .A1(net1012),
    .A2(_04389_));
 sg13g2_a22oi_1 _21667_ (.Y(_04391_),
    .B1(net142),
    .B2(net189),
    .A2(net140),
    .A1(_04025_));
 sg13g2_a22oi_1 _21668_ (.Y(_04392_),
    .B1(net168),
    .B2(_03498_),
    .A2(net117),
    .A1(net193));
 sg13g2_a221oi_1 _21669_ (.B2(_03968_),
    .C1(_04073_),
    .B1(net141),
    .A1(net194),
    .Y(_04393_),
    .A2(net144));
 sg13g2_and3_1 _21670_ (.X(_04394_),
    .A(_04391_),
    .B(_04392_),
    .C(_04393_));
 sg13g2_nand2_1 _21671_ (.Y(_04395_),
    .A(net237),
    .B(_11132_));
 sg13g2_a21oi_1 _21672_ (.A1(_11183_),
    .A2(_04395_),
    .Y(_04396_),
    .B1(_04196_));
 sg13g2_a221oi_1 _21673_ (.B2(net221),
    .C1(_04396_),
    .B1(net118),
    .A1(_04169_),
    .Y(_04397_),
    .A2(net147));
 sg13g2_a221oi_1 _21674_ (.B2(_04397_),
    .C1(_03977_),
    .B1(_04394_),
    .A1(net148),
    .Y(_04398_),
    .A2(net145));
 sg13g2_a22oi_1 _21675_ (.Y(_04399_),
    .B1(net118),
    .B2(net229),
    .A2(net141),
    .A1(net188));
 sg13g2_a22oi_1 _21676_ (.Y(_04400_),
    .B1(net140),
    .B2(net222),
    .A2(net170),
    .A1(net167));
 sg13g2_nand3_1 _21677_ (.B(_04399_),
    .C(_04400_),
    .A(net143),
    .Y(_04401_));
 sg13g2_nor2_1 _21678_ (.A(_09662_),
    .B(_04315_),
    .Y(_04402_));
 sg13g2_a221oi_1 _21679_ (.B2(_04402_),
    .C1(net223),
    .B1(_04401_),
    .A1(net1088),
    .Y(_04403_),
    .A2(_11472_));
 sg13g2_nor2b_1 _21680_ (.A(_04398_),
    .B_N(_04403_),
    .Y(_04404_));
 sg13g2_and2_1 _21681_ (.A(_03530_),
    .B(_03531_),
    .X(_04405_));
 sg13g2_xnor2_1 _21682_ (.Y(_04406_),
    .A(_03528_),
    .B(_04405_));
 sg13g2_nand2_1 _21683_ (.Y(_04407_),
    .A(_03995_),
    .B(_04406_));
 sg13g2_xnor2_1 _21684_ (.Y(_04408_),
    .A(net102),
    .B(_04405_));
 sg13g2_nand2b_1 _21685_ (.Y(_04409_),
    .B(net1086),
    .A_N(_04408_));
 sg13g2_nand4_1 _21686_ (.B(_04404_),
    .C(_04407_),
    .A(_04390_),
    .Y(_04410_),
    .D(_04409_));
 sg13g2_o21ai_1 _21687_ (.B1(_04410_),
    .Y(_04411_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[5] ));
 sg13g2_buf_1 _21688_ (.A(_08482_),
    .X(_04412_));
 sg13g2_nand2_1 _21689_ (.Y(_04413_),
    .A(net1038),
    .B(_04097_));
 sg13g2_xnor2_1 _21690_ (.Y(_04414_),
    .A(_10929_),
    .B(_04413_));
 sg13g2_a22oi_1 _21691_ (.Y(_04415_),
    .B1(_04414_),
    .B2(net32),
    .A2(net28),
    .A1(net948));
 sg13g2_o21ai_1 _21692_ (.B1(_04415_),
    .Y(_00991_),
    .A1(net30),
    .A2(_04411_));
 sg13g2_a21oi_1 _21693_ (.A1(_03528_),
    .A2(_03530_),
    .Y(_04416_),
    .B1(_03532_));
 sg13g2_nand2_1 _21694_ (.Y(_04417_),
    .A(net204),
    .B(net148));
 sg13g2_inv_1 _21695_ (.Y(_04418_),
    .A(_04417_));
 sg13g2_nor2_1 _21696_ (.A(_04418_),
    .B(_03507_),
    .Y(_04419_));
 sg13g2_xnor2_1 _21697_ (.Y(_04420_),
    .A(_04416_),
    .B(_04419_));
 sg13g2_nor2_1 _21698_ (.A(net191),
    .B(net236),
    .Y(_04421_));
 sg13g2_nand2_1 _21699_ (.Y(_04422_),
    .A(net191),
    .B(net236));
 sg13g2_o21ai_1 _21700_ (.B1(_04422_),
    .Y(_04423_),
    .A1(net102),
    .A2(_04421_));
 sg13g2_xnor2_1 _21701_ (.Y(_04424_),
    .A(_04419_),
    .B(_04423_));
 sg13g2_nand2_1 _21702_ (.Y(_04425_),
    .A(_03456_),
    .B(net145));
 sg13g2_a21oi_1 _21703_ (.A1(net228),
    .A2(_04066_),
    .Y(_04426_),
    .B1(_03974_));
 sg13g2_nand2_1 _21704_ (.Y(_04427_),
    .A(net172),
    .B(net170));
 sg13g2_o21ai_1 _21705_ (.B1(_04427_),
    .Y(_04428_),
    .A1(net171),
    .A2(_04207_));
 sg13g2_a221oi_1 _21706_ (.B2(net189),
    .C1(_04428_),
    .B1(_04128_),
    .A1(net239),
    .Y(_04429_),
    .A2(_04064_));
 sg13g2_a22oi_1 _21707_ (.Y(_04430_),
    .B1(net147),
    .B2(net194),
    .A2(_04076_),
    .A1(_03489_));
 sg13g2_nand4_1 _21708_ (.B(_04426_),
    .C(_04429_),
    .A(_04211_),
    .Y(_04431_),
    .D(_04430_));
 sg13g2_a21o_1 _21709_ (.A2(_04431_),
    .A1(_04293_),
    .B1(_04396_),
    .X(_04432_));
 sg13g2_a22oi_1 _21710_ (.Y(_04433_),
    .B1(net118),
    .B2(net225),
    .A2(_04076_),
    .A1(net222));
 sg13g2_a21oi_1 _21711_ (.A1(net167),
    .A2(_04081_),
    .Y(_04434_),
    .B1(_03974_));
 sg13g2_nor2_1 _21712_ (.A(_03513_),
    .B(_04069_),
    .Y(_04435_));
 sg13g2_a21oi_1 _21713_ (.A1(net188),
    .A2(_04128_),
    .Y(_04436_),
    .B1(_04435_));
 sg13g2_nand3_1 _21714_ (.B(_04434_),
    .C(_04436_),
    .A(_04433_),
    .Y(_04437_));
 sg13g2_nand3_1 _21715_ (.B(_04368_),
    .C(_04437_),
    .A(net1080),
    .Y(_04438_));
 sg13g2_nand2_1 _21716_ (.Y(_04439_),
    .A(net1079),
    .B(_03507_));
 sg13g2_o21ai_1 _21717_ (.B1(_04439_),
    .Y(_04440_),
    .A1(_08840_),
    .A2(_03507_));
 sg13g2_o21ai_1 _21718_ (.B1(_04417_),
    .Y(_04441_),
    .A1(net1012),
    .A2(_04440_));
 sg13g2_a21oi_1 _21719_ (.A1(net1088),
    .A2(_11497_),
    .Y(_04442_),
    .B1(net223));
 sg13g2_nand3_1 _21720_ (.B(_04441_),
    .C(_04442_),
    .A(_04438_),
    .Y(_04443_));
 sg13g2_a221oi_1 _21721_ (.B2(_04432_),
    .C1(_04443_),
    .B1(_04425_),
    .A1(net1086),
    .Y(_04444_),
    .A2(_04424_));
 sg13g2_o21ai_1 _21722_ (.B1(_04444_),
    .Y(_04445_),
    .A1(_03992_),
    .A2(_04420_));
 sg13g2_o21ai_1 _21723_ (.B1(_04445_),
    .Y(_04446_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[6] ));
 sg13g2_buf_1 _21724_ (.A(_08435_),
    .X(_04447_));
 sg13g2_nand3_1 _21725_ (.B(_08482_),
    .C(_04097_),
    .A(net1038),
    .Y(_04448_));
 sg13g2_xnor2_1 _21726_ (.Y(_04449_),
    .A(_10982_),
    .B(_04448_));
 sg13g2_a22oi_1 _21727_ (.Y(_04450_),
    .B1(_04449_),
    .B2(net32),
    .A2(net28),
    .A1(net947));
 sg13g2_o21ai_1 _21728_ (.B1(_04450_),
    .Y(_00992_),
    .A1(net30),
    .A2(_04446_));
 sg13g2_nand2_1 _21729_ (.Y(_04451_),
    .A(_03995_),
    .B(_04048_));
 sg13g2_a22oi_1 _21730_ (.Y(_04452_),
    .B1(_03440_),
    .B2(_03443_),
    .A2(_03435_),
    .A1(net102));
 sg13g2_xor2_1 _21731_ (.B(_04047_),
    .A(_04452_),
    .X(_04453_));
 sg13g2_nand2_1 _21732_ (.Y(_04454_),
    .A(net949),
    .B(_04453_));
 sg13g2_and4_1 _21733_ (.A(_10859_),
    .B(net332),
    .C(net235),
    .D(_03523_),
    .X(_04455_));
 sg13g2_a21o_1 _21734_ (.A2(_04128_),
    .A1(_10877_),
    .B1(_04455_),
    .X(_04456_));
 sg13g2_nor2_1 _21735_ (.A(_03493_),
    .B(_03956_),
    .Y(_04457_));
 sg13g2_and4_1 _21736_ (.A(net290),
    .B(_11272_),
    .C(_03473_),
    .D(_03954_),
    .X(_04458_));
 sg13g2_a21o_1 _21737_ (.A2(_04081_),
    .A1(_03561_),
    .B1(_04458_),
    .X(_04459_));
 sg13g2_nor4_1 _21738_ (.A(_04147_),
    .B(_04456_),
    .C(_04457_),
    .D(_04459_),
    .Y(_04460_));
 sg13g2_o21ai_1 _21739_ (.B1(_04460_),
    .Y(_04461_),
    .A1(net231),
    .A2(_04203_));
 sg13g2_a21oi_1 _21740_ (.A1(net290),
    .A2(_11175_),
    .Y(_04462_),
    .B1(net201));
 sg13g2_o21ai_1 _21741_ (.B1(_04460_),
    .Y(_04463_),
    .A1(net231),
    .A2(_04462_));
 sg13g2_a22oi_1 _21742_ (.Y(_04464_),
    .B1(_04463_),
    .B2(net1043),
    .A2(_04461_),
    .A1(net1081));
 sg13g2_a21o_1 _21743_ (.A2(net145),
    .A1(_03537_),
    .B1(_04464_),
    .X(_04465_));
 sg13g2_mux2_1 _21744_ (.A0(net1087),
    .A1(net1011),
    .S(_03568_),
    .X(_04466_));
 sg13g2_o21ai_1 _21745_ (.B1(_03552_),
    .Y(_04467_),
    .A1(net1012),
    .A2(_04466_));
 sg13g2_a22oi_1 _21746_ (.Y(_04468_),
    .B1(net142),
    .B2(net188),
    .A2(net140),
    .A1(net167));
 sg13g2_a21oi_1 _21747_ (.A1(net229),
    .A2(net141),
    .Y(_04469_),
    .B1(net145));
 sg13g2_a22oi_1 _21748_ (.Y(_04470_),
    .B1(net118),
    .B2(net191),
    .A2(net117),
    .A1(net222));
 sg13g2_nand4_1 _21749_ (.B(_04468_),
    .C(_04469_),
    .A(_03929_),
    .Y(_04471_),
    .D(_04470_));
 sg13g2_a21oi_1 _21750_ (.A1(net148),
    .A2(net145),
    .Y(_04472_),
    .B1(_09662_));
 sg13g2_a221oi_1 _21751_ (.B2(_04472_),
    .C1(net223),
    .B1(_04471_),
    .A1(net1088),
    .Y(_04473_),
    .A2(_10230_));
 sg13g2_and3_1 _21752_ (.X(_04474_),
    .A(_04465_),
    .B(_04467_),
    .C(_04473_));
 sg13g2_nand3_1 _21753_ (.B(_04454_),
    .C(_04474_),
    .A(_04451_),
    .Y(_04475_));
 sg13g2_o21ai_1 _21754_ (.B1(_04475_),
    .Y(_04476_),
    .A1(net226),
    .A2(\cpu.ex.c_mult[7] ));
 sg13g2_xnor2_1 _21755_ (.Y(_04477_),
    .A(_10945_),
    .B(_04098_));
 sg13g2_a22oi_1 _21756_ (.Y(_04478_),
    .B1(_04477_),
    .B2(net32),
    .A2(net28),
    .A1(\cpu.ex.pc[7] ));
 sg13g2_o21ai_1 _21757_ (.B1(_04478_),
    .Y(_00993_),
    .A1(net30),
    .A2(_04476_));
 sg13g2_a21oi_1 _21758_ (.A1(_09652_),
    .A2(_04048_),
    .Y(_04479_),
    .B1(net630));
 sg13g2_a22oi_1 _21759_ (.Y(_04480_),
    .B1(net142),
    .B2(_03402_),
    .A2(net170),
    .A1(net189));
 sg13g2_a22oi_1 _21760_ (.Y(_04481_),
    .B1(net141),
    .B2(net193),
    .A2(net140),
    .A1(net166));
 sg13g2_nor2b_1 _21761_ (.A(_04462_),
    .B_N(net1043),
    .Y(_04482_));
 sg13g2_o21ai_1 _21762_ (.B1(net192),
    .Y(_04483_),
    .A1(net117),
    .A2(_04482_));
 sg13g2_nand4_1 _21763_ (.B(_04480_),
    .C(_04481_),
    .A(_04126_),
    .Y(_04484_),
    .D(_04483_));
 sg13g2_a21oi_1 _21764_ (.A1(_03474_),
    .A2(net120),
    .Y(_04485_),
    .B1(_03977_));
 sg13g2_nor2_1 _21765_ (.A(_04286_),
    .B(_04360_),
    .Y(_04486_));
 sg13g2_a22oi_1 _21766_ (.Y(_04487_),
    .B1(net142),
    .B2(net167),
    .A2(net117),
    .A1(net188));
 sg13g2_a21oi_1 _21767_ (.A1(_03926_),
    .A2(_04081_),
    .Y(_04488_),
    .B1(_03974_));
 sg13g2_a22oi_1 _21768_ (.Y(_04489_),
    .B1(net147),
    .B2(net222),
    .A2(_04128_),
    .A1(net229));
 sg13g2_nand4_1 _21769_ (.B(_04487_),
    .C(_04488_),
    .A(_04486_),
    .Y(_04490_),
    .D(_04489_));
 sg13g2_nand3_1 _21770_ (.B(_04425_),
    .C(_04490_),
    .A(net1080),
    .Y(_04491_));
 sg13g2_nand2_1 _21771_ (.Y(_04492_),
    .A(net1079),
    .B(_03539_));
 sg13g2_o21ai_1 _21772_ (.B1(_04492_),
    .Y(_04493_),
    .A1(net883),
    .A2(_03539_));
 sg13g2_o21ai_1 _21773_ (.B1(_03545_),
    .Y(_04494_),
    .A1(net1012),
    .A2(_04493_));
 sg13g2_nand2_1 _21774_ (.Y(_04495_),
    .A(_04491_),
    .B(_04494_));
 sg13g2_a221oi_1 _21775_ (.B2(_04485_),
    .C1(_04495_),
    .B1(_04484_),
    .A1(net1024),
    .Y(_04496_),
    .A2(_11193_));
 sg13g2_and2_1 _21776_ (.A(_04479_),
    .B(_04496_),
    .X(_04497_));
 sg13g2_or3_1 _21777_ (.A(_04027_),
    .B(_03457_),
    .C(_04029_),
    .X(_04498_));
 sg13g2_nand2b_1 _21778_ (.Y(_04499_),
    .B(_03545_),
    .A_N(_03539_));
 sg13g2_o21ai_1 _21779_ (.B1(net1086),
    .Y(_04500_),
    .A1(_04498_),
    .A2(_04499_));
 sg13g2_a21o_1 _21780_ (.A2(_04499_),
    .A1(_04498_),
    .B1(_04500_),
    .X(_04501_));
 sg13g2_nor3_1 _21781_ (.A(_10962_),
    .B(_03507_),
    .C(_03534_),
    .Y(_04502_));
 sg13g2_o21ai_1 _21782_ (.B1(net221),
    .Y(_04503_),
    .A1(_03507_),
    .A2(_03534_));
 sg13g2_o21ai_1 _21783_ (.B1(_04503_),
    .Y(_04504_),
    .A1(_11166_),
    .A2(_04502_));
 sg13g2_buf_1 _21784_ (.A(_04504_),
    .X(_04505_));
 sg13g2_xor2_1 _21785_ (.B(_04505_),
    .A(_04499_),
    .X(_04506_));
 sg13g2_a221oi_1 _21786_ (.B2(net630),
    .C1(net187),
    .B1(_04506_),
    .A1(_04497_),
    .Y(_04507_),
    .A2(_04501_));
 sg13g2_a21oi_1 _21787_ (.A1(net187),
    .A2(\cpu.ex.c_mult[8] ),
    .Y(_04508_),
    .B1(_04507_));
 sg13g2_xnor2_1 _21788_ (.Y(_04509_),
    .A(_10681_),
    .B(_04100_));
 sg13g2_a22oi_1 _21789_ (.Y(_04510_),
    .B1(_04509_),
    .B2(_04104_),
    .A2(_04020_),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_o21ai_1 _21790_ (.B1(_04510_),
    .Y(_00994_),
    .A1(net30),
    .A2(_04508_));
 sg13g2_xor2_1 _21791_ (.B(net146),
    .A(_11373_),
    .X(_04511_));
 sg13g2_a21oi_1 _21792_ (.A1(_03545_),
    .A2(_04505_),
    .Y(_04512_),
    .B1(_03539_));
 sg13g2_xnor2_1 _21793_ (.Y(_04513_),
    .A(_04511_),
    .B(_04512_));
 sg13g2_and2_1 _21794_ (.A(_03452_),
    .B(_03460_),
    .X(_04514_));
 sg13g2_xor2_1 _21795_ (.B(_04511_),
    .A(_04514_),
    .X(_04515_));
 sg13g2_a22oi_1 _21796_ (.Y(_04516_),
    .B1(_04066_),
    .B2(_03561_),
    .A2(_04076_),
    .A1(net239));
 sg13g2_a22oi_1 _21797_ (.Y(_04517_),
    .B1(_04081_),
    .B2(net166),
    .A2(_04128_),
    .A1(_10859_));
 sg13g2_nand4_1 _21798_ (.B(_04255_),
    .C(_04516_),
    .A(net143),
    .Y(_04518_),
    .D(_04517_));
 sg13g2_a21oi_1 _21799_ (.A1(_04207_),
    .A2(_04462_),
    .Y(_04519_),
    .B1(_03398_));
 sg13g2_o21ai_1 _21800_ (.B1(net1043),
    .Y(_04520_),
    .A1(_04518_),
    .A2(_04519_));
 sg13g2_nand2_1 _21801_ (.Y(_04521_),
    .A(net1081),
    .B(_04518_));
 sg13g2_nand2_1 _21802_ (.Y(_04522_),
    .A(_04520_),
    .B(_04521_));
 sg13g2_nand2_1 _21803_ (.Y(_04523_),
    .A(_04090_),
    .B(_04522_));
 sg13g2_nand3_1 _21804_ (.B(_11373_),
    .C(net146),
    .A(net1011),
    .Y(_04524_));
 sg13g2_o21ai_1 _21805_ (.B1(net1087),
    .Y(_04525_),
    .A1(_10365_),
    .A2(_03474_));
 sg13g2_nand3_1 _21806_ (.B(_04524_),
    .C(_04525_),
    .A(_04060_),
    .Y(_04526_));
 sg13g2_a22oi_1 _21807_ (.Y(_04527_),
    .B1(_03543_),
    .B2(_04526_),
    .A2(_11173_),
    .A1(net1024));
 sg13g2_a22oi_1 _21808_ (.Y(_04528_),
    .B1(net147),
    .B2(net188),
    .A2(net142),
    .A1(net190));
 sg13g2_a221oi_1 _21809_ (.B2(net225),
    .C1(_04319_),
    .B1(net140),
    .A1(net167),
    .Y(_04529_),
    .A2(net117));
 sg13g2_a221oi_1 _21810_ (.B2(net221),
    .C1(_03949_),
    .B1(net118),
    .A1(net222),
    .Y(_04530_),
    .A2(net144));
 sg13g2_nand3_1 _21811_ (.B(_04529_),
    .C(_04530_),
    .A(_04528_),
    .Y(_04531_));
 sg13g2_a21oi_1 _21812_ (.A1(_03537_),
    .A2(net120),
    .Y(_04532_),
    .B1(_09662_));
 sg13g2_nand2_1 _21813_ (.Y(_04533_),
    .A(_04531_),
    .B(_04532_));
 sg13g2_nand4_1 _21814_ (.B(_04523_),
    .C(_04527_),
    .A(_04050_),
    .Y(_04534_),
    .D(_04533_));
 sg13g2_a221oi_1 _21815_ (.B2(net949),
    .C1(_04534_),
    .B1(_04515_),
    .A1(net630),
    .Y(_04535_),
    .A2(_04513_));
 sg13g2_a21oi_1 _21816_ (.A1(net187),
    .A2(_11390_),
    .Y(_04536_),
    .B1(_04535_));
 sg13g2_nand2_1 _21817_ (.Y(_04537_),
    .A(_04227_),
    .B(_04536_));
 sg13g2_xnor2_1 _21818_ (.Y(_04538_),
    .A(_00292_),
    .B(_04101_));
 sg13g2_a22oi_1 _21819_ (.Y(_04539_),
    .B1(_04538_),
    .B2(net32),
    .A2(net28),
    .A1(_08460_));
 sg13g2_nand2_1 _21820_ (.Y(_00995_),
    .A(_04537_),
    .B(_04539_));
 sg13g2_nand2_1 _21821_ (.Y(_04540_),
    .A(_10184_),
    .B(net119));
 sg13g2_and2_1 _21822_ (.A(_04540_),
    .B(_03554_),
    .X(_04541_));
 sg13g2_and2_1 _21823_ (.A(_03543_),
    .B(_03545_),
    .X(_04542_));
 sg13g2_nor2_1 _21824_ (.A(_03562_),
    .B(_03563_),
    .Y(_04543_));
 sg13g2_a21oi_1 _21825_ (.A1(_04542_),
    .A2(_04505_),
    .Y(_04544_),
    .B1(_04543_));
 sg13g2_xnor2_1 _21826_ (.Y(_04545_),
    .A(_04541_),
    .B(_04544_));
 sg13g2_xnor2_1 _21827_ (.Y(_04546_),
    .A(_04037_),
    .B(_04541_));
 sg13g2_nand3_1 _21828_ (.B(net208),
    .C(net119),
    .A(net1011),
    .Y(_04547_));
 sg13g2_nand2_1 _21829_ (.Y(_04548_),
    .A(net1087),
    .B(_04540_));
 sg13g2_nand3_1 _21830_ (.B(_04547_),
    .C(_04548_),
    .A(_04060_),
    .Y(_04549_));
 sg13g2_a21oi_1 _21831_ (.A1(net190),
    .A2(_04087_),
    .Y(_04550_),
    .B1(_04288_));
 sg13g2_nor2_1 _21832_ (.A(_03432_),
    .B(_03946_),
    .Y(_04551_));
 sg13g2_a21oi_1 _21833_ (.A1(net221),
    .A2(net170),
    .Y(_04552_),
    .B1(_04551_));
 sg13g2_a22oi_1 _21834_ (.Y(_04553_),
    .B1(_03967_),
    .B2(_03425_),
    .A2(_04076_),
    .A1(net225));
 sg13g2_a22oi_1 _21835_ (.Y(_04554_),
    .B1(_03964_),
    .B2(net222),
    .A2(net144),
    .A1(_03420_));
 sg13g2_and4_1 _21836_ (.A(_04426_),
    .B(_04552_),
    .C(_04553_),
    .D(_04554_),
    .X(_04555_));
 sg13g2_a221oi_1 _21837_ (.B2(_04555_),
    .C1(_09662_),
    .B1(_04550_),
    .A1(_03474_),
    .Y(_04556_),
    .A2(net145));
 sg13g2_a221oi_1 _21838_ (.B2(_04549_),
    .C1(_04556_),
    .B1(_03554_),
    .A1(net1024),
    .Y(_04557_),
    .A2(_11258_));
 sg13g2_nor2_1 _21839_ (.A(net362),
    .B(_11258_),
    .Y(_04558_));
 sg13g2_nor2_1 _21840_ (.A(net334),
    .B(net290),
    .Y(_04559_));
 sg13g2_a221oi_1 _21841_ (.B2(net283),
    .C1(_04559_),
    .B1(_04558_),
    .A1(_11111_),
    .Y(_04560_),
    .A2(_11115_));
 sg13g2_a22oi_1 _21842_ (.Y(_04561_),
    .B1(_04082_),
    .B2(_03400_),
    .A2(_04204_),
    .A1(net239));
 sg13g2_a21oi_1 _21843_ (.A1(net166),
    .A2(net170),
    .Y(_04562_),
    .B1(_03974_));
 sg13g2_nand3_1 _21844_ (.B(_04561_),
    .C(_04562_),
    .A(_04210_),
    .Y(_04563_));
 sg13g2_nand2_1 _21845_ (.Y(_04564_),
    .A(_04293_),
    .B(_04563_));
 sg13g2_o21ai_1 _21846_ (.B1(_04564_),
    .Y(_04565_),
    .A1(_04196_),
    .A2(_04560_));
 sg13g2_nand2_1 _21847_ (.Y(_04566_),
    .A(_04132_),
    .B(_04565_));
 sg13g2_nand3_1 _21848_ (.B(_04557_),
    .C(_04566_),
    .A(_04050_),
    .Y(_04567_));
 sg13g2_a221oi_1 _21849_ (.B2(net949),
    .C1(_04567_),
    .B1(_04546_),
    .A1(net630),
    .Y(_04568_),
    .A2(_04545_));
 sg13g2_a21o_1 _21850_ (.A2(_11423_),
    .A1(_04141_),
    .B1(_04568_),
    .X(_04569_));
 sg13g2_buf_1 _21851_ (.A(_08490_),
    .X(_04570_));
 sg13g2_nand2_1 _21852_ (.Y(_04571_),
    .A(_08460_),
    .B(_04101_));
 sg13g2_xnor2_1 _21853_ (.Y(_04572_),
    .A(_10527_),
    .B(_04571_));
 sg13g2_a22oi_1 _21854_ (.Y(_04573_),
    .B1(_04572_),
    .B2(net35),
    .A2(_04020_),
    .A1(net946));
 sg13g2_o21ai_1 _21855_ (.B1(_04573_),
    .Y(_00996_),
    .A1(_03913_),
    .A2(_04569_));
 sg13g2_mux2_1 _21856_ (.A0(\cpu.dec.r_set_cc ),
    .A1(\cpu.ex.r_set_cc ),
    .S(_03396_),
    .X(_00999_));
 sg13g2_buf_1 _21857_ (.A(_00256_),
    .X(_04574_));
 sg13g2_nor4_1 _21858_ (.A(net1076),
    .B(_09967_),
    .C(_04574_),
    .D(_03341_),
    .Y(_04575_));
 sg13g2_buf_2 _21859_ (.A(_04575_),
    .X(_04576_));
 sg13g2_buf_1 _21860_ (.A(_04576_),
    .X(_04577_));
 sg13g2_mux2_1 _21861_ (.A0(_10810_),
    .A1(net441),
    .S(net495),
    .X(_01000_));
 sg13g2_buf_1 _21862_ (.A(net952),
    .X(_04578_));
 sg13g2_mux2_1 _21863_ (.A0(\cpu.ex.r_sp[11] ),
    .A1(_04578_),
    .S(net495),
    .X(_01001_));
 sg13g2_mux2_1 _21864_ (.A0(_10332_),
    .A1(net497),
    .S(net495),
    .X(_01002_));
 sg13g2_mux2_1 _21865_ (.A0(_10287_),
    .A1(net498),
    .S(_04577_),
    .X(_01003_));
 sg13g2_mux2_1 _21866_ (.A0(_10250_),
    .A1(net438),
    .S(net495),
    .X(_01004_));
 sg13g2_mux2_1 _21867_ (.A0(_10209_),
    .A1(_03354_),
    .S(_04577_),
    .X(_01005_));
 sg13g2_mux2_1 _21868_ (.A0(_10554_),
    .A1(net505),
    .S(net495),
    .X(_01006_));
 sg13g2_mux2_1 _21869_ (.A0(_10781_),
    .A1(net440),
    .S(net495),
    .X(_01007_));
 sg13g2_mux2_1 _21870_ (.A0(_10474_),
    .A1(net504),
    .S(net495),
    .X(_01008_));
 sg13g2_mux2_1 _21871_ (.A0(_10436_),
    .A1(net501),
    .S(net495),
    .X(_01009_));
 sg13g2_mux2_1 _21872_ (.A0(_10421_),
    .A1(net827),
    .S(_04576_),
    .X(_01010_));
 sg13g2_buf_1 _21873_ (.A(net956),
    .X(_04579_));
 sg13g2_mux2_1 _21874_ (.A0(_10390_),
    .A1(_04579_),
    .S(_04576_),
    .X(_01011_));
 sg13g2_buf_1 _21875_ (.A(_02869_),
    .X(_04580_));
 sg13g2_mux2_1 _21876_ (.A0(_10096_),
    .A1(_04580_),
    .S(_04576_),
    .X(_01012_));
 sg13g2_mux2_1 _21877_ (.A0(_10030_),
    .A1(net828),
    .S(_04576_),
    .X(_01013_));
 sg13g2_mux2_1 _21878_ (.A0(_10161_),
    .A1(net830),
    .S(_04576_),
    .X(_01014_));
 sg13g2_or2_1 _21879_ (.X(_04581_),
    .B(_03341_),
    .A(_09970_));
 sg13g2_buf_1 _21880_ (.A(_04581_),
    .X(_04582_));
 sg13g2_buf_1 _21881_ (.A(_04582_),
    .X(_04583_));
 sg13g2_nor2b_1 _21882_ (.A(_04574_),
    .B_N(net896),
    .Y(_04584_));
 sg13g2_nand2_1 _21883_ (.Y(_04585_),
    .A(_03339_),
    .B(_04584_));
 sg13g2_and2_1 _21884_ (.A(net896),
    .B(_09967_),
    .X(_04586_));
 sg13g2_a21oi_1 _21885_ (.A1(_09968_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04587_),
    .B1(_04586_));
 sg13g2_or4_1 _21886_ (.A(net1076),
    .B(_04574_),
    .C(_03341_),
    .D(_04587_),
    .X(_04588_));
 sg13g2_buf_1 _21887_ (.A(_04588_),
    .X(_04589_));
 sg13g2_buf_1 _21888_ (.A(_04589_),
    .X(_04590_));
 sg13g2_nand2_1 _21889_ (.Y(_04591_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net434));
 sg13g2_o21ai_1 _21890_ (.B1(_04591_),
    .Y(_01015_),
    .A1(net494),
    .A2(_04585_));
 sg13g2_mux2_1 _21891_ (.A0(net1075),
    .A1(_10161_),
    .S(net494),
    .X(_04592_));
 sg13g2_buf_1 _21892_ (.A(_04589_),
    .X(_04593_));
 sg13g2_mux2_1 _21893_ (.A0(_04592_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net433),
    .X(_01016_));
 sg13g2_mux2_1 _21894_ (.A0(_10147_),
    .A1(\cpu.ex.r_sp[11] ),
    .S(_04583_),
    .X(_04594_));
 sg13g2_mux2_1 _21895_ (.A0(_04594_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net433),
    .X(_01017_));
 sg13g2_buf_1 _21896_ (.A(_04582_),
    .X(_04595_));
 sg13g2_mux2_1 _21897_ (.A0(net576),
    .A1(_10332_),
    .S(net493),
    .X(_04596_));
 sg13g2_mux2_1 _21898_ (.A0(_04596_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net434),
    .X(_01018_));
 sg13g2_mux2_1 _21899_ (.A0(net577),
    .A1(_10287_),
    .S(_04595_),
    .X(_04597_));
 sg13g2_mux2_1 _21900_ (.A0(_04597_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(_04590_),
    .X(_01019_));
 sg13g2_mux2_1 _21901_ (.A0(net578),
    .A1(_10250_),
    .S(net493),
    .X(_04598_));
 sg13g2_mux2_1 _21902_ (.A0(_04598_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net434),
    .X(_01020_));
 sg13g2_nor2_1 _21903_ (.A(net679),
    .B(net493),
    .Y(_04599_));
 sg13g2_a21oi_1 _21904_ (.A1(_10209_),
    .A2(net494),
    .Y(_04600_),
    .B1(_04599_));
 sg13g2_nand2_1 _21905_ (.Y(_04601_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(_04590_));
 sg13g2_o21ai_1 _21906_ (.B1(_04601_),
    .Y(_01021_),
    .A1(_04593_),
    .A2(_04600_));
 sg13g2_nor2_1 _21907_ (.A(net464),
    .B(net493),
    .Y(_04602_));
 sg13g2_a21oi_1 _21908_ (.A1(_10810_),
    .A2(net494),
    .Y(_04603_),
    .B1(_04602_));
 sg13g2_nand2_1 _21909_ (.Y(_04604_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net434));
 sg13g2_o21ai_1 _21910_ (.B1(_04604_),
    .Y(_01022_),
    .A1(net433),
    .A2(_04603_));
 sg13g2_nor2_1 _21911_ (.A(_03609_),
    .B(net493),
    .Y(_04605_));
 sg13g2_a21oi_1 _21912_ (.A1(_10554_),
    .A2(net494),
    .Y(_04606_),
    .B1(_04605_));
 sg13g2_nand2_1 _21913_ (.Y(_04607_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net434));
 sg13g2_o21ai_1 _21914_ (.B1(_04607_),
    .Y(_01023_),
    .A1(_04593_),
    .A2(_04606_));
 sg13g2_nor2_1 _21915_ (.A(_09041_),
    .B(_04595_),
    .Y(_04608_));
 sg13g2_a21oi_1 _21916_ (.A1(_10781_),
    .A2(_04583_),
    .Y(_04609_),
    .B1(_04608_));
 sg13g2_nand2_1 _21917_ (.Y(_04610_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(net434));
 sg13g2_o21ai_1 _21918_ (.B1(_04610_),
    .Y(_01024_),
    .A1(net433),
    .A2(_04609_));
 sg13g2_nor2_1 _21919_ (.A(net708),
    .B(net493),
    .Y(_04611_));
 sg13g2_a21oi_1 _21920_ (.A1(_10474_),
    .A2(net494),
    .Y(_04612_),
    .B1(_04611_));
 sg13g2_nand2_1 _21921_ (.Y(_04613_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04589_));
 sg13g2_o21ai_1 _21922_ (.B1(_04613_),
    .Y(_01025_),
    .A1(net433),
    .A2(_04612_));
 sg13g2_nor2_1 _21923_ (.A(_02855_),
    .B(_04582_),
    .Y(_04614_));
 sg13g2_a21oi_1 _21924_ (.A1(_10436_),
    .A2(net494),
    .Y(_04615_),
    .B1(_04614_));
 sg13g2_nand2_1 _21925_ (.Y(_04616_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04589_));
 sg13g2_o21ai_1 _21926_ (.B1(_04616_),
    .Y(_01026_),
    .A1(net433),
    .A2(_04615_));
 sg13g2_nor2_1 _21927_ (.A(net715),
    .B(_04582_),
    .Y(_04617_));
 sg13g2_a21oi_1 _21928_ (.A1(_10421_),
    .A2(net494),
    .Y(_04618_),
    .B1(_04617_));
 sg13g2_nand2_1 _21929_ (.Y(_04619_),
    .A(\cpu.ex.r_stmp[6] ),
    .B(_04589_));
 sg13g2_o21ai_1 _21930_ (.B1(_04619_),
    .Y(_01027_),
    .A1(net433),
    .A2(_04618_));
 sg13g2_mux2_1 _21931_ (.A0(net956),
    .A1(_10390_),
    .S(net493),
    .X(_04620_));
 sg13g2_mux2_1 _21932_ (.A0(_04620_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net434),
    .X(_01028_));
 sg13g2_mux2_1 _21933_ (.A0(net1085),
    .A1(_10096_),
    .S(net493),
    .X(_04621_));
 sg13g2_mux2_1 _21934_ (.A0(_04621_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net434),
    .X(_01029_));
 sg13g2_mux2_1 _21935_ (.A0(_09985_),
    .A1(_10030_),
    .S(_04582_),
    .X(_04622_));
 sg13g2_nor2_1 _21936_ (.A(_04589_),
    .B(_04622_),
    .Y(_04623_));
 sg13g2_a21oi_1 _21937_ (.A1(_10048_),
    .A2(net433),
    .Y(_01030_),
    .B1(_04623_));
 sg13g2_buf_1 _21938_ (.A(_11226_),
    .X(_04624_));
 sg13g2_buf_1 _21939_ (.A(net101),
    .X(_04625_));
 sg13g2_buf_1 _21940_ (.A(_03394_),
    .X(_04626_));
 sg13g2_buf_1 _21941_ (.A(net986),
    .X(_04627_));
 sg13g2_buf_1 _21942_ (.A(_11668_),
    .X(_04628_));
 sg13g2_inv_1 _21943_ (.Y(_04629_),
    .A(_00311_));
 sg13g2_a22oi_1 _21944_ (.Y(_04630_),
    .B1(net513),
    .B2(\cpu.dcache.r_data[7][24] ),
    .A2(net536),
    .A1(_04629_));
 sg13g2_a22oi_1 _21945_ (.Y(_04631_),
    .B1(_11884_),
    .B2(\cpu.dcache.r_data[1][24] ),
    .A2(net456),
    .A1(\cpu.dcache.r_data[3][24] ));
 sg13g2_a22oi_1 _21946_ (.Y(_04632_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][24] ),
    .A2(net515),
    .A1(\cpu.dcache.r_data[5][24] ));
 sg13g2_a22oi_1 _21947_ (.Y(_04633_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_and4_1 _21948_ (.A(_04630_),
    .B(_04631_),
    .C(_04632_),
    .D(_04633_),
    .X(_04634_));
 sg13g2_buf_1 _21949_ (.A(_04634_),
    .X(_04635_));
 sg13g2_nand2_1 _21950_ (.Y(_04636_),
    .A(\cpu.dcache.r_data[3][16] ),
    .B(net393));
 sg13g2_buf_1 _21951_ (.A(net536),
    .X(_04637_));
 sg13g2_buf_1 _21952_ (.A(net432),
    .X(_04638_));
 sg13g2_a22oi_1 _21953_ (.Y(_04639_),
    .B1(net452),
    .B2(\cpu.dcache.r_data[7][16] ),
    .A2(net384),
    .A1(\cpu.dcache.r_data[0][16] ));
 sg13g2_a22oi_1 _21954_ (.Y(_04640_),
    .B1(net354),
    .B2(\cpu.dcache.r_data[1][16] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][16] ));
 sg13g2_mux2_1 _21955_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(\cpu.dcache.r_data[6][16] ),
    .S(net594),
    .X(_04641_));
 sg13g2_a22oi_1 _21956_ (.Y(_04642_),
    .B1(_04641_),
    .B2(net632),
    .A2(_09151_),
    .A1(\cpu.dcache.r_data[5][16] ));
 sg13g2_nand2b_1 _21957_ (.Y(_04643_),
    .B(_11604_),
    .A_N(_04642_));
 sg13g2_nand4_1 _21958_ (.B(_04639_),
    .C(_04640_),
    .A(_04636_),
    .Y(_04644_),
    .D(_04643_));
 sg13g2_nand2_1 _21959_ (.Y(_04645_),
    .A(net665),
    .B(_04644_));
 sg13g2_or3_1 _21960_ (.A(_10512_),
    .B(_08534_),
    .C(_08593_),
    .X(_04646_));
 sg13g2_buf_2 _21961_ (.A(_04646_),
    .X(_04647_));
 sg13g2_buf_1 _21962_ (.A(_04647_),
    .X(_04648_));
 sg13g2_mux2_1 _21963_ (.A0(_04635_),
    .A1(_04645_),
    .S(net629),
    .X(_04649_));
 sg13g2_a22oi_1 _21964_ (.Y(_04650_),
    .B1(net456),
    .B2(\cpu.dcache.r_data[3][0] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][0] ));
 sg13g2_a22oi_1 _21965_ (.Y(_04651_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][0] ),
    .A2(net458),
    .A1(\cpu.dcache.r_data[1][0] ));
 sg13g2_mux2_1 _21966_ (.A0(\cpu.dcache.r_data[5][0] ),
    .A1(\cpu.dcache.r_data[7][0] ),
    .S(net594),
    .X(_04652_));
 sg13g2_a22oi_1 _21967_ (.Y(_04653_),
    .B1(_04652_),
    .B2(net692),
    .A2(_09260_),
    .A1(\cpu.dcache.r_data[4][0] ));
 sg13g2_nand2b_1 _21968_ (.Y(_04654_),
    .B(net726),
    .A_N(_04653_));
 sg13g2_nand3_1 _21969_ (.B(_04651_),
    .C(_04654_),
    .A(_04650_),
    .Y(_04655_));
 sg13g2_mux2_1 _21970_ (.A0(\cpu.dcache.r_data[0][0] ),
    .A1(_04655_),
    .S(net532),
    .X(_04656_));
 sg13g2_and2_1 _21971_ (.A(net945),
    .B(_04647_),
    .X(_04657_));
 sg13g2_a22oi_1 _21972_ (.Y(_04658_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][8] ),
    .A2(net456),
    .A1(\cpu.dcache.r_data[3][8] ));
 sg13g2_a22oi_1 _21973_ (.Y(_04659_),
    .B1(net458),
    .B2(\cpu.dcache.r_data[1][8] ),
    .A2(net515),
    .A1(\cpu.dcache.r_data[5][8] ));
 sg13g2_inv_1 _21974_ (.Y(_04660_),
    .A(_00312_));
 sg13g2_a22oi_1 _21975_ (.Y(_04661_),
    .B1(net513),
    .B2(\cpu.dcache.r_data[7][8] ),
    .A2(net536),
    .A1(_04660_));
 sg13g2_a22oi_1 _21976_ (.Y(_04662_),
    .B1(net589),
    .B2(\cpu.dcache.r_data[4][8] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_nand4_1 _21977_ (.B(_04659_),
    .C(_04661_),
    .A(_04658_),
    .Y(_04663_),
    .D(_04662_));
 sg13g2_buf_1 _21978_ (.A(_04663_),
    .X(_04664_));
 sg13g2_nor2_1 _21979_ (.A(net582),
    .B(net629),
    .Y(_04665_));
 sg13g2_a22oi_1 _21980_ (.Y(_04666_),
    .B1(_04664_),
    .B2(_04665_),
    .A2(_04657_),
    .A1(_04656_));
 sg13g2_o21ai_1 _21981_ (.B1(_04666_),
    .Y(_04667_),
    .A1(net945),
    .A2(_04649_));
 sg13g2_nor4_2 _21982_ (.A(net1090),
    .B(_08589_),
    .C(_10512_),
    .Y(_04668_),
    .D(_08534_));
 sg13g2_buf_1 _21983_ (.A(_04668_),
    .X(_04669_));
 sg13g2_buf_1 _21984_ (.A(net707),
    .X(_04670_));
 sg13g2_nand2_1 _21985_ (.Y(_04671_),
    .A(net581),
    .B(_04656_));
 sg13g2_nand3_1 _21986_ (.B(net628),
    .C(_04671_),
    .A(_04645_),
    .Y(_04672_));
 sg13g2_o21ai_1 _21987_ (.B1(_04672_),
    .Y(_04673_),
    .A1(_04667_),
    .A2(net628));
 sg13g2_nand2b_1 _21988_ (.Y(_04674_),
    .B(_08950_),
    .A_N(_08954_));
 sg13g2_buf_1 _21989_ (.A(_04674_),
    .X(_04675_));
 sg13g2_buf_1 _21990_ (.A(_09476_),
    .X(_04676_));
 sg13g2_o21ai_1 _21991_ (.B1(_04676_),
    .Y(_04677_),
    .A1(net1020),
    .A2(net875));
 sg13g2_nor2_1 _21992_ (.A(_09732_),
    .B(net693),
    .Y(_04678_));
 sg13g2_nor2_1 _21993_ (.A(_02855_),
    .B(net760),
    .Y(_04679_));
 sg13g2_a21oi_1 _21994_ (.A1(_04677_),
    .A2(_04678_),
    .Y(_04680_),
    .B1(_04679_));
 sg13g2_inv_2 _21995_ (.Y(_04681_),
    .A(_09476_));
 sg13g2_nand2_1 _21996_ (.Y(_04682_),
    .A(net875),
    .B(_04681_));
 sg13g2_o21ai_1 _21997_ (.B1(_04682_),
    .Y(_04683_),
    .A1(_09040_),
    .A2(_04681_));
 sg13g2_nand2_1 _21998_ (.Y(_04684_),
    .A(net762),
    .B(net873));
 sg13g2_buf_1 _21999_ (.A(_04684_),
    .X(_04685_));
 sg13g2_nand2_1 _22000_ (.Y(_04686_),
    .A(net851),
    .B(_04676_));
 sg13g2_o21ai_1 _22001_ (.B1(_04682_),
    .Y(_04687_),
    .A1(_04685_),
    .A2(_04686_));
 sg13g2_a22oi_1 _22002_ (.Y(_04688_),
    .B1(_04681_),
    .B2(_04678_),
    .A2(net693),
    .A1(net875));
 sg13g2_nor2_1 _22003_ (.A(net873),
    .B(_04688_),
    .Y(_04689_));
 sg13g2_a221oi_1 _22004_ (.B2(net1010),
    .C1(_04689_),
    .B1(_04687_),
    .A1(net692),
    .Y(_04690_),
    .A2(_04683_));
 sg13g2_o21ai_1 _22005_ (.B1(_04690_),
    .Y(_04691_),
    .A1(_08961_),
    .A2(_04680_));
 sg13g2_buf_2 _22006_ (.A(_04691_),
    .X(_04692_));
 sg13g2_nand2_1 _22007_ (.Y(_04693_),
    .A(net632),
    .B(net873));
 sg13g2_nor2_1 _22008_ (.A(net875),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_buf_1 _22009_ (.A(_04694_),
    .X(_04695_));
 sg13g2_nand2_1 _22010_ (.Y(_04696_),
    .A(net693),
    .B(_04695_));
 sg13g2_buf_2 _22011_ (.A(_04696_),
    .X(_04697_));
 sg13g2_nor2_1 _22012_ (.A(net1010),
    .B(_04697_),
    .Y(_04698_));
 sg13g2_buf_1 _22013_ (.A(_04698_),
    .X(_04699_));
 sg13g2_a21o_1 _22014_ (.A2(_04692_),
    .A1(_08980_),
    .B1(net281),
    .X(_04700_));
 sg13g2_buf_1 _22015_ (.A(_09136_),
    .X(_04701_));
 sg13g2_nor3_1 _22016_ (.A(net1010),
    .B(net627),
    .C(net558),
    .Y(_04702_));
 sg13g2_buf_2 _22017_ (.A(_04702_),
    .X(_04703_));
 sg13g2_nor3_1 _22018_ (.A(net944),
    .B(net627),
    .C(net558),
    .Y(_04704_));
 sg13g2_buf_2 _22019_ (.A(_04704_),
    .X(_04705_));
 sg13g2_buf_2 _22020_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04706_));
 sg13g2_a22oi_1 _22021_ (.Y(_04707_),
    .B1(_04705_),
    .B2(_04706_),
    .A2(_04703_),
    .A1(_08980_));
 sg13g2_nor3_1 _22022_ (.A(net875),
    .B(net944),
    .C(_09164_),
    .Y(_04708_));
 sg13g2_buf_1 _22023_ (.A(_04708_),
    .X(_04709_));
 sg13g2_buf_2 _22024_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04710_));
 sg13g2_buf_2 _22025_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04711_));
 sg13g2_mux2_1 _22026_ (.A0(_04710_),
    .A1(_04711_),
    .S(_11687_),
    .X(_04712_));
 sg13g2_nand2_1 _22027_ (.Y(_04713_),
    .A(net762),
    .B(_08962_));
 sg13g2_buf_2 _22028_ (.A(_04713_),
    .X(_04714_));
 sg13g2_nor2_1 _22029_ (.A(net627),
    .B(_04714_),
    .Y(_04715_));
 sg13g2_buf_2 _22030_ (.A(_04715_),
    .X(_04716_));
 sg13g2_nand2_1 _22031_ (.Y(_04717_),
    .A(net1010),
    .B(_04716_));
 sg13g2_buf_1 _22032_ (.A(_04717_),
    .X(_04718_));
 sg13g2_inv_1 _22033_ (.Y(_04719_),
    .A(_04718_));
 sg13g2_buf_2 _22034_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04720_));
 sg13g2_a22oi_1 _22035_ (.Y(_04721_),
    .B1(_04719_),
    .B2(_04720_),
    .A2(_04712_),
    .A1(net626));
 sg13g2_buf_2 _22036_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04722_));
 sg13g2_nor3_2 _22037_ (.A(net746),
    .B(_04681_),
    .C(net748),
    .Y(_04723_));
 sg13g2_nor3_2 _22038_ (.A(net1010),
    .B(net1020),
    .C(_09433_),
    .Y(_04724_));
 sg13g2_buf_2 _22039_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04725_));
 sg13g2_a22oi_1 _22040_ (.Y(_04726_),
    .B1(_04724_),
    .B2(_04725_),
    .A2(_04723_),
    .A1(_04722_));
 sg13g2_nand3_1 _22041_ (.B(_04721_),
    .C(_04726_),
    .A(_04707_),
    .Y(_04727_));
 sg13g2_a21oi_1 _22042_ (.A1(\cpu.gpio.r_enable_in[0] ),
    .A2(_04700_),
    .Y(_04728_),
    .B1(_04727_));
 sg13g2_nor2_1 _22043_ (.A(_04675_),
    .B(_04728_),
    .Y(_04729_));
 sg13g2_mux2_1 _22044_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(net744),
    .X(_04730_));
 sg13g2_nand2_1 _22045_ (.Y(_04731_),
    .A(net744),
    .B(_09743_));
 sg13g2_o21ai_1 _22046_ (.B1(_04731_),
    .Y(_04732_),
    .A1(net642),
    .A2(_00285_));
 sg13g2_a22oi_1 _22047_ (.Y(_04733_),
    .B1(_04732_),
    .B2(net353),
    .A2(_04730_),
    .A1(net392));
 sg13g2_nor2_2 _22048_ (.A(net627),
    .B(net558),
    .Y(_04734_));
 sg13g2_buf_1 _22049_ (.A(_04734_),
    .X(_04735_));
 sg13g2_nand2_1 _22050_ (.Y(_04736_),
    .A(_09470_),
    .B(_08962_));
 sg13g2_buf_1 _22051_ (.A(_04736_),
    .X(_04737_));
 sg13g2_nor3_2 _22052_ (.A(net851),
    .B(net594),
    .C(net557),
    .Y(_04738_));
 sg13g2_buf_1 _22053_ (.A(_04738_),
    .X(_04739_));
 sg13g2_buf_1 _22054_ (.A(net430),
    .X(_04740_));
 sg13g2_buf_1 _22055_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04741_));
 sg13g2_a22oi_1 _22056_ (.Y(_04742_),
    .B1(net383),
    .B2(_04741_),
    .A2(net431),
    .A1(_09003_));
 sg13g2_nand2_1 _22057_ (.Y(_04743_),
    .A(_04733_),
    .B(_04742_));
 sg13g2_a22oi_1 _22058_ (.Y(_04744_),
    .B1(net400),
    .B2(_09876_),
    .A2(net390),
    .A1(\cpu.intr.r_timer_reload[0] ));
 sg13g2_nand3_1 _22059_ (.B(\cpu.intr.r_timer_reload[16] ),
    .C(net390),
    .A(net665),
    .Y(_04745_));
 sg13g2_o21ai_1 _22060_ (.B1(_04745_),
    .Y(_04746_),
    .A1(net582),
    .A2(_04744_));
 sg13g2_nor2_1 _22061_ (.A(_09001_),
    .B(_09002_),
    .Y(_04747_));
 sg13g2_and2_1 _22062_ (.A(net558),
    .B(_04737_),
    .X(_04748_));
 sg13g2_buf_1 _22063_ (.A(_04748_),
    .X(_04749_));
 sg13g2_nor2_1 _22064_ (.A(net594),
    .B(_04749_),
    .Y(_04750_));
 sg13g2_nor2_1 _22065_ (.A(net726),
    .B(_04750_),
    .Y(_04751_));
 sg13g2_buf_2 _22066_ (.A(_04751_),
    .X(_04752_));
 sg13g2_nor2_1 _22067_ (.A(_04701_),
    .B(net557),
    .Y(_04753_));
 sg13g2_buf_1 _22068_ (.A(_04753_),
    .X(_04754_));
 sg13g2_buf_1 _22069_ (.A(_04754_),
    .X(_04755_));
 sg13g2_a21oi_1 _22070_ (.A1(_09003_),
    .A2(_04752_),
    .Y(_04756_),
    .B1(net382));
 sg13g2_nor2_1 _22071_ (.A(_04747_),
    .B(_04756_),
    .Y(_04757_));
 sg13g2_nor3_1 _22072_ (.A(_04743_),
    .B(_04746_),
    .C(_04757_),
    .Y(_04758_));
 sg13g2_and2_1 _22073_ (.A(_08954_),
    .B(_09736_),
    .X(_04759_));
 sg13g2_buf_1 _22074_ (.A(_04759_),
    .X(_04760_));
 sg13g2_nor3_1 _22075_ (.A(net726),
    .B(net760),
    .C(_04693_),
    .Y(_04761_));
 sg13g2_buf_1 _22076_ (.A(_04761_),
    .X(_04762_));
 sg13g2_nand2_1 _22077_ (.Y(_04763_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(net429));
 sg13g2_a22oi_1 _22078_ (.Y(_04764_),
    .B1(_04716_),
    .B2(\cpu.uart.r_x_invert ),
    .A2(net431),
    .A1(_09001_));
 sg13g2_nor3_1 _22079_ (.A(_09262_),
    .B(_09040_),
    .C(_04736_),
    .Y(_04765_));
 sg13g2_buf_2 _22080_ (.A(_04765_),
    .X(_04766_));
 sg13g2_o21ai_1 _22081_ (.B1(net851),
    .Y(_04767_),
    .A1(_09151_),
    .A2(net749));
 sg13g2_buf_2 _22082_ (.A(_04767_),
    .X(_04768_));
 sg13g2_a22oi_1 _22083_ (.Y(_04769_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[0] ),
    .A2(_04766_),
    .A1(\cpu.uart.r_div_value[8] ));
 sg13g2_nand3_1 _22084_ (.B(_04764_),
    .C(_04769_),
    .A(_04763_),
    .Y(_04770_));
 sg13g2_nand2_1 _22085_ (.Y(_04771_),
    .A(net852),
    .B(\cpu.spi.r_mode[2][0] ));
 sg13g2_o21ai_1 _22086_ (.B1(_04771_),
    .Y(_04772_),
    .A1(net852),
    .A2(_00224_));
 sg13g2_nand3_1 _22087_ (.B(net944),
    .C(net533),
    .A(net1020),
    .Y(_04773_));
 sg13g2_buf_2 _22088_ (.A(_04773_),
    .X(_04774_));
 sg13g2_nor2_1 _22089_ (.A(_00313_),
    .B(_04774_),
    .Y(_04775_));
 sg13g2_a221oi_1 _22090_ (.B2(_04772_),
    .C1(_04775_),
    .B1(net429),
    .A1(\cpu.spi.r_mode[1][0] ),
    .Y(_04776_),
    .A2(_04724_));
 sg13g2_nand2_1 _22091_ (.Y(_04777_),
    .A(net693),
    .B(_04682_));
 sg13g2_buf_1 _22092_ (.A(_00228_),
    .X(_04778_));
 sg13g2_or2_1 _22093_ (.X(_04779_),
    .B(_04778_),
    .A(net693));
 sg13g2_o21ai_1 _22094_ (.B1(_04779_),
    .Y(_04780_),
    .A1(_08961_),
    .A2(_04686_));
 sg13g2_a21oi_1 _22095_ (.A1(_09164_),
    .A2(_09167_),
    .Y(_04781_),
    .B1(_08963_));
 sg13g2_a221oi_1 _22096_ (.B2(_08963_),
    .C1(_04781_),
    .B1(_04780_),
    .A1(net632),
    .Y(_04782_),
    .A2(_04777_));
 sg13g2_nor2_2 _22097_ (.A(net875),
    .B(_04736_),
    .Y(_04783_));
 sg13g2_nand2_1 _22098_ (.Y(_04784_),
    .A(net693),
    .B(_04783_));
 sg13g2_buf_1 _22099_ (.A(_04784_),
    .X(_04785_));
 sg13g2_nor2_2 _22100_ (.A(net1010),
    .B(net428),
    .Y(_04786_));
 sg13g2_nor3_1 _22101_ (.A(_04724_),
    .B(_04782_),
    .C(_04786_),
    .Y(_04787_));
 sg13g2_buf_2 _22102_ (.A(_04787_),
    .X(_04788_));
 sg13g2_a22oi_1 _22103_ (.Y(_04789_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net538),
    .A2(_04778_),
    .A1(_08998_));
 sg13g2_nand3_1 _22104_ (.B(net760),
    .C(\cpu.spi.r_ready ),
    .A(net746),
    .Y(_04790_));
 sg13g2_o21ai_1 _22105_ (.B1(_04790_),
    .Y(_04791_),
    .A1(net666),
    .A2(_04789_));
 sg13g2_nand2_1 _22106_ (.Y(_04792_),
    .A(_02855_),
    .B(_04766_));
 sg13g2_buf_1 _22107_ (.A(_04792_),
    .X(_04793_));
 sg13g2_buf_1 _22108_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04794_));
 sg13g2_nor2_1 _22109_ (.A(net944),
    .B(_04785_),
    .Y(_04795_));
 sg13g2_buf_2 _22110_ (.A(_04795_),
    .X(_04796_));
 sg13g2_nand2_1 _22111_ (.Y(_04797_),
    .A(_04794_),
    .B(_04796_));
 sg13g2_o21ai_1 _22112_ (.B1(_04797_),
    .Y(_04798_),
    .A1(_00314_),
    .A2(net381));
 sg13g2_a221oi_1 _22113_ (.B2(net565),
    .C1(_04798_),
    .B1(_04791_),
    .A1(_09072_),
    .Y(_04799_),
    .A2(_04788_));
 sg13g2_a21oi_1 _22114_ (.A1(_04776_),
    .A2(_04799_),
    .Y(_04800_),
    .B1(_08956_));
 sg13g2_a21oi_1 _22115_ (.A1(_04760_),
    .A2(_04770_),
    .Y(_04801_),
    .B1(_04800_));
 sg13g2_o21ai_1 _22116_ (.B1(_04801_),
    .Y(_04802_),
    .A1(net583),
    .A2(_04758_));
 sg13g2_o21ai_1 _22117_ (.B1(net823),
    .Y(_04803_),
    .A1(_04729_),
    .A2(_04802_));
 sg13g2_o21ai_1 _22118_ (.B1(_04803_),
    .Y(_04804_),
    .A1(_04627_),
    .A2(_04673_));
 sg13g2_buf_1 _22119_ (.A(_03394_),
    .X(_04805_));
 sg13g2_nor2b_1 _22120_ (.A(net74),
    .B_N(net831),
    .Y(_04806_));
 sg13g2_a21oi_1 _22121_ (.A1(net75),
    .A2(_04804_),
    .Y(_04807_),
    .B1(_04806_));
 sg13g2_nand2_1 _22122_ (.Y(_04808_),
    .A(_11216_),
    .B(_03911_));
 sg13g2_a221oi_1 _22123_ (.B2(_11203_),
    .C1(net226),
    .B1(net291),
    .A1(net463),
    .Y(_04809_),
    .A2(_11195_));
 sg13g2_a22oi_1 _22124_ (.Y(_04810_),
    .B1(_04558_),
    .B2(_03473_),
    .A2(_04559_),
    .A1(_10903_));
 sg13g2_nor3_1 _22125_ (.A(_03617_),
    .B(_11273_),
    .C(_04810_),
    .Y(_04811_));
 sg13g2_a22oi_1 _22126_ (.Y(_04812_),
    .B1(_03954_),
    .B2(net194),
    .A2(_11175_),
    .A1(_10877_));
 sg13g2_nor2_1 _22127_ (.A(_03932_),
    .B(_04812_),
    .Y(_04813_));
 sg13g2_nand2_1 _22128_ (.Y(_04814_),
    .A(net228),
    .B(_03966_));
 sg13g2_nand3_1 _22129_ (.B(_04488_),
    .C(_04814_),
    .A(_04370_),
    .Y(_04815_));
 sg13g2_nand3_1 _22130_ (.B(_03916_),
    .C(net224),
    .A(net166),
    .Y(_04816_));
 sg13g2_nand2_1 _22131_ (.Y(_04817_),
    .A(net149),
    .B(net168));
 sg13g2_a21oi_1 _22132_ (.A1(net189),
    .A2(_03952_),
    .Y(_04818_),
    .B1(_04123_));
 sg13g2_nor3_1 _22133_ (.A(_04208_),
    .B(_04435_),
    .C(_04551_),
    .Y(_04819_));
 sg13g2_nand4_1 _22134_ (.B(_04817_),
    .C(_04818_),
    .A(_04816_),
    .Y(_04820_),
    .D(_04819_));
 sg13g2_nor4_1 _22135_ (.A(_04811_),
    .B(_04813_),
    .C(_04815_),
    .D(_04820_),
    .Y(_04821_));
 sg13g2_nor2b_1 _22136_ (.A(_04821_),
    .B_N(net1081),
    .Y(_04822_));
 sg13g2_nor2_1 _22137_ (.A(net1043),
    .B(_04822_),
    .Y(_04823_));
 sg13g2_o21ai_1 _22138_ (.B1(_04821_),
    .Y(_04824_),
    .A1(net231),
    .A2(_11183_));
 sg13g2_o21ai_1 _22139_ (.B1(_04824_),
    .Y(_04825_),
    .A1(_04085_),
    .A2(_04072_));
 sg13g2_nor3_1 _22140_ (.A(_09673_),
    .B(net293),
    .C(net283),
    .Y(_04826_));
 sg13g2_nor4_1 _22141_ (.A(net1087),
    .B(net1086),
    .C(_11193_),
    .D(_03995_),
    .Y(_04827_));
 sg13g2_o21ai_1 _22142_ (.B1(_04060_),
    .Y(_04828_),
    .A1(_04826_),
    .A2(_04827_));
 sg13g2_nor4_1 _22143_ (.A(net1087),
    .B(_08921_),
    .C(_09654_),
    .D(_03995_),
    .Y(_04829_));
 sg13g2_o21ai_1 _22144_ (.B1(net293),
    .Y(_04830_),
    .A1(net283),
    .A2(_04829_));
 sg13g2_a221oi_1 _22145_ (.B2(_04830_),
    .C1(net223),
    .B1(_04828_),
    .A1(_08763_),
    .Y(_04831_),
    .A2(_10368_));
 sg13g2_o21ai_1 _22146_ (.B1(_04831_),
    .Y(_04832_),
    .A1(_04823_),
    .A2(_04825_));
 sg13g2_nor2b_1 _22147_ (.A(_04809_),
    .B_N(_04832_),
    .Y(_04833_));
 sg13g2_nand2b_1 _22148_ (.Y(_04834_),
    .B(_04833_),
    .A_N(_04808_));
 sg13g2_a21oi_1 _22149_ (.A1(net710),
    .A2(_04808_),
    .Y(_04835_),
    .B1(net101));
 sg13g2_a22oi_1 _22150_ (.Y(_01031_),
    .B1(_04834_),
    .B2(_04835_),
    .A2(_04807_),
    .A1(_04625_));
 sg13g2_buf_1 _22151_ (.A(_11226_),
    .X(_04836_));
 sg13g2_nor2_1 _22152_ (.A(net1020),
    .B(_09871_),
    .Y(_04837_));
 sg13g2_buf_1 _22153_ (.A(_04837_),
    .X(_04838_));
 sg13g2_nand2b_1 _22154_ (.Y(_04839_),
    .B(net1020),
    .A_N(_00162_));
 sg13g2_nand2_1 _22155_ (.Y(_04840_),
    .A(net873),
    .B(net10));
 sg13g2_a21oi_1 _22156_ (.A1(_04839_),
    .A2(_04840_),
    .Y(_04841_),
    .B1(net748));
 sg13g2_a221oi_1 _22157_ (.B2(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .C1(_04841_),
    .B1(_04838_),
    .A1(_08971_),
    .Y(_04842_),
    .A2(_04716_));
 sg13g2_inv_1 _22158_ (.Y(_04843_),
    .A(_04842_));
 sg13g2_a21o_1 _22159_ (.A2(_04692_),
    .A1(_08976_),
    .B1(net281),
    .X(_04844_));
 sg13g2_nor2_1 _22160_ (.A(_00159_),
    .B(net352),
    .Y(_04845_));
 sg13g2_a221oi_1 _22161_ (.B2(_08970_),
    .C1(_04845_),
    .B1(_04786_),
    .A1(_08976_),
    .Y(_04846_),
    .A2(_04703_));
 sg13g2_nand3_1 _22162_ (.B(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .C(_04738_),
    .A(net944),
    .Y(_04847_));
 sg13g2_nor2_1 _22163_ (.A(net873),
    .B(_00158_),
    .Y(_04848_));
 sg13g2_buf_1 _22164_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_04849_));
 sg13g2_nor2b_1 _22165_ (.A(net880),
    .B_N(_04849_),
    .Y(_04850_));
 sg13g2_o21ai_1 _22166_ (.B1(net626),
    .Y(_04851_),
    .A1(_04848_),
    .A2(_04850_));
 sg13g2_inv_1 _22167_ (.Y(_04852_),
    .A(_00160_));
 sg13g2_nand3_1 _22168_ (.B(_08971_),
    .C(net944),
    .A(_08970_),
    .Y(_04853_));
 sg13g2_o21ai_1 _22169_ (.B1(_04853_),
    .Y(_04854_),
    .A1(_02855_),
    .A2(_00161_));
 sg13g2_a22oi_1 _22170_ (.Y(_04855_),
    .B1(_04754_),
    .B2(_04854_),
    .A2(_04705_),
    .A1(_04852_));
 sg13g2_nand4_1 _22171_ (.B(_04847_),
    .C(_04851_),
    .A(_04846_),
    .Y(_04856_),
    .D(_04855_));
 sg13g2_a221oi_1 _22172_ (.B2(\cpu.gpio.r_enable_in[7] ),
    .C1(_04856_),
    .B1(_04844_),
    .A1(net944),
    .Y(_04857_),
    .A2(_04843_));
 sg13g2_nor2_1 _22173_ (.A(_09736_),
    .B(_04752_),
    .Y(_04858_));
 sg13g2_buf_1 _22174_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_04859_));
 sg13g2_mux2_1 _22175_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net880),
    .X(_04860_));
 sg13g2_a22oi_1 _22176_ (.Y(_04861_),
    .B1(_04860_),
    .B2(net515),
    .A2(_04738_),
    .A1(_04859_));
 sg13g2_nor2_1 _22177_ (.A(net1020),
    .B(_09731_),
    .Y(_04862_));
 sg13g2_buf_2 _22178_ (.A(_04862_),
    .X(_04863_));
 sg13g2_nand2_1 _22179_ (.Y(_04864_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_04863_));
 sg13g2_a22oi_1 _22180_ (.Y(_04865_),
    .B1(net533),
    .B2(_09766_),
    .A2(net585),
    .A1(\cpu.intr.r_timer_reload[23] ));
 sg13g2_nand2b_1 _22181_ (.Y(_04866_),
    .B(net880),
    .A_N(_04865_));
 sg13g2_nor2_1 _22182_ (.A(net1020),
    .B(_09433_),
    .Y(_04867_));
 sg13g2_buf_2 _22183_ (.A(_04867_),
    .X(_04868_));
 sg13g2_a22oi_1 _22184_ (.Y(_04869_),
    .B1(net556),
    .B2(_09911_),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[7] ));
 sg13g2_nand4_1 _22185_ (.B(_04864_),
    .C(_04866_),
    .A(_04861_),
    .Y(_04870_),
    .D(_04869_));
 sg13g2_buf_1 _22186_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_04871_));
 sg13g2_nor2_1 _22187_ (.A(net760),
    .B(_04714_),
    .Y(_04872_));
 sg13g2_buf_2 _22188_ (.A(_04872_),
    .X(_04873_));
 sg13g2_or2_1 _22189_ (.X(_04874_),
    .B(_04774_),
    .A(_00156_));
 sg13g2_o21ai_1 _22190_ (.B1(_04874_),
    .Y(_04875_),
    .A1(_00157_),
    .A2(_04792_));
 sg13g2_a221oi_1 _22191_ (.B2(\cpu.spi.r_timeout[7] ),
    .C1(_04875_),
    .B1(_04873_),
    .A1(_04871_),
    .Y(_04876_),
    .A2(_04796_));
 sg13g2_nand2b_1 _22192_ (.Y(_04877_),
    .B(_04788_),
    .A_N(_00222_));
 sg13g2_a21oi_1 _22193_ (.A1(_04876_),
    .A2(_04877_),
    .Y(_04878_),
    .B1(_08956_));
 sg13g2_a21oi_1 _22194_ (.A1(_04858_),
    .A2(_04870_),
    .Y(_04879_),
    .B1(_04878_));
 sg13g2_o21ai_1 _22195_ (.B1(_04879_),
    .Y(_04880_),
    .A1(_04675_),
    .A2(_04857_));
 sg13g2_a22oi_1 _22196_ (.Y(_04881_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04761_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_nand2_1 _22197_ (.Y(_04882_),
    .A(_04760_),
    .B(_04881_));
 sg13g2_o21ai_1 _22198_ (.B1(_04882_),
    .Y(_04883_),
    .A1(_04760_),
    .A2(_04880_));
 sg13g2_a22oi_1 _22199_ (.Y(_04884_),
    .B1(net534),
    .B2(\cpu.dcache.r_data[1][7] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][7] ));
 sg13g2_o21ai_1 _22200_ (.B1(_04884_),
    .Y(_04885_),
    .A1(_00152_),
    .A2(net532));
 sg13g2_a221oi_1 _22201_ (.B2(\cpu.dcache.r_data[7][7] ),
    .C1(_04885_),
    .B1(net585),
    .A1(\cpu.dcache.r_data[2][7] ),
    .Y(_04886_),
    .A2(net592));
 sg13g2_mux2_1 _22202_ (.A0(\cpu.dcache.r_data[4][7] ),
    .A1(\cpu.dcache.r_data[6][7] ),
    .S(net693),
    .X(_04887_));
 sg13g2_a22oi_1 _22203_ (.Y(_04888_),
    .B1(_04887_),
    .B2(net632),
    .A2(_09151_),
    .A1(\cpu.dcache.r_data[5][7] ));
 sg13g2_nand2b_1 _22204_ (.Y(_04889_),
    .B(_11603_),
    .A_N(_04888_));
 sg13g2_and2_1 _22205_ (.A(_04886_),
    .B(_04889_),
    .X(_04890_));
 sg13g2_buf_1 _22206_ (.A(_04890_),
    .X(_04891_));
 sg13g2_inv_1 _22207_ (.Y(_04892_),
    .A(_04891_));
 sg13g2_inv_1 _22208_ (.Y(_04893_),
    .A(_00153_));
 sg13g2_a22oi_1 _22209_ (.Y(_04894_),
    .B1(net585),
    .B2(\cpu.dcache.r_data[7][23] ),
    .A2(net536),
    .A1(_04893_));
 sg13g2_a22oi_1 _22210_ (.Y(_04895_),
    .B1(net534),
    .B2(\cpu.dcache.r_data[1][23] ),
    .A2(net592),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_a22oi_1 _22211_ (.Y(_04896_),
    .B1(net533),
    .B2(\cpu.dcache.r_data[6][23] ),
    .A2(net591),
    .A1(\cpu.dcache.r_data[5][23] ));
 sg13g2_a22oi_1 _22212_ (.Y(_04897_),
    .B1(net589),
    .B2(\cpu.dcache.r_data[4][23] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_nand4_1 _22213_ (.B(_04895_),
    .C(_04896_),
    .A(_04894_),
    .Y(_04898_),
    .D(_04897_));
 sg13g2_buf_1 _22214_ (.A(_04898_),
    .X(_04899_));
 sg13g2_nor2_1 _22215_ (.A(net873),
    .B(_11668_),
    .Y(_04900_));
 sg13g2_buf_2 _22216_ (.A(_04900_),
    .X(_04901_));
 sg13g2_a22oi_1 _22217_ (.Y(_04902_),
    .B1(_04899_),
    .B2(_04901_),
    .A2(_04892_),
    .A1(_11668_));
 sg13g2_inv_1 _22218_ (.Y(_04903_),
    .A(_00155_));
 sg13g2_a22oi_1 _22219_ (.Y(_04904_),
    .B1(net585),
    .B2(\cpu.dcache.r_data[7][15] ),
    .A2(net536),
    .A1(_04903_));
 sg13g2_a22oi_1 _22220_ (.Y(_04905_),
    .B1(net534),
    .B2(\cpu.dcache.r_data[1][15] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][15] ));
 sg13g2_a22oi_1 _22221_ (.Y(_04906_),
    .B1(net533),
    .B2(\cpu.dcache.r_data[6][15] ),
    .A2(net591),
    .A1(\cpu.dcache.r_data[5][15] ));
 sg13g2_a22oi_1 _22222_ (.Y(_04907_),
    .B1(net589),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(net592),
    .A1(\cpu.dcache.r_data[2][15] ));
 sg13g2_nand4_1 _22223_ (.B(_04905_),
    .C(_04906_),
    .A(_04904_),
    .Y(_04908_),
    .D(_04907_));
 sg13g2_inv_1 _22224_ (.Y(_04909_),
    .A(_00154_));
 sg13g2_a22oi_1 _22225_ (.Y(_04910_),
    .B1(net591),
    .B2(\cpu.dcache.r_data[5][31] ),
    .A2(net536),
    .A1(_04909_));
 sg13g2_a22oi_1 _22226_ (.Y(_04911_),
    .B1(net589),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(net585),
    .A1(\cpu.dcache.r_data[7][31] ));
 sg13g2_a22oi_1 _22227_ (.Y(_04912_),
    .B1(net534),
    .B2(\cpu.dcache.r_data[1][31] ),
    .A2(net592),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_a22oi_1 _22228_ (.Y(_04913_),
    .B1(net533),
    .B2(\cpu.dcache.r_data[6][31] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_nand4_1 _22229_ (.B(_04911_),
    .C(_04912_),
    .A(_04910_),
    .Y(_04914_),
    .D(_04913_));
 sg13g2_a221oi_1 _22230_ (.B2(net983),
    .C1(_04647_),
    .B1(_04914_),
    .A1(net873),
    .Y(_04915_),
    .A2(_04908_));
 sg13g2_a21oi_1 _22231_ (.A1(_04647_),
    .A2(_04902_),
    .Y(_04916_),
    .B1(_04915_));
 sg13g2_nand2_1 _22232_ (.Y(_04917_),
    .A(_08964_),
    .B(_04899_));
 sg13g2_o21ai_1 _22233_ (.B1(_04917_),
    .Y(_04918_),
    .A1(_08964_),
    .A2(_04891_));
 sg13g2_mux2_1 _22234_ (.A0(_04916_),
    .A1(_04918_),
    .S(_04668_),
    .X(_04919_));
 sg13g2_nor2_1 _22235_ (.A(net986),
    .B(_04919_),
    .Y(_04920_));
 sg13g2_a21oi_2 _22236_ (.B1(_04920_),
    .Y(_04921_),
    .A2(_04883_),
    .A1(net986));
 sg13g2_a21oi_1 _22237_ (.A1(net1090),
    .A2(_04921_),
    .Y(_04922_),
    .B1(_11222_));
 sg13g2_buf_2 _22238_ (.A(_04922_),
    .X(_04923_));
 sg13g2_buf_1 _22239_ (.A(net1090),
    .X(_04924_));
 sg13g2_and2_1 _22240_ (.A(_11665_),
    .B(_04858_),
    .X(_04925_));
 sg13g2_buf_2 _22241_ (.A(_04925_),
    .X(_04926_));
 sg13g2_buf_1 _22242_ (.A(_04838_),
    .X(_04927_));
 sg13g2_buf_1 _22243_ (.A(_04863_),
    .X(_04928_));
 sg13g2_a22oi_1 _22244_ (.Y(_04929_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[10] ),
    .A2(net492),
    .A1(_09928_));
 sg13g2_buf_2 _22245_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_04930_));
 sg13g2_mux2_1 _22246_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(\cpu.intr.r_clock_cmp[26] ),
    .S(net642),
    .X(_04931_));
 sg13g2_a22oi_1 _22247_ (.Y(_04932_),
    .B1(_04931_),
    .B2(net392),
    .A2(net383),
    .A1(_04930_));
 sg13g2_buf_1 _22248_ (.A(_04868_),
    .X(_04933_));
 sg13g2_nand2_1 _22249_ (.Y(_04934_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(net555));
 sg13g2_nand3_1 _22250_ (.B(_04932_),
    .C(_04934_),
    .A(_04929_),
    .Y(_04935_));
 sg13g2_inv_1 _22251_ (.Y(_04936_),
    .A(_00102_));
 sg13g2_buf_1 _22252_ (.A(net515),
    .X(_04937_));
 sg13g2_a22oi_1 _22253_ (.Y(_04938_),
    .B1(net426),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(_04638_),
    .A1(_04936_));
 sg13g2_a22oi_1 _22254_ (.Y(_04939_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][26] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[7][26] ));
 sg13g2_buf_1 _22255_ (.A(net456),
    .X(_04940_));
 sg13g2_a22oi_1 _22256_ (.Y(_04941_),
    .B1(net380),
    .B2(\cpu.dcache.r_data[3][26] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][26] ));
 sg13g2_a22oi_1 _22257_ (.Y(_04942_),
    .B1(net391),
    .B2(\cpu.dcache.r_data[6][26] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[1][26] ));
 sg13g2_nand4_1 _22258_ (.B(_04939_),
    .C(_04941_),
    .A(_04938_),
    .Y(_04943_),
    .D(_04942_));
 sg13g2_inv_1 _22259_ (.Y(_04944_),
    .A(_00103_));
 sg13g2_a22oi_1 _22260_ (.Y(_04945_),
    .B1(net452),
    .B2(\cpu.dcache.r_data[7][10] ),
    .A2(net432),
    .A1(_04944_));
 sg13g2_a22oi_1 _22261_ (.Y(_04946_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][10] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][10] ));
 sg13g2_a22oi_1 _22262_ (.Y(_04947_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net426),
    .A1(\cpu.dcache.r_data[5][10] ));
 sg13g2_a22oi_1 _22263_ (.Y(_04948_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_nand4_1 _22264_ (.B(_04946_),
    .C(_04947_),
    .A(_04945_),
    .Y(_04949_),
    .D(_04948_));
 sg13g2_buf_1 _22265_ (.A(_04949_),
    .X(_04950_));
 sg13g2_mux2_1 _22266_ (.A0(_04943_),
    .A1(_04950_),
    .S(net581),
    .X(_04951_));
 sg13g2_a22oi_1 _22267_ (.Y(_04952_),
    .B1(_04951_),
    .B2(_04669_),
    .A2(_04935_),
    .A1(_04926_));
 sg13g2_or2_1 _22268_ (.X(_04953_),
    .B(_04952_),
    .A(net943));
 sg13g2_nand3_1 _22269_ (.B(_04923_),
    .C(_04953_),
    .A(_04805_),
    .Y(_04954_));
 sg13g2_o21ai_1 _22270_ (.B1(_04954_),
    .Y(_04955_),
    .A1(net1075),
    .A2(net75));
 sg13g2_a21oi_1 _22271_ (.A1(_00258_),
    .A2(_11213_),
    .Y(_04956_),
    .B1(_11553_));
 sg13g2_buf_1 _22272_ (.A(_04956_),
    .X(_04957_));
 sg13g2_buf_1 _22273_ (.A(_04957_),
    .X(_04958_));
 sg13g2_a221oi_1 _22274_ (.B2(net187),
    .C1(_04568_),
    .B1(_11423_),
    .A1(_04924_),
    .Y(_04959_),
    .A2(_11214_));
 sg13g2_a21oi_1 _22275_ (.A1(_04958_),
    .A2(_04572_),
    .Y(_04960_),
    .B1(_04959_));
 sg13g2_nand2_1 _22276_ (.Y(_04961_),
    .A(_08619_),
    .B(_10654_));
 sg13g2_buf_1 _22277_ (.A(_04961_),
    .X(_04962_));
 sg13g2_nor2_1 _22278_ (.A(_11226_),
    .B(_04962_),
    .Y(_04963_));
 sg13g2_buf_1 _22279_ (.A(_03911_),
    .X(_04964_));
 sg13g2_buf_1 _22280_ (.A(net165),
    .X(_04965_));
 sg13g2_nor3_1 _22281_ (.A(net946),
    .B(net101),
    .C(net139),
    .Y(_04966_));
 sg13g2_a221oi_1 _22282_ (.B2(_04963_),
    .C1(_04966_),
    .B1(_04960_),
    .A1(net100),
    .Y(_01032_),
    .A2(_04955_));
 sg13g2_buf_1 _22283_ (.A(_11223_),
    .X(_04967_));
 sg13g2_buf_1 _22284_ (.A(_04957_),
    .X(_04968_));
 sg13g2_nand3b_1 _22285_ (.B(net165),
    .C(net624),
    .Y(_04969_),
    .A_N(_04103_));
 sg13g2_o21ai_1 _22286_ (.B1(_04969_),
    .Y(_04970_),
    .A1(\cpu.ex.pc[11] ),
    .A2(net165));
 sg13g2_nor2_1 _22287_ (.A(_11226_),
    .B(_04808_),
    .Y(_04971_));
 sg13g2_nor2_1 _22288_ (.A(net880),
    .B(net748),
    .Y(_04972_));
 sg13g2_buf_1 _22289_ (.A(_04972_),
    .X(_04973_));
 sg13g2_a22oi_1 _22290_ (.Y(_04974_),
    .B1(net554),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net555),
    .A1(_09744_));
 sg13g2_a22oi_1 _22291_ (.Y(_04975_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[11] ),
    .A2(net492),
    .A1(_09932_));
 sg13g2_nor2_1 _22292_ (.A(net746),
    .B(net748),
    .Y(_04976_));
 sg13g2_buf_1 _22293_ (.A(_04976_),
    .X(_04977_));
 sg13g2_buf_2 _22294_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_04978_));
 sg13g2_a22oi_1 _22295_ (.Y(_04979_),
    .B1(net383),
    .B2(_04978_),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_nand3_1 _22296_ (.B(_04975_),
    .C(_04979_),
    .A(_04974_),
    .Y(_04980_));
 sg13g2_inv_1 _22297_ (.Y(_04981_),
    .A(_00112_));
 sg13g2_a22oi_1 _22298_ (.Y(_04982_),
    .B1(_04937_),
    .B2(\cpu.dcache.r_data[5][27] ),
    .A2(_04638_),
    .A1(_04981_));
 sg13g2_a22oi_1 _22299_ (.Y(_04983_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][27] ),
    .A2(_02743_),
    .A1(\cpu.dcache.r_data[7][27] ));
 sg13g2_a22oi_1 _22300_ (.Y(_04984_),
    .B1(_11885_),
    .B2(\cpu.dcache.r_data[1][27] ),
    .A2(_12009_),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_a22oi_1 _22301_ (.Y(_04985_),
    .B1(net391),
    .B2(\cpu.dcache.r_data[6][27] ),
    .A2(_04940_),
    .A1(\cpu.dcache.r_data[3][27] ));
 sg13g2_nand4_1 _22302_ (.B(_04983_),
    .C(_04984_),
    .A(_04982_),
    .Y(_04986_),
    .D(_04985_));
 sg13g2_a22oi_1 _22303_ (.Y(_04987_),
    .B1(_12439_),
    .B2(\cpu.dcache.r_data[6][11] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][11] ));
 sg13g2_a22oi_1 _22304_ (.Y(_04988_),
    .B1(_02743_),
    .B2(\cpu.dcache.r_data[7][11] ),
    .A2(net515),
    .A1(\cpu.dcache.r_data[5][11] ));
 sg13g2_a22oi_1 _22305_ (.Y(_04989_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][11] ),
    .A2(_12121_),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_nand3_1 _22306_ (.B(_04988_),
    .C(_04989_),
    .A(_04987_),
    .Y(_04990_));
 sg13g2_nand2_1 _22307_ (.Y(_04991_),
    .A(_00113_),
    .B(_09454_));
 sg13g2_o21ai_1 _22308_ (.B1(_04991_),
    .Y(_04992_),
    .A1(_09454_),
    .A2(_04990_));
 sg13g2_o21ai_1 _22309_ (.B1(_11886_),
    .Y(_04993_),
    .A1(\cpu.dcache.r_data[1][11] ),
    .A2(_04990_));
 sg13g2_o21ai_1 _22310_ (.B1(_04993_),
    .Y(_04994_),
    .A1(_11886_),
    .A2(_04992_));
 sg13g2_mux2_1 _22311_ (.A0(_04986_),
    .A1(_04994_),
    .S(net529),
    .X(_04995_));
 sg13g2_a22oi_1 _22312_ (.Y(_04996_),
    .B1(_04995_),
    .B2(net628),
    .A2(_04980_),
    .A1(_04926_));
 sg13g2_o21ai_1 _22313_ (.B1(_04923_),
    .Y(_04997_),
    .A1(net943),
    .A2(_04996_));
 sg13g2_nand2b_1 _22314_ (.Y(_04998_),
    .B(net36),
    .A_N(_10147_));
 sg13g2_o21ai_1 _22315_ (.B1(_04998_),
    .Y(_04999_),
    .A1(net36),
    .A2(_04997_));
 sg13g2_a221oi_1 _22316_ (.B2(_04095_),
    .C1(_04999_),
    .B1(_04971_),
    .A1(net85),
    .Y(_01033_),
    .A2(_04970_));
 sg13g2_nand3b_1 _22317_ (.B(_04964_),
    .C(net625),
    .Y(_05000_),
    .A_N(_04139_));
 sg13g2_o21ai_1 _22318_ (.B1(_05000_),
    .Y(_05001_),
    .A1(net769),
    .A2(_04965_));
 sg13g2_buf_1 _22319_ (.A(_11223_),
    .X(_05002_));
 sg13g2_a22oi_1 _22320_ (.Y(_05003_),
    .B1(net554),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net555),
    .A1(\cpu.intr.r_timer_count[12] ));
 sg13g2_a22oi_1 _22321_ (.Y(_05004_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[12] ),
    .A2(net492),
    .A1(_09939_));
 sg13g2_buf_2 _22322_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05005_));
 sg13g2_a22oi_1 _22323_ (.Y(_05006_),
    .B1(net383),
    .B2(_05005_),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_nand3_1 _22324_ (.B(_05004_),
    .C(_05006_),
    .A(_05003_),
    .Y(_05007_));
 sg13g2_inv_1 _22325_ (.Y(_05008_),
    .A(_00123_));
 sg13g2_a22oi_1 _22326_ (.Y(_05009_),
    .B1(net515),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(net432),
    .A1(_05008_));
 sg13g2_a22oi_1 _22327_ (.Y(_05010_),
    .B1(_09858_),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(net585),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_a22oi_1 _22328_ (.Y(_05011_),
    .B1(net456),
    .B2(\cpu.dcache.r_data[3][28] ),
    .A2(_12008_),
    .A1(\cpu.dcache.r_data[2][28] ));
 sg13g2_a22oi_1 _22329_ (.Y(_05012_),
    .B1(_12439_),
    .B2(\cpu.dcache.r_data[6][28] ),
    .A2(net458),
    .A1(\cpu.dcache.r_data[1][28] ));
 sg13g2_nand4_1 _22330_ (.B(_05010_),
    .C(_05011_),
    .A(_05009_),
    .Y(_05013_),
    .D(_05012_));
 sg13g2_a22oi_1 _22331_ (.Y(_05014_),
    .B1(net534),
    .B2(\cpu.dcache.r_data[1][12] ),
    .A2(_12008_),
    .A1(\cpu.dcache.r_data[2][12] ));
 sg13g2_a22oi_1 _22332_ (.Y(_05015_),
    .B1(_09208_),
    .B2(\cpu.dcache.r_data[6][12] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][12] ));
 sg13g2_mux2_1 _22333_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(\cpu.dcache.r_data[7][12] ),
    .S(_08946_),
    .X(_05016_));
 sg13g2_a22oi_1 _22334_ (.Y(_05017_),
    .B1(_05016_),
    .B2(net692),
    .A2(_09260_),
    .A1(\cpu.dcache.r_data[4][12] ));
 sg13g2_nand2b_1 _22335_ (.Y(_05018_),
    .B(_11603_),
    .A_N(_05017_));
 sg13g2_and4_1 _22336_ (.A(net532),
    .B(_05014_),
    .C(_05015_),
    .D(_05018_),
    .X(_05019_));
 sg13g2_a21oi_1 _22337_ (.A1(_00124_),
    .A2(net432),
    .Y(_05020_),
    .B1(_05019_));
 sg13g2_mux2_1 _22338_ (.A0(_05013_),
    .A1(_05020_),
    .S(net581),
    .X(_05021_));
 sg13g2_a22oi_1 _22339_ (.Y(_05022_),
    .B1(_05021_),
    .B2(net628),
    .A2(_05007_),
    .A1(_04926_));
 sg13g2_o21ai_1 _22340_ (.B1(_04923_),
    .Y(_05023_),
    .A1(net943),
    .A2(_05022_));
 sg13g2_nand2b_1 _22341_ (.Y(_05024_),
    .B(net36),
    .A_N(net576));
 sg13g2_o21ai_1 _22342_ (.B1(_05024_),
    .Y(_05025_),
    .A1(net36),
    .A2(_05023_));
 sg13g2_a221oi_1 _22343_ (.B2(net84),
    .C1(_05025_),
    .B1(_05001_),
    .A1(_04137_),
    .Y(_01034_),
    .A2(_04971_));
 sg13g2_nand3b_1 _22344_ (.B(net165),
    .C(net625),
    .Y(_05026_),
    .A_N(_04188_));
 sg13g2_o21ai_1 _22345_ (.B1(_05026_),
    .Y(_05027_),
    .A1(net768),
    .A2(_04964_));
 sg13g2_a22oi_1 _22346_ (.Y(_05028_),
    .B1(net554),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net427),
    .A1(\cpu.intr.r_timer_reload[13] ));
 sg13g2_a22oi_1 _22347_ (.Y(_05029_),
    .B1(net492),
    .B2(_09944_),
    .A2(net555),
    .A1(\cpu.intr.r_timer_count[13] ));
 sg13g2_buf_1 _22348_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05030_));
 sg13g2_a22oi_1 _22349_ (.Y(_05031_),
    .B1(net383),
    .B2(_05030_),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_nand3_1 _22350_ (.B(_05029_),
    .C(_05031_),
    .A(_05028_),
    .Y(_05032_));
 sg13g2_inv_1 _22351_ (.Y(_05033_),
    .A(_00130_));
 sg13g2_a22oi_1 _22352_ (.Y(_05034_),
    .B1(net455),
    .B2(\cpu.dcache.r_data[5][29] ),
    .A2(net384),
    .A1(_05033_));
 sg13g2_a22oi_1 _22353_ (.Y(_05035_),
    .B1(_09860_),
    .B2(\cpu.dcache.r_data[4][29] ),
    .A2(net390),
    .A1(\cpu.dcache.r_data[7][29] ));
 sg13g2_a22oi_1 _22354_ (.Y(_05036_),
    .B1(_12122_),
    .B2(\cpu.dcache.r_data[3][29] ),
    .A2(_12010_),
    .A1(\cpu.dcache.r_data[2][29] ));
 sg13g2_a22oi_1 _22355_ (.Y(_05037_),
    .B1(_12441_),
    .B2(\cpu.dcache.r_data[6][29] ),
    .A2(net354),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_nand4_1 _22356_ (.B(_05035_),
    .C(_05036_),
    .A(_05034_),
    .Y(_05038_),
    .D(_05037_));
 sg13g2_a22oi_1 _22357_ (.Y(_05039_),
    .B1(net354),
    .B2(\cpu.dcache.r_data[1][13] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[5][13] ));
 sg13g2_a22oi_1 _22358_ (.Y(_05040_),
    .B1(_12440_),
    .B2(\cpu.dcache.r_data[6][13] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_inv_1 _22359_ (.Y(_05041_),
    .A(_00131_));
 sg13g2_a22oi_1 _22360_ (.Y(_05042_),
    .B1(_02745_),
    .B2(\cpu.dcache.r_data[7][13] ),
    .A2(net384),
    .A1(_05041_));
 sg13g2_a22oi_1 _22361_ (.Y(_05043_),
    .B1(_09859_),
    .B2(\cpu.dcache.r_data[4][13] ),
    .A2(_12010_),
    .A1(\cpu.dcache.r_data[2][13] ));
 sg13g2_nand4_1 _22362_ (.B(_05040_),
    .C(_05042_),
    .A(_05039_),
    .Y(_05044_),
    .D(_05043_));
 sg13g2_mux2_1 _22363_ (.A0(_05038_),
    .A1(_05044_),
    .S(net581),
    .X(_05045_));
 sg13g2_a22oi_1 _22364_ (.Y(_05046_),
    .B1(_05045_),
    .B2(net628),
    .A2(_05032_),
    .A1(_04926_));
 sg13g2_or2_1 _22365_ (.X(_05047_),
    .B(_05046_),
    .A(net943));
 sg13g2_a21oi_1 _22366_ (.A1(_04923_),
    .A2(_05047_),
    .Y(_05048_),
    .B1(_03395_));
 sg13g2_a21oi_1 _22367_ (.A1(_03350_),
    .A2(net36),
    .Y(_05049_),
    .B1(_05048_));
 sg13g2_a221oi_1 _22368_ (.B2(net85),
    .C1(_05049_),
    .B1(_05027_),
    .A1(_04186_),
    .Y(_01035_),
    .A2(_04971_));
 sg13g2_a22oi_1 _22369_ (.Y(_05050_),
    .B1(_04863_),
    .B2(\cpu.intr.r_timer_reload[14] ),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[14] ));
 sg13g2_buf_1 _22370_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05051_));
 sg13g2_mux2_1 _22371_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(\cpu.intr.r_clock_cmp[30] ),
    .S(net744),
    .X(_05052_));
 sg13g2_a22oi_1 _22372_ (.Y(_05053_),
    .B1(_05052_),
    .B2(net392),
    .A2(net430),
    .A1(_05051_));
 sg13g2_nand2_1 _22373_ (.Y(_05054_),
    .A(_09950_),
    .B(net556));
 sg13g2_nand3_1 _22374_ (.B(_05053_),
    .C(_05054_),
    .A(_05050_),
    .Y(_05055_));
 sg13g2_a22oi_1 _22375_ (.Y(_05056_),
    .B1(net533),
    .B2(\cpu.dcache.r_data[6][30] ),
    .A2(net592),
    .A1(\cpu.dcache.r_data[2][30] ));
 sg13g2_a22oi_1 _22376_ (.Y(_05057_),
    .B1(net585),
    .B2(\cpu.dcache.r_data[7][30] ),
    .A2(net591),
    .A1(\cpu.dcache.r_data[5][30] ));
 sg13g2_a22oi_1 _22377_ (.Y(_05058_),
    .B1(net589),
    .B2(\cpu.dcache.r_data[4][30] ),
    .A2(net535),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_nand3_1 _22378_ (.B(_05057_),
    .C(_05058_),
    .A(_05056_),
    .Y(_05059_));
 sg13g2_nand2_1 _22379_ (.Y(_05060_),
    .A(_00142_),
    .B(_09454_));
 sg13g2_o21ai_1 _22380_ (.B1(_05060_),
    .Y(_05061_),
    .A1(_09454_),
    .A2(_05059_));
 sg13g2_nor3_1 _22381_ (.A(\cpu.dcache.r_data[1][30] ),
    .B(net668),
    .C(_05059_),
    .Y(_05062_));
 sg13g2_a21o_1 _22382_ (.A2(_05061_),
    .A1(net668),
    .B1(_05062_),
    .X(_05063_));
 sg13g2_buf_1 _22383_ (.A(_05063_),
    .X(_05064_));
 sg13g2_inv_1 _22384_ (.Y(_05065_),
    .A(_00143_));
 sg13g2_a22oi_1 _22385_ (.Y(_05066_),
    .B1(net515),
    .B2(\cpu.dcache.r_data[5][14] ),
    .A2(_04637_),
    .A1(_05065_));
 sg13g2_a22oi_1 _22386_ (.Y(_05067_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[7][14] ));
 sg13g2_a22oi_1 _22387_ (.Y(_05068_),
    .B1(net456),
    .B2(\cpu.dcache.r_data[3][14] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_a22oi_1 _22388_ (.Y(_05069_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][14] ),
    .A2(net458),
    .A1(\cpu.dcache.r_data[1][14] ));
 sg13g2_nand4_1 _22389_ (.B(_05067_),
    .C(_05068_),
    .A(_05066_),
    .Y(_05070_),
    .D(_05069_));
 sg13g2_nand2_1 _22390_ (.Y(_05071_),
    .A(_09728_),
    .B(_05070_));
 sg13g2_o21ai_1 _22391_ (.B1(_05071_),
    .Y(_05072_),
    .A1(net666),
    .A2(_05064_));
 sg13g2_a22oi_1 _22392_ (.Y(_05073_),
    .B1(_05072_),
    .B2(net707),
    .A2(_05055_),
    .A1(_04926_));
 sg13g2_nand2_1 _22393_ (.Y(_05074_),
    .A(net1090),
    .B(_04921_));
 sg13g2_o21ai_1 _22394_ (.B1(_05074_),
    .Y(_05075_),
    .A1(net1090),
    .A2(_05073_));
 sg13g2_mux2_1 _22395_ (.A0(net578),
    .A1(_05075_),
    .S(_03394_),
    .X(_05076_));
 sg13g2_nand3_1 _22396_ (.B(_11222_),
    .C(_04962_),
    .A(_08344_),
    .Y(_05077_));
 sg13g2_o21ai_1 _22397_ (.B1(_05077_),
    .Y(_05078_),
    .A1(net106),
    .A2(_05076_));
 sg13g2_nor2_1 _22398_ (.A(net625),
    .B(_05078_),
    .Y(_05079_));
 sg13g2_o21ai_1 _22399_ (.B1(_05079_),
    .Y(_05080_),
    .A1(_03915_),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_nand2_1 _22400_ (.Y(_05081_),
    .A(_04958_),
    .B(_04230_));
 sg13g2_a21o_1 _22401_ (.A2(_05081_),
    .A1(_04963_),
    .B1(_05078_),
    .X(_05082_));
 sg13g2_o21ai_1 _22402_ (.B1(_05082_),
    .Y(_01036_),
    .A1(_04226_),
    .A2(_05080_));
 sg13g2_a22oi_1 _22403_ (.Y(_05083_),
    .B1(net554),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net555),
    .A1(\cpu.intr.r_timer_count[15] ));
 sg13g2_a22oi_1 _22404_ (.Y(_05084_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[15] ),
    .A2(net556),
    .A1(_09955_));
 sg13g2_buf_1 _22405_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05085_));
 sg13g2_a22oi_1 _22406_ (.Y(_05086_),
    .B1(net430),
    .B2(_05085_),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_nand3_1 _22407_ (.B(_05084_),
    .C(_05086_),
    .A(_05083_),
    .Y(_05087_));
 sg13g2_mux2_1 _22408_ (.A0(_04908_),
    .A1(_04914_),
    .S(_09867_),
    .X(_05088_));
 sg13g2_a22oi_1 _22409_ (.Y(_05089_),
    .B1(_05088_),
    .B2(net707),
    .A2(_05087_),
    .A1(_04926_));
 sg13g2_o21ai_1 _22410_ (.B1(_04923_),
    .Y(_05090_),
    .A1(net1090),
    .A2(_05089_));
 sg13g2_inv_1 _22411_ (.Y(_05091_),
    .A(_05090_));
 sg13g2_nor2_1 _22412_ (.A(net1094),
    .B(_03911_),
    .Y(_05092_));
 sg13g2_nor3_1 _22413_ (.A(_11216_),
    .B(_04962_),
    .C(_04272_),
    .Y(_05093_));
 sg13g2_nor4_1 _22414_ (.A(_03395_),
    .B(_05091_),
    .C(_05092_),
    .D(_05093_),
    .Y(_05094_));
 sg13g2_nand2_1 _22415_ (.Y(_05095_),
    .A(_04269_),
    .B(_05094_));
 sg13g2_nand2_1 _22416_ (.Y(_05096_),
    .A(net74),
    .B(_05090_));
 sg13g2_o21ai_1 _22417_ (.B1(_05096_),
    .Y(_05097_),
    .A1(net679),
    .A2(net74));
 sg13g2_buf_1 _22418_ (.A(_04962_),
    .X(_05098_));
 sg13g2_a21o_1 _22419_ (.A2(_04272_),
    .A1(net625),
    .B1(net164),
    .X(_05099_));
 sg13g2_a22oi_1 _22420_ (.Y(_05100_),
    .B1(_05094_),
    .B2(_05099_),
    .A2(_05097_),
    .A1(_04624_));
 sg13g2_o21ai_1 _22421_ (.B1(_05100_),
    .Y(_01037_),
    .A1(_04268_),
    .A2(_05095_));
 sg13g2_nand2_1 _22422_ (.Y(_05101_),
    .A(_10771_),
    .B(_04957_));
 sg13g2_o21ai_1 _22423_ (.B1(_05101_),
    .Y(_05102_),
    .A1(net624),
    .A2(_04007_));
 sg13g2_nor2_1 _22424_ (.A(net764),
    .B(net165),
    .Y(_05103_));
 sg13g2_a21oi_1 _22425_ (.A1(net139),
    .A2(_05102_),
    .Y(_05104_),
    .B1(_05103_));
 sg13g2_a22oi_1 _22426_ (.Y(_05105_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][1] ),
    .A2(net456),
    .A1(\cpu.dcache.r_data[3][1] ));
 sg13g2_a22oi_1 _22427_ (.Y(_05106_),
    .B1(net458),
    .B2(\cpu.dcache.r_data[1][1] ),
    .A2(net518),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_mux2_1 _22428_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(\cpu.dcache.r_data[7][1] ),
    .S(net594),
    .X(_05107_));
 sg13g2_a22oi_1 _22429_ (.Y(_05108_),
    .B1(_05107_),
    .B2(net692),
    .A2(net749),
    .A1(\cpu.dcache.r_data[6][1] ));
 sg13g2_nand2b_1 _22430_ (.Y(_05109_),
    .B(net726),
    .A_N(_05108_));
 sg13g2_nand3_1 _22431_ (.B(_05106_),
    .C(_05109_),
    .A(_05105_),
    .Y(_05110_));
 sg13g2_mux2_1 _22432_ (.A0(\cpu.dcache.r_data[0][1] ),
    .A1(_05110_),
    .S(net532),
    .X(_05111_));
 sg13g2_a22oi_1 _22433_ (.Y(_05112_),
    .B1(net391),
    .B2(\cpu.dcache.r_data[6][17] ),
    .A2(net458),
    .A1(\cpu.dcache.r_data[1][17] ));
 sg13g2_a22oi_1 _22434_ (.Y(_05113_),
    .B1(net513),
    .B2(\cpu.dcache.r_data[7][17] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][17] ));
 sg13g2_inv_1 _22435_ (.Y(_05114_),
    .A(_00091_));
 sg13g2_a22oi_1 _22436_ (.Y(_05115_),
    .B1(net426),
    .B2(\cpu.dcache.r_data[5][17] ),
    .A2(net432),
    .A1(_05114_));
 sg13g2_a22oi_1 _22437_ (.Y(_05116_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][17] ));
 sg13g2_nand4_1 _22438_ (.B(_05113_),
    .C(_05115_),
    .A(_05112_),
    .Y(_05117_),
    .D(_05116_));
 sg13g2_buf_1 _22439_ (.A(_05117_),
    .X(_05118_));
 sg13g2_and2_1 _22440_ (.A(net582),
    .B(_05118_),
    .X(_05119_));
 sg13g2_a21oi_1 _22441_ (.A1(net581),
    .A2(_05111_),
    .Y(_05120_),
    .B1(_05119_));
 sg13g2_a22oi_1 _22442_ (.Y(_05121_),
    .B1(_05118_),
    .B2(_04901_),
    .A2(_05111_),
    .A1(_11668_));
 sg13g2_a22oi_1 _22443_ (.Y(_05122_),
    .B1(net533),
    .B2(\cpu.dcache.r_data[6][9] ),
    .A2(_12326_),
    .A1(\cpu.dcache.r_data[5][9] ));
 sg13g2_a22oi_1 _22444_ (.Y(_05123_),
    .B1(net585),
    .B2(\cpu.dcache.r_data[7][9] ),
    .A2(net592),
    .A1(\cpu.dcache.r_data[2][9] ));
 sg13g2_nand2_1 _22445_ (.Y(_05124_),
    .A(_05122_),
    .B(_05123_));
 sg13g2_a221oi_1 _22446_ (.B2(\cpu.dcache.r_data[4][9] ),
    .C1(_05124_),
    .B1(net589),
    .A1(\cpu.dcache.r_data[3][9] ),
    .Y(_05125_),
    .A2(_12121_));
 sg13g2_mux2_1 _22447_ (.A0(_00093_),
    .A1(_05125_),
    .S(net627),
    .X(_05126_));
 sg13g2_nor2_1 _22448_ (.A(\cpu.dcache.r_data[1][9] ),
    .B(net668),
    .Y(_05127_));
 sg13g2_a22oi_1 _22449_ (.Y(_05128_),
    .B1(_05127_),
    .B2(_05125_),
    .A2(_05126_),
    .A1(net668));
 sg13g2_a22oi_1 _22450_ (.Y(_05129_),
    .B1(_12440_),
    .B2(\cpu.dcache.r_data[6][25] ),
    .A2(_04940_),
    .A1(\cpu.dcache.r_data[3][25] ));
 sg13g2_a22oi_1 _22451_ (.Y(_05130_),
    .B1(_11885_),
    .B2(\cpu.dcache.r_data[1][25] ),
    .A2(_04937_),
    .A1(\cpu.dcache.r_data[5][25] ));
 sg13g2_inv_1 _22452_ (.Y(_05131_),
    .A(_00092_));
 sg13g2_a22oi_1 _22453_ (.Y(_05132_),
    .B1(net452),
    .B2(\cpu.dcache.r_data[7][25] ),
    .A2(_04637_),
    .A1(_05131_));
 sg13g2_a22oi_1 _22454_ (.Y(_05133_),
    .B1(_09859_),
    .B2(\cpu.dcache.r_data[4][25] ),
    .A2(_12009_),
    .A1(\cpu.dcache.r_data[2][25] ));
 sg13g2_nand4_1 _22455_ (.B(_05130_),
    .C(_05132_),
    .A(_05129_),
    .Y(_05134_),
    .D(_05133_));
 sg13g2_a221oi_1 _22456_ (.B2(net983),
    .C1(_04647_),
    .B1(_05134_),
    .A1(_09729_),
    .Y(_05135_),
    .A2(_05128_));
 sg13g2_a21oi_1 _22457_ (.A1(net629),
    .A2(_05121_),
    .Y(_05136_),
    .B1(_05135_));
 sg13g2_nor2_1 _22458_ (.A(net707),
    .B(_05136_),
    .Y(_05137_));
 sg13g2_a21oi_1 _22459_ (.A1(net707),
    .A2(_05120_),
    .Y(_05138_),
    .B1(_05137_));
 sg13g2_nor2_1 _22460_ (.A(_00095_),
    .B(net428),
    .Y(_05139_));
 sg13g2_a221oi_1 _22461_ (.B2(_11595_),
    .C1(_05139_),
    .B1(_04762_),
    .A1(_11596_),
    .Y(_05140_),
    .A2(_04868_));
 sg13g2_buf_1 _22462_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05141_));
 sg13g2_nor2_1 _22463_ (.A(_02855_),
    .B(_04697_),
    .Y(_05142_));
 sg13g2_nand2_1 _22464_ (.Y(_05143_),
    .A(\cpu.spi.r_timeout[1] ),
    .B(_04873_));
 sg13g2_o21ai_1 _22465_ (.B1(_05143_),
    .Y(_05144_),
    .A1(_00094_),
    .A2(_04774_));
 sg13g2_a221oi_1 _22466_ (.B2(_11599_),
    .C1(_05144_),
    .B1(_05142_),
    .A1(_05141_),
    .Y(_05145_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22467_ (.B1(_05145_),
    .Y(_05146_),
    .A1(net852),
    .A2(_05140_));
 sg13g2_mux2_1 _22468_ (.A0(_05146_),
    .A1(_09071_),
    .S(_04788_),
    .X(_05147_));
 sg13g2_nand2b_1 _22469_ (.Y(_05148_),
    .B(_04723_),
    .A_N(_00100_));
 sg13g2_nand2b_1 _22470_ (.Y(_05149_),
    .B(_04724_),
    .A_N(_00099_));
 sg13g2_inv_1 _22471_ (.Y(_05150_),
    .A(_00098_));
 sg13g2_buf_2 _22472_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05151_));
 sg13g2_nand2_1 _22473_ (.Y(_05152_),
    .A(net746),
    .B(_05151_));
 sg13g2_o21ai_1 _22474_ (.B1(_05152_),
    .Y(_05153_),
    .A1(net746),
    .A2(_00096_));
 sg13g2_a21oi_1 _22475_ (.A1(_04709_),
    .A2(_05153_),
    .Y(_05154_),
    .B1(net1022));
 sg13g2_o21ai_1 _22476_ (.B1(_05154_),
    .Y(_05155_),
    .A1(_00097_),
    .A2(net352));
 sg13g2_a221oi_1 _22477_ (.B2(_05150_),
    .C1(_05155_),
    .B1(_04705_),
    .A1(_08973_),
    .Y(_05156_),
    .A2(_04703_));
 sg13g2_a21oi_1 _22478_ (.A1(_08973_),
    .A2(_04692_),
    .Y(_05157_),
    .B1(net281));
 sg13g2_nand2b_1 _22479_ (.Y(_05158_),
    .B(\cpu.gpio.r_enable_in[1] ),
    .A_N(_05157_));
 sg13g2_nand4_1 _22480_ (.B(_05149_),
    .C(_05156_),
    .A(_05148_),
    .Y(_05159_),
    .D(_05158_));
 sg13g2_o21ai_1 _22481_ (.B1(_05159_),
    .Y(_05160_),
    .A1(_08950_),
    .A2(_05147_));
 sg13g2_nand2_1 _22482_ (.Y(_05161_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(net429));
 sg13g2_a22oi_1 _22483_ (.Y(_05162_),
    .B1(_04716_),
    .B2(\cpu.uart.r_r_invert ),
    .A2(net431),
    .A1(_09002_));
 sg13g2_a22oi_1 _22484_ (.Y(_05163_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[1] ),
    .A2(_04766_),
    .A1(\cpu.uart.r_div_value[9] ));
 sg13g2_nand3_1 _22485_ (.B(_05162_),
    .C(_05163_),
    .A(_05161_),
    .Y(_05164_));
 sg13g2_a22oi_1 _22486_ (.Y(_05165_),
    .B1(net353),
    .B2(_09742_),
    .A2(net452),
    .A1(\cpu.intr.r_timer_reload[17] ));
 sg13g2_a221oi_1 _22487_ (.B2(_09746_),
    .C1(net744),
    .B1(net391),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .Y(_05166_),
    .A2(net455));
 sg13g2_a21oi_1 _22488_ (.A1(net642),
    .A2(_05165_),
    .Y(_05167_),
    .B1(_05166_));
 sg13g2_nand2_1 _22489_ (.Y(_05168_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(_04863_));
 sg13g2_buf_2 _22490_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05169_));
 sg13g2_a22oi_1 _22491_ (.Y(_05170_),
    .B1(_04739_),
    .B2(_05169_),
    .A2(_04734_),
    .A1(_08997_));
 sg13g2_a22oi_1 _22492_ (.Y(_05171_),
    .B1(net556),
    .B2(_09877_),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_nand3_1 _22493_ (.B(_05170_),
    .C(_05171_),
    .A(_05168_),
    .Y(_05172_));
 sg13g2_nor2_1 _22494_ (.A(_05167_),
    .B(_05172_),
    .Y(_05173_));
 sg13g2_a21oi_1 _22495_ (.A1(_08997_),
    .A2(_04752_),
    .Y(_05174_),
    .B1(net382));
 sg13g2_nand2b_1 _22496_ (.Y(_05175_),
    .B(\cpu.intr.r_clock ),
    .A_N(_05174_));
 sg13g2_a21oi_1 _22497_ (.A1(_05173_),
    .A2(_05175_),
    .Y(_05176_),
    .B1(net583));
 sg13g2_a21oi_1 _22498_ (.A1(_04760_),
    .A2(_05164_),
    .Y(_05177_),
    .B1(_05176_));
 sg13g2_o21ai_1 _22499_ (.B1(_05177_),
    .Y(_05178_),
    .A1(_08954_),
    .A2(_05160_));
 sg13g2_mux2_1 _22500_ (.A0(_05138_),
    .A1(_05178_),
    .S(net986),
    .X(_05179_));
 sg13g2_nand2_1 _22501_ (.Y(_05180_),
    .A(net74),
    .B(_05179_));
 sg13g2_o21ai_1 _22502_ (.B1(_05180_),
    .Y(_05181_),
    .A1(_09881_),
    .A2(net74));
 sg13g2_nand2_1 _22503_ (.Y(_05182_),
    .A(net100),
    .B(_05181_));
 sg13g2_o21ai_1 _22504_ (.B1(_05182_),
    .Y(_01038_),
    .A1(net86),
    .A2(_05104_));
 sg13g2_nor2_1 _22505_ (.A(\cpu.dcache.r_data[0][2] ),
    .B(net532),
    .Y(_05183_));
 sg13g2_a22oi_1 _22506_ (.Y(_05184_),
    .B1(net455),
    .B2(\cpu.dcache.r_data[5][2] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_a22oi_1 _22507_ (.Y(_05185_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][2] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][2] ));
 sg13g2_mux2_1 _22508_ (.A0(\cpu.dcache.r_data[4][2] ),
    .A1(\cpu.dcache.r_data[6][2] ),
    .S(_08946_),
    .X(_05186_));
 sg13g2_a22oi_1 _22509_ (.Y(_05187_),
    .B1(_05186_),
    .B2(net632),
    .A2(_09157_),
    .A1(\cpu.dcache.r_data[7][2] ));
 sg13g2_nand2b_1 _22510_ (.Y(_05188_),
    .B(net726),
    .A_N(_05187_));
 sg13g2_nand4_1 _22511_ (.B(_05184_),
    .C(_05185_),
    .A(net532),
    .Y(_05189_),
    .D(_05188_));
 sg13g2_nor2b_1 _22512_ (.A(_05183_),
    .B_N(_05189_),
    .Y(_05190_));
 sg13g2_a22oi_1 _22513_ (.Y(_05191_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][18] ),
    .A2(net426),
    .A1(\cpu.dcache.r_data[5][18] ));
 sg13g2_a22oi_1 _22514_ (.Y(_05192_),
    .B1(net391),
    .B2(\cpu.dcache.r_data[6][18] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][18] ));
 sg13g2_inv_1 _22515_ (.Y(_05193_),
    .A(_00101_));
 sg13g2_a22oi_1 _22516_ (.Y(_05194_),
    .B1(net452),
    .B2(\cpu.dcache.r_data[7][18] ),
    .A2(net384),
    .A1(_05193_));
 sg13g2_a22oi_1 _22517_ (.Y(_05195_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][18] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][18] ));
 sg13g2_nand4_1 _22518_ (.B(_05192_),
    .C(_05194_),
    .A(_05191_),
    .Y(_05196_),
    .D(_05195_));
 sg13g2_and2_1 _22519_ (.A(net582),
    .B(_05196_),
    .X(_05197_));
 sg13g2_a21oi_1 _22520_ (.A1(net529),
    .A2(_05190_),
    .Y(_05198_),
    .B1(_05197_));
 sg13g2_a22oi_1 _22521_ (.Y(_05199_),
    .B1(_05190_),
    .B2(net945),
    .A2(_05196_),
    .A1(_04901_));
 sg13g2_a221oi_1 _22522_ (.B2(_09879_),
    .C1(net629),
    .B1(_04950_),
    .A1(net983),
    .Y(_05200_),
    .A2(_04943_));
 sg13g2_a21oi_1 _22523_ (.A1(_04648_),
    .A2(_05199_),
    .Y(_05201_),
    .B1(_05200_));
 sg13g2_nor2_1 _22524_ (.A(net707),
    .B(_05201_),
    .Y(_05202_));
 sg13g2_a21oi_1 _22525_ (.A1(_04670_),
    .A2(_05198_),
    .Y(_05203_),
    .B1(_05202_));
 sg13g2_nand2b_1 _22526_ (.Y(_05204_),
    .B(_04868_),
    .A_N(_00283_));
 sg13g2_o21ai_1 _22527_ (.B1(_05204_),
    .Y(_05205_),
    .A1(_00105_),
    .A2(net428));
 sg13g2_a21oi_1 _22528_ (.A1(_11581_),
    .A2(_04762_),
    .Y(_05206_),
    .B1(_05205_));
 sg13g2_buf_1 _22529_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05207_));
 sg13g2_a21oi_1 _22530_ (.A1(\cpu.spi.r_timeout[2] ),
    .A2(_04873_),
    .Y(_05208_),
    .B1(_08950_));
 sg13g2_o21ai_1 _22531_ (.B1(_05208_),
    .Y(_05209_),
    .A1(_00104_),
    .A2(_04774_));
 sg13g2_a221oi_1 _22532_ (.B2(_11582_),
    .C1(_05209_),
    .B1(_05142_),
    .A1(_05207_),
    .Y(_05210_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22533_ (.B1(_05210_),
    .Y(_05211_),
    .A1(net852),
    .A2(_05206_));
 sg13g2_a21oi_1 _22534_ (.A1(_09075_),
    .A2(_04788_),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_nor2_1 _22535_ (.A(_08954_),
    .B(_05212_),
    .Y(_05213_));
 sg13g2_nand2b_1 _22536_ (.Y(_05214_),
    .B(_04723_),
    .A_N(_00110_));
 sg13g2_nand2b_1 _22537_ (.Y(_05215_),
    .B(_04724_),
    .A_N(_00109_));
 sg13g2_inv_1 _22538_ (.Y(_05216_),
    .A(_00108_));
 sg13g2_buf_1 _22539_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05217_));
 sg13g2_nand2_1 _22540_ (.Y(_05218_),
    .A(net746),
    .B(_05217_));
 sg13g2_o21ai_1 _22541_ (.B1(_05218_),
    .Y(_05219_),
    .A1(net746),
    .A2(_00106_));
 sg13g2_a21oi_1 _22542_ (.A1(_04709_),
    .A2(_05219_),
    .Y(_05220_),
    .B1(net1022));
 sg13g2_o21ai_1 _22543_ (.B1(_05220_),
    .Y(_05221_),
    .A1(_00107_),
    .A2(_04718_));
 sg13g2_a221oi_1 _22544_ (.B2(_05216_),
    .C1(_05221_),
    .B1(_04705_),
    .A1(_08984_),
    .Y(_05222_),
    .A2(_04703_));
 sg13g2_a21oi_1 _22545_ (.A1(_08984_),
    .A2(_04692_),
    .Y(_05223_),
    .B1(net281));
 sg13g2_nand2b_1 _22546_ (.Y(_05224_),
    .B(\cpu.gpio.r_enable_in[2] ),
    .A_N(_05223_));
 sg13g2_nand4_1 _22547_ (.B(_05215_),
    .C(_05222_),
    .A(_05214_),
    .Y(_05225_),
    .D(_05224_));
 sg13g2_inv_1 _22548_ (.Y(_05226_),
    .A(\cpu.uart.r_div_value[2] ));
 sg13g2_a22oi_1 _22549_ (.Y(_05227_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[2] ),
    .A2(_04766_),
    .A1(_09717_));
 sg13g2_o21ai_1 _22550_ (.B1(_05227_),
    .Y(_05228_),
    .A1(_05226_),
    .A2(_04697_));
 sg13g2_a22oi_1 _22551_ (.Y(_05229_),
    .B1(net353),
    .B2(_09741_),
    .A2(net390),
    .A1(\cpu.intr.r_timer_reload[18] ));
 sg13g2_a221oi_1 _22552_ (.B2(\cpu.intr.r_timer_reload[2] ),
    .C1(net642),
    .B1(net390),
    .A1(\cpu.intr.r_clock_cmp[2] ),
    .Y(_05230_),
    .A2(net392));
 sg13g2_a21oi_1 _22553_ (.A1(net665),
    .A2(_05229_),
    .Y(_05231_),
    .B1(_05230_));
 sg13g2_nand2_1 _22554_ (.Y(_05232_),
    .A(_09886_),
    .B(net556));
 sg13g2_buf_1 _22555_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05233_));
 sg13g2_a22oi_1 _22556_ (.Y(_05234_),
    .B1(net382),
    .B2(_08994_),
    .A2(net430),
    .A1(_05233_));
 sg13g2_a22oi_1 _22557_ (.Y(_05235_),
    .B1(net555),
    .B2(\cpu.intr.r_timer_count[2] ),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_nand3_1 _22558_ (.B(_05234_),
    .C(_05235_),
    .A(_05232_),
    .Y(_05236_));
 sg13g2_nor2_1 _22559_ (.A(_05231_),
    .B(_05236_),
    .Y(_05237_));
 sg13g2_a21oi_1 _22560_ (.A1(_08994_),
    .A2(_04752_),
    .Y(_05238_),
    .B1(_04735_));
 sg13g2_nand2b_1 _22561_ (.Y(_05239_),
    .B(\cpu.intr.r_enable[2] ),
    .A_N(_05238_));
 sg13g2_a21oi_1 _22562_ (.A1(_05237_),
    .A2(_05239_),
    .Y(_05240_),
    .B1(_09737_));
 sg13g2_a221oi_1 _22563_ (.B2(_04760_),
    .C1(_05240_),
    .B1(_05228_),
    .A1(_05213_),
    .Y(_05241_),
    .A2(_05225_));
 sg13g2_nand2_1 _22564_ (.Y(_05242_),
    .A(net823),
    .B(_05241_));
 sg13g2_o21ai_1 _22565_ (.B1(_05242_),
    .Y(_05243_),
    .A1(net823),
    .A2(_05203_));
 sg13g2_mux2_1 _22566_ (.A0(net632),
    .A1(_05243_),
    .S(net75),
    .X(_05244_));
 sg13g2_o21ai_1 _22567_ (.B1(net165),
    .Y(_05245_),
    .A1(net885),
    .A2(_11216_));
 sg13g2_nand3_1 _22568_ (.B(net885),
    .C(_04957_),
    .A(net771),
    .Y(_05246_));
 sg13g2_o21ai_1 _22569_ (.B1(_05246_),
    .Y(_05247_),
    .A1(net625),
    .A2(_04313_));
 sg13g2_a221oi_1 _22570_ (.B2(net139),
    .C1(_04624_),
    .B1(_05247_),
    .A1(net770),
    .Y(_05248_),
    .A2(_05245_));
 sg13g2_a21oi_1 _22571_ (.A1(net86),
    .A2(_05244_),
    .Y(_01039_),
    .B1(_05248_));
 sg13g2_nand2_1 _22572_ (.Y(_05249_),
    .A(net624),
    .B(_04097_));
 sg13g2_o21ai_1 _22573_ (.B1(_05249_),
    .Y(_05250_),
    .A1(net624),
    .A2(_04346_));
 sg13g2_nand2_1 _22574_ (.Y(_05251_),
    .A(net624),
    .B(_04347_));
 sg13g2_a21oi_1 _22575_ (.A1(net165),
    .A2(_05251_),
    .Y(_05252_),
    .B1(net703));
 sg13g2_a21oi_1 _22576_ (.A1(net139),
    .A2(_05250_),
    .Y(_05253_),
    .B1(_05252_));
 sg13g2_nand2_1 _22577_ (.Y(_05254_),
    .A(\cpu.dcache.r_data[3][3] ),
    .B(net393));
 sg13g2_a22oi_1 _22578_ (.Y(_05255_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][3] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[0][3] ));
 sg13g2_a22oi_1 _22579_ (.Y(_05256_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][3] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][3] ));
 sg13g2_mux2_1 _22580_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(\cpu.dcache.r_data[7][3] ),
    .S(net594),
    .X(_05257_));
 sg13g2_a22oi_1 _22581_ (.Y(_05258_),
    .B1(_05257_),
    .B2(net692),
    .A2(net749),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_nand2b_1 _22582_ (.Y(_05259_),
    .B(net726),
    .A_N(_05258_));
 sg13g2_nand4_1 _22583_ (.B(_05255_),
    .C(_05256_),
    .A(_05254_),
    .Y(_05260_),
    .D(_05259_));
 sg13g2_inv_1 _22584_ (.Y(_05261_),
    .A(_00111_));
 sg13g2_a22oi_1 _22585_ (.Y(_05262_),
    .B1(net426),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net432),
    .A1(_05261_));
 sg13g2_a22oi_1 _22586_ (.Y(_05263_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][19] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_a22oi_1 _22587_ (.Y(_05264_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][19] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[7][19] ));
 sg13g2_a22oi_1 _22588_ (.Y(_05265_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][19] ));
 sg13g2_nand4_1 _22589_ (.B(_05263_),
    .C(_05264_),
    .A(_05262_),
    .Y(_05266_),
    .D(_05265_));
 sg13g2_buf_1 _22590_ (.A(_05266_),
    .X(_05267_));
 sg13g2_a22oi_1 _22591_ (.Y(_05268_),
    .B1(_05267_),
    .B2(_04901_),
    .A2(_05260_),
    .A1(net945));
 sg13g2_a221oi_1 _22592_ (.B2(_09729_),
    .C1(_04647_),
    .B1(_04994_),
    .A1(net983),
    .Y(_05269_),
    .A2(_04986_));
 sg13g2_a21oi_1 _22593_ (.A1(_04648_),
    .A2(_05268_),
    .Y(_05270_),
    .B1(_05269_));
 sg13g2_mux2_1 _22594_ (.A0(_05260_),
    .A1(_05267_),
    .S(net582),
    .X(_05271_));
 sg13g2_mux2_1 _22595_ (.A0(_05270_),
    .A1(_05271_),
    .S(_04669_),
    .X(_05272_));
 sg13g2_or2_1 _22596_ (.X(_05273_),
    .B(_05272_),
    .A(_11665_));
 sg13g2_a21o_1 _22597_ (.A2(_04692_),
    .A1(_08988_),
    .B1(net281),
    .X(_05274_));
 sg13g2_inv_1 _22598_ (.Y(_05275_),
    .A(_00119_));
 sg13g2_a22oi_1 _22599_ (.Y(_05276_),
    .B1(net492),
    .B2(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A2(_04977_),
    .A1(_05275_));
 sg13g2_inv_1 _22600_ (.Y(_05277_),
    .A(_00118_));
 sg13g2_nor2_1 _22601_ (.A(net666),
    .B(_00116_),
    .Y(_05278_));
 sg13g2_buf_1 _22602_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05279_));
 sg13g2_nor2b_1 _22603_ (.A(_09866_),
    .B_N(_05279_),
    .Y(_05280_));
 sg13g2_o21ai_1 _22604_ (.B1(net626),
    .Y(_05281_),
    .A1(_05278_),
    .A2(_05280_));
 sg13g2_o21ai_1 _22605_ (.B1(_05281_),
    .Y(_05282_),
    .A1(_00117_),
    .A2(net352));
 sg13g2_a221oi_1 _22606_ (.B2(_05277_),
    .C1(_05282_),
    .B1(_04705_),
    .A1(_08988_),
    .Y(_05283_),
    .A2(_04703_));
 sg13g2_o21ai_1 _22607_ (.B1(_05283_),
    .Y(_05284_),
    .A1(_04681_),
    .A2(_05276_));
 sg13g2_a21oi_1 _22608_ (.A1(\cpu.gpio.r_enable_in[3] ),
    .A2(_05274_),
    .Y(_05285_),
    .B1(_05284_));
 sg13g2_buf_1 _22609_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05286_));
 sg13g2_nor2_1 _22610_ (.A(_00114_),
    .B(_04774_),
    .Y(_05287_));
 sg13g2_a221oi_1 _22611_ (.B2(\cpu.spi.r_timeout[3] ),
    .C1(_05287_),
    .B1(_04873_),
    .A1(_05286_),
    .Y(_05288_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22612_ (.B1(_05288_),
    .Y(_05289_),
    .A1(_00115_),
    .A2(net381));
 sg13g2_a21oi_1 _22613_ (.A1(_09069_),
    .A2(_04788_),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_nor2_1 _22614_ (.A(_08956_),
    .B(_05290_),
    .Y(_05291_));
 sg13g2_a21o_1 _22615_ (.A2(_04752_),
    .A1(_08995_),
    .B1(net431),
    .X(_05292_));
 sg13g2_a22oi_1 _22616_ (.Y(_05293_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[3] ),
    .A2(_04933_),
    .A1(\cpu.intr.r_timer_count[3] ));
 sg13g2_nand2_1 _22617_ (.Y(_05294_),
    .A(_09891_),
    .B(net556));
 sg13g2_buf_2 _22618_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05295_));
 sg13g2_a22oi_1 _22619_ (.Y(_05296_),
    .B1(net382),
    .B2(_08995_),
    .A2(net430),
    .A1(_05295_));
 sg13g2_nand2_1 _22620_ (.Y(_05297_),
    .A(net880),
    .B(net726));
 sg13g2_mux2_1 _22621_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .S(net538),
    .X(_05298_));
 sg13g2_a22oi_1 _22622_ (.Y(_05299_),
    .B1(_05298_),
    .B2(net565),
    .A2(net749),
    .A1(_09740_));
 sg13g2_nor2_1 _22623_ (.A(_05297_),
    .B(_05299_),
    .Y(_05300_));
 sg13g2_a21oi_1 _22624_ (.A1(\cpu.intr.r_clock_cmp[3] ),
    .A2(net554),
    .Y(_05301_),
    .B1(_05300_));
 sg13g2_nand4_1 _22625_ (.B(_05294_),
    .C(_05296_),
    .A(_05293_),
    .Y(_05302_),
    .D(_05301_));
 sg13g2_a21oi_1 _22626_ (.A1(\cpu.intr.r_enable[3] ),
    .A2(_05292_),
    .Y(_05303_),
    .B1(_05302_));
 sg13g2_nor2_1 _22627_ (.A(net583),
    .B(_05303_),
    .Y(_05304_));
 sg13g2_nand2_1 _22628_ (.Y(_05305_),
    .A(_08954_),
    .B(_09737_));
 sg13g2_and2_1 _22629_ (.A(\cpu.uart.r_in[3] ),
    .B(_04768_),
    .X(_05306_));
 sg13g2_a221oi_1 _22630_ (.B2(\cpu.uart.r_div_value[11] ),
    .C1(_05306_),
    .B1(_04766_),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05307_),
    .A2(net429));
 sg13g2_o21ai_1 _22631_ (.B1(net986),
    .Y(_05308_),
    .A1(_05305_),
    .A2(_05307_));
 sg13g2_nor3_1 _22632_ (.A(_05291_),
    .B(_05304_),
    .C(_05308_),
    .Y(_05309_));
 sg13g2_o21ai_1 _22633_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_04675_),
    .A2(_05285_));
 sg13g2_nand3_1 _22634_ (.B(_05273_),
    .C(_05310_),
    .A(net74),
    .Y(_05311_));
 sg13g2_o21ai_1 _22635_ (.B1(_05311_),
    .Y(_05312_),
    .A1(net760),
    .A2(net75));
 sg13g2_mux2_1 _22636_ (.A0(_05253_),
    .A1(_05312_),
    .S(net100),
    .X(_01040_));
 sg13g2_o21ai_1 _22637_ (.B1(net165),
    .Y(_05313_),
    .A1(_11216_),
    .A2(_04097_));
 sg13g2_nand2_1 _22638_ (.Y(_05314_),
    .A(_04968_),
    .B(_04385_));
 sg13g2_o21ai_1 _22639_ (.B1(_05314_),
    .Y(_05315_),
    .A1(net625),
    .A2(_04382_));
 sg13g2_a22oi_1 _22640_ (.Y(_05316_),
    .B1(_05315_),
    .B2(net139),
    .A2(_05313_),
    .A1(net1038));
 sg13g2_o21ai_1 _22641_ (.B1(net708),
    .Y(_05317_),
    .A1(_10512_),
    .A2(_03392_));
 sg13g2_mux2_1 _22642_ (.A0(\cpu.dcache.r_data[4][4] ),
    .A1(\cpu.dcache.r_data[6][4] ),
    .S(net538),
    .X(_05318_));
 sg13g2_a22oi_1 _22643_ (.Y(_05319_),
    .B1(_05318_),
    .B2(net632),
    .A2(_09157_),
    .A1(\cpu.dcache.r_data[7][4] ));
 sg13g2_a22oi_1 _22644_ (.Y(_05320_),
    .B1(net458),
    .B2(\cpu.dcache.r_data[1][4] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_o21ai_1 _22645_ (.B1(_05320_),
    .Y(_05321_),
    .A1(_00121_),
    .A2(net532));
 sg13g2_a221oi_1 _22646_ (.B2(\cpu.dcache.r_data[5][4] ),
    .C1(_05321_),
    .B1(net455),
    .A1(\cpu.dcache.r_data[2][4] ),
    .Y(_05322_),
    .A2(net394));
 sg13g2_o21ai_1 _22647_ (.B1(_05322_),
    .Y(_05323_),
    .A1(net851),
    .A2(_05319_));
 sg13g2_inv_1 _22648_ (.Y(_05324_),
    .A(_00122_));
 sg13g2_a22oi_1 _22649_ (.Y(_05325_),
    .B1(net518),
    .B2(\cpu.dcache.r_data[2][20] ),
    .A2(net432),
    .A1(_05324_));
 sg13g2_a22oi_1 _22650_ (.Y(_05326_),
    .B1(net380),
    .B2(\cpu.dcache.r_data[3][20] ),
    .A2(_12326_),
    .A1(\cpu.dcache.r_data[5][20] ));
 sg13g2_a22oi_1 _22651_ (.Y(_05327_),
    .B1(_09858_),
    .B2(\cpu.dcache.r_data[4][20] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_a22oi_1 _22652_ (.Y(_05328_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[6][20] ),
    .A2(_11884_),
    .A1(\cpu.dcache.r_data[1][20] ));
 sg13g2_nand4_1 _22653_ (.B(_05326_),
    .C(_05327_),
    .A(_05325_),
    .Y(_05329_),
    .D(_05328_));
 sg13g2_buf_1 _22654_ (.A(_05329_),
    .X(_05330_));
 sg13g2_a22oi_1 _22655_ (.Y(_05331_),
    .B1(_05330_),
    .B2(_04901_),
    .A2(_05323_),
    .A1(net945));
 sg13g2_a221oi_1 _22656_ (.B2(net581),
    .C1(net629),
    .B1(_05020_),
    .A1(net983),
    .Y(_05332_),
    .A2(_05013_));
 sg13g2_a21oi_1 _22657_ (.A1(net629),
    .A2(_05331_),
    .Y(_05333_),
    .B1(_05332_));
 sg13g2_mux2_1 _22658_ (.A0(_05323_),
    .A1(_05330_),
    .S(net582),
    .X(_05334_));
 sg13g2_mux2_1 _22659_ (.A0(_05333_),
    .A1(_05334_),
    .S(net707),
    .X(_05335_));
 sg13g2_buf_1 _22660_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05336_));
 sg13g2_nor2_1 _22661_ (.A(_00125_),
    .B(_04774_),
    .Y(_05337_));
 sg13g2_a221oi_1 _22662_ (.B2(\cpu.spi.r_timeout[4] ),
    .C1(_05337_),
    .B1(_04873_),
    .A1(_05336_),
    .Y(_05338_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22663_ (.B1(_05338_),
    .Y(_05339_),
    .A1(_00126_),
    .A2(_04793_));
 sg13g2_a21oi_1 _22664_ (.A1(_09077_),
    .A2(_04788_),
    .Y(_05340_),
    .B1(_05339_));
 sg13g2_a22oi_1 _22665_ (.Y(_05341_),
    .B1(_04863_),
    .B2(\cpu.intr.r_timer_reload[4] ),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[4] ));
 sg13g2_nand2_1 _22666_ (.Y(_05342_),
    .A(_09896_),
    .B(net556));
 sg13g2_buf_2 _22667_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05343_));
 sg13g2_a22oi_1 _22668_ (.Y(_05344_),
    .B1(net430),
    .B2(_05343_),
    .A2(_04734_),
    .A1(_08992_));
 sg13g2_mux2_1 _22669_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net594),
    .X(_05345_));
 sg13g2_a22oi_1 _22670_ (.Y(_05346_),
    .B1(_05345_),
    .B2(net692),
    .A2(net749),
    .A1(_09763_));
 sg13g2_nor2_1 _22671_ (.A(_05297_),
    .B(_05346_),
    .Y(_05347_));
 sg13g2_a21oi_1 _22672_ (.A1(\cpu.intr.r_clock_cmp[4] ),
    .A2(net554),
    .Y(_05348_),
    .B1(_05347_));
 sg13g2_nand4_1 _22673_ (.B(_05342_),
    .C(_05344_),
    .A(_05341_),
    .Y(_05349_),
    .D(_05348_));
 sg13g2_o21ai_1 _22674_ (.B1(net851),
    .Y(_05350_),
    .A1(net538),
    .A2(net558));
 sg13g2_nor2_1 _22675_ (.A(_10514_),
    .B(_05350_),
    .Y(_05351_));
 sg13g2_inv_1 _22676_ (.Y(_05352_),
    .A(_08992_));
 sg13g2_a21oi_1 _22677_ (.A1(_05352_),
    .A2(_04752_),
    .Y(_05353_),
    .B1(net583));
 sg13g2_o21ai_1 _22678_ (.B1(_05353_),
    .Y(_05354_),
    .A1(_05349_),
    .A2(_05351_));
 sg13g2_o21ai_1 _22679_ (.B1(_05354_),
    .Y(_05355_),
    .A1(_08956_),
    .A2(_05340_));
 sg13g2_a21o_1 _22680_ (.A2(_04692_),
    .A1(_08974_),
    .B1(net281),
    .X(_05356_));
 sg13g2_a21oi_1 _22681_ (.A1(_08977_),
    .A2(_04754_),
    .Y(_05357_),
    .B1(_04716_));
 sg13g2_nor2b_1 _22682_ (.A(_05357_),
    .B_N(_08978_),
    .Y(_05358_));
 sg13g2_a22oi_1 _22683_ (.Y(_05359_),
    .B1(net465),
    .B2(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A2(net426),
    .A1(net7));
 sg13g2_buf_2 _22684_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05360_));
 sg13g2_nand3_1 _22685_ (.B(_05360_),
    .C(net426),
    .A(_09866_),
    .Y(_05361_));
 sg13g2_o21ai_1 _22686_ (.B1(_05361_),
    .Y(_05362_),
    .A1(net744),
    .A2(_05359_));
 sg13g2_buf_1 _22687_ (.A(net944),
    .X(_05363_));
 sg13g2_o21ai_1 _22688_ (.B1(net822),
    .Y(_05364_),
    .A1(_05358_),
    .A2(_05362_));
 sg13g2_nand3_1 _22689_ (.B(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .C(_04739_),
    .A(net822),
    .Y(_05365_));
 sg13g2_buf_2 _22690_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05366_));
 sg13g2_a22oi_1 _22691_ (.Y(_05367_),
    .B1(_04786_),
    .B2(_08977_),
    .A2(_04705_),
    .A1(_05366_));
 sg13g2_buf_2 _22692_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05368_));
 sg13g2_buf_2 _22693_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05369_));
 sg13g2_mux2_1 _22694_ (.A0(_05368_),
    .A1(_05369_),
    .S(net880),
    .X(_05370_));
 sg13g2_buf_2 _22695_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05371_));
 sg13g2_buf_2 _22696_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05372_));
 sg13g2_a22oi_1 _22697_ (.Y(_05373_),
    .B1(_04754_),
    .B2(_05372_),
    .A2(_04716_),
    .A1(_05371_));
 sg13g2_nor2_1 _22698_ (.A(_02855_),
    .B(_05373_),
    .Y(_05374_));
 sg13g2_a221oi_1 _22699_ (.B2(_05370_),
    .C1(_05374_),
    .B1(net626),
    .A1(_08974_),
    .Y(_05375_),
    .A2(_04703_));
 sg13g2_nand4_1 _22700_ (.B(_05365_),
    .C(_05367_),
    .A(_05364_),
    .Y(_05376_),
    .D(_05375_));
 sg13g2_a21oi_1 _22701_ (.A1(\cpu.gpio.r_enable_in[4] ),
    .A2(_05356_),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_nor2_1 _22702_ (.A(_04675_),
    .B(_05377_),
    .Y(_05378_));
 sg13g2_nor3_1 _22703_ (.A(_04760_),
    .B(_05355_),
    .C(_05378_),
    .Y(_05379_));
 sg13g2_a221oi_1 _22704_ (.B2(\cpu.uart.r_in[4] ),
    .C1(_05305_),
    .B1(_04768_),
    .A1(\cpu.uart.r_div_value[4] ),
    .Y(_05380_),
    .A2(net429));
 sg13g2_o21ai_1 _22705_ (.B1(net986),
    .Y(_05381_),
    .A1(_05379_),
    .A2(_05380_));
 sg13g2_o21ai_1 _22706_ (.B1(_05381_),
    .Y(_05382_),
    .A1(net823),
    .A2(_05335_));
 sg13g2_nand2_1 _22707_ (.Y(_05383_),
    .A(net75),
    .B(_05382_));
 sg13g2_nand3_1 _22708_ (.B(_05317_),
    .C(_05383_),
    .A(net101),
    .Y(_05384_));
 sg13g2_o21ai_1 _22709_ (.B1(_05384_),
    .Y(_01041_),
    .A1(net86),
    .A2(_05316_));
 sg13g2_nand2_1 _22710_ (.Y(_05385_),
    .A(net624),
    .B(_04414_));
 sg13g2_o21ai_1 _22711_ (.B1(_05385_),
    .Y(_05386_),
    .A1(net625),
    .A2(_04411_));
 sg13g2_and2_1 _22712_ (.A(net948),
    .B(net164),
    .X(_05387_));
 sg13g2_a21oi_1 _22713_ (.A1(net139),
    .A2(_05386_),
    .Y(_05388_),
    .B1(_05387_));
 sg13g2_a22oi_1 _22714_ (.Y(_05389_),
    .B1(net353),
    .B2(\cpu.dcache.r_data[6][5] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_a22oi_1 _22715_ (.Y(_05390_),
    .B1(net354),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[5][5] ));
 sg13g2_inv_1 _22716_ (.Y(_05391_),
    .A(_00128_));
 sg13g2_a22oi_1 _22717_ (.Y(_05392_),
    .B1(_02745_),
    .B2(\cpu.dcache.r_data[7][5] ),
    .A2(net384),
    .A1(_05391_));
 sg13g2_a22oi_1 _22718_ (.Y(_05393_),
    .B1(net400),
    .B2(\cpu.dcache.r_data[4][5] ),
    .A2(_12122_),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_nand4_1 _22719_ (.B(_05390_),
    .C(_05392_),
    .A(_05389_),
    .Y(_05394_),
    .D(_05393_));
 sg13g2_buf_1 _22720_ (.A(_05394_),
    .X(_05395_));
 sg13g2_inv_1 _22721_ (.Y(_05396_),
    .A(_00129_));
 sg13g2_a22oi_1 _22722_ (.Y(_05397_),
    .B1(_12327_),
    .B2(\cpu.dcache.r_data[5][21] ),
    .A2(net384),
    .A1(_05396_));
 sg13g2_a22oi_1 _22723_ (.Y(_05398_),
    .B1(net354),
    .B2(\cpu.dcache.r_data[1][21] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][21] ));
 sg13g2_a22oi_1 _22724_ (.Y(_05399_),
    .B1(_12441_),
    .B2(\cpu.dcache.r_data[6][21] ),
    .A2(_02744_),
    .A1(\cpu.dcache.r_data[7][21] ));
 sg13g2_a22oi_1 _22725_ (.Y(_05400_),
    .B1(net400),
    .B2(\cpu.dcache.r_data[4][21] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_nand4_1 _22726_ (.B(_05398_),
    .C(_05399_),
    .A(_05397_),
    .Y(_05401_),
    .D(_05400_));
 sg13g2_buf_1 _22727_ (.A(_05401_),
    .X(_05402_));
 sg13g2_a22oi_1 _22728_ (.Y(_05403_),
    .B1(_05402_),
    .B2(_04901_),
    .A2(_05395_),
    .A1(net945));
 sg13g2_a221oi_1 _22729_ (.B2(net581),
    .C1(net629),
    .B1(_05044_),
    .A1(net983),
    .Y(_05404_),
    .A2(_05038_));
 sg13g2_a21o_1 _22730_ (.A2(_05403_),
    .A1(net629),
    .B1(_05404_),
    .X(_05405_));
 sg13g2_and2_1 _22731_ (.A(_09868_),
    .B(_05402_),
    .X(_05406_));
 sg13g2_a21oi_1 _22732_ (.A1(net529),
    .A2(_05395_),
    .Y(_05407_),
    .B1(_05406_));
 sg13g2_mux2_1 _22733_ (.A0(_05405_),
    .A1(_05407_),
    .S(net628),
    .X(_05408_));
 sg13g2_a21o_1 _22734_ (.A2(_04692_),
    .A1(_08981_),
    .B1(net281),
    .X(_05409_));
 sg13g2_nor3_1 _22735_ (.A(net666),
    .B(_00138_),
    .C(net748),
    .Y(_05410_));
 sg13g2_a22oi_1 _22736_ (.Y(_05411_),
    .B1(net400),
    .B2(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A2(_12327_),
    .A1(net8));
 sg13g2_a21oi_1 _22737_ (.A1(_08985_),
    .A2(net382),
    .Y(_05412_),
    .B1(_04716_));
 sg13g2_nand2b_1 _22738_ (.Y(_05413_),
    .B(_08986_),
    .A_N(_05412_));
 sg13g2_o21ai_1 _22739_ (.B1(_05413_),
    .Y(_05414_),
    .A1(_09867_),
    .A2(_05411_));
 sg13g2_or2_1 _22740_ (.X(_05415_),
    .B(_05414_),
    .A(_05410_));
 sg13g2_nand2_1 _22741_ (.Y(_05416_),
    .A(_04681_),
    .B(_04734_));
 sg13g2_nor2_1 _22742_ (.A(_00136_),
    .B(_05416_),
    .Y(_05417_));
 sg13g2_a221oi_1 _22743_ (.B2(_08985_),
    .C1(_05417_),
    .B1(_04786_),
    .A1(_08981_),
    .Y(_05418_),
    .A2(_04703_));
 sg13g2_or2_1 _22744_ (.X(_05419_),
    .B(_04714_),
    .A(net627));
 sg13g2_buf_1 _22745_ (.A(_05419_),
    .X(_05420_));
 sg13g2_nor2_1 _22746_ (.A(_00135_),
    .B(_05420_),
    .Y(_05421_));
 sg13g2_nor3_1 _22747_ (.A(_00137_),
    .B(_04701_),
    .C(net557),
    .Y(_05422_));
 sg13g2_o21ai_1 _22748_ (.B1(_11602_),
    .Y(_05423_),
    .A1(_05421_),
    .A2(_05422_));
 sg13g2_nor2_1 _22749_ (.A(net666),
    .B(_00134_),
    .Y(_05424_));
 sg13g2_buf_2 _22750_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05425_));
 sg13g2_nor2b_1 _22751_ (.A(_11687_),
    .B_N(_05425_),
    .Y(_05426_));
 sg13g2_o21ai_1 _22752_ (.B1(net626),
    .Y(_05427_),
    .A1(_05424_),
    .A2(_05426_));
 sg13g2_nand3_1 _22753_ (.B(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .C(net383),
    .A(net822),
    .Y(_05428_));
 sg13g2_nand4_1 _22754_ (.B(_05423_),
    .C(_05427_),
    .A(_05418_),
    .Y(_05429_),
    .D(_05428_));
 sg13g2_a221oi_1 _22755_ (.B2(net822),
    .C1(_05429_),
    .B1(_05415_),
    .A1(\cpu.gpio.r_enable_in[5] ),
    .Y(_05430_),
    .A2(_05409_));
 sg13g2_buf_1 _22756_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05431_));
 sg13g2_nor2_1 _22757_ (.A(_00132_),
    .B(_04774_),
    .Y(_05432_));
 sg13g2_a221oi_1 _22758_ (.B2(\cpu.spi.r_timeout[5] ),
    .C1(_05432_),
    .B1(_04873_),
    .A1(_05431_),
    .Y(_05433_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22759_ (.B1(_05433_),
    .Y(_05434_),
    .A1(_00133_),
    .A2(_04793_));
 sg13g2_a21oi_1 _22760_ (.A1(_09076_),
    .A2(_04788_),
    .Y(_05435_),
    .B1(_05434_));
 sg13g2_nor2_1 _22761_ (.A(_08956_),
    .B(_05435_),
    .Y(_05436_));
 sg13g2_a22oi_1 _22762_ (.Y(_05437_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_nor2_1 _22763_ (.A(_05305_),
    .B(_05437_),
    .Y(_05438_));
 sg13g2_a21o_1 _22764_ (.A2(_04752_),
    .A1(_08999_),
    .B1(net382),
    .X(_05439_));
 sg13g2_a22oi_1 _22765_ (.Y(_05440_),
    .B1(net556),
    .B2(_09901_),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[5] ));
 sg13g2_nand2_1 _22766_ (.Y(_05441_),
    .A(_08999_),
    .B(net431));
 sg13g2_buf_1 _22767_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05442_));
 sg13g2_mux2_1 _22768_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .S(net744),
    .X(_05443_));
 sg13g2_a22oi_1 _22769_ (.Y(_05444_),
    .B1(_05443_),
    .B2(net392),
    .A2(net430),
    .A1(_05442_));
 sg13g2_a22oi_1 _22770_ (.Y(_05445_),
    .B1(net391),
    .B2(_09764_),
    .A2(net452),
    .A1(\cpu.intr.r_timer_reload[21] ));
 sg13g2_inv_1 _22771_ (.Y(_05446_),
    .A(_05445_));
 sg13g2_a22oi_1 _22772_ (.Y(_05447_),
    .B1(_05446_),
    .B2(net642),
    .A2(_04863_),
    .A1(\cpu.intr.r_timer_reload[5] ));
 sg13g2_nand4_1 _22773_ (.B(_05441_),
    .C(_05444_),
    .A(_05440_),
    .Y(_05448_),
    .D(_05447_));
 sg13g2_a21oi_1 _22774_ (.A1(_08998_),
    .A2(_05439_),
    .Y(_05449_),
    .B1(_05448_));
 sg13g2_nor2_1 _22775_ (.A(net583),
    .B(_05449_),
    .Y(_05450_));
 sg13g2_nor3_1 _22776_ (.A(_05436_),
    .B(_05438_),
    .C(_05450_),
    .Y(_05451_));
 sg13g2_o21ai_1 _22777_ (.B1(_05451_),
    .Y(_05452_),
    .A1(_04675_),
    .A2(_05430_));
 sg13g2_nand2_1 _22778_ (.Y(_05453_),
    .A(net823),
    .B(_05452_));
 sg13g2_o21ai_1 _22779_ (.B1(_05453_),
    .Y(_05454_),
    .A1(net823),
    .A2(_05408_));
 sg13g2_nor2_1 _22780_ (.A(net716),
    .B(net75),
    .Y(_05455_));
 sg13g2_a221oi_1 _22781_ (.B2(_05454_),
    .C1(_05455_),
    .B1(net75),
    .A1(net761),
    .Y(_05456_),
    .A2(_11220_));
 sg13g2_a21oi_1 _22782_ (.A1(net84),
    .A2(_05388_),
    .Y(_01042_),
    .B1(_05456_));
 sg13g2_nand2_1 _22783_ (.Y(_05457_),
    .A(net624),
    .B(_04449_));
 sg13g2_o21ai_1 _22784_ (.B1(_05457_),
    .Y(_05458_),
    .A1(net624),
    .A2(_04446_));
 sg13g2_nand2b_1 _22785_ (.Y(_05459_),
    .B(net164),
    .A_N(net947));
 sg13g2_o21ai_1 _22786_ (.B1(_05459_),
    .Y(_05460_),
    .A1(net164),
    .A2(_05458_));
 sg13g2_a22oi_1 _22787_ (.Y(_05461_),
    .B1(_04768_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_nor2_1 _22788_ (.A(_05305_),
    .B(_05461_),
    .Y(_05462_));
 sg13g2_buf_1 _22789_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05463_));
 sg13g2_nor2_1 _22790_ (.A(_00144_),
    .B(_04774_),
    .Y(_05464_));
 sg13g2_a221oi_1 _22791_ (.B2(\cpu.spi.r_timeout[6] ),
    .C1(_05464_),
    .B1(_04873_),
    .A1(_05463_),
    .Y(_05465_),
    .A2(_04796_));
 sg13g2_o21ai_1 _22792_ (.B1(_05465_),
    .Y(_05466_),
    .A1(_00145_),
    .A2(net381));
 sg13g2_a21oi_1 _22793_ (.A1(_09070_),
    .A2(_04788_),
    .Y(_05467_),
    .B1(_05466_));
 sg13g2_nand2_1 _22794_ (.Y(_05468_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_04933_));
 sg13g2_a22oi_1 _22795_ (.Y(_05469_),
    .B1(_04928_),
    .B2(\cpu.intr.r_timer_reload[6] ),
    .A2(net553),
    .A1(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_buf_1 _22796_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05470_));
 sg13g2_a22oi_1 _22797_ (.Y(_05471_),
    .B1(net492),
    .B2(_09906_),
    .A2(net430),
    .A1(_05470_));
 sg13g2_nand3_1 _22798_ (.B(_05469_),
    .C(_05471_),
    .A(_05468_),
    .Y(_05472_));
 sg13g2_a22oi_1 _22799_ (.Y(_05473_),
    .B1(net353),
    .B2(_09765_),
    .A2(net390),
    .A1(\cpu.intr.r_timer_reload[22] ));
 sg13g2_a21oi_1 _22800_ (.A1(\cpu.intr.r_clock_cmp[6] ),
    .A2(net392),
    .Y(_05474_),
    .B1(net665));
 sg13g2_a21oi_1 _22801_ (.A1(net582),
    .A2(_05473_),
    .Y(_05475_),
    .B1(_05474_));
 sg13g2_o21ai_1 _22802_ (.B1(_04858_),
    .Y(_05476_),
    .A1(_05472_),
    .A2(_05475_));
 sg13g2_o21ai_1 _22803_ (.B1(_05476_),
    .Y(_05477_),
    .A1(_08956_),
    .A2(_05467_));
 sg13g2_nand3_1 _22804_ (.B(_08969_),
    .C(_04692_),
    .A(_08968_),
    .Y(_05478_));
 sg13g2_nand2_1 _22805_ (.Y(_05479_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_04927_));
 sg13g2_a22oi_1 _22806_ (.Y(_05480_),
    .B1(_04740_),
    .B2(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A2(_04716_),
    .A1(_08989_));
 sg13g2_nand2_1 _22807_ (.Y(_05481_),
    .A(net9),
    .B(net554));
 sg13g2_nand3_1 _22808_ (.B(_05480_),
    .C(_05481_),
    .A(_05479_),
    .Y(_05482_));
 sg13g2_nand2b_1 _22809_ (.Y(_05483_),
    .B(_04723_),
    .A_N(_00150_));
 sg13g2_buf_1 _22810_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05484_));
 sg13g2_nand2_1 _22811_ (.Y(_05485_),
    .A(net746),
    .B(_05484_));
 sg13g2_o21ai_1 _22812_ (.B1(_05485_),
    .Y(_05486_),
    .A1(net666),
    .A2(_00146_));
 sg13g2_nor2_1 _22813_ (.A(_00148_),
    .B(_05416_),
    .Y(_05487_));
 sg13g2_a221oi_1 _22814_ (.B2(_05486_),
    .C1(_05487_),
    .B1(net626),
    .A1(_08969_),
    .Y(_05488_),
    .A2(_04703_));
 sg13g2_and3_1 _22815_ (.X(_05489_),
    .A(_08989_),
    .B(net822),
    .C(net382));
 sg13g2_o21ai_1 _22816_ (.B1(\cpu.gpio.r_enable_io[6] ),
    .Y(_05490_),
    .A1(_04786_),
    .A2(_05489_));
 sg13g2_nand2b_1 _22817_ (.Y(_05491_),
    .B(_04755_),
    .A_N(_00149_));
 sg13g2_o21ai_1 _22818_ (.B1(_05491_),
    .Y(_05492_),
    .A1(_00147_),
    .A2(_05420_));
 sg13g2_a22oi_1 _22819_ (.Y(_05493_),
    .B1(_05492_),
    .B2(_11602_),
    .A2(net281),
    .A1(_08968_));
 sg13g2_nand4_1 _22820_ (.B(_05488_),
    .C(_05490_),
    .A(_05483_),
    .Y(_05494_),
    .D(_05493_));
 sg13g2_a21oi_1 _22821_ (.A1(net822),
    .A2(_05482_),
    .Y(_05495_),
    .B1(_05494_));
 sg13g2_a21oi_1 _22822_ (.A1(_05478_),
    .A2(_05495_),
    .Y(_05496_),
    .B1(_04675_));
 sg13g2_nor3_1 _22823_ (.A(_05462_),
    .B(_05477_),
    .C(_05496_),
    .Y(_05497_));
 sg13g2_o21ai_1 _22824_ (.B1(_05071_),
    .Y(_05498_),
    .A1(_11668_),
    .A2(_05064_));
 sg13g2_inv_1 _22825_ (.Y(_05499_),
    .A(_05498_));
 sg13g2_a22oi_1 _22826_ (.Y(_05500_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net426),
    .A1(\cpu.dcache.r_data[5][22] ));
 sg13g2_a22oi_1 _22827_ (.Y(_05501_),
    .B1(net391),
    .B2(\cpu.dcache.r_data[6][22] ),
    .A2(net457),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_inv_1 _22828_ (.Y(_05502_),
    .A(_00141_));
 sg13g2_a22oi_1 _22829_ (.Y(_05503_),
    .B1(_02744_),
    .B2(\cpu.dcache.r_data[7][22] ),
    .A2(net384),
    .A1(_05502_));
 sg13g2_a22oi_1 _22830_ (.Y(_05504_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][22] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_nand4_1 _22831_ (.B(_05501_),
    .C(_05503_),
    .A(_05500_),
    .Y(_05505_),
    .D(_05504_));
 sg13g2_nand2_1 _22832_ (.Y(_05506_),
    .A(net665),
    .B(_05505_));
 sg13g2_mux2_1 _22833_ (.A0(_05499_),
    .A1(_05506_),
    .S(_04647_),
    .X(_05507_));
 sg13g2_a22oi_1 _22834_ (.Y(_05508_),
    .B1(net353),
    .B2(\cpu.dcache.r_data[6][6] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_a22oi_1 _22835_ (.Y(_05509_),
    .B1(net354),
    .B2(\cpu.dcache.r_data[1][6] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[5][6] ));
 sg13g2_inv_1 _22836_ (.Y(_05510_),
    .A(_00140_));
 sg13g2_a22oi_1 _22837_ (.Y(_05511_),
    .B1(net452),
    .B2(\cpu.dcache.r_data[7][6] ),
    .A2(net384),
    .A1(_05510_));
 sg13g2_a22oi_1 _22838_ (.Y(_05512_),
    .B1(net465),
    .B2(\cpu.dcache.r_data[4][6] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][6] ));
 sg13g2_and4_1 _22839_ (.A(_05508_),
    .B(_05509_),
    .C(_05511_),
    .D(_05512_),
    .X(_05513_));
 sg13g2_buf_1 _22840_ (.A(_05513_),
    .X(_05514_));
 sg13g2_mux2_1 _22841_ (.A0(_05507_),
    .A1(_05514_),
    .S(_04657_),
    .X(_05515_));
 sg13g2_o21ai_1 _22842_ (.B1(_05506_),
    .Y(_05516_),
    .A1(_09868_),
    .A2(_05514_));
 sg13g2_nand2_1 _22843_ (.Y(_05517_),
    .A(net707),
    .B(_05516_));
 sg13g2_o21ai_1 _22844_ (.B1(_05517_),
    .Y(_05518_),
    .A1(net628),
    .A2(_05515_));
 sg13g2_nor2_1 _22845_ (.A(net823),
    .B(_05518_),
    .Y(_05519_));
 sg13g2_a21oi_1 _22846_ (.A1(net823),
    .A2(_05497_),
    .Y(_05520_),
    .B1(_05519_));
 sg13g2_nor2_1 _22847_ (.A(net715),
    .B(net74),
    .Y(_05521_));
 sg13g2_a221oi_1 _22848_ (.B2(_05520_),
    .C1(_05521_),
    .B1(net75),
    .A1(net761),
    .Y(_05522_),
    .A2(_11220_));
 sg13g2_a21oi_1 _22849_ (.A1(net84),
    .A2(_05460_),
    .Y(_01043_),
    .B1(_05522_));
 sg13g2_a21oi_1 _22850_ (.A1(_04957_),
    .A2(_04477_),
    .Y(_05523_),
    .B1(net164));
 sg13g2_o21ai_1 _22851_ (.B1(_05523_),
    .Y(_05524_),
    .A1(net625),
    .A2(_04476_));
 sg13g2_o21ai_1 _22852_ (.B1(_05524_),
    .Y(_05525_),
    .A1(\cpu.ex.pc[7] ),
    .A2(net139));
 sg13g2_mux2_1 _22853_ (.A0(net956),
    .A1(_04921_),
    .S(_04805_),
    .X(_05526_));
 sg13g2_nand2_1 _22854_ (.Y(_05527_),
    .A(_04836_),
    .B(_05526_));
 sg13g2_o21ai_1 _22855_ (.B1(_05527_),
    .Y(_01044_),
    .A1(_04625_),
    .A2(_05525_));
 sg13g2_nor3_1 _22856_ (.A(_11216_),
    .B(net164),
    .C(_04509_),
    .Y(_05528_));
 sg13g2_a21o_1 _22857_ (.A2(net164),
    .A1(net950),
    .B1(_05528_),
    .X(_05529_));
 sg13g2_a22oi_1 _22858_ (.Y(_05530_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[8] ),
    .A2(net492),
    .A1(_09916_));
 sg13g2_buf_1 _22859_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05531_));
 sg13g2_mux2_1 _22860_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(\cpu.intr.r_clock_cmp[24] ),
    .S(net665),
    .X(_05532_));
 sg13g2_a22oi_1 _22861_ (.Y(_05533_),
    .B1(_05532_),
    .B2(net392),
    .A2(net383),
    .A1(_05531_));
 sg13g2_nand2_1 _22862_ (.Y(_05534_),
    .A(_09745_),
    .B(net555));
 sg13g2_nand3_1 _22863_ (.B(_05533_),
    .C(_05534_),
    .A(_05530_),
    .Y(_05535_));
 sg13g2_nand2_1 _22864_ (.Y(_05536_),
    .A(_09879_),
    .B(_04664_));
 sg13g2_o21ai_1 _22865_ (.B1(_05536_),
    .Y(_05537_),
    .A1(net529),
    .A2(_04635_));
 sg13g2_a22oi_1 _22866_ (.Y(_05538_),
    .B1(_05537_),
    .B2(net628),
    .A2(_05535_),
    .A1(_04926_));
 sg13g2_o21ai_1 _22867_ (.B1(_04923_),
    .Y(_05539_),
    .A1(net943),
    .A2(_05538_));
 sg13g2_nor2b_1 _22868_ (.A(net74),
    .B_N(net1085),
    .Y(_05540_));
 sg13g2_a221oi_1 _22869_ (.B2(_05539_),
    .C1(_05540_),
    .B1(_04626_),
    .A1(_09037_),
    .Y(_05541_),
    .A2(_11220_));
 sg13g2_a221oi_1 _22870_ (.B2(_04967_),
    .C1(_05541_),
    .B1(_05529_),
    .A1(_04508_),
    .Y(_01045_),
    .A2(_04971_));
 sg13g2_nor2_1 _22871_ (.A(_11226_),
    .B(net139),
    .Y(_05542_));
 sg13g2_and2_1 _22872_ (.A(_04968_),
    .B(_04538_),
    .X(_05543_));
 sg13g2_a21oi_1 _22873_ (.A1(_11216_),
    .A2(_04536_),
    .Y(_05544_),
    .B1(_05543_));
 sg13g2_a22oi_1 _22874_ (.Y(_05545_),
    .B1(net427),
    .B2(\cpu.intr.r_timer_reload[9] ),
    .A2(net492),
    .A1(_09923_));
 sg13g2_buf_1 _22875_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05546_));
 sg13g2_mux2_1 _22876_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(\cpu.intr.r_clock_cmp[25] ),
    .S(net665),
    .X(_05547_));
 sg13g2_a22oi_1 _22877_ (.Y(_05548_),
    .B1(_05547_),
    .B2(net392),
    .A2(net383),
    .A1(_05546_));
 sg13g2_nand2_1 _22878_ (.Y(_05549_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(net555));
 sg13g2_nand3_1 _22879_ (.B(_05548_),
    .C(_05549_),
    .A(_05545_),
    .Y(_05550_));
 sg13g2_mux2_1 _22880_ (.A0(_05128_),
    .A1(_05134_),
    .S(net530),
    .X(_05551_));
 sg13g2_a22oi_1 _22881_ (.Y(_05552_),
    .B1(_05551_),
    .B2(_04670_),
    .A2(_05550_),
    .A1(_04926_));
 sg13g2_o21ai_1 _22882_ (.B1(_04923_),
    .Y(_05553_),
    .A1(net943),
    .A2(_05552_));
 sg13g2_nand2b_1 _22883_ (.Y(_05554_),
    .B(_03396_),
    .A_N(_09985_));
 sg13g2_o21ai_1 _22884_ (.B1(_05554_),
    .Y(_05555_),
    .A1(net36),
    .A2(_05553_));
 sg13g2_a221oi_1 _22885_ (.B2(_04963_),
    .C1(_05555_),
    .B1(_05544_),
    .A1(_08462_),
    .Y(_01046_),
    .A2(_05542_));
 sg13g2_inv_1 _22886_ (.Y(_05556_),
    .A(\cpu.dec.r_rd[0] ));
 sg13g2_o21ai_1 _22887_ (.B1(_04965_),
    .Y(_05557_),
    .A1(_03294_),
    .A2(_05556_));
 sg13g2_mux2_1 _22888_ (.A0(_09964_),
    .A1(_05557_),
    .S(_04967_),
    .X(_01047_));
 sg13g2_nor2b_1 _22889_ (.A(_03294_),
    .B_N(\cpu.dec.r_rd[1] ),
    .Y(_05558_));
 sg13g2_o21ai_1 _22890_ (.B1(net106),
    .Y(_05559_),
    .A1(_05098_),
    .A2(_05558_));
 sg13g2_o21ai_1 _22891_ (.B1(_05559_),
    .Y(_01048_),
    .A1(_03370_),
    .A2(net84));
 sg13g2_nor3_1 _22892_ (.A(_03294_),
    .B(_09095_),
    .C(net164),
    .Y(_05560_));
 sg13g2_nand3_1 _22893_ (.B(net106),
    .C(_05560_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05561_));
 sg13g2_o21ai_1 _22894_ (.B1(_05561_),
    .Y(_01049_),
    .A1(_09968_),
    .A2(_05002_));
 sg13g2_inv_1 _22895_ (.Y(_05562_),
    .A(net1076));
 sg13g2_nand3_1 _22896_ (.B(net106),
    .C(_05560_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05563_));
 sg13g2_o21ai_1 _22897_ (.B1(_05563_),
    .Y(_01050_),
    .A1(_05562_),
    .A2(_05002_));
 sg13g2_mux2_1 _22898_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_04836_),
    .X(_01051_));
 sg13g2_buf_1 _22899_ (.A(_09808_),
    .X(_05564_));
 sg13g2_buf_1 _22900_ (.A(net942),
    .X(_05565_));
 sg13g2_nand2_1 _22901_ (.Y(_05566_),
    .A(net821),
    .B(net100));
 sg13g2_o21ai_1 _22902_ (.B1(_05566_),
    .Y(_01052_),
    .A1(_11019_),
    .A2(net86));
 sg13g2_buf_1 _22903_ (.A(net943),
    .X(_05567_));
 sg13g2_nand2_1 _22904_ (.Y(_05568_),
    .A(_11068_),
    .B(_11074_));
 sg13g2_a22oi_1 _22905_ (.Y(_05569_),
    .B1(net527),
    .B2(_10178_),
    .A2(net528),
    .A1(net1075));
 sg13g2_nor2_1 _22906_ (.A(net820),
    .B(_05569_),
    .Y(_05570_));
 sg13g2_a21oi_1 _22907_ (.A1(net820),
    .A2(_05568_),
    .Y(_05571_),
    .B1(_05570_));
 sg13g2_nand2_1 _22908_ (.Y(_05572_),
    .A(\cpu.dcache.wdata[10] ),
    .B(net100));
 sg13g2_o21ai_1 _22909_ (.B1(_05572_),
    .Y(_01053_),
    .A1(net86),
    .A2(_05571_));
 sg13g2_nand2b_1 _22910_ (.Y(_05573_),
    .B(_11109_),
    .A_N(_11103_));
 sg13g2_mux2_1 _22911_ (.A0(_10149_),
    .A1(_05573_),
    .S(net820),
    .X(_05574_));
 sg13g2_mux2_1 _22912_ (.A0(_09937_),
    .A1(_05574_),
    .S(net85),
    .X(_01054_));
 sg13g2_nor2_1 _22913_ (.A(net820),
    .B(_10338_),
    .Y(_05575_));
 sg13g2_a21oi_1 _22914_ (.A1(net820),
    .A2(_10482_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_nand2_1 _22915_ (.Y(_05577_),
    .A(_09942_),
    .B(net100));
 sg13g2_o21ai_1 _22916_ (.B1(_05577_),
    .Y(_01055_),
    .A1(net86),
    .A2(_05576_));
 sg13g2_nand2_1 _22917_ (.Y(_05578_),
    .A(_10453_),
    .B(_10454_));
 sg13g2_nand2_1 _22918_ (.Y(_05579_),
    .A(_04924_),
    .B(_05578_));
 sg13g2_o21ai_1 _22919_ (.B1(_05579_),
    .Y(_05580_),
    .A1(_05567_),
    .A2(_10310_));
 sg13g2_nand2_1 _22920_ (.Y(_05581_),
    .A(net85),
    .B(_05580_));
 sg13g2_o21ai_1 _22921_ (.B1(_05581_),
    .Y(_01056_),
    .A1(_11737_),
    .A2(net84));
 sg13g2_nand2_1 _22922_ (.Y(_05582_),
    .A(_10429_),
    .B(_10430_));
 sg13g2_mux2_1 _22923_ (.A0(_10264_),
    .A1(_05582_),
    .S(net943),
    .X(_05583_));
 sg13g2_nand2_1 _22924_ (.Y(_05584_),
    .A(net106),
    .B(_05583_));
 sg13g2_o21ai_1 _22925_ (.B1(_05584_),
    .Y(_01057_),
    .A1(_11747_),
    .A2(net84));
 sg13g2_mux2_1 _22926_ (.A0(_10225_),
    .A1(_10397_),
    .S(net820),
    .X(_05585_));
 sg13g2_nand2_1 _22927_ (.Y(_05586_),
    .A(_09958_),
    .B(net101));
 sg13g2_o21ai_1 _22928_ (.B1(_05586_),
    .Y(_01058_),
    .A1(net86),
    .A2(_05585_));
 sg13g2_o21ai_1 _22929_ (.B1(net527),
    .Y(_05587_),
    .A1(_11032_),
    .A2(_11045_));
 sg13g2_nand2_1 _22930_ (.Y(_05588_),
    .A(_09869_),
    .B(net528));
 sg13g2_nand2_1 _22931_ (.Y(_05589_),
    .A(_05587_),
    .B(_05588_));
 sg13g2_mux2_1 _22932_ (.A0(net871),
    .A1(_05589_),
    .S(net85),
    .X(_01059_));
 sg13g2_mux2_1 _22933_ (.A0(_09827_),
    .A1(_05568_),
    .S(net85),
    .X(_01060_));
 sg13g2_nand2_1 _22934_ (.Y(_05590_),
    .A(_05573_),
    .B(net106));
 sg13g2_o21ai_1 _22935_ (.B1(_05590_),
    .Y(_01061_),
    .A1(net720),
    .A2(net84));
 sg13g2_buf_1 _22936_ (.A(net1007),
    .X(_05591_));
 sg13g2_mux2_1 _22937_ (.A0(net819),
    .A1(_10482_),
    .S(net85),
    .X(_01062_));
 sg13g2_buf_1 _22938_ (.A(net1006),
    .X(_05592_));
 sg13g2_mux2_1 _22939_ (.A0(net818),
    .A1(_05578_),
    .S(net85),
    .X(_01063_));
 sg13g2_nand2_1 _22940_ (.Y(_05593_),
    .A(_05582_),
    .B(net106));
 sg13g2_o21ai_1 _22941_ (.B1(_05593_),
    .Y(_01064_),
    .A1(net719),
    .A2(net84));
 sg13g2_nand2_1 _22942_ (.Y(_05594_),
    .A(net1005),
    .B(net101));
 sg13g2_o21ai_1 _22943_ (.B1(_05594_),
    .Y(_01065_),
    .A1(_10397_),
    .A2(net86));
 sg13g2_nor2_1 _22944_ (.A(_11553_),
    .B(_11019_),
    .Y(_05595_));
 sg13g2_a21oi_1 _22945_ (.A1(_10068_),
    .A2(_10102_),
    .Y(_05596_),
    .B1(_05567_));
 sg13g2_nor2_1 _22946_ (.A(_05595_),
    .B(_05596_),
    .Y(_05597_));
 sg13g2_nand2_1 _22947_ (.Y(_05598_),
    .A(_09921_),
    .B(net101));
 sg13g2_o21ai_1 _22948_ (.B1(_05598_),
    .Y(_01066_),
    .A1(net100),
    .A2(_05597_));
 sg13g2_nor2_1 _22949_ (.A(net820),
    .B(_10061_),
    .Y(_05599_));
 sg13g2_a21oi_1 _22950_ (.A1(net820),
    .A2(_05589_),
    .Y(_05600_),
    .B1(_05599_));
 sg13g2_nand2_1 _22951_ (.Y(_05601_),
    .A(_09926_),
    .B(net101));
 sg13g2_o21ai_1 _22952_ (.B1(_05601_),
    .Y(_01067_),
    .A1(net100),
    .A2(_05600_));
 sg13g2_buf_1 _22953_ (.A(net253),
    .X(_05602_));
 sg13g2_nand2_1 _22954_ (.Y(_05603_),
    .A(_08582_),
    .B(_08587_));
 sg13g2_buf_2 _22955_ (.A(_05603_),
    .X(_05604_));
 sg13g2_nand2_1 _22956_ (.Y(_05605_),
    .A(_10316_),
    .B(_05604_));
 sg13g2_o21ai_1 _22957_ (.B1(_05605_),
    .Y(_05606_),
    .A1(_08149_),
    .A2(_05604_));
 sg13g2_or3_1 _22958_ (.A(_11021_),
    .B(_11078_),
    .C(_11112_),
    .X(_05607_));
 sg13g2_o21ai_1 _22959_ (.B1(_03171_),
    .Y(_05608_),
    .A1(_11048_),
    .A2(_05607_));
 sg13g2_nor4_2 _22960_ (.A(_08514_),
    .B(_04574_),
    .C(_09970_),
    .Y(_05609_),
    .D(_03371_));
 sg13g2_and2_1 _22961_ (.A(_05608_),
    .B(_05609_),
    .X(_05610_));
 sg13g2_buf_2 _22962_ (.A(_05610_),
    .X(_05611_));
 sg13g2_buf_1 _22963_ (.A(_00288_),
    .X(_05612_));
 sg13g2_nand2b_1 _22964_ (.Y(_05613_),
    .B(net951),
    .A_N(net1052));
 sg13g2_o21ai_1 _22965_ (.B1(_05613_),
    .Y(_05614_),
    .A1(net831),
    .A2(_10316_));
 sg13g2_nand3_1 _22966_ (.B(_05611_),
    .C(_05614_),
    .A(_08620_),
    .Y(_05615_));
 sg13g2_o21ai_1 _22967_ (.B1(_05615_),
    .Y(_05616_),
    .A1(net186),
    .A2(_05606_));
 sg13g2_nand2b_1 _22968_ (.Y(_05617_),
    .B(net253),
    .A_N(_05611_));
 sg13g2_nand2_2 _22969_ (.Y(_05618_),
    .A(_09037_),
    .B(_05617_));
 sg13g2_inv_1 _22970_ (.Y(_05619_),
    .A(_10317_));
 sg13g2_a22oi_1 _22971_ (.Y(_01070_),
    .B1(_05618_),
    .B2(_05619_),
    .A2(_05616_),
    .A1(_09039_));
 sg13g2_inv_1 _22972_ (.Y(_05620_),
    .A(net1072));
 sg13g2_nand2_1 _22973_ (.Y(_05621_),
    .A(net577),
    .B(_05604_));
 sg13g2_o21ai_1 _22974_ (.B1(_05621_),
    .Y(_05622_),
    .A1(_08084_),
    .A2(_05604_));
 sg13g2_nor2_1 _22975_ (.A(_05619_),
    .B(_05620_),
    .Y(_05623_));
 sg13g2_buf_2 _22976_ (.A(_05623_),
    .X(_05624_));
 sg13g2_buf_1 _22977_ (.A(_10317_),
    .X(_05625_));
 sg13g2_nor2_1 _22978_ (.A(_05625_),
    .B(net1072),
    .Y(_05626_));
 sg13g2_o21ai_1 _22979_ (.B1(net831),
    .Y(_05627_),
    .A1(_05624_),
    .A2(_05626_));
 sg13g2_o21ai_1 _22980_ (.B1(_05627_),
    .Y(_05628_),
    .A1(net831),
    .A2(_10286_));
 sg13g2_nand3_1 _22981_ (.B(_05611_),
    .C(_05628_),
    .A(net186),
    .Y(_05629_));
 sg13g2_o21ai_1 _22982_ (.B1(_05629_),
    .Y(_05630_),
    .A1(net186),
    .A2(_05622_));
 sg13g2_buf_1 _22983_ (.A(_09038_),
    .X(_05631_));
 sg13g2_a22oi_1 _22984_ (.Y(_01071_),
    .B1(_05630_),
    .B2(_05631_),
    .A2(_05618_),
    .A1(_05620_));
 sg13g2_buf_1 _22985_ (.A(_10241_),
    .X(_05632_));
 sg13g2_nand2_1 _22986_ (.Y(_05633_),
    .A(_10262_),
    .B(_05604_));
 sg13g2_o21ai_1 _22987_ (.B1(_05633_),
    .Y(_05634_),
    .A1(_08344_),
    .A2(_05604_));
 sg13g2_nand2_1 _22988_ (.Y(_05635_),
    .A(_10317_),
    .B(net1072));
 sg13g2_buf_1 _22989_ (.A(_05635_),
    .X(_05636_));
 sg13g2_nor2_2 _22990_ (.A(net817),
    .B(net816),
    .Y(_05637_));
 sg13g2_buf_1 _22991_ (.A(_10240_),
    .X(_05638_));
 sg13g2_nor2_1 _22992_ (.A(net940),
    .B(_05624_),
    .Y(_05639_));
 sg13g2_o21ai_1 _22993_ (.B1(net951),
    .Y(_05640_),
    .A1(_05637_),
    .A2(_05639_));
 sg13g2_o21ai_1 _22994_ (.B1(_05640_),
    .Y(_05641_),
    .A1(net831),
    .A2(_10262_));
 sg13g2_nand3_1 _22995_ (.B(_05611_),
    .C(_05641_),
    .A(net186),
    .Y(_05642_));
 sg13g2_o21ai_1 _22996_ (.B1(_05642_),
    .Y(_05643_),
    .A1(net186),
    .A2(_05634_));
 sg13g2_buf_2 _22997_ (.A(net761),
    .X(_05644_));
 sg13g2_a22oi_1 _22998_ (.Y(_01072_),
    .B1(_05643_),
    .B2(net622),
    .A2(_05618_),
    .A1(net817));
 sg13g2_nor2_1 _22999_ (.A(_08069_),
    .B(_05604_),
    .Y(_05645_));
 sg13g2_a21oi_1 _23000_ (.A1(_09220_),
    .A2(_05604_),
    .Y(_05646_),
    .B1(_05645_));
 sg13g2_buf_1 _23001_ (.A(_10220_),
    .X(_05647_));
 sg13g2_xnor2_1 _23002_ (.Y(_05648_),
    .A(net939),
    .B(_05637_));
 sg13g2_nand2_1 _23003_ (.Y(_05649_),
    .A(_03338_),
    .B(_05648_));
 sg13g2_o21ai_1 _23004_ (.B1(_05649_),
    .Y(_05650_),
    .A1(_03338_),
    .A2(_10200_));
 sg13g2_nand3_1 _23005_ (.B(_05611_),
    .C(_05650_),
    .A(_08620_),
    .Y(_05651_));
 sg13g2_o21ai_1 _23006_ (.B1(_05651_),
    .Y(_05652_),
    .A1(net186),
    .A2(_05646_));
 sg13g2_a22oi_1 _23007_ (.Y(_01073_),
    .B1(_05652_),
    .B2(_05644_),
    .A2(_05618_),
    .A1(_10892_));
 sg13g2_buf_1 _23008_ (.A(net573),
    .X(_05653_));
 sg13g2_buf_2 _23009_ (.A(_00188_),
    .X(_05654_));
 sg13g2_nor2_1 _23010_ (.A(_10576_),
    .B(_10220_),
    .Y(_05655_));
 sg13g2_buf_2 _23011_ (.A(_05655_),
    .X(_05656_));
 sg13g2_nand2_1 _23012_ (.Y(_05657_),
    .A(_05654_),
    .B(_05656_));
 sg13g2_nand4_1 _23013_ (.B(_11095_),
    .C(_05609_),
    .A(net951),
    .Y(_05658_),
    .D(_05626_));
 sg13g2_buf_1 _23014_ (.A(_05658_),
    .X(_05659_));
 sg13g2_nor2_1 _23015_ (.A(_05657_),
    .B(_05659_),
    .Y(_05660_));
 sg13g2_buf_1 _23016_ (.A(_05660_),
    .X(_05661_));
 sg13g2_buf_1 _23017_ (.A(_05661_),
    .X(_05662_));
 sg13g2_mux2_1 _23018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(net491),
    .S(net351),
    .X(_01141_));
 sg13g2_mux2_1 _23019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net438),
    .S(net351),
    .X(_01142_));
 sg13g2_buf_1 _23020_ (.A(net994),
    .X(_05663_));
 sg13g2_mux2_1 _23021_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(net815),
    .S(net351),
    .X(_01143_));
 sg13g2_mux2_1 _23022_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net501),
    .S(net351),
    .X(_01144_));
 sg13g2_mux2_1 _23023_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net827),
    .S(net351),
    .X(_01145_));
 sg13g2_mux2_1 _23024_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net825),
    .S(net351),
    .X(_01146_));
 sg13g2_mux2_1 _23025_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net824),
    .S(_05662_),
    .X(_01147_));
 sg13g2_mux2_1 _23026_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(_03369_),
    .S(net351),
    .X(_01148_));
 sg13g2_buf_1 _23027_ (.A(net953),
    .X(_05664_));
 sg13g2_mux2_1 _23028_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net814),
    .S(net351),
    .X(_01149_));
 sg13g2_mux2_1 _23029_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net826),
    .S(_05662_),
    .X(_01150_));
 sg13g2_mux2_1 _23030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(net497),
    .S(_05661_),
    .X(_01151_));
 sg13g2_mux2_1 _23031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net498),
    .S(_05661_),
    .X(_01152_));
 sg13g2_nand3_1 _23032_ (.B(_11095_),
    .C(_05609_),
    .A(_03337_),
    .Y(_05665_));
 sg13g2_buf_1 _23033_ (.A(_05665_),
    .X(_05666_));
 sg13g2_buf_1 _23034_ (.A(_05666_),
    .X(_05667_));
 sg13g2_nand2_1 _23035_ (.Y(_05668_),
    .A(_05619_),
    .B(_10302_));
 sg13g2_buf_1 _23036_ (.A(_05668_),
    .X(_05669_));
 sg13g2_inv_1 _23037_ (.Y(_05670_),
    .A(_10576_));
 sg13g2_nand2_1 _23038_ (.Y(_05671_),
    .A(_05670_),
    .B(_05647_));
 sg13g2_buf_1 _23039_ (.A(_05671_),
    .X(_05672_));
 sg13g2_nor3_2 _23040_ (.A(_05638_),
    .B(_05669_),
    .C(_05672_),
    .Y(_05673_));
 sg13g2_nor2b_1 _23041_ (.A(net425),
    .B_N(_05673_),
    .Y(_05674_));
 sg13g2_buf_1 _23042_ (.A(_05674_),
    .X(_05675_));
 sg13g2_buf_1 _23043_ (.A(_05675_),
    .X(_05676_));
 sg13g2_mux2_1 _23044_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net491),
    .S(net330),
    .X(_01153_));
 sg13g2_mux2_1 _23045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net438),
    .S(net330),
    .X(_01154_));
 sg13g2_mux2_1 _23046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net815),
    .S(net330),
    .X(_01155_));
 sg13g2_mux2_1 _23047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net501),
    .S(_05676_),
    .X(_01156_));
 sg13g2_mux2_1 _23048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net827),
    .S(net330),
    .X(_01157_));
 sg13g2_mux2_1 _23049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net825),
    .S(net330),
    .X(_01158_));
 sg13g2_mux2_1 _23050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net824),
    .S(net330),
    .X(_01159_));
 sg13g2_mux2_1 _23051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(_03369_),
    .S(net330),
    .X(_01160_));
 sg13g2_mux2_1 _23052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net814),
    .S(net330),
    .X(_01161_));
 sg13g2_mux2_1 _23053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net826),
    .S(_05676_),
    .X(_01162_));
 sg13g2_mux2_1 _23054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net497),
    .S(_05675_),
    .X(_01163_));
 sg13g2_mux2_1 _23055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net498),
    .S(_05675_),
    .X(_01164_));
 sg13g2_nor3_1 _23056_ (.A(net1073),
    .B(net816),
    .C(_05672_),
    .Y(_05677_));
 sg13g2_buf_2 _23057_ (.A(_05677_),
    .X(_05678_));
 sg13g2_nor2b_1 _23058_ (.A(net425),
    .B_N(_05678_),
    .Y(_05679_));
 sg13g2_buf_1 _23059_ (.A(_05679_),
    .X(_05680_));
 sg13g2_buf_1 _23060_ (.A(_05680_),
    .X(_05681_));
 sg13g2_mux2_1 _23061_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net491),
    .S(net329),
    .X(_01165_));
 sg13g2_mux2_1 _23062_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net438),
    .S(net329),
    .X(_01166_));
 sg13g2_mux2_1 _23063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net815),
    .S(net329),
    .X(_01167_));
 sg13g2_mux2_1 _23064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(_03378_),
    .S(_05681_),
    .X(_01168_));
 sg13g2_mux2_1 _23065_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(_03379_),
    .S(net329),
    .X(_01169_));
 sg13g2_mux2_1 _23066_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net825),
    .S(net329),
    .X(_01170_));
 sg13g2_mux2_1 _23067_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net824),
    .S(net329),
    .X(_01171_));
 sg13g2_buf_1 _23068_ (.A(net954),
    .X(_05682_));
 sg13g2_mux2_1 _23069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(net813),
    .S(net329),
    .X(_01172_));
 sg13g2_mux2_1 _23070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net814),
    .S(net329),
    .X(_01173_));
 sg13g2_mux2_1 _23071_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net826),
    .S(_05681_),
    .X(_01174_));
 sg13g2_mux2_1 _23072_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net497),
    .S(_05680_),
    .X(_01175_));
 sg13g2_mux2_1 _23073_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net498),
    .S(_05680_),
    .X(_01176_));
 sg13g2_nor2_2 _23074_ (.A(_10576_),
    .B(_10892_),
    .Y(_05683_));
 sg13g2_nand2b_1 _23075_ (.Y(_05684_),
    .B(_05683_),
    .A_N(_05654_));
 sg13g2_buf_1 _23076_ (.A(_05684_),
    .X(_05685_));
 sg13g2_nor2_1 _23077_ (.A(_05659_),
    .B(_05685_),
    .Y(_05686_));
 sg13g2_buf_1 _23078_ (.A(_05686_),
    .X(_05687_));
 sg13g2_buf_1 _23079_ (.A(_05687_),
    .X(_05688_));
 sg13g2_mux2_1 _23080_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net491),
    .S(net350),
    .X(_01177_));
 sg13g2_mux2_1 _23081_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net438),
    .S(net350),
    .X(_01178_));
 sg13g2_mux2_1 _23082_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net815),
    .S(net350),
    .X(_01179_));
 sg13g2_mux2_1 _23083_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(_03378_),
    .S(net350),
    .X(_01180_));
 sg13g2_mux2_1 _23084_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(_03379_),
    .S(net350),
    .X(_01181_));
 sg13g2_mux2_1 _23085_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net825),
    .S(net350),
    .X(_01182_));
 sg13g2_mux2_1 _23086_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net824),
    .S(_05688_),
    .X(_01183_));
 sg13g2_mux2_1 _23087_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(net813),
    .S(net350),
    .X(_01184_));
 sg13g2_mux2_1 _23088_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net814),
    .S(net350),
    .X(_01185_));
 sg13g2_mux2_1 _23089_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net826),
    .S(_05688_),
    .X(_01186_));
 sg13g2_mux2_1 _23090_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net497),
    .S(_05687_),
    .X(_01187_));
 sg13g2_mux2_1 _23091_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net498),
    .S(_05687_),
    .X(_01188_));
 sg13g2_nand2_2 _23092_ (.Y(_05689_),
    .A(net941),
    .B(_05620_));
 sg13g2_or2_1 _23093_ (.X(_05690_),
    .B(_05666_),
    .A(_05689_));
 sg13g2_buf_2 _23094_ (.A(_05690_),
    .X(_05691_));
 sg13g2_nor2_1 _23095_ (.A(_05685_),
    .B(_05691_),
    .Y(_05692_));
 sg13g2_buf_1 _23096_ (.A(_05692_),
    .X(_05693_));
 sg13g2_buf_1 _23097_ (.A(_05693_),
    .X(_05694_));
 sg13g2_mux2_1 _23098_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net491),
    .S(net280),
    .X(_01189_));
 sg13g2_mux2_1 _23099_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net438),
    .S(net280),
    .X(_01190_));
 sg13g2_mux2_1 _23100_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net815),
    .S(net280),
    .X(_01191_));
 sg13g2_buf_1 _23101_ (.A(_02877_),
    .X(_05695_));
 sg13g2_mux2_1 _23102_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(net552),
    .S(net280),
    .X(_01192_));
 sg13g2_buf_1 _23103_ (.A(_08949_),
    .X(_05696_));
 sg13g2_mux2_1 _23104_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net812),
    .S(net280),
    .X(_01193_));
 sg13g2_mux2_1 _23105_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net825),
    .S(_05694_),
    .X(_01194_));
 sg13g2_mux2_1 _23106_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net824),
    .S(net280),
    .X(_01195_));
 sg13g2_mux2_1 _23107_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net813),
    .S(net280),
    .X(_01196_));
 sg13g2_mux2_1 _23108_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net814),
    .S(net280),
    .X(_01197_));
 sg13g2_mux2_1 _23109_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net826),
    .S(_05694_),
    .X(_01198_));
 sg13g2_mux2_1 _23110_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net497),
    .S(_05693_),
    .X(_01199_));
 sg13g2_mux2_1 _23111_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net498),
    .S(_05693_),
    .X(_01200_));
 sg13g2_buf_1 _23112_ (.A(_05666_),
    .X(_05697_));
 sg13g2_nor3_1 _23113_ (.A(net706),
    .B(_05697_),
    .C(_05685_),
    .Y(_05698_));
 sg13g2_buf_1 _23114_ (.A(_05698_),
    .X(_05699_));
 sg13g2_buf_1 _23115_ (.A(_05699_),
    .X(_05700_));
 sg13g2_mux2_1 _23116_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(net491),
    .S(net328),
    .X(_01201_));
 sg13g2_mux2_1 _23117_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(_03390_),
    .S(net328),
    .X(_01202_));
 sg13g2_mux2_1 _23118_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net815),
    .S(net328),
    .X(_01203_));
 sg13g2_mux2_1 _23119_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(net552),
    .S(net328),
    .X(_01204_));
 sg13g2_mux2_1 _23120_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(net812),
    .S(net328),
    .X(_01205_));
 sg13g2_mux2_1 _23121_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net825),
    .S(_05700_),
    .X(_01206_));
 sg13g2_mux2_1 _23122_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net824),
    .S(net328),
    .X(_01207_));
 sg13g2_mux2_1 _23123_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net813),
    .S(net328),
    .X(_01208_));
 sg13g2_mux2_1 _23124_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(_05664_),
    .S(net328),
    .X(_01209_));
 sg13g2_mux2_1 _23125_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net826),
    .S(_05700_),
    .X(_01210_));
 sg13g2_mux2_1 _23126_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(net497),
    .S(_05699_),
    .X(_01211_));
 sg13g2_mux2_1 _23127_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03389_),
    .S(_05699_),
    .X(_01212_));
 sg13g2_nor3_1 _23128_ (.A(net816),
    .B(net424),
    .C(_05685_),
    .Y(_05701_));
 sg13g2_buf_1 _23129_ (.A(_05701_),
    .X(_05702_));
 sg13g2_buf_1 _23130_ (.A(_05702_),
    .X(_05703_));
 sg13g2_mux2_1 _23131_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(net491),
    .S(net327),
    .X(_01213_));
 sg13g2_mux2_1 _23132_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(_03390_),
    .S(net327),
    .X(_01214_));
 sg13g2_mux2_1 _23133_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(_05663_),
    .S(net327),
    .X(_01215_));
 sg13g2_mux2_1 _23134_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(net552),
    .S(net327),
    .X(_01216_));
 sg13g2_mux2_1 _23135_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(net812),
    .S(net327),
    .X(_01217_));
 sg13g2_mux2_1 _23136_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(net825),
    .S(_05703_),
    .X(_01218_));
 sg13g2_mux2_1 _23137_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(net824),
    .S(_05703_),
    .X(_01219_));
 sg13g2_mux2_1 _23138_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(net813),
    .S(net327),
    .X(_01220_));
 sg13g2_mux2_1 _23139_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(_05664_),
    .S(net327),
    .X(_01221_));
 sg13g2_mux2_1 _23140_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(_04578_),
    .S(net327),
    .X(_01222_));
 sg13g2_mux2_1 _23141_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_03598_),
    .S(_05702_),
    .X(_01223_));
 sg13g2_mux2_1 _23142_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03389_),
    .S(_05702_),
    .X(_01224_));
 sg13g2_buf_1 _23143_ (.A(_10576_),
    .X(_05704_));
 sg13g2_nand2_1 _23144_ (.Y(_05705_),
    .A(_05704_),
    .B(_10892_));
 sg13g2_buf_1 _23145_ (.A(_05705_),
    .X(_05706_));
 sg13g2_nand2_1 _23146_ (.Y(_05707_),
    .A(_05632_),
    .B(_05626_));
 sg13g2_nor3_1 _23147_ (.A(net424),
    .B(_05706_),
    .C(_05707_),
    .Y(_05708_));
 sg13g2_buf_1 _23148_ (.A(_05708_),
    .X(_05709_));
 sg13g2_buf_1 _23149_ (.A(_05709_),
    .X(_05710_));
 sg13g2_mux2_1 _23150_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net491),
    .S(net326),
    .X(_01225_));
 sg13g2_buf_1 _23151_ (.A(net578),
    .X(_05711_));
 sg13g2_mux2_1 _23152_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net490),
    .S(net326),
    .X(_01226_));
 sg13g2_mux2_1 _23153_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net815),
    .S(net326),
    .X(_01227_));
 sg13g2_mux2_1 _23154_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net552),
    .S(net326),
    .X(_01228_));
 sg13g2_mux2_1 _23155_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net812),
    .S(net326),
    .X(_01229_));
 sg13g2_mux2_1 _23156_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net825),
    .S(_05710_),
    .X(_01230_));
 sg13g2_mux2_1 _23157_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net824),
    .S(net326),
    .X(_01231_));
 sg13g2_mux2_1 _23158_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net813),
    .S(net326),
    .X(_01232_));
 sg13g2_mux2_1 _23159_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net814),
    .S(net326),
    .X(_01233_));
 sg13g2_mux2_1 _23160_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net826),
    .S(_05710_),
    .X(_01234_));
 sg13g2_mux2_1 _23161_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(_03598_),
    .S(_05709_),
    .X(_01235_));
 sg13g2_buf_1 _23162_ (.A(net577),
    .X(_05712_));
 sg13g2_mux2_1 _23163_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net489),
    .S(_05709_),
    .X(_01236_));
 sg13g2_nor3_1 _23164_ (.A(net940),
    .B(_05691_),
    .C(_05706_),
    .Y(_05713_));
 sg13g2_buf_1 _23165_ (.A(_05713_),
    .X(_05714_));
 sg13g2_buf_1 _23166_ (.A(_05714_),
    .X(_05715_));
 sg13g2_mux2_1 _23167_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(_05653_),
    .S(net279),
    .X(_01237_));
 sg13g2_mux2_1 _23168_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net490),
    .S(net279),
    .X(_01238_));
 sg13g2_mux2_1 _23169_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(_05663_),
    .S(net279),
    .X(_01239_));
 sg13g2_mux2_1 _23170_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net552),
    .S(net279),
    .X(_01240_));
 sg13g2_mux2_1 _23171_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net812),
    .S(net279),
    .X(_01241_));
 sg13g2_mux2_1 _23172_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(_04579_),
    .S(_05715_),
    .X(_01242_));
 sg13g2_mux2_1 _23173_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(_04580_),
    .S(net279),
    .X(_01243_));
 sg13g2_mux2_1 _23174_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net813),
    .S(net279),
    .X(_01244_));
 sg13g2_mux2_1 _23175_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net814),
    .S(net279),
    .X(_01245_));
 sg13g2_mux2_1 _23176_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net826),
    .S(_05715_),
    .X(_01246_));
 sg13g2_buf_1 _23177_ (.A(net576),
    .X(_05716_));
 sg13g2_mux2_1 _23178_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net488),
    .S(_05714_),
    .X(_01247_));
 sg13g2_mux2_1 _23179_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net489),
    .S(_05714_),
    .X(_01248_));
 sg13g2_nor2_1 _23180_ (.A(_05670_),
    .B(_05625_),
    .Y(_05717_));
 sg13g2_nand3_1 _23181_ (.B(net817),
    .C(_05717_),
    .A(net1072),
    .Y(_05718_));
 sg13g2_nor2_2 _23182_ (.A(net939),
    .B(_05718_),
    .Y(_05719_));
 sg13g2_nor2b_1 _23183_ (.A(net425),
    .B_N(_05719_),
    .Y(_05720_));
 sg13g2_buf_1 _23184_ (.A(_05720_),
    .X(_05721_));
 sg13g2_buf_1 _23185_ (.A(_05721_),
    .X(_05722_));
 sg13g2_mux2_1 _23186_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(_05653_),
    .S(net325),
    .X(_01249_));
 sg13g2_mux2_1 _23187_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net490),
    .S(net325),
    .X(_01250_));
 sg13g2_mux2_1 _23188_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net815),
    .S(net325),
    .X(_01251_));
 sg13g2_mux2_1 _23189_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net552),
    .S(net325),
    .X(_01252_));
 sg13g2_mux2_1 _23190_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net812),
    .S(net325),
    .X(_01253_));
 sg13g2_buf_1 _23191_ (.A(_02866_),
    .X(_05723_));
 sg13g2_mux2_1 _23192_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net811),
    .S(_05722_),
    .X(_01254_));
 sg13g2_buf_1 _23193_ (.A(_08951_),
    .X(_05724_));
 sg13g2_mux2_1 _23194_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net937),
    .S(net325),
    .X(_01255_));
 sg13g2_mux2_1 _23195_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(_05682_),
    .S(net325),
    .X(_01256_));
 sg13g2_mux2_1 _23196_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net814),
    .S(net325),
    .X(_01257_));
 sg13g2_buf_1 _23197_ (.A(_10147_),
    .X(_05725_));
 sg13g2_mux2_1 _23198_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(_05725_),
    .S(_05722_),
    .X(_01258_));
 sg13g2_mux2_1 _23199_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net488),
    .S(_05721_),
    .X(_01259_));
 sg13g2_mux2_1 _23200_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net489),
    .S(_05721_),
    .X(_01260_));
 sg13g2_buf_1 _23201_ (.A(net573),
    .X(_05726_));
 sg13g2_nor3_1 _23202_ (.A(net1073),
    .B(net816),
    .C(_05706_),
    .Y(_05727_));
 sg13g2_buf_2 _23203_ (.A(_05727_),
    .X(_05728_));
 sg13g2_nor2b_1 _23204_ (.A(net425),
    .B_N(_05728_),
    .Y(_05729_));
 sg13g2_buf_1 _23205_ (.A(_05729_),
    .X(_05730_));
 sg13g2_buf_1 _23206_ (.A(_05730_),
    .X(_05731_));
 sg13g2_mux2_1 _23207_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(_05726_),
    .S(net324),
    .X(_01261_));
 sg13g2_mux2_1 _23208_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(net490),
    .S(net324),
    .X(_01262_));
 sg13g2_buf_1 _23209_ (.A(net994),
    .X(_05732_));
 sg13g2_mux2_1 _23210_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net810),
    .S(net324),
    .X(_01263_));
 sg13g2_mux2_1 _23211_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net552),
    .S(net324),
    .X(_01264_));
 sg13g2_mux2_1 _23212_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(_05696_),
    .S(net324),
    .X(_01265_));
 sg13g2_mux2_1 _23213_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(net811),
    .S(net324),
    .X(_01266_));
 sg13g2_mux2_1 _23214_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(_05724_),
    .S(_05731_),
    .X(_01267_));
 sg13g2_mux2_1 _23215_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(_05682_),
    .S(net324),
    .X(_01268_));
 sg13g2_buf_1 _23216_ (.A(net1075),
    .X(_05733_));
 sg13g2_mux2_1 _23217_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net935),
    .S(net324),
    .X(_01269_));
 sg13g2_mux2_1 _23218_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(_05725_),
    .S(_05731_),
    .X(_01270_));
 sg13g2_mux2_1 _23219_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net488),
    .S(_05730_),
    .X(_01271_));
 sg13g2_mux2_1 _23220_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net489),
    .S(_05730_),
    .X(_01272_));
 sg13g2_nor2_1 _23221_ (.A(_05657_),
    .B(_05691_),
    .Y(_05734_));
 sg13g2_buf_1 _23222_ (.A(_05734_),
    .X(_05735_));
 sg13g2_buf_1 _23223_ (.A(_05735_),
    .X(_05736_));
 sg13g2_mux2_1 _23224_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(_05726_),
    .S(net278),
    .X(_01273_));
 sg13g2_mux2_1 _23225_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(net490),
    .S(net278),
    .X(_01274_));
 sg13g2_mux2_1 _23226_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(net810),
    .S(net278),
    .X(_01275_));
 sg13g2_mux2_1 _23227_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(net552),
    .S(net278),
    .X(_01276_));
 sg13g2_mux2_1 _23228_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(_05696_),
    .S(net278),
    .X(_01277_));
 sg13g2_mux2_1 _23229_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(net811),
    .S(net278),
    .X(_01278_));
 sg13g2_mux2_1 _23230_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(net937),
    .S(_05736_),
    .X(_01279_));
 sg13g2_mux2_1 _23231_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(net813),
    .S(net278),
    .X(_01280_));
 sg13g2_mux2_1 _23232_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(net935),
    .S(net278),
    .X(_01281_));
 sg13g2_mux2_1 _23233_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(net936),
    .S(_05736_),
    .X(_01282_));
 sg13g2_mux2_1 _23234_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net488),
    .S(_05735_),
    .X(_01283_));
 sg13g2_mux2_1 _23235_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05712_),
    .S(_05735_),
    .X(_01284_));
 sg13g2_or2_1 _23236_ (.X(_05737_),
    .B(_05706_),
    .A(_05654_));
 sg13g2_buf_1 _23237_ (.A(_05737_),
    .X(_05738_));
 sg13g2_nor2_1 _23238_ (.A(_05659_),
    .B(_05738_),
    .Y(_05739_));
 sg13g2_buf_1 _23239_ (.A(_05739_),
    .X(_05740_));
 sg13g2_buf_1 _23240_ (.A(_05740_),
    .X(_05741_));
 sg13g2_mux2_1 _23241_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net487),
    .S(net349),
    .X(_01285_));
 sg13g2_mux2_1 _23242_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net490),
    .S(net349),
    .X(_01286_));
 sg13g2_mux2_1 _23243_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net810),
    .S(net349),
    .X(_01287_));
 sg13g2_mux2_1 _23244_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(_05695_),
    .S(net349),
    .X(_01288_));
 sg13g2_mux2_1 _23245_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net812),
    .S(net349),
    .X(_01289_));
 sg13g2_mux2_1 _23246_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net811),
    .S(_05741_),
    .X(_01290_));
 sg13g2_mux2_1 _23247_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net937),
    .S(net349),
    .X(_01291_));
 sg13g2_buf_1 _23248_ (.A(_09985_),
    .X(_05742_));
 sg13g2_mux2_1 _23249_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(_05742_),
    .S(net349),
    .X(_01292_));
 sg13g2_mux2_1 _23250_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net935),
    .S(net349),
    .X(_01293_));
 sg13g2_mux2_1 _23251_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net936),
    .S(_05741_),
    .X(_01294_));
 sg13g2_mux2_1 _23252_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net488),
    .S(_05740_),
    .X(_01295_));
 sg13g2_mux2_1 _23253_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net489),
    .S(_05740_),
    .X(_01296_));
 sg13g2_nor2_1 _23254_ (.A(_05691_),
    .B(_05738_),
    .Y(_05743_));
 sg13g2_buf_1 _23255_ (.A(_05743_),
    .X(_05744_));
 sg13g2_buf_1 _23256_ (.A(_05744_),
    .X(_05745_));
 sg13g2_mux2_1 _23257_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net487),
    .S(net277),
    .X(_01297_));
 sg13g2_mux2_1 _23258_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net490),
    .S(net277),
    .X(_01298_));
 sg13g2_mux2_1 _23259_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(_05732_),
    .S(net277),
    .X(_01299_));
 sg13g2_mux2_1 _23260_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(_05695_),
    .S(net277),
    .X(_01300_));
 sg13g2_mux2_1 _23261_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net812),
    .S(net277),
    .X(_01301_));
 sg13g2_mux2_1 _23262_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net811),
    .S(_05745_),
    .X(_01302_));
 sg13g2_mux2_1 _23263_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(_05724_),
    .S(net277),
    .X(_01303_));
 sg13g2_mux2_1 _23264_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net934),
    .S(net277),
    .X(_01304_));
 sg13g2_mux2_1 _23265_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net935),
    .S(net277),
    .X(_01305_));
 sg13g2_mux2_1 _23266_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net936),
    .S(_05745_),
    .X(_01306_));
 sg13g2_mux2_1 _23267_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net488),
    .S(_05744_),
    .X(_01307_));
 sg13g2_mux2_1 _23268_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net489),
    .S(_05744_),
    .X(_01308_));
 sg13g2_nor3_1 _23269_ (.A(net706),
    .B(net424),
    .C(_05738_),
    .Y(_05746_));
 sg13g2_buf_1 _23270_ (.A(_05746_),
    .X(_05747_));
 sg13g2_buf_1 _23271_ (.A(_05747_),
    .X(_05748_));
 sg13g2_mux2_1 _23272_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net487),
    .S(net323),
    .X(_01309_));
 sg13g2_mux2_1 _23273_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(_05711_),
    .S(net323),
    .X(_01310_));
 sg13g2_mux2_1 _23274_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net810),
    .S(net323),
    .X(_01311_));
 sg13g2_buf_1 _23275_ (.A(_02877_),
    .X(_05749_));
 sg13g2_mux2_1 _23276_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net551),
    .S(net323),
    .X(_01312_));
 sg13g2_buf_1 _23277_ (.A(_08949_),
    .X(_05750_));
 sg13g2_mux2_1 _23278_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net809),
    .S(net323),
    .X(_01313_));
 sg13g2_mux2_1 _23279_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(_05723_),
    .S(_05748_),
    .X(_01314_));
 sg13g2_mux2_1 _23280_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net937),
    .S(net323),
    .X(_01315_));
 sg13g2_mux2_1 _23281_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net934),
    .S(net323),
    .X(_01316_));
 sg13g2_mux2_1 _23282_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net935),
    .S(net323),
    .X(_01317_));
 sg13g2_mux2_1 _23283_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net936),
    .S(_05748_),
    .X(_01318_));
 sg13g2_mux2_1 _23284_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net488),
    .S(_05747_),
    .X(_01319_));
 sg13g2_mux2_1 _23285_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net489),
    .S(_05747_),
    .X(_01320_));
 sg13g2_nor3_1 _23286_ (.A(net816),
    .B(net424),
    .C(_05738_),
    .Y(_05751_));
 sg13g2_buf_1 _23287_ (.A(_05751_),
    .X(_05752_));
 sg13g2_buf_1 _23288_ (.A(_05752_),
    .X(_05753_));
 sg13g2_mux2_1 _23289_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net487),
    .S(net322),
    .X(_01321_));
 sg13g2_mux2_1 _23290_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(_05711_),
    .S(net322),
    .X(_01322_));
 sg13g2_mux2_1 _23291_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net810),
    .S(net322),
    .X(_01323_));
 sg13g2_mux2_1 _23292_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net551),
    .S(net322),
    .X(_01324_));
 sg13g2_mux2_1 _23293_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net809),
    .S(net322),
    .X(_01325_));
 sg13g2_mux2_1 _23294_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(_05723_),
    .S(_05753_),
    .X(_01326_));
 sg13g2_mux2_1 _23295_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net937),
    .S(net322),
    .X(_01327_));
 sg13g2_mux2_1 _23296_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net934),
    .S(net322),
    .X(_01328_));
 sg13g2_mux2_1 _23297_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net935),
    .S(net322),
    .X(_01329_));
 sg13g2_mux2_1 _23298_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net936),
    .S(_05753_),
    .X(_01330_));
 sg13g2_mux2_1 _23299_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net488),
    .S(_05752_),
    .X(_01331_));
 sg13g2_mux2_1 _23300_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(_05712_),
    .S(_05752_),
    .X(_01332_));
 sg13g2_nand2_2 _23301_ (.Y(_05754_),
    .A(net938),
    .B(net939));
 sg13g2_nor3_1 _23302_ (.A(net424),
    .B(_05707_),
    .C(_05754_),
    .Y(_05755_));
 sg13g2_buf_1 _23303_ (.A(_05755_),
    .X(_05756_));
 sg13g2_buf_1 _23304_ (.A(_05756_),
    .X(_05757_));
 sg13g2_mux2_1 _23305_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net487),
    .S(net321),
    .X(_01333_));
 sg13g2_mux2_1 _23306_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net490),
    .S(net321),
    .X(_01334_));
 sg13g2_mux2_1 _23307_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net810),
    .S(net321),
    .X(_01335_));
 sg13g2_mux2_1 _23308_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net551),
    .S(net321),
    .X(_01336_));
 sg13g2_mux2_1 _23309_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net809),
    .S(net321),
    .X(_01337_));
 sg13g2_mux2_1 _23310_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net811),
    .S(net321),
    .X(_01338_));
 sg13g2_mux2_1 _23311_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net937),
    .S(_05757_),
    .X(_01339_));
 sg13g2_mux2_1 _23312_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net934),
    .S(net321),
    .X(_01340_));
 sg13g2_mux2_1 _23313_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net935),
    .S(net321),
    .X(_01341_));
 sg13g2_mux2_1 _23314_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net936),
    .S(_05757_),
    .X(_01342_));
 sg13g2_mux2_1 _23315_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(_05716_),
    .S(_05756_),
    .X(_01343_));
 sg13g2_mux2_1 _23316_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net489),
    .S(_05756_),
    .X(_01344_));
 sg13g2_nor3_1 _23317_ (.A(_05638_),
    .B(_05691_),
    .C(_05754_),
    .Y(_05758_));
 sg13g2_buf_1 _23318_ (.A(_05758_),
    .X(_05759_));
 sg13g2_buf_1 _23319_ (.A(_05759_),
    .X(_05760_));
 sg13g2_mux2_1 _23320_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net487),
    .S(net276),
    .X(_01345_));
 sg13g2_buf_1 _23321_ (.A(net578),
    .X(_05761_));
 sg13g2_mux2_1 _23322_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(_05761_),
    .S(net276),
    .X(_01346_));
 sg13g2_mux2_1 _23323_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net810),
    .S(net276),
    .X(_01347_));
 sg13g2_mux2_1 _23324_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net551),
    .S(net276),
    .X(_01348_));
 sg13g2_mux2_1 _23325_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net809),
    .S(net276),
    .X(_01349_));
 sg13g2_mux2_1 _23326_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net811),
    .S(net276),
    .X(_01350_));
 sg13g2_mux2_1 _23327_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net937),
    .S(_05760_),
    .X(_01351_));
 sg13g2_mux2_1 _23328_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net934),
    .S(net276),
    .X(_01352_));
 sg13g2_mux2_1 _23329_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net935),
    .S(net276),
    .X(_01353_));
 sg13g2_mux2_1 _23330_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net936),
    .S(_05760_),
    .X(_01354_));
 sg13g2_mux2_1 _23331_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(_05716_),
    .S(_05759_),
    .X(_01355_));
 sg13g2_buf_1 _23332_ (.A(net577),
    .X(_05762_));
 sg13g2_mux2_1 _23333_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net485),
    .S(_05759_),
    .X(_01356_));
 sg13g2_nor2_2 _23334_ (.A(_10892_),
    .B(_05718_),
    .Y(_05763_));
 sg13g2_nor2b_1 _23335_ (.A(net425),
    .B_N(_05763_),
    .Y(_05764_));
 sg13g2_buf_1 _23336_ (.A(_05764_),
    .X(_05765_));
 sg13g2_buf_1 _23337_ (.A(_05765_),
    .X(_05766_));
 sg13g2_mux2_1 _23338_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net487),
    .S(net320),
    .X(_01357_));
 sg13g2_mux2_1 _23339_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(_05761_),
    .S(net320),
    .X(_01358_));
 sg13g2_mux2_1 _23340_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net810),
    .S(net320),
    .X(_01359_));
 sg13g2_mux2_1 _23341_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net551),
    .S(net320),
    .X(_01360_));
 sg13g2_mux2_1 _23342_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(_05750_),
    .S(net320),
    .X(_01361_));
 sg13g2_mux2_1 _23343_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net811),
    .S(net320),
    .X(_01362_));
 sg13g2_mux2_1 _23344_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net937),
    .S(_05766_),
    .X(_01363_));
 sg13g2_mux2_1 _23345_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(_05742_),
    .S(net320),
    .X(_01364_));
 sg13g2_mux2_1 _23346_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(_05733_),
    .S(net320),
    .X(_01365_));
 sg13g2_mux2_1 _23347_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net936),
    .S(_05766_),
    .X(_01366_));
 sg13g2_buf_1 _23348_ (.A(net576),
    .X(_05767_));
 sg13g2_mux2_1 _23349_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net484),
    .S(_05765_),
    .X(_01367_));
 sg13g2_mux2_1 _23350_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net485),
    .S(_05765_),
    .X(_01368_));
 sg13g2_nor3_1 _23351_ (.A(net1073),
    .B(net816),
    .C(_05754_),
    .Y(_05768_));
 sg13g2_buf_2 _23352_ (.A(_05768_),
    .X(_05769_));
 sg13g2_nor2b_1 _23353_ (.A(net425),
    .B_N(_05769_),
    .Y(_05770_));
 sg13g2_buf_1 _23354_ (.A(_05770_),
    .X(_05771_));
 sg13g2_buf_1 _23355_ (.A(_05771_),
    .X(_05772_));
 sg13g2_mux2_1 _23356_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net487),
    .S(net319),
    .X(_01369_));
 sg13g2_mux2_1 _23357_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net486),
    .S(net319),
    .X(_01370_));
 sg13g2_mux2_1 _23358_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(_05732_),
    .S(net319),
    .X(_01371_));
 sg13g2_mux2_1 _23359_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net551),
    .S(net319),
    .X(_01372_));
 sg13g2_mux2_1 _23360_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(_05750_),
    .S(net319),
    .X(_01373_));
 sg13g2_buf_1 _23361_ (.A(_02866_),
    .X(_05773_));
 sg13g2_mux2_1 _23362_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net808),
    .S(net319),
    .X(_01374_));
 sg13g2_buf_1 _23363_ (.A(_08951_),
    .X(_05774_));
 sg13g2_mux2_1 _23364_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net933),
    .S(_05772_),
    .X(_01375_));
 sg13g2_mux2_1 _23365_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net934),
    .S(net319),
    .X(_01376_));
 sg13g2_mux2_1 _23366_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(_05733_),
    .S(net319),
    .X(_01377_));
 sg13g2_buf_1 _23367_ (.A(_10147_),
    .X(_05775_));
 sg13g2_mux2_1 _23368_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(_05775_),
    .S(_05772_),
    .X(_01378_));
 sg13g2_mux2_1 _23369_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net484),
    .S(_05771_),
    .X(_01379_));
 sg13g2_mux2_1 _23370_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net485),
    .S(_05771_),
    .X(_01380_));
 sg13g2_buf_1 _23371_ (.A(net573),
    .X(_05776_));
 sg13g2_or2_1 _23372_ (.X(_05777_),
    .B(_05754_),
    .A(_05654_));
 sg13g2_buf_1 _23373_ (.A(_05777_),
    .X(_05778_));
 sg13g2_nor2_1 _23374_ (.A(_05659_),
    .B(_05778_),
    .Y(_05779_));
 sg13g2_buf_1 _23375_ (.A(_05779_),
    .X(_05780_));
 sg13g2_buf_1 _23376_ (.A(_05780_),
    .X(_05781_));
 sg13g2_mux2_1 _23377_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net483),
    .S(net348),
    .X(_01381_));
 sg13g2_mux2_1 _23378_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net486),
    .S(net348),
    .X(_01382_));
 sg13g2_buf_1 _23379_ (.A(net994),
    .X(_05782_));
 sg13g2_mux2_1 _23380_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net807),
    .S(net348),
    .X(_01383_));
 sg13g2_mux2_1 _23381_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net551),
    .S(net348),
    .X(_01384_));
 sg13g2_mux2_1 _23382_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net809),
    .S(net348),
    .X(_01385_));
 sg13g2_mux2_1 _23383_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net808),
    .S(_05781_),
    .X(_01386_));
 sg13g2_mux2_1 _23384_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net933),
    .S(net348),
    .X(_01387_));
 sg13g2_mux2_1 _23385_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net934),
    .S(net348),
    .X(_01388_));
 sg13g2_buf_1 _23386_ (.A(_10156_),
    .X(_05783_));
 sg13g2_mux2_1 _23387_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net931),
    .S(net348),
    .X(_01389_));
 sg13g2_mux2_1 _23388_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net932),
    .S(_05781_),
    .X(_01390_));
 sg13g2_mux2_1 _23389_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net484),
    .S(_05780_),
    .X(_01391_));
 sg13g2_mux2_1 _23390_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net485),
    .S(_05780_),
    .X(_01392_));
 sg13g2_nor2_1 _23391_ (.A(_05691_),
    .B(_05778_),
    .Y(_05784_));
 sg13g2_buf_1 _23392_ (.A(_05784_),
    .X(_05785_));
 sg13g2_buf_1 _23393_ (.A(_05785_),
    .X(_05786_));
 sg13g2_mux2_1 _23394_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net483),
    .S(net275),
    .X(_01393_));
 sg13g2_mux2_1 _23395_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net486),
    .S(net275),
    .X(_01394_));
 sg13g2_mux2_1 _23396_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net807),
    .S(net275),
    .X(_01395_));
 sg13g2_mux2_1 _23397_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net551),
    .S(net275),
    .X(_01396_));
 sg13g2_mux2_1 _23398_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net809),
    .S(net275),
    .X(_01397_));
 sg13g2_mux2_1 _23399_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net808),
    .S(_05786_),
    .X(_01398_));
 sg13g2_mux2_1 _23400_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net933),
    .S(net275),
    .X(_01399_));
 sg13g2_mux2_1 _23401_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net934),
    .S(net275),
    .X(_01400_));
 sg13g2_mux2_1 _23402_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net931),
    .S(net275),
    .X(_01401_));
 sg13g2_mux2_1 _23403_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net932),
    .S(_05786_),
    .X(_01402_));
 sg13g2_mux2_1 _23404_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net484),
    .S(_05785_),
    .X(_01403_));
 sg13g2_mux2_1 _23405_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net485),
    .S(_05785_),
    .X(_01404_));
 sg13g2_nor3_1 _23406_ (.A(net706),
    .B(_05657_),
    .C(net425),
    .Y(_05787_));
 sg13g2_buf_1 _23407_ (.A(_05787_),
    .X(_05788_));
 sg13g2_buf_1 _23408_ (.A(_05788_),
    .X(_05789_));
 sg13g2_mux2_1 _23409_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net483),
    .S(net318),
    .X(_01405_));
 sg13g2_mux2_1 _23410_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net486),
    .S(net318),
    .X(_01406_));
 sg13g2_mux2_1 _23411_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(net807),
    .S(net318),
    .X(_01407_));
 sg13g2_mux2_1 _23412_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05749_),
    .S(net318),
    .X(_01408_));
 sg13g2_mux2_1 _23413_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net809),
    .S(net318),
    .X(_01409_));
 sg13g2_mux2_1 _23414_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net808),
    .S(_05789_),
    .X(_01410_));
 sg13g2_mux2_1 _23415_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net933),
    .S(net318),
    .X(_01411_));
 sg13g2_buf_1 _23416_ (.A(_09985_),
    .X(_05790_));
 sg13g2_mux2_1 _23417_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(net930),
    .S(net318),
    .X(_01412_));
 sg13g2_mux2_1 _23418_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(net931),
    .S(net318),
    .X(_01413_));
 sg13g2_mux2_1 _23419_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net932),
    .S(_05789_),
    .X(_01414_));
 sg13g2_mux2_1 _23420_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(net484),
    .S(_05788_),
    .X(_01415_));
 sg13g2_mux2_1 _23421_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(_05762_),
    .S(_05788_),
    .X(_01416_));
 sg13g2_nor3_1 _23422_ (.A(net706),
    .B(net424),
    .C(_05778_),
    .Y(_05791_));
 sg13g2_buf_1 _23423_ (.A(_05791_),
    .X(_05792_));
 sg13g2_buf_1 _23424_ (.A(_05792_),
    .X(_05793_));
 sg13g2_mux2_1 _23425_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(_05776_),
    .S(net317),
    .X(_01417_));
 sg13g2_mux2_1 _23426_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net486),
    .S(net317),
    .X(_01418_));
 sg13g2_mux2_1 _23427_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(_05782_),
    .S(net317),
    .X(_01419_));
 sg13g2_mux2_1 _23428_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(_05749_),
    .S(net317),
    .X(_01420_));
 sg13g2_mux2_1 _23429_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net809),
    .S(net317),
    .X(_01421_));
 sg13g2_mux2_1 _23430_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(_05773_),
    .S(_05793_),
    .X(_01422_));
 sg13g2_mux2_1 _23431_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(_05774_),
    .S(net317),
    .X(_01423_));
 sg13g2_mux2_1 _23432_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(_05790_),
    .S(net317),
    .X(_01424_));
 sg13g2_mux2_1 _23433_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(_05783_),
    .S(net317),
    .X(_01425_));
 sg13g2_mux2_1 _23434_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net932),
    .S(_05793_),
    .X(_01426_));
 sg13g2_mux2_1 _23435_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net484),
    .S(_05792_),
    .X(_01427_));
 sg13g2_mux2_1 _23436_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net485),
    .S(_05792_),
    .X(_01428_));
 sg13g2_nor3_1 _23437_ (.A(net816),
    .B(net424),
    .C(_05778_),
    .Y(_05794_));
 sg13g2_buf_1 _23438_ (.A(_05794_),
    .X(_05795_));
 sg13g2_buf_1 _23439_ (.A(_05795_),
    .X(_05796_));
 sg13g2_mux2_1 _23440_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(_05776_),
    .S(net316),
    .X(_01429_));
 sg13g2_mux2_1 _23441_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net486),
    .S(net316),
    .X(_01430_));
 sg13g2_mux2_1 _23442_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(_05782_),
    .S(net316),
    .X(_01431_));
 sg13g2_mux2_1 _23443_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(_02878_),
    .S(net316),
    .X(_01432_));
 sg13g2_mux2_1 _23444_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net838),
    .S(net316),
    .X(_01433_));
 sg13g2_mux2_1 _23445_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(_05773_),
    .S(_05796_),
    .X(_01434_));
 sg13g2_mux2_1 _23446_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(_05774_),
    .S(net316),
    .X(_01435_));
 sg13g2_mux2_1 _23447_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(_05790_),
    .S(net316),
    .X(_01436_));
 sg13g2_mux2_1 _23448_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(_05783_),
    .S(net316),
    .X(_01437_));
 sg13g2_mux2_1 _23449_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net932),
    .S(_05796_),
    .X(_01438_));
 sg13g2_mux2_1 _23450_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net484),
    .S(_05795_),
    .X(_01439_));
 sg13g2_mux2_1 _23451_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net485),
    .S(_05795_),
    .X(_01440_));
 sg13g2_nor3_1 _23452_ (.A(_05636_),
    .B(_05657_),
    .C(_05697_),
    .Y(_05797_));
 sg13g2_buf_1 _23453_ (.A(_05797_),
    .X(_05798_));
 sg13g2_buf_1 _23454_ (.A(_05798_),
    .X(_05799_));
 sg13g2_mux2_1 _23455_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net483),
    .S(net315),
    .X(_01441_));
 sg13g2_mux2_1 _23456_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net486),
    .S(net315),
    .X(_01442_));
 sg13g2_mux2_1 _23457_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(net807),
    .S(net315),
    .X(_01443_));
 sg13g2_mux2_1 _23458_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net566),
    .S(net315),
    .X(_01444_));
 sg13g2_mux2_1 _23459_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(net838),
    .S(net315),
    .X(_01445_));
 sg13g2_mux2_1 _23460_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net808),
    .S(net315),
    .X(_01446_));
 sg13g2_mux2_1 _23461_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net933),
    .S(_05799_),
    .X(_01447_));
 sg13g2_mux2_1 _23462_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net930),
    .S(net315),
    .X(_01448_));
 sg13g2_mux2_1 _23463_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net931),
    .S(net315),
    .X(_01449_));
 sg13g2_mux2_1 _23464_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net932),
    .S(_05799_),
    .X(_01450_));
 sg13g2_mux2_1 _23465_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net484),
    .S(_05798_),
    .X(_01451_));
 sg13g2_mux2_1 _23466_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(net485),
    .S(_05798_),
    .X(_01452_));
 sg13g2_nand2_1 _23467_ (.Y(_05800_),
    .A(net1073),
    .B(_05656_));
 sg13g2_nor2_1 _23468_ (.A(_05659_),
    .B(_05800_),
    .Y(_05801_));
 sg13g2_buf_1 _23469_ (.A(_05801_),
    .X(_05802_));
 sg13g2_buf_1 _23470_ (.A(_05802_),
    .X(_05803_));
 sg13g2_mux2_1 _23471_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net483),
    .S(net347),
    .X(_01453_));
 sg13g2_mux2_1 _23472_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net486),
    .S(net347),
    .X(_01454_));
 sg13g2_mux2_1 _23473_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net807),
    .S(net347),
    .X(_01455_));
 sg13g2_mux2_1 _23474_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net566),
    .S(net347),
    .X(_01456_));
 sg13g2_mux2_1 _23475_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net838),
    .S(net347),
    .X(_01457_));
 sg13g2_mux2_1 _23476_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net808),
    .S(_05803_),
    .X(_01458_));
 sg13g2_mux2_1 _23477_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net933),
    .S(net347),
    .X(_01459_));
 sg13g2_mux2_1 _23478_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net930),
    .S(net347),
    .X(_01460_));
 sg13g2_mux2_1 _23479_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net931),
    .S(net347),
    .X(_01461_));
 sg13g2_mux2_1 _23480_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net932),
    .S(_05803_),
    .X(_01462_));
 sg13g2_mux2_1 _23481_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(_05767_),
    .S(_05802_),
    .X(_01463_));
 sg13g2_mux2_1 _23482_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05762_),
    .S(_05802_),
    .X(_01464_));
 sg13g2_nor2_1 _23483_ (.A(_05689_),
    .B(_05800_),
    .Y(_05804_));
 sg13g2_buf_2 _23484_ (.A(_05804_),
    .X(_05805_));
 sg13g2_nor2b_1 _23485_ (.A(net425),
    .B_N(_05805_),
    .Y(_05806_));
 sg13g2_buf_1 _23486_ (.A(_05806_),
    .X(_05807_));
 sg13g2_buf_1 _23487_ (.A(_05807_),
    .X(_05808_));
 sg13g2_mux2_1 _23488_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net483),
    .S(net314),
    .X(_01465_));
 sg13g2_mux2_1 _23489_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net506),
    .S(net314),
    .X(_01466_));
 sg13g2_mux2_1 _23490_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net807),
    .S(net314),
    .X(_01467_));
 sg13g2_mux2_1 _23491_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net566),
    .S(net314),
    .X(_01468_));
 sg13g2_mux2_1 _23492_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net838),
    .S(net314),
    .X(_01469_));
 sg13g2_mux2_1 _23493_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net808),
    .S(_05808_),
    .X(_01470_));
 sg13g2_mux2_1 _23494_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(net933),
    .S(net314),
    .X(_01471_));
 sg13g2_mux2_1 _23495_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net930),
    .S(net314),
    .X(_01472_));
 sg13g2_mux2_1 _23496_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net931),
    .S(net314),
    .X(_01473_));
 sg13g2_mux2_1 _23497_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net932),
    .S(_05808_),
    .X(_01474_));
 sg13g2_mux2_1 _23498_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(_05767_),
    .S(_05807_),
    .X(_01475_));
 sg13g2_mux2_1 _23499_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net507),
    .S(_05807_),
    .X(_01476_));
 sg13g2_nor2_1 _23500_ (.A(net817),
    .B(net706),
    .Y(_05809_));
 sg13g2_and2_1 _23501_ (.A(_05656_),
    .B(_05809_),
    .X(_05810_));
 sg13g2_buf_1 _23502_ (.A(_05810_),
    .X(_05811_));
 sg13g2_nor2b_1 _23503_ (.A(_05667_),
    .B_N(_05811_),
    .Y(_05812_));
 sg13g2_buf_1 _23504_ (.A(_05812_),
    .X(_05813_));
 sg13g2_buf_1 _23505_ (.A(_05813_),
    .X(_05814_));
 sg13g2_mux2_1 _23506_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net483),
    .S(net313),
    .X(_01477_));
 sg13g2_mux2_1 _23507_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(net506),
    .S(net313),
    .X(_01478_));
 sg13g2_mux2_1 _23508_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net807),
    .S(net313),
    .X(_01479_));
 sg13g2_mux2_1 _23509_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net566),
    .S(net313),
    .X(_01480_));
 sg13g2_mux2_1 _23510_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net838),
    .S(net313),
    .X(_01481_));
 sg13g2_mux2_1 _23511_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net808),
    .S(_05814_),
    .X(_01482_));
 sg13g2_mux2_1 _23512_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net933),
    .S(net313),
    .X(_01483_));
 sg13g2_mux2_1 _23513_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(net930),
    .S(net313),
    .X(_01484_));
 sg13g2_mux2_1 _23514_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(net931),
    .S(net313),
    .X(_01485_));
 sg13g2_mux2_1 _23515_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(_05775_),
    .S(_05814_),
    .X(_01486_));
 sg13g2_mux2_1 _23516_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net508),
    .S(_05813_),
    .X(_01487_));
 sg13g2_mux2_1 _23517_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net507),
    .S(_05813_),
    .X(_01488_));
 sg13g2_and2_1 _23518_ (.A(_05637_),
    .B(_05656_),
    .X(_05815_));
 sg13g2_buf_2 _23519_ (.A(_05815_),
    .X(_05816_));
 sg13g2_nor2b_1 _23520_ (.A(_05667_),
    .B_N(_05816_),
    .Y(_05817_));
 sg13g2_buf_1 _23521_ (.A(_05817_),
    .X(_05818_));
 sg13g2_buf_1 _23522_ (.A(_05818_),
    .X(_05819_));
 sg13g2_mux2_1 _23523_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(net483),
    .S(_05819_),
    .X(_01489_));
 sg13g2_mux2_1 _23524_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net506),
    .S(net312),
    .X(_01490_));
 sg13g2_mux2_1 _23525_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net807),
    .S(net312),
    .X(_01491_));
 sg13g2_mux2_1 _23526_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net566),
    .S(net312),
    .X(_01492_));
 sg13g2_mux2_1 _23527_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net838),
    .S(net312),
    .X(_01493_));
 sg13g2_mux2_1 _23528_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net843),
    .S(net312),
    .X(_01494_));
 sg13g2_mux2_1 _23529_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net955),
    .S(net312),
    .X(_01495_));
 sg13g2_mux2_1 _23530_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net930),
    .S(net312),
    .X(_01496_));
 sg13g2_mux2_1 _23531_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net931),
    .S(net312),
    .X(_01497_));
 sg13g2_mux2_1 _23532_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net952),
    .S(_05819_),
    .X(_01498_));
 sg13g2_mux2_1 _23533_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net508),
    .S(_05818_),
    .X(_01499_));
 sg13g2_mux2_1 _23534_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net507),
    .S(_05818_),
    .X(_01500_));
 sg13g2_nor3_1 _23535_ (.A(net424),
    .B(_05672_),
    .C(_05707_),
    .Y(_05820_));
 sg13g2_buf_1 _23536_ (.A(_05820_),
    .X(_05821_));
 sg13g2_buf_1 _23537_ (.A(_05821_),
    .X(_05822_));
 sg13g2_mux2_1 _23538_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_11613_),
    .S(_05822_),
    .X(_01501_));
 sg13g2_mux2_1 _23539_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(_03352_),
    .S(net311),
    .X(_01502_));
 sg13g2_mux2_1 _23540_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_10200_),
    .S(net311),
    .X(_01503_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(net566),
    .S(_05822_),
    .X(_01504_));
 sg13g2_mux2_1 _23542_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(_02881_),
    .S(net311),
    .X(_01505_));
 sg13g2_mux2_1 _23543_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(net843),
    .S(net311),
    .X(_01506_));
 sg13g2_mux2_1 _23544_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net955),
    .S(net311),
    .X(_01507_));
 sg13g2_mux2_1 _23545_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net930),
    .S(net311),
    .X(_01508_));
 sg13g2_mux2_1 _23546_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net953),
    .S(net311),
    .X(_01509_));
 sg13g2_mux2_1 _23547_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net952),
    .S(net311),
    .X(_01510_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net508),
    .S(_05821_),
    .X(_01511_));
 sg13g2_mux2_1 _23549_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(net507),
    .S(_05821_),
    .X(_01512_));
 sg13g2_nor3_1 _23550_ (.A(net940),
    .B(_05672_),
    .C(_05691_),
    .Y(_05823_));
 sg13g2_buf_1 _23551_ (.A(_05823_),
    .X(_05824_));
 sg13g2_buf_1 _23552_ (.A(_05824_),
    .X(_05825_));
 sg13g2_mux2_1 _23553_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(_11613_),
    .S(_05825_),
    .X(_01513_));
 sg13g2_mux2_1 _23554_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_03352_),
    .S(net274),
    .X(_01514_));
 sg13g2_mux2_1 _23555_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(net994),
    .S(net274),
    .X(_01515_));
 sg13g2_mux2_1 _23556_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(net566),
    .S(_05825_),
    .X(_01516_));
 sg13g2_mux2_1 _23557_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(_02881_),
    .S(net274),
    .X(_01517_));
 sg13g2_mux2_1 _23558_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_02867_),
    .S(net274),
    .X(_01518_));
 sg13g2_mux2_1 _23559_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(net955),
    .S(net274),
    .X(_01519_));
 sg13g2_mux2_1 _23560_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(net930),
    .S(net274),
    .X(_01520_));
 sg13g2_mux2_1 _23561_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(net953),
    .S(net274),
    .X(_01521_));
 sg13g2_mux2_1 _23562_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_02875_),
    .S(net274),
    .X(_01522_));
 sg13g2_mux2_1 _23563_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_03348_),
    .S(_05824_),
    .X(_01523_));
 sg13g2_mux2_1 _23564_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03350_),
    .S(_05824_),
    .X(_01524_));
 sg13g2_and2_1 _23565_ (.A(_05654_),
    .B(_05656_),
    .X(_05826_));
 sg13g2_buf_1 _23566_ (.A(_05826_),
    .X(_05827_));
 sg13g2_nand2_1 _23567_ (.Y(_05828_),
    .A(_03337_),
    .B(_05609_));
 sg13g2_nor2_1 _23568_ (.A(_11095_),
    .B(_05828_),
    .Y(_05829_));
 sg13g2_buf_1 _23569_ (.A(_05829_),
    .X(_05830_));
 sg13g2_and2_1 _23570_ (.A(_05626_),
    .B(_05830_),
    .X(_05831_));
 sg13g2_buf_1 _23571_ (.A(_05831_),
    .X(_05832_));
 sg13g2_nand2_1 _23572_ (.Y(_05833_),
    .A(_05827_),
    .B(_05832_));
 sg13g2_buf_2 _23573_ (.A(_05833_),
    .X(_05834_));
 sg13g2_buf_1 _23574_ (.A(_05834_),
    .X(_05835_));
 sg13g2_nand2_1 _23575_ (.Y(_05836_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(_05834_));
 sg13g2_o21ai_1 _23576_ (.B1(_05836_),
    .Y(_01525_),
    .A1(net631),
    .A2(net220));
 sg13g2_mux2_1 _23577_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(_05835_),
    .X(_01526_));
 sg13g2_nand2_1 _23578_ (.Y(_05837_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(_05834_));
 sg13g2_o21ai_1 _23579_ (.B1(_05837_),
    .Y(_01527_),
    .A1(net560),
    .A2(_05835_));
 sg13g2_nand2_1 _23580_ (.Y(_05838_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(_05834_));
 sg13g2_o21ai_1 _23581_ (.B1(_05838_),
    .Y(_01528_),
    .A1(net637),
    .A2(net220));
 sg13g2_nand2_1 _23582_ (.Y(_05839_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .B(_05834_));
 sg13g2_o21ai_1 _23583_ (.B1(_05839_),
    .Y(_01529_),
    .A1(net636),
    .A2(net220));
 sg13g2_mux2_1 _23584_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .S(net220),
    .X(_01530_));
 sg13g2_mux2_1 _23585_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net220),
    .X(_01531_));
 sg13g2_mux2_1 _23586_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net220),
    .X(_01532_));
 sg13g2_mux2_1 _23587_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(net220),
    .X(_01533_));
 sg13g2_mux2_1 _23588_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net220),
    .X(_01534_));
 sg13g2_mux2_1 _23589_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(_05834_),
    .X(_01535_));
 sg13g2_mux2_1 _23590_ (.A0(_03605_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_05834_),
    .X(_01536_));
 sg13g2_buf_1 _23591_ (.A(_05830_),
    .X(_05840_));
 sg13g2_nand2_1 _23592_ (.Y(_05841_),
    .A(_05673_),
    .B(net379));
 sg13g2_buf_2 _23593_ (.A(_05841_),
    .X(_05842_));
 sg13g2_buf_1 _23594_ (.A(_05842_),
    .X(_05843_));
 sg13g2_nand2_1 _23595_ (.Y(_05844_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(_05842_));
 sg13g2_o21ai_1 _23596_ (.B1(_05844_),
    .Y(_01537_),
    .A1(net631),
    .A2(net273));
 sg13g2_mux2_1 _23597_ (.A0(_03606_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(net273),
    .X(_01538_));
 sg13g2_nand2_1 _23598_ (.Y(_05845_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(_05842_));
 sg13g2_o21ai_1 _23599_ (.B1(_05845_),
    .Y(_01539_),
    .A1(_03607_),
    .A2(_05843_));
 sg13g2_nand2_1 _23600_ (.Y(_05846_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(_05842_));
 sg13g2_o21ai_1 _23601_ (.B1(_05846_),
    .Y(_01540_),
    .A1(net637),
    .A2(net273));
 sg13g2_nand2_1 _23602_ (.Y(_05847_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .B(_05842_));
 sg13g2_o21ai_1 _23603_ (.B1(_05847_),
    .Y(_01541_),
    .A1(net636),
    .A2(net273));
 sg13g2_mux2_1 _23604_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .S(net273),
    .X(_01542_));
 sg13g2_mux2_1 _23605_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net273),
    .X(_01543_));
 sg13g2_mux2_1 _23606_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net273),
    .X(_01544_));
 sg13g2_mux2_1 _23607_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(_05843_),
    .X(_01545_));
 sg13g2_mux2_1 _23608_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net273),
    .X(_01546_));
 sg13g2_mux2_1 _23609_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(_05842_),
    .X(_01547_));
 sg13g2_mux2_1 _23610_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(_05842_),
    .X(_01548_));
 sg13g2_nand2_1 _23611_ (.Y(_05848_),
    .A(_05678_),
    .B(net379));
 sg13g2_buf_2 _23612_ (.A(_05848_),
    .X(_05849_));
 sg13g2_buf_1 _23613_ (.A(_05849_),
    .X(_05850_));
 sg13g2_nand2_1 _23614_ (.Y(_05851_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(_05849_));
 sg13g2_o21ai_1 _23615_ (.B1(_05851_),
    .Y(_01549_),
    .A1(net631),
    .A2(net272));
 sg13g2_mux2_1 _23616_ (.A0(_03606_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(net272),
    .X(_01550_));
 sg13g2_nand2_1 _23617_ (.Y(_05852_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(_05849_));
 sg13g2_o21ai_1 _23618_ (.B1(_05852_),
    .Y(_01551_),
    .A1(_03607_),
    .A2(_05850_));
 sg13g2_nand2_1 _23619_ (.Y(_05853_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(_05849_));
 sg13g2_o21ai_1 _23620_ (.B1(_05853_),
    .Y(_01552_),
    .A1(net637),
    .A2(net272));
 sg13g2_nand2_1 _23621_ (.Y(_05854_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .B(_05849_));
 sg13g2_o21ai_1 _23622_ (.B1(_05854_),
    .Y(_01553_),
    .A1(net636),
    .A2(net272));
 sg13g2_mux2_1 _23623_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S(net272),
    .X(_01554_));
 sg13g2_mux2_1 _23624_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net272),
    .X(_01555_));
 sg13g2_mux2_1 _23625_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net272),
    .X(_01556_));
 sg13g2_mux2_1 _23626_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(_05850_),
    .X(_01557_));
 sg13g2_mux2_1 _23627_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net272),
    .X(_01558_));
 sg13g2_mux2_1 _23628_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(_05849_),
    .X(_01559_));
 sg13g2_mux2_1 _23629_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(_05849_),
    .X(_01560_));
 sg13g2_nor2_1 _23630_ (.A(_05654_),
    .B(_05672_),
    .Y(_05855_));
 sg13g2_nand2_1 _23631_ (.Y(_05856_),
    .A(_05855_),
    .B(_05832_));
 sg13g2_buf_2 _23632_ (.A(_05856_),
    .X(_05857_));
 sg13g2_buf_1 _23633_ (.A(_05857_),
    .X(_05858_));
 sg13g2_nand2_1 _23634_ (.Y(_05859_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(_05857_));
 sg13g2_o21ai_1 _23635_ (.B1(_05859_),
    .Y(_01561_),
    .A1(net631),
    .A2(net219));
 sg13g2_mux2_1 _23636_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net219),
    .X(_01562_));
 sg13g2_nand2_1 _23637_ (.Y(_05860_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(_05857_));
 sg13g2_o21ai_1 _23638_ (.B1(_05860_),
    .Y(_01563_),
    .A1(net560),
    .A2(_05858_));
 sg13g2_nand2_1 _23639_ (.Y(_05861_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(_05857_));
 sg13g2_o21ai_1 _23640_ (.B1(_05861_),
    .Y(_01564_),
    .A1(net637),
    .A2(net219));
 sg13g2_nand2_1 _23641_ (.Y(_05862_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .B(_05857_));
 sg13g2_o21ai_1 _23642_ (.B1(_05862_),
    .Y(_01565_),
    .A1(net636),
    .A2(_05858_));
 sg13g2_mux2_1 _23643_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .S(net219),
    .X(_01566_));
 sg13g2_mux2_1 _23644_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net219),
    .X(_01567_));
 sg13g2_mux2_1 _23645_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net219),
    .X(_01568_));
 sg13g2_mux2_1 _23646_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net219),
    .X(_01569_));
 sg13g2_mux2_1 _23647_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net219),
    .X(_01570_));
 sg13g2_mux2_1 _23648_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_05857_),
    .X(_01571_));
 sg13g2_mux2_1 _23649_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_05857_),
    .X(_01572_));
 sg13g2_nor3_1 _23650_ (.A(_11095_),
    .B(_05689_),
    .C(_05828_),
    .Y(_05863_));
 sg13g2_buf_2 _23651_ (.A(_05863_),
    .X(_05864_));
 sg13g2_nand2_1 _23652_ (.Y(_05865_),
    .A(_05855_),
    .B(_05864_));
 sg13g2_buf_2 _23653_ (.A(_05865_),
    .X(_05866_));
 sg13g2_buf_1 _23654_ (.A(_05866_),
    .X(_05867_));
 sg13g2_nand2_1 _23655_ (.Y(_05868_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(_05866_));
 sg13g2_o21ai_1 _23656_ (.B1(_05868_),
    .Y(_01573_),
    .A1(net631),
    .A2(net310));
 sg13g2_mux2_1 _23657_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net310),
    .X(_01574_));
 sg13g2_nand2_1 _23658_ (.Y(_05869_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(_05866_));
 sg13g2_o21ai_1 _23659_ (.B1(_05869_),
    .Y(_01575_),
    .A1(net560),
    .A2(_05867_));
 sg13g2_nand2_1 _23660_ (.Y(_05870_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(_05866_));
 sg13g2_o21ai_1 _23661_ (.B1(_05870_),
    .Y(_01576_),
    .A1(net637),
    .A2(net310));
 sg13g2_nand2_1 _23662_ (.Y(_05871_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .B(_05866_));
 sg13g2_o21ai_1 _23663_ (.B1(_05871_),
    .Y(_01577_),
    .A1(net636),
    .A2(net310));
 sg13g2_mux2_1 _23664_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .S(net310),
    .X(_01578_));
 sg13g2_mux2_1 _23665_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net310),
    .X(_01579_));
 sg13g2_mux2_1 _23666_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net310),
    .X(_01580_));
 sg13g2_mux2_1 _23667_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(_05867_),
    .X(_01581_));
 sg13g2_mux2_1 _23668_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net310),
    .X(_01582_));
 sg13g2_mux2_1 _23669_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_05866_),
    .X(_01583_));
 sg13g2_mux2_1 _23670_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_05866_),
    .X(_01584_));
 sg13g2_nor2_1 _23671_ (.A(net941),
    .B(_05620_),
    .Y(_05872_));
 sg13g2_nand3_1 _23672_ (.B(_05855_),
    .C(net379),
    .A(_05872_),
    .Y(_05873_));
 sg13g2_buf_2 _23673_ (.A(_05873_),
    .X(_05874_));
 sg13g2_buf_1 _23674_ (.A(_05874_),
    .X(_05875_));
 sg13g2_nand2_1 _23675_ (.Y(_05876_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(_05874_));
 sg13g2_o21ai_1 _23676_ (.B1(_05876_),
    .Y(_01585_),
    .A1(net631),
    .A2(net271));
 sg13g2_mux2_1 _23677_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net271),
    .X(_01586_));
 sg13g2_nand2_1 _23678_ (.Y(_05877_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(_05874_));
 sg13g2_o21ai_1 _23679_ (.B1(_05877_),
    .Y(_01587_),
    .A1(net560),
    .A2(_05875_));
 sg13g2_nand2_1 _23680_ (.Y(_05878_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(_05874_));
 sg13g2_o21ai_1 _23681_ (.B1(_05878_),
    .Y(_01588_),
    .A1(_02857_),
    .A2(net271));
 sg13g2_nand2_1 _23682_ (.Y(_05879_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .B(_05874_));
 sg13g2_o21ai_1 _23683_ (.B1(_05879_),
    .Y(_01589_),
    .A1(_02864_),
    .A2(net271));
 sg13g2_mux2_1 _23684_ (.A0(_02868_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .S(net271),
    .X(_01590_));
 sg13g2_mux2_1 _23685_ (.A0(_02870_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net271),
    .X(_01591_));
 sg13g2_mux2_1 _23686_ (.A0(_02872_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net271),
    .X(_01592_));
 sg13g2_mux2_1 _23687_ (.A0(_02874_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(_05875_),
    .X(_01593_));
 sg13g2_mux2_1 _23688_ (.A0(_02876_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net271),
    .X(_01594_));
 sg13g2_mux2_1 _23689_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_05874_),
    .X(_01595_));
 sg13g2_mux2_1 _23690_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_05874_),
    .X(_01596_));
 sg13g2_buf_1 _23691_ (.A(_05830_),
    .X(_05880_));
 sg13g2_nand3_1 _23692_ (.B(_05855_),
    .C(net378),
    .A(_05624_),
    .Y(_05881_));
 sg13g2_buf_2 _23693_ (.A(_05881_),
    .X(_05882_));
 sg13g2_buf_1 _23694_ (.A(_05882_),
    .X(_05883_));
 sg13g2_nand2_1 _23695_ (.Y(_05884_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(_05882_));
 sg13g2_o21ai_1 _23696_ (.B1(_05884_),
    .Y(_01597_),
    .A1(net631),
    .A2(net270));
 sg13g2_mux2_1 _23697_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net270),
    .X(_01598_));
 sg13g2_nand2_1 _23698_ (.Y(_05885_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(_05882_));
 sg13g2_o21ai_1 _23699_ (.B1(_05885_),
    .Y(_01599_),
    .A1(net560),
    .A2(_05883_));
 sg13g2_nand2_1 _23700_ (.Y(_05886_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(_05882_));
 sg13g2_o21ai_1 _23701_ (.B1(_05886_),
    .Y(_01600_),
    .A1(_02857_),
    .A2(net270));
 sg13g2_nand2_1 _23702_ (.Y(_05887_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .B(_05882_));
 sg13g2_o21ai_1 _23703_ (.B1(_05887_),
    .Y(_01601_),
    .A1(_02864_),
    .A2(net270));
 sg13g2_mux2_1 _23704_ (.A0(_02868_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S(net270),
    .X(_01602_));
 sg13g2_mux2_1 _23705_ (.A0(_02870_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net270),
    .X(_01603_));
 sg13g2_mux2_1 _23706_ (.A0(_02872_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net270),
    .X(_01604_));
 sg13g2_mux2_1 _23707_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(_05883_),
    .X(_01605_));
 sg13g2_mux2_1 _23708_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net270),
    .X(_01606_));
 sg13g2_mux2_1 _23709_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_05882_),
    .X(_01607_));
 sg13g2_mux2_1 _23710_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_05882_),
    .X(_01608_));
 sg13g2_nor3_2 _23711_ (.A(net941),
    .B(net1072),
    .C(net940),
    .Y(_05888_));
 sg13g2_nand4_1 _23712_ (.B(_10892_),
    .C(_05888_),
    .A(net938),
    .Y(_05889_),
    .D(net378));
 sg13g2_buf_2 _23713_ (.A(_05889_),
    .X(_05890_));
 sg13g2_buf_1 _23714_ (.A(_05890_),
    .X(_05891_));
 sg13g2_nand2_1 _23715_ (.Y(_05892_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(_05890_));
 sg13g2_o21ai_1 _23716_ (.B1(_05892_),
    .Y(_01609_),
    .A1(_03613_),
    .A2(net269));
 sg13g2_mux2_1 _23717_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net269),
    .X(_01610_));
 sg13g2_nand2_1 _23718_ (.Y(_05893_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(_05890_));
 sg13g2_o21ai_1 _23719_ (.B1(_05893_),
    .Y(_01611_),
    .A1(net560),
    .A2(net269));
 sg13g2_buf_1 _23720_ (.A(net716),
    .X(_05894_));
 sg13g2_nand2_1 _23721_ (.Y(_05895_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(_05890_));
 sg13g2_o21ai_1 _23722_ (.B1(_05895_),
    .Y(_01612_),
    .A1(net621),
    .A2(_05891_));
 sg13g2_buf_1 _23723_ (.A(net715),
    .X(_05896_));
 sg13g2_nand2_1 _23724_ (.Y(_05897_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .B(_05890_));
 sg13g2_o21ai_1 _23725_ (.B1(_05897_),
    .Y(_01613_),
    .A1(net620),
    .A2(net269));
 sg13g2_buf_1 _23726_ (.A(net843),
    .X(_05898_));
 sg13g2_mux2_1 _23727_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .S(net269),
    .X(_01614_));
 sg13g2_buf_1 _23728_ (.A(net955),
    .X(_05899_));
 sg13g2_mux2_1 _23729_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net269),
    .X(_01615_));
 sg13g2_buf_1 _23730_ (.A(net954),
    .X(_05900_));
 sg13g2_mux2_1 _23731_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net269),
    .X(_01616_));
 sg13g2_buf_1 _23732_ (.A(net953),
    .X(_05901_));
 sg13g2_mux2_1 _23733_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net269),
    .X(_01617_));
 sg13g2_buf_1 _23734_ (.A(net952),
    .X(_05902_));
 sg13g2_mux2_1 _23735_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(_05891_),
    .X(_01618_));
 sg13g2_mux2_1 _23736_ (.A0(net437),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_05890_),
    .X(_01619_));
 sg13g2_mux2_1 _23737_ (.A0(_03605_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_05890_),
    .X(_01620_));
 sg13g2_nand4_1 _23738_ (.B(net817),
    .C(_10892_),
    .A(net938),
    .Y(_05903_),
    .D(_05864_));
 sg13g2_buf_2 _23739_ (.A(_05903_),
    .X(_05904_));
 sg13g2_buf_1 _23740_ (.A(_05904_),
    .X(_05905_));
 sg13g2_nand2_1 _23741_ (.Y(_05906_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(_05904_));
 sg13g2_o21ai_1 _23742_ (.B1(_05906_),
    .Y(_01621_),
    .A1(_03613_),
    .A2(net309));
 sg13g2_mux2_1 _23743_ (.A0(net435),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(net309),
    .X(_01622_));
 sg13g2_nand2_1 _23744_ (.Y(_05907_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(_05904_));
 sg13g2_o21ai_1 _23745_ (.B1(_05907_),
    .Y(_01623_),
    .A1(net560),
    .A2(net309));
 sg13g2_nand2_1 _23746_ (.Y(_05908_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_05904_));
 sg13g2_o21ai_1 _23747_ (.B1(_05908_),
    .Y(_01624_),
    .A1(net621),
    .A2(_05905_));
 sg13g2_nand2_1 _23748_ (.Y(_05909_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .B(_05904_));
 sg13g2_o21ai_1 _23749_ (.B1(_05909_),
    .Y(_01625_),
    .A1(_05896_),
    .A2(net309));
 sg13g2_mux2_1 _23750_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .S(net309),
    .X(_01626_));
 sg13g2_mux2_1 _23751_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net309),
    .X(_01627_));
 sg13g2_mux2_1 _23752_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net309),
    .X(_01628_));
 sg13g2_mux2_1 _23753_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net309),
    .X(_01629_));
 sg13g2_mux2_1 _23754_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(_05905_),
    .X(_01630_));
 sg13g2_mux2_1 _23755_ (.A0(_03604_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(_05904_),
    .X(_01631_));
 sg13g2_mux2_1 _23756_ (.A0(net436),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_05904_),
    .X(_01632_));
 sg13g2_buf_1 _23757_ (.A(net708),
    .X(_05910_));
 sg13g2_nand2_1 _23758_ (.Y(_05911_),
    .A(_05719_),
    .B(net379));
 sg13g2_buf_2 _23759_ (.A(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _23760_ (.A(_05912_),
    .X(_05913_));
 sg13g2_nand2_1 _23761_ (.Y(_05914_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(_05912_));
 sg13g2_o21ai_1 _23762_ (.B1(_05914_),
    .Y(_01633_),
    .A1(net619),
    .A2(net268));
 sg13g2_buf_1 _23763_ (.A(net506),
    .X(_05915_));
 sg13g2_mux2_1 _23764_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(net268),
    .X(_01634_));
 sg13g2_buf_1 _23765_ (.A(net679),
    .X(_05916_));
 sg13g2_nand2_1 _23766_ (.Y(_05917_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(_05912_));
 sg13g2_o21ai_1 _23767_ (.B1(_05917_),
    .Y(_01635_),
    .A1(_05916_),
    .A2(net268));
 sg13g2_nand2_1 _23768_ (.Y(_05918_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_05912_));
 sg13g2_o21ai_1 _23769_ (.B1(_05918_),
    .Y(_01636_),
    .A1(_05894_),
    .A2(_05913_));
 sg13g2_nand2_1 _23770_ (.Y(_05919_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .B(_05912_));
 sg13g2_o21ai_1 _23771_ (.B1(_05919_),
    .Y(_01637_),
    .A1(net620),
    .A2(net268));
 sg13g2_mux2_1 _23772_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .S(net268),
    .X(_01638_));
 sg13g2_mux2_1 _23773_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net268),
    .X(_01639_));
 sg13g2_mux2_1 _23774_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net268),
    .X(_01640_));
 sg13g2_mux2_1 _23775_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net268),
    .X(_01641_));
 sg13g2_mux2_1 _23776_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(_05913_),
    .X(_01642_));
 sg13g2_buf_1 _23777_ (.A(net508),
    .X(_05920_));
 sg13g2_mux2_1 _23778_ (.A0(_05920_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_05912_),
    .X(_01643_));
 sg13g2_buf_1 _23779_ (.A(net507),
    .X(_05921_));
 sg13g2_mux2_1 _23780_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_05912_),
    .X(_01644_));
 sg13g2_nand2_1 _23781_ (.Y(_05922_),
    .A(_05728_),
    .B(net379));
 sg13g2_buf_2 _23782_ (.A(_05922_),
    .X(_05923_));
 sg13g2_buf_1 _23783_ (.A(_05923_),
    .X(_05924_));
 sg13g2_nand2_1 _23784_ (.Y(_05925_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(_05923_));
 sg13g2_o21ai_1 _23785_ (.B1(_05925_),
    .Y(_01645_),
    .A1(net619),
    .A2(net267));
 sg13g2_mux2_1 _23786_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(net267),
    .X(_01646_));
 sg13g2_nand2_1 _23787_ (.Y(_05926_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(_05923_));
 sg13g2_o21ai_1 _23788_ (.B1(_05926_),
    .Y(_01647_),
    .A1(net550),
    .A2(net267));
 sg13g2_nand2_1 _23789_ (.Y(_05927_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_05923_));
 sg13g2_o21ai_1 _23790_ (.B1(_05927_),
    .Y(_01648_),
    .A1(net621),
    .A2(_05924_));
 sg13g2_nand2_1 _23791_ (.Y(_05928_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .B(_05923_));
 sg13g2_o21ai_1 _23792_ (.B1(_05928_),
    .Y(_01649_),
    .A1(net620),
    .A2(net267));
 sg13g2_mux2_1 _23793_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S(net267),
    .X(_01650_));
 sg13g2_mux2_1 _23794_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net267),
    .X(_01651_));
 sg13g2_mux2_1 _23795_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net267),
    .X(_01652_));
 sg13g2_mux2_1 _23796_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net267),
    .X(_01653_));
 sg13g2_mux2_1 _23797_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(_05924_),
    .X(_01654_));
 sg13g2_mux2_1 _23798_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(_05923_),
    .X(_01655_));
 sg13g2_mux2_1 _23799_ (.A0(_05921_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_05923_),
    .X(_01656_));
 sg13g2_nand2_1 _23800_ (.Y(_05929_),
    .A(_05827_),
    .B(_05864_));
 sg13g2_buf_2 _23801_ (.A(_05929_),
    .X(_05930_));
 sg13g2_buf_1 _23802_ (.A(_05930_),
    .X(_05931_));
 sg13g2_nand2_1 _23803_ (.Y(_05932_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(_05930_));
 sg13g2_o21ai_1 _23804_ (.B1(_05932_),
    .Y(_01657_),
    .A1(_05910_),
    .A2(net308));
 sg13g2_mux2_1 _23805_ (.A0(_05915_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net308),
    .X(_01658_));
 sg13g2_nand2_1 _23806_ (.Y(_05933_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(_05930_));
 sg13g2_o21ai_1 _23807_ (.B1(_05933_),
    .Y(_01659_),
    .A1(net550),
    .A2(net308));
 sg13g2_nand2_1 _23808_ (.Y(_05934_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(_05930_));
 sg13g2_o21ai_1 _23809_ (.B1(_05934_),
    .Y(_01660_),
    .A1(_05894_),
    .A2(_05931_));
 sg13g2_nand2_1 _23810_ (.Y(_05935_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .B(_05930_));
 sg13g2_o21ai_1 _23811_ (.B1(_05935_),
    .Y(_01661_),
    .A1(net620),
    .A2(_05931_));
 sg13g2_mux2_1 _23812_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .S(net308),
    .X(_01662_));
 sg13g2_mux2_1 _23813_ (.A0(_05899_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net308),
    .X(_01663_));
 sg13g2_mux2_1 _23814_ (.A0(_05900_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net308),
    .X(_01664_));
 sg13g2_mux2_1 _23815_ (.A0(_05901_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net308),
    .X(_01665_));
 sg13g2_mux2_1 _23816_ (.A0(_05902_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net308),
    .X(_01666_));
 sg13g2_mux2_1 _23817_ (.A0(_05920_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_05930_),
    .X(_01667_));
 sg13g2_mux2_1 _23818_ (.A0(_05921_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_05930_),
    .X(_01668_));
 sg13g2_nor2_1 _23819_ (.A(_05654_),
    .B(_05706_),
    .Y(_05936_));
 sg13g2_nand2_1 _23820_ (.Y(_05937_),
    .A(_05936_),
    .B(_05832_));
 sg13g2_buf_2 _23821_ (.A(_05937_),
    .X(_05938_));
 sg13g2_buf_1 _23822_ (.A(_05938_),
    .X(_05939_));
 sg13g2_nand2_1 _23823_ (.Y(_05940_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(_05938_));
 sg13g2_o21ai_1 _23824_ (.B1(_05940_),
    .Y(_01669_),
    .A1(net619),
    .A2(_05939_));
 sg13g2_mux2_1 _23825_ (.A0(_05915_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net218),
    .X(_01670_));
 sg13g2_nand2_1 _23826_ (.Y(_05941_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(_05938_));
 sg13g2_o21ai_1 _23827_ (.B1(_05941_),
    .Y(_01671_),
    .A1(net550),
    .A2(net218));
 sg13g2_nand2_1 _23828_ (.Y(_05942_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(_05938_));
 sg13g2_o21ai_1 _23829_ (.B1(_05942_),
    .Y(_01672_),
    .A1(net621),
    .A2(_05939_));
 sg13g2_nand2_1 _23830_ (.Y(_05943_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .B(_05938_));
 sg13g2_o21ai_1 _23831_ (.B1(_05943_),
    .Y(_01673_),
    .A1(net620),
    .A2(net218));
 sg13g2_mux2_1 _23832_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .S(net218),
    .X(_01674_));
 sg13g2_mux2_1 _23833_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net218),
    .X(_01675_));
 sg13g2_mux2_1 _23834_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(net218),
    .X(_01676_));
 sg13g2_mux2_1 _23835_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net218),
    .X(_01677_));
 sg13g2_mux2_1 _23836_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(net218),
    .X(_01678_));
 sg13g2_mux2_1 _23837_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(_05938_),
    .X(_01679_));
 sg13g2_mux2_1 _23838_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(_05938_),
    .X(_01680_));
 sg13g2_nand2_1 _23839_ (.Y(_05944_),
    .A(_05936_),
    .B(_05864_));
 sg13g2_buf_2 _23840_ (.A(_05944_),
    .X(_05945_));
 sg13g2_buf_1 _23841_ (.A(_05945_),
    .X(_05946_));
 sg13g2_nand2_1 _23842_ (.Y(_05947_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(_05945_));
 sg13g2_o21ai_1 _23843_ (.B1(_05947_),
    .Y(_01681_),
    .A1(net619),
    .A2(_05946_));
 sg13g2_mux2_1 _23844_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net307),
    .X(_01682_));
 sg13g2_nand2_1 _23845_ (.Y(_05948_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(_05945_));
 sg13g2_o21ai_1 _23846_ (.B1(_05948_),
    .Y(_01683_),
    .A1(net550),
    .A2(net307));
 sg13g2_nand2_1 _23847_ (.Y(_05949_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(_05945_));
 sg13g2_o21ai_1 _23848_ (.B1(_05949_),
    .Y(_01684_),
    .A1(net621),
    .A2(_05946_));
 sg13g2_nand2_1 _23849_ (.Y(_05950_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .B(_05945_));
 sg13g2_o21ai_1 _23850_ (.B1(_05950_),
    .Y(_01685_),
    .A1(net620),
    .A2(net307));
 sg13g2_mux2_1 _23851_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .S(net307),
    .X(_01686_));
 sg13g2_mux2_1 _23852_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net307),
    .X(_01687_));
 sg13g2_mux2_1 _23853_ (.A0(_05900_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(net307),
    .X(_01688_));
 sg13g2_mux2_1 _23854_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net307),
    .X(_01689_));
 sg13g2_mux2_1 _23855_ (.A0(_05902_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(net307),
    .X(_01690_));
 sg13g2_mux2_1 _23856_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(_05945_),
    .X(_01691_));
 sg13g2_mux2_1 _23857_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(_05945_),
    .X(_01692_));
 sg13g2_nand3_1 _23858_ (.B(_05936_),
    .C(_05880_),
    .A(_05872_),
    .Y(_05951_));
 sg13g2_buf_2 _23859_ (.A(_05951_),
    .X(_05952_));
 sg13g2_buf_1 _23860_ (.A(_05952_),
    .X(_05953_));
 sg13g2_nand2_1 _23861_ (.Y(_05954_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(_05952_));
 sg13g2_o21ai_1 _23862_ (.B1(_05954_),
    .Y(_01693_),
    .A1(net619),
    .A2(_05953_));
 sg13g2_mux2_1 _23863_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net266),
    .X(_01694_));
 sg13g2_nand2_1 _23864_ (.Y(_05955_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(_05952_));
 sg13g2_o21ai_1 _23865_ (.B1(_05955_),
    .Y(_01695_),
    .A1(net550),
    .A2(net266));
 sg13g2_nand2_1 _23866_ (.Y(_05956_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(_05952_));
 sg13g2_o21ai_1 _23867_ (.B1(_05956_),
    .Y(_01696_),
    .A1(net621),
    .A2(_05953_));
 sg13g2_nand2_1 _23868_ (.Y(_05957_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .B(_05952_));
 sg13g2_o21ai_1 _23869_ (.B1(_05957_),
    .Y(_01697_),
    .A1(net620),
    .A2(net266));
 sg13g2_mux2_1 _23870_ (.A0(_05898_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .S(net266),
    .X(_01698_));
 sg13g2_mux2_1 _23871_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net266),
    .X(_01699_));
 sg13g2_mux2_1 _23872_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(net266),
    .X(_01700_));
 sg13g2_mux2_1 _23873_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net266),
    .X(_01701_));
 sg13g2_mux2_1 _23874_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(net266),
    .X(_01702_));
 sg13g2_mux2_1 _23875_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(_05952_),
    .X(_01703_));
 sg13g2_mux2_1 _23876_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_05952_),
    .X(_01704_));
 sg13g2_nand3_1 _23877_ (.B(_05936_),
    .C(net378),
    .A(_05624_),
    .Y(_05958_));
 sg13g2_buf_2 _23878_ (.A(_05958_),
    .X(_05959_));
 sg13g2_buf_1 _23879_ (.A(_05959_),
    .X(_05960_));
 sg13g2_nand2_1 _23880_ (.Y(_05961_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(_05959_));
 sg13g2_o21ai_1 _23881_ (.B1(_05961_),
    .Y(_01705_),
    .A1(_05910_),
    .A2(_05960_));
 sg13g2_mux2_1 _23882_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net265),
    .X(_01706_));
 sg13g2_nand2_1 _23883_ (.Y(_05962_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(_05959_));
 sg13g2_o21ai_1 _23884_ (.B1(_05962_),
    .Y(_01707_),
    .A1(net550),
    .A2(net265));
 sg13g2_nand2_1 _23885_ (.Y(_05963_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(_05959_));
 sg13g2_o21ai_1 _23886_ (.B1(_05963_),
    .Y(_01708_),
    .A1(net621),
    .A2(_05960_));
 sg13g2_nand2_1 _23887_ (.Y(_05964_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .B(_05959_));
 sg13g2_o21ai_1 _23888_ (.B1(_05964_),
    .Y(_01709_),
    .A1(_05896_),
    .A2(net265));
 sg13g2_mux2_1 _23889_ (.A0(_05898_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S(net265),
    .X(_01710_));
 sg13g2_mux2_1 _23890_ (.A0(_05899_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net265),
    .X(_01711_));
 sg13g2_mux2_1 _23891_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(net265),
    .X(_01712_));
 sg13g2_mux2_1 _23892_ (.A0(_05901_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net265),
    .X(_01713_));
 sg13g2_mux2_1 _23893_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net265),
    .X(_01714_));
 sg13g2_mux2_1 _23894_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(_05959_),
    .X(_01715_));
 sg13g2_mux2_1 _23895_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_05959_),
    .X(_01716_));
 sg13g2_nand4_1 _23896_ (.B(net939),
    .C(_05888_),
    .A(net938),
    .Y(_05965_),
    .D(net378));
 sg13g2_buf_2 _23897_ (.A(_05965_),
    .X(_05966_));
 sg13g2_buf_1 _23898_ (.A(_05966_),
    .X(_05967_));
 sg13g2_nand2_1 _23899_ (.Y(_05968_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(_05966_));
 sg13g2_o21ai_1 _23900_ (.B1(_05968_),
    .Y(_01717_),
    .A1(net619),
    .A2(_05967_));
 sg13g2_mux2_1 _23901_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(_05967_),
    .X(_01718_));
 sg13g2_nand2_1 _23902_ (.Y(_05969_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(_05966_));
 sg13g2_o21ai_1 _23903_ (.B1(_05969_),
    .Y(_01719_),
    .A1(net550),
    .A2(net264));
 sg13g2_nand2_1 _23904_ (.Y(_05970_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(_05966_));
 sg13g2_o21ai_1 _23905_ (.B1(_05970_),
    .Y(_01720_),
    .A1(net621),
    .A2(net264));
 sg13g2_nand2_1 _23906_ (.Y(_05971_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .B(_05966_));
 sg13g2_o21ai_1 _23907_ (.B1(_05971_),
    .Y(_01721_),
    .A1(net620),
    .A2(net264));
 sg13g2_mux2_1 _23908_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .S(net264),
    .X(_01722_));
 sg13g2_mux2_1 _23909_ (.A0(net806),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net264),
    .X(_01723_));
 sg13g2_mux2_1 _23910_ (.A0(net805),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(net264),
    .X(_01724_));
 sg13g2_mux2_1 _23911_ (.A0(net804),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net264),
    .X(_01725_));
 sg13g2_mux2_1 _23912_ (.A0(net803),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net264),
    .X(_01726_));
 sg13g2_mux2_1 _23913_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_05966_),
    .X(_01727_));
 sg13g2_mux2_1 _23914_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(_05966_),
    .X(_01728_));
 sg13g2_nand4_1 _23915_ (.B(net817),
    .C(net939),
    .A(net938),
    .Y(_05972_),
    .D(_05864_));
 sg13g2_buf_2 _23916_ (.A(_05972_),
    .X(_05973_));
 sg13g2_buf_1 _23917_ (.A(_05973_),
    .X(_05974_));
 sg13g2_nand2_1 _23918_ (.Y(_05975_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(_05973_));
 sg13g2_o21ai_1 _23919_ (.B1(_05975_),
    .Y(_01729_),
    .A1(net619),
    .A2(_05974_));
 sg13g2_mux2_1 _23920_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(_05974_),
    .X(_01730_));
 sg13g2_nand2_1 _23921_ (.Y(_05976_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(_05973_));
 sg13g2_o21ai_1 _23922_ (.B1(_05976_),
    .Y(_01731_),
    .A1(net550),
    .A2(net306));
 sg13g2_buf_1 _23923_ (.A(net716),
    .X(_05977_));
 sg13g2_nand2_1 _23924_ (.Y(_05978_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(_05973_));
 sg13g2_o21ai_1 _23925_ (.B1(_05978_),
    .Y(_01732_),
    .A1(net618),
    .A2(net306));
 sg13g2_buf_1 _23926_ (.A(net715),
    .X(_05979_));
 sg13g2_nand2_1 _23927_ (.Y(_05980_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .B(_05973_));
 sg13g2_o21ai_1 _23928_ (.B1(_05980_),
    .Y(_01733_),
    .A1(net617),
    .A2(net306));
 sg13g2_buf_1 _23929_ (.A(net843),
    .X(_05981_));
 sg13g2_mux2_1 _23930_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .S(net306),
    .X(_01734_));
 sg13g2_buf_1 _23931_ (.A(net955),
    .X(_05982_));
 sg13g2_mux2_1 _23932_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net306),
    .X(_01735_));
 sg13g2_buf_1 _23933_ (.A(_02871_),
    .X(_05983_));
 sg13g2_mux2_1 _23934_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(net306),
    .X(_01736_));
 sg13g2_buf_1 _23935_ (.A(_02873_),
    .X(_05984_));
 sg13g2_mux2_1 _23936_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net306),
    .X(_01737_));
 sg13g2_buf_1 _23937_ (.A(net952),
    .X(_05985_));
 sg13g2_mux2_1 _23938_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net306),
    .X(_01738_));
 sg13g2_mux2_1 _23939_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(_05973_),
    .X(_01739_));
 sg13g2_mux2_1 _23940_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(_05973_),
    .X(_01740_));
 sg13g2_nand2_1 _23941_ (.Y(_05986_),
    .A(_05763_),
    .B(_05840_));
 sg13g2_buf_2 _23942_ (.A(_05986_),
    .X(_05987_));
 sg13g2_buf_1 _23943_ (.A(_05987_),
    .X(_05988_));
 sg13g2_nand2_1 _23944_ (.Y(_05989_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(_05987_));
 sg13g2_o21ai_1 _23945_ (.B1(_05989_),
    .Y(_01741_),
    .A1(net619),
    .A2(net263));
 sg13g2_mux2_1 _23946_ (.A0(net423),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(_05988_),
    .X(_01742_));
 sg13g2_nand2_1 _23947_ (.Y(_05990_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(_05987_));
 sg13g2_o21ai_1 _23948_ (.B1(_05990_),
    .Y(_01743_),
    .A1(_05916_),
    .A2(net263));
 sg13g2_nand2_1 _23949_ (.Y(_05991_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(_05987_));
 sg13g2_o21ai_1 _23950_ (.B1(_05991_),
    .Y(_01744_),
    .A1(net618),
    .A2(net263));
 sg13g2_nand2_1 _23951_ (.Y(_05992_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .B(_05987_));
 sg13g2_o21ai_1 _23952_ (.B1(_05992_),
    .Y(_01745_),
    .A1(net617),
    .A2(net263));
 sg13g2_mux2_1 _23953_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .S(net263),
    .X(_01746_));
 sg13g2_mux2_1 _23954_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net263),
    .X(_01747_));
 sg13g2_mux2_1 _23955_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(net263),
    .X(_01748_));
 sg13g2_mux2_1 _23956_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(_05988_),
    .X(_01749_));
 sg13g2_mux2_1 _23957_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net263),
    .X(_01750_));
 sg13g2_mux2_1 _23958_ (.A0(net422),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_05987_),
    .X(_01751_));
 sg13g2_mux2_1 _23959_ (.A0(net421),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_05987_),
    .X(_01752_));
 sg13g2_buf_1 _23960_ (.A(net708),
    .X(_05993_));
 sg13g2_nand2_1 _23961_ (.Y(_05994_),
    .A(_05769_),
    .B(net379));
 sg13g2_buf_2 _23962_ (.A(_05994_),
    .X(_05995_));
 sg13g2_buf_1 _23963_ (.A(_05995_),
    .X(_05996_));
 sg13g2_nand2_1 _23964_ (.Y(_05997_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(_05995_));
 sg13g2_o21ai_1 _23965_ (.B1(_05997_),
    .Y(_01753_),
    .A1(net616),
    .A2(_05996_));
 sg13g2_buf_1 _23966_ (.A(net506),
    .X(_05998_));
 sg13g2_mux2_1 _23967_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net262),
    .X(_01754_));
 sg13g2_buf_1 _23968_ (.A(net679),
    .X(_05999_));
 sg13g2_nand2_1 _23969_ (.Y(_06000_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(_05995_));
 sg13g2_o21ai_1 _23970_ (.B1(_06000_),
    .Y(_01755_),
    .A1(net549),
    .A2(net262));
 sg13g2_nand2_1 _23971_ (.Y(_06001_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(_05995_));
 sg13g2_o21ai_1 _23972_ (.B1(_06001_),
    .Y(_01756_),
    .A1(net618),
    .A2(net262));
 sg13g2_nand2_1 _23973_ (.Y(_06002_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .B(_05995_));
 sg13g2_o21ai_1 _23974_ (.B1(_06002_),
    .Y(_01757_),
    .A1(_05979_),
    .A2(net262));
 sg13g2_mux2_1 _23975_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S(net262),
    .X(_01758_));
 sg13g2_mux2_1 _23976_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net262),
    .X(_01759_));
 sg13g2_mux2_1 _23977_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(net262),
    .X(_01760_));
 sg13g2_mux2_1 _23978_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(_05996_),
    .X(_01761_));
 sg13g2_mux2_1 _23979_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net262),
    .X(_01762_));
 sg13g2_buf_1 _23980_ (.A(net508),
    .X(_06003_));
 sg13g2_mux2_1 _23981_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(_05995_),
    .X(_01763_));
 sg13g2_buf_1 _23982_ (.A(net507),
    .X(_06004_));
 sg13g2_mux2_1 _23983_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(_05995_),
    .X(_01764_));
 sg13g2_nor2_1 _23984_ (.A(_05654_),
    .B(_05754_),
    .Y(_06005_));
 sg13g2_nand2_1 _23985_ (.Y(_06006_),
    .A(_06005_),
    .B(_05832_));
 sg13g2_buf_2 _23986_ (.A(_06006_),
    .X(_06007_));
 sg13g2_buf_1 _23987_ (.A(_06007_),
    .X(_06008_));
 sg13g2_nand2_1 _23988_ (.Y(_06009_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(_06007_));
 sg13g2_o21ai_1 _23989_ (.B1(_06009_),
    .Y(_01765_),
    .A1(net616),
    .A2(net217));
 sg13g2_mux2_1 _23990_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net217),
    .X(_01766_));
 sg13g2_nand2_1 _23991_ (.Y(_06010_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(_06007_));
 sg13g2_o21ai_1 _23992_ (.B1(_06010_),
    .Y(_01767_),
    .A1(net549),
    .A2(net217));
 sg13g2_nand2_1 _23993_ (.Y(_06011_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(_06007_));
 sg13g2_o21ai_1 _23994_ (.B1(_06011_),
    .Y(_01768_),
    .A1(net618),
    .A2(net217));
 sg13g2_nand2_1 _23995_ (.Y(_06012_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .B(_06007_));
 sg13g2_o21ai_1 _23996_ (.B1(_06012_),
    .Y(_01769_),
    .A1(net617),
    .A2(net217));
 sg13g2_mux2_1 _23997_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .S(net217),
    .X(_01770_));
 sg13g2_mux2_1 _23998_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net217),
    .X(_01771_));
 sg13g2_mux2_1 _23999_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(net217),
    .X(_01772_));
 sg13g2_mux2_1 _24000_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(_06008_),
    .X(_01773_));
 sg13g2_mux2_1 _24001_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(_06008_),
    .X(_01774_));
 sg13g2_mux2_1 _24002_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06007_),
    .X(_01775_));
 sg13g2_mux2_1 _24003_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(_06007_),
    .X(_01776_));
 sg13g2_nand2_1 _24004_ (.Y(_06013_),
    .A(_06005_),
    .B(_05864_));
 sg13g2_buf_2 _24005_ (.A(_06013_),
    .X(_06014_));
 sg13g2_buf_1 _24006_ (.A(_06014_),
    .X(_06015_));
 sg13g2_nand2_1 _24007_ (.Y(_06016_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(_06014_));
 sg13g2_o21ai_1 _24008_ (.B1(_06016_),
    .Y(_01777_),
    .A1(net616),
    .A2(net305));
 sg13g2_mux2_1 _24009_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net305),
    .X(_01778_));
 sg13g2_nand2_1 _24010_ (.Y(_06017_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(_06014_));
 sg13g2_o21ai_1 _24011_ (.B1(_06017_),
    .Y(_01779_),
    .A1(net549),
    .A2(net305));
 sg13g2_nand2_1 _24012_ (.Y(_06018_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(_06014_));
 sg13g2_o21ai_1 _24013_ (.B1(_06018_),
    .Y(_01780_),
    .A1(net618),
    .A2(net305));
 sg13g2_nand2_1 _24014_ (.Y(_06019_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .B(_06014_));
 sg13g2_o21ai_1 _24015_ (.B1(_06019_),
    .Y(_01781_),
    .A1(net617),
    .A2(net305));
 sg13g2_mux2_1 _24016_ (.A0(_05981_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .S(net305),
    .X(_01782_));
 sg13g2_mux2_1 _24017_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net305),
    .X(_01783_));
 sg13g2_mux2_1 _24018_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(net305),
    .X(_01784_));
 sg13g2_mux2_1 _24019_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(_06015_),
    .X(_01785_));
 sg13g2_mux2_1 _24020_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(_06015_),
    .X(_01786_));
 sg13g2_mux2_1 _24021_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06014_),
    .X(_01787_));
 sg13g2_mux2_1 _24022_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(_06014_),
    .X(_01788_));
 sg13g2_nand3_1 _24023_ (.B(_05827_),
    .C(net378),
    .A(_05872_),
    .Y(_06020_));
 sg13g2_buf_2 _24024_ (.A(_06020_),
    .X(_06021_));
 sg13g2_buf_1 _24025_ (.A(_06021_),
    .X(_06022_));
 sg13g2_nand2_1 _24026_ (.Y(_06023_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24027_ (.B1(_06023_),
    .Y(_01789_),
    .A1(net616),
    .A2(net261));
 sg13g2_mux2_1 _24028_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(net261),
    .X(_01790_));
 sg13g2_nand2_1 _24029_ (.Y(_06024_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24030_ (.B1(_06024_),
    .Y(_01791_),
    .A1(net549),
    .A2(net261));
 sg13g2_nand2_1 _24031_ (.Y(_06025_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24032_ (.B1(_06025_),
    .Y(_01792_),
    .A1(net618),
    .A2(_06022_));
 sg13g2_nand2_1 _24033_ (.Y(_06026_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24034_ (.B1(_06026_),
    .Y(_01793_),
    .A1(net617),
    .A2(net261));
 sg13g2_mux2_1 _24035_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .S(_06022_),
    .X(_01794_));
 sg13g2_mux2_1 _24036_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net261),
    .X(_01795_));
 sg13g2_mux2_1 _24037_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(net261),
    .X(_01796_));
 sg13g2_mux2_1 _24038_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net261),
    .X(_01797_));
 sg13g2_mux2_1 _24039_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net261),
    .X(_01798_));
 sg13g2_mux2_1 _24040_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(_06021_),
    .X(_01799_));
 sg13g2_mux2_1 _24041_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(_06021_),
    .X(_01800_));
 sg13g2_nand3_1 _24042_ (.B(_06005_),
    .C(net378),
    .A(_05872_),
    .Y(_06027_));
 sg13g2_buf_2 _24043_ (.A(_06027_),
    .X(_06028_));
 sg13g2_buf_1 _24044_ (.A(_06028_),
    .X(_06029_));
 sg13g2_nand2_1 _24045_ (.Y(_06030_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(_06028_));
 sg13g2_o21ai_1 _24046_ (.B1(_06030_),
    .Y(_01801_),
    .A1(_05993_),
    .A2(net260));
 sg13g2_mux2_1 _24047_ (.A0(_05998_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net260),
    .X(_01802_));
 sg13g2_nand2_1 _24048_ (.Y(_06031_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(_06028_));
 sg13g2_o21ai_1 _24049_ (.B1(_06031_),
    .Y(_01803_),
    .A1(_05999_),
    .A2(net260));
 sg13g2_nand2_1 _24050_ (.Y(_06032_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(_06028_));
 sg13g2_o21ai_1 _24051_ (.B1(_06032_),
    .Y(_01804_),
    .A1(_05977_),
    .A2(net260));
 sg13g2_nand2_1 _24052_ (.Y(_06033_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .B(_06028_));
 sg13g2_o21ai_1 _24053_ (.B1(_06033_),
    .Y(_01805_),
    .A1(net617),
    .A2(net260));
 sg13g2_mux2_1 _24054_ (.A0(_05981_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .S(net260),
    .X(_01806_));
 sg13g2_mux2_1 _24055_ (.A0(_05982_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net260),
    .X(_01807_));
 sg13g2_mux2_1 _24056_ (.A0(_05983_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(net260),
    .X(_01808_));
 sg13g2_mux2_1 _24057_ (.A0(_05984_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(_06029_),
    .X(_01809_));
 sg13g2_mux2_1 _24058_ (.A0(_05985_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(_06029_),
    .X(_01810_));
 sg13g2_mux2_1 _24059_ (.A0(_06003_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06028_),
    .X(_01811_));
 sg13g2_mux2_1 _24060_ (.A0(_06004_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(_06028_),
    .X(_01812_));
 sg13g2_nand3_1 _24061_ (.B(_06005_),
    .C(_05880_),
    .A(_05624_),
    .Y(_06034_));
 sg13g2_buf_2 _24062_ (.A(_06034_),
    .X(_06035_));
 sg13g2_buf_1 _24063_ (.A(_06035_),
    .X(_06036_));
 sg13g2_nand2_1 _24064_ (.Y(_06037_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(_06035_));
 sg13g2_o21ai_1 _24065_ (.B1(_06037_),
    .Y(_01813_),
    .A1(_05993_),
    .A2(net259));
 sg13g2_mux2_1 _24066_ (.A0(_05998_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net259),
    .X(_01814_));
 sg13g2_nand2_1 _24067_ (.Y(_06038_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(_06035_));
 sg13g2_o21ai_1 _24068_ (.B1(_06038_),
    .Y(_01815_),
    .A1(_05999_),
    .A2(net259));
 sg13g2_nand2_1 _24069_ (.Y(_06039_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(_06035_));
 sg13g2_o21ai_1 _24070_ (.B1(_06039_),
    .Y(_01816_),
    .A1(_05977_),
    .A2(net259));
 sg13g2_nand2_1 _24071_ (.Y(_06040_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .B(_06035_));
 sg13g2_o21ai_1 _24072_ (.B1(_06040_),
    .Y(_01817_),
    .A1(net617),
    .A2(net259));
 sg13g2_mux2_1 _24073_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S(net259),
    .X(_01818_));
 sg13g2_mux2_1 _24074_ (.A0(_05982_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net259),
    .X(_01819_));
 sg13g2_mux2_1 _24075_ (.A0(_05983_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(net259),
    .X(_01820_));
 sg13g2_mux2_1 _24076_ (.A0(_05984_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(_06036_),
    .X(_01821_));
 sg13g2_mux2_1 _24077_ (.A0(_05985_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(_06036_),
    .X(_01822_));
 sg13g2_mux2_1 _24078_ (.A0(_06003_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06035_),
    .X(_01823_));
 sg13g2_mux2_1 _24079_ (.A0(_06004_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(_06035_),
    .X(_01824_));
 sg13g2_nand3_1 _24080_ (.B(_05827_),
    .C(net378),
    .A(_05624_),
    .Y(_06041_));
 sg13g2_buf_2 _24081_ (.A(_06041_),
    .X(_06042_));
 sg13g2_buf_1 _24082_ (.A(_06042_),
    .X(_06043_));
 sg13g2_nand2_1 _24083_ (.Y(_06044_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(_06042_));
 sg13g2_o21ai_1 _24084_ (.B1(_06044_),
    .Y(_01825_),
    .A1(net616),
    .A2(net258));
 sg13g2_mux2_1 _24085_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net258),
    .X(_01826_));
 sg13g2_nand2_1 _24086_ (.Y(_06045_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(_06042_));
 sg13g2_o21ai_1 _24087_ (.B1(_06045_),
    .Y(_01827_),
    .A1(net549),
    .A2(net258));
 sg13g2_nand2_1 _24088_ (.Y(_06046_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(_06042_));
 sg13g2_o21ai_1 _24089_ (.B1(_06046_),
    .Y(_01828_),
    .A1(net618),
    .A2(_06043_));
 sg13g2_nand2_1 _24090_ (.Y(_06047_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .B(_06042_));
 sg13g2_o21ai_1 _24091_ (.B1(_06047_),
    .Y(_01829_),
    .A1(net617),
    .A2(net258));
 sg13g2_mux2_1 _24092_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S(_06043_),
    .X(_01830_));
 sg13g2_mux2_1 _24093_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net258),
    .X(_01831_));
 sg13g2_mux2_1 _24094_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(net258),
    .X(_01832_));
 sg13g2_mux2_1 _24095_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net258),
    .X(_01833_));
 sg13g2_mux2_1 _24096_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net258),
    .X(_01834_));
 sg13g2_mux2_1 _24097_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(_06042_),
    .X(_01835_));
 sg13g2_mux2_1 _24098_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06042_),
    .X(_01836_));
 sg13g2_nand2b_1 _24099_ (.Y(_06048_),
    .B(_05832_),
    .A_N(_05800_));
 sg13g2_buf_2 _24100_ (.A(_06048_),
    .X(_06049_));
 sg13g2_buf_1 _24101_ (.A(_06049_),
    .X(_06050_));
 sg13g2_nand2_1 _24102_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24103_ (.B1(_06051_),
    .Y(_01837_),
    .A1(net616),
    .A2(net216));
 sg13g2_mux2_1 _24104_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net216),
    .X(_01838_));
 sg13g2_nand2_1 _24105_ (.Y(_06052_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24106_ (.B1(_06052_),
    .Y(_01839_),
    .A1(net549),
    .A2(net216));
 sg13g2_nand2_1 _24107_ (.Y(_06053_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24108_ (.B1(_06053_),
    .Y(_01840_),
    .A1(net618),
    .A2(_06050_));
 sg13g2_nand2_1 _24109_ (.Y(_06054_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24110_ (.B1(_06054_),
    .Y(_01841_),
    .A1(_05979_),
    .A2(_06050_));
 sg13g2_mux2_1 _24111_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .S(net216),
    .X(_01842_));
 sg13g2_mux2_1 _24112_ (.A0(net802),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net216),
    .X(_01843_));
 sg13g2_mux2_1 _24113_ (.A0(net801),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net216),
    .X(_01844_));
 sg13g2_mux2_1 _24114_ (.A0(net800),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net216),
    .X(_01845_));
 sg13g2_mux2_1 _24115_ (.A0(net799),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(net216),
    .X(_01846_));
 sg13g2_mux2_1 _24116_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(_06049_),
    .X(_01847_));
 sg13g2_mux2_1 _24117_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(_06049_),
    .X(_01848_));
 sg13g2_nand2_1 _24118_ (.Y(_06055_),
    .A(_05805_),
    .B(net379));
 sg13g2_buf_2 _24119_ (.A(_06055_),
    .X(_06056_));
 sg13g2_buf_1 _24120_ (.A(_06056_),
    .X(_06057_));
 sg13g2_nand2_1 _24121_ (.Y(_06058_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(_06056_));
 sg13g2_o21ai_1 _24122_ (.B1(_06058_),
    .Y(_01849_),
    .A1(net616),
    .A2(_06057_));
 sg13g2_mux2_1 _24123_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net257),
    .X(_01850_));
 sg13g2_nand2_1 _24124_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(_06056_));
 sg13g2_o21ai_1 _24125_ (.B1(_06059_),
    .Y(_01851_),
    .A1(net549),
    .A2(_06057_));
 sg13g2_nand2_1 _24126_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(_06056_));
 sg13g2_o21ai_1 _24127_ (.B1(_06060_),
    .Y(_01852_),
    .A1(net716),
    .A2(net257));
 sg13g2_nand2_1 _24128_ (.Y(_06061_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .B(_06056_));
 sg13g2_o21ai_1 _24129_ (.B1(_06061_),
    .Y(_01853_),
    .A1(net715),
    .A2(net257));
 sg13g2_mux2_1 _24130_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .S(net257),
    .X(_01854_));
 sg13g2_mux2_1 _24131_ (.A0(net837),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net257),
    .X(_01855_));
 sg13g2_mux2_1 _24132_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net257),
    .X(_01856_));
 sg13g2_mux2_1 _24133_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net257),
    .X(_01857_));
 sg13g2_mux2_1 _24134_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net257),
    .X(_01858_));
 sg13g2_mux2_1 _24135_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(_06056_),
    .X(_01859_));
 sg13g2_mux2_1 _24136_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06056_),
    .X(_01860_));
 sg13g2_nand2_1 _24137_ (.Y(_06062_),
    .A(_05811_),
    .B(_05840_));
 sg13g2_buf_2 _24138_ (.A(_06062_),
    .X(_06063_));
 sg13g2_buf_1 _24139_ (.A(_06063_),
    .X(_06064_));
 sg13g2_nand2_1 _24140_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24141_ (.B1(_06065_),
    .Y(_01861_),
    .A1(net616),
    .A2(_06064_));
 sg13g2_mux2_1 _24142_ (.A0(net420),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net256),
    .X(_01862_));
 sg13g2_nand2_1 _24143_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24144_ (.B1(_06066_),
    .Y(_01863_),
    .A1(net549),
    .A2(_06064_));
 sg13g2_nand2_1 _24145_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24146_ (.B1(_06067_),
    .Y(_01864_),
    .A1(net716),
    .A2(net256));
 sg13g2_nand2_1 _24147_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24148_ (.B1(_06068_),
    .Y(_01865_),
    .A1(net715),
    .A2(net256));
 sg13g2_mux2_1 _24149_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .S(net256),
    .X(_01866_));
 sg13g2_mux2_1 _24150_ (.A0(net837),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net256),
    .X(_01867_));
 sg13g2_mux2_1 _24151_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net256),
    .X(_01868_));
 sg13g2_mux2_1 _24152_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net256),
    .X(_01869_));
 sg13g2_mux2_1 _24153_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(net256),
    .X(_01870_));
 sg13g2_mux2_1 _24154_ (.A0(net419),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(_06063_),
    .X(_01871_));
 sg13g2_mux2_1 _24155_ (.A0(net418),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06063_),
    .X(_01872_));
 sg13g2_nand2_1 _24156_ (.Y(_06069_),
    .A(_05816_),
    .B(net379));
 sg13g2_buf_2 _24157_ (.A(_06069_),
    .X(_06070_));
 sg13g2_buf_1 _24158_ (.A(_06070_),
    .X(_06071_));
 sg13g2_nand2_1 _24159_ (.Y(_06072_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24160_ (.B1(_06072_),
    .Y(_01873_),
    .A1(net708),
    .A2(net255));
 sg13g2_mux2_1 _24161_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net255),
    .X(_01874_));
 sg13g2_nand2_1 _24162_ (.Y(_06073_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24163_ (.B1(_06073_),
    .Y(_01875_),
    .A1(net679),
    .A2(_06071_));
 sg13g2_nand2_1 _24164_ (.Y(_06074_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24165_ (.B1(_06074_),
    .Y(_01876_),
    .A1(net716),
    .A2(net255));
 sg13g2_nand2_1 _24166_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24167_ (.B1(_06075_),
    .Y(_01877_),
    .A1(net715),
    .A2(_06071_));
 sg13g2_mux2_1 _24168_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S(net255),
    .X(_01878_));
 sg13g2_mux2_1 _24169_ (.A0(net837),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net255),
    .X(_01879_));
 sg13g2_mux2_1 _24170_ (.A0(net836),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net255),
    .X(_01880_));
 sg13g2_mux2_1 _24171_ (.A0(net835),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net255),
    .X(_01881_));
 sg13g2_mux2_1 _24172_ (.A0(net834),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(net255),
    .X(_01882_));
 sg13g2_mux2_1 _24173_ (.A0(net439),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(_06070_),
    .X(_01883_));
 sg13g2_mux2_1 _24174_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06070_),
    .X(_01884_));
 sg13g2_nand3_1 _24175_ (.B(_05888_),
    .C(net378),
    .A(_05683_),
    .Y(_06076_));
 sg13g2_buf_2 _24176_ (.A(_06076_),
    .X(_06077_));
 sg13g2_buf_1 _24177_ (.A(_06077_),
    .X(_06078_));
 sg13g2_nand2_1 _24178_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24179_ (.B1(_06079_),
    .Y(_01885_),
    .A1(net708),
    .A2(net254));
 sg13g2_mux2_1 _24180_ (.A0(_03353_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(net254),
    .X(_01886_));
 sg13g2_nand2_1 _24181_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24182_ (.B1(_06080_),
    .Y(_01887_),
    .A1(net679),
    .A2(_06078_));
 sg13g2_nand2_1 _24183_ (.Y(_06081_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24184_ (.B1(_06081_),
    .Y(_01888_),
    .A1(_02856_),
    .A2(net254));
 sg13g2_nand2_1 _24185_ (.Y(_06082_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24186_ (.B1(_06082_),
    .Y(_01889_),
    .A1(_02863_),
    .A2(_06078_));
 sg13g2_mux2_1 _24187_ (.A0(_02884_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .S(net254),
    .X(_01890_));
 sg13g2_mux2_1 _24188_ (.A0(_02885_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net254),
    .X(_01891_));
 sg13g2_mux2_1 _24189_ (.A0(_02886_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net254),
    .X(_01892_));
 sg13g2_mux2_1 _24190_ (.A0(_02887_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net254),
    .X(_01893_));
 sg13g2_mux2_1 _24191_ (.A0(_02888_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net254),
    .X(_01894_));
 sg13g2_mux2_1 _24192_ (.A0(_03363_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(_06077_),
    .X(_01895_));
 sg13g2_mux2_1 _24193_ (.A0(_03351_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06077_),
    .X(_01896_));
 sg13g2_nand3_1 _24194_ (.B(_05683_),
    .C(_05864_),
    .A(net817),
    .Y(_06083_));
 sg13g2_buf_2 _24195_ (.A(_06083_),
    .X(_06084_));
 sg13g2_buf_1 _24196_ (.A(_06084_),
    .X(_06085_));
 sg13g2_nand2_1 _24197_ (.Y(_06086_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(_06084_));
 sg13g2_o21ai_1 _24198_ (.B1(_06086_),
    .Y(_01897_),
    .A1(_03612_),
    .A2(net304));
 sg13g2_mux2_1 _24199_ (.A0(_03353_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(net304),
    .X(_01898_));
 sg13g2_nand2_1 _24200_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(_06084_));
 sg13g2_o21ai_1 _24201_ (.B1(_06087_),
    .Y(_01899_),
    .A1(_09220_),
    .A2(_06085_));
 sg13g2_nand2_1 _24202_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(_06084_));
 sg13g2_o21ai_1 _24203_ (.B1(_06088_),
    .Y(_01900_),
    .A1(net716),
    .A2(net304));
 sg13g2_nand2_1 _24204_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .B(_06084_));
 sg13g2_o21ai_1 _24205_ (.B1(_06089_),
    .Y(_01901_),
    .A1(_02863_),
    .A2(_06085_));
 sg13g2_mux2_1 _24206_ (.A0(_02884_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .S(net304),
    .X(_01902_));
 sg13g2_mux2_1 _24207_ (.A0(_02885_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net304),
    .X(_01903_));
 sg13g2_mux2_1 _24208_ (.A0(_02886_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net304),
    .X(_01904_));
 sg13g2_mux2_1 _24209_ (.A0(_02887_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net304),
    .X(_01905_));
 sg13g2_mux2_1 _24210_ (.A0(_02888_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net304),
    .X(_01906_));
 sg13g2_mux2_1 _24211_ (.A0(_03363_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(_06084_),
    .X(_01907_));
 sg13g2_mux2_1 _24212_ (.A0(_03351_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06084_),
    .X(_01908_));
 sg13g2_buf_1 _24213_ (.A(net565),
    .X(_06090_));
 sg13g2_mux2_1 _24214_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(net482),
    .S(_05661_),
    .X(_01909_));
 sg13g2_mux2_1 _24215_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net482),
    .S(_05675_),
    .X(_01910_));
 sg13g2_mux2_1 _24216_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net482),
    .S(_05680_),
    .X(_01911_));
 sg13g2_mux2_1 _24217_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net482),
    .S(_05687_),
    .X(_01912_));
 sg13g2_mux2_1 _24218_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net482),
    .S(_05693_),
    .X(_01913_));
 sg13g2_mux2_1 _24219_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06090_),
    .S(_05699_),
    .X(_01914_));
 sg13g2_mux2_1 _24220_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06090_),
    .S(_05702_),
    .X(_01915_));
 sg13g2_mux2_1 _24221_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net482),
    .S(_05709_),
    .X(_01916_));
 sg13g2_mux2_1 _24222_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net482),
    .S(_05714_),
    .X(_01917_));
 sg13g2_mux2_1 _24223_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net482),
    .S(_05721_),
    .X(_01918_));
 sg13g2_buf_1 _24224_ (.A(net565),
    .X(_06091_));
 sg13g2_mux2_1 _24225_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net481),
    .S(_05730_),
    .X(_01919_));
 sg13g2_mux2_1 _24226_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(net481),
    .S(_05735_),
    .X(_01920_));
 sg13g2_mux2_1 _24227_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net481),
    .S(_05740_),
    .X(_01921_));
 sg13g2_mux2_1 _24228_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net481),
    .S(_05744_),
    .X(_01922_));
 sg13g2_mux2_1 _24229_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net481),
    .S(_05747_),
    .X(_01923_));
 sg13g2_mux2_1 _24230_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net481),
    .S(_05752_),
    .X(_01924_));
 sg13g2_mux2_1 _24231_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net481),
    .S(_05756_),
    .X(_01925_));
 sg13g2_mux2_1 _24232_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(_06091_),
    .S(_05759_),
    .X(_01926_));
 sg13g2_mux2_1 _24233_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net481),
    .S(_05765_),
    .X(_01927_));
 sg13g2_mux2_1 _24234_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(_06091_),
    .S(_05771_),
    .X(_01928_));
 sg13g2_buf_1 _24235_ (.A(net565),
    .X(_06092_));
 sg13g2_mux2_1 _24236_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net480),
    .S(_05780_),
    .X(_01929_));
 sg13g2_mux2_1 _24237_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net480),
    .S(_05785_),
    .X(_01930_));
 sg13g2_mux2_1 _24238_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(net480),
    .S(_05788_),
    .X(_01931_));
 sg13g2_mux2_1 _24239_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net480),
    .S(_05792_),
    .X(_01932_));
 sg13g2_mux2_1 _24240_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net480),
    .S(_05795_),
    .X(_01933_));
 sg13g2_mux2_1 _24241_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(_06092_),
    .S(_05798_),
    .X(_01934_));
 sg13g2_mux2_1 _24242_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net480),
    .S(_05802_),
    .X(_01935_));
 sg13g2_mux2_1 _24243_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net480),
    .S(_05807_),
    .X(_01936_));
 sg13g2_mux2_1 _24244_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net480),
    .S(_05813_),
    .X(_01937_));
 sg13g2_mux2_1 _24245_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(_06092_),
    .S(_05818_),
    .X(_01938_));
 sg13g2_mux2_1 _24246_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(net565),
    .S(_05821_),
    .X(_01939_));
 sg13g2_mux2_1 _24247_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_03356_),
    .S(_05824_),
    .X(_01940_));
 sg13g2_nor2_2 _24248_ (.A(net1022),
    .B(_09022_),
    .Y(_06093_));
 sg13g2_nand3_1 _24249_ (.B(_09497_),
    .C(_06093_),
    .A(net956),
    .Y(_06094_));
 sg13g2_buf_1 _24250_ (.A(_06094_),
    .X(_06095_));
 sg13g2_nor2_1 _24251_ (.A(net1019),
    .B(net138),
    .Y(_06096_));
 sg13g2_buf_2 _24252_ (.A(_06096_),
    .X(_06097_));
 sg13g2_and3_1 _24253_ (.X(_06098_),
    .A(_05363_),
    .B(_04740_),
    .C(_06097_));
 sg13g2_buf_1 _24254_ (.A(_06098_),
    .X(_06099_));
 sg13g2_mux2_1 _24255_ (.A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net971),
    .S(_06099_),
    .X(_01957_));
 sg13g2_mux2_1 _24256_ (.A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net969),
    .S(_06099_),
    .X(_01958_));
 sg13g2_buf_1 _24257_ (.A(_09851_),
    .X(_06100_));
 sg13g2_mux2_1 _24258_ (.A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net929),
    .S(_06099_),
    .X(_01959_));
 sg13g2_mux2_1 _24259_ (.A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1005),
    .S(_06099_),
    .X(_01960_));
 sg13g2_nand3_1 _24260_ (.B(_04927_),
    .C(_06097_),
    .A(net822),
    .Y(_06101_));
 sg13g2_buf_2 _24261_ (.A(_06101_),
    .X(_06102_));
 sg13g2_nand2_1 _24262_ (.Y(_06103_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24263_ (.B1(_06103_),
    .Y(_01961_),
    .A1(net720),
    .A2(_06102_));
 sg13g2_mux2_1 _24264_ (.A0(net819),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06102_),
    .X(_01962_));
 sg13g2_mux2_1 _24265_ (.A0(net818),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06102_),
    .X(_01963_));
 sg13g2_nand2_1 _24266_ (.Y(_06104_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24267_ (.B1(_06104_),
    .Y(_01964_),
    .A1(net719),
    .A2(_06102_));
 sg13g2_nand2_1 _24268_ (.Y(_06105_),
    .A(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24269_ (.B1(_06105_),
    .Y(_01965_),
    .A1(net718),
    .A2(_06102_));
 sg13g2_nand2_1 _24270_ (.Y(_06106_),
    .A(_04723_),
    .B(_06097_));
 sg13g2_buf_1 _24271_ (.A(_06106_),
    .X(_06107_));
 sg13g2_nand2_1 _24272_ (.Y(_06108_),
    .A(_04722_),
    .B(_06107_));
 sg13g2_o21ai_1 _24273_ (.B1(_06108_),
    .Y(_01966_),
    .A1(_12245_),
    .A2(_06107_));
 sg13g2_buf_1 _24274_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06109_));
 sg13g2_mux2_1 _24275_ (.A0(_09820_),
    .A1(_06109_),
    .S(net79),
    .X(_01967_));
 sg13g2_mux2_1 _24276_ (.A0(net870),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(net79),
    .X(_01968_));
 sg13g2_nand2_1 _24277_ (.Y(_06110_),
    .A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .B(net79));
 sg13g2_o21ai_1 _24278_ (.B1(_06110_),
    .Y(_01969_),
    .A1(_12362_),
    .A2(net79));
 sg13g2_mux2_1 _24279_ (.A0(_05591_),
    .A1(_05360_),
    .S(net79),
    .X(_01970_));
 sg13g2_buf_1 _24280_ (.A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .X(_06111_));
 sg13g2_mux2_1 _24281_ (.A0(net818),
    .A1(_06111_),
    .S(net79),
    .X(_01971_));
 sg13g2_nand2_1 _24282_ (.Y(_06112_),
    .A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B(_06106_));
 sg13g2_o21ai_1 _24283_ (.B1(_06112_),
    .Y(_01972_),
    .A1(_12376_),
    .A2(net79));
 sg13g2_nand2_1 _24284_ (.Y(_06113_),
    .A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .B(_06106_));
 sg13g2_o21ai_1 _24285_ (.B1(_06113_),
    .Y(_01973_),
    .A1(net718),
    .A2(net79));
 sg13g2_and3_1 _24286_ (.X(_06114_),
    .A(net529),
    .B(net626),
    .C(_06097_));
 sg13g2_buf_4 _24287_ (.X(_06115_),
    .A(_06114_));
 sg13g2_mux2_1 _24288_ (.A0(_04710_),
    .A1(net821),
    .S(_06115_),
    .X(_01974_));
 sg13g2_mux2_1 _24289_ (.A0(_05151_),
    .A1(net871),
    .S(_06115_),
    .X(_01975_));
 sg13g2_mux2_1 _24290_ (.A0(_05217_),
    .A1(net870),
    .S(_06115_),
    .X(_01976_));
 sg13g2_buf_1 _24291_ (.A(net1078),
    .X(_06116_));
 sg13g2_mux2_1 _24292_ (.A0(_05279_),
    .A1(net928),
    .S(_06115_),
    .X(_01977_));
 sg13g2_mux2_1 _24293_ (.A0(_05368_),
    .A1(_11801_),
    .S(_06115_),
    .X(_01978_));
 sg13g2_mux2_1 _24294_ (.A0(_05425_),
    .A1(_11806_),
    .S(_06115_),
    .X(_01979_));
 sg13g2_mux2_1 _24295_ (.A0(_05484_),
    .A1(net929),
    .S(_06115_),
    .X(_01980_));
 sg13g2_mux2_1 _24296_ (.A0(_04849_),
    .A1(_09857_),
    .S(_06115_),
    .X(_01981_));
 sg13g2_nand3_1 _24297_ (.B(net626),
    .C(_06097_),
    .A(net530),
    .Y(_06117_));
 sg13g2_buf_1 _24298_ (.A(_06117_),
    .X(_06118_));
 sg13g2_buf_1 _24299_ (.A(_06118_),
    .X(_06119_));
 sg13g2_nand2_1 _24300_ (.Y(_06120_),
    .A(_04711_),
    .B(net73));
 sg13g2_o21ai_1 _24301_ (.B1(_06120_),
    .Y(_01982_),
    .A1(_12245_),
    .A2(net73));
 sg13g2_buf_1 _24302_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06121_));
 sg13g2_mux2_1 _24303_ (.A0(_09820_),
    .A1(_06121_),
    .S(net73),
    .X(_01983_));
 sg13g2_mux2_1 _24304_ (.A0(net870),
    .A1(\cpu.gpio.r_src_io[6][2] ),
    .S(_06119_),
    .X(_01984_));
 sg13g2_nand2_1 _24305_ (.Y(_06122_),
    .A(\cpu.gpio.r_src_io[6][3] ),
    .B(net73));
 sg13g2_o21ai_1 _24306_ (.B1(_06122_),
    .Y(_01985_),
    .A1(net720),
    .A2(net73));
 sg13g2_mux2_1 _24307_ (.A0(net819),
    .A1(_05369_),
    .S(_06119_),
    .X(_01986_));
 sg13g2_buf_1 _24308_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06123_));
 sg13g2_mux2_1 _24309_ (.A0(net818),
    .A1(_06123_),
    .S(net73),
    .X(_01987_));
 sg13g2_nand2_1 _24310_ (.Y(_06124_),
    .A(\cpu.gpio.r_src_io[7][2] ),
    .B(_06118_));
 sg13g2_o21ai_1 _24311_ (.B1(_06124_),
    .Y(_01988_),
    .A1(net719),
    .A2(net73));
 sg13g2_nand2_1 _24312_ (.Y(_06125_),
    .A(\cpu.gpio.r_src_io[7][3] ),
    .B(_06118_));
 sg13g2_o21ai_1 _24313_ (.B1(_06125_),
    .Y(_01989_),
    .A1(net718),
    .A2(net73));
 sg13g2_and3_1 _24314_ (.X(_06126_),
    .A(net635),
    .B(_04755_),
    .C(_06097_));
 sg13g2_buf_1 _24315_ (.A(_06126_),
    .X(_06127_));
 sg13g2_mux2_1 _24316_ (.A0(_05372_),
    .A1(net971),
    .S(_06127_),
    .X(_01990_));
 sg13g2_buf_1 _24317_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06128_));
 sg13g2_mux2_1 _24318_ (.A0(_06128_),
    .A1(_11806_),
    .S(_06127_),
    .X(_01991_));
 sg13g2_mux2_1 _24319_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(net929),
    .S(_06127_),
    .X(_01992_));
 sg13g2_mux2_1 _24320_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net1005),
    .S(_06127_),
    .X(_01993_));
 sg13g2_nand2_1 _24321_ (.Y(_06129_),
    .A(_04705_),
    .B(_06097_));
 sg13g2_buf_1 _24322_ (.A(_06129_),
    .X(_06130_));
 sg13g2_nand2_1 _24323_ (.Y(_06131_),
    .A(_04706_),
    .B(net78));
 sg13g2_o21ai_1 _24324_ (.B1(_06131_),
    .Y(_01994_),
    .A1(net721),
    .A2(_06130_));
 sg13g2_buf_1 _24325_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06132_));
 sg13g2_mux2_1 _24326_ (.A0(net871),
    .A1(_06132_),
    .S(_06130_),
    .X(_01995_));
 sg13g2_mux2_1 _24327_ (.A0(_09827_),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(net78),
    .X(_01996_));
 sg13g2_nand2_1 _24328_ (.Y(_06133_),
    .A(\cpu.gpio.r_src_o[4][3] ),
    .B(net78));
 sg13g2_o21ai_1 _24329_ (.B1(_06133_),
    .Y(_01997_),
    .A1(_11716_),
    .A2(net78));
 sg13g2_mux2_1 _24330_ (.A0(net819),
    .A1(_05366_),
    .S(net78),
    .X(_01998_));
 sg13g2_buf_1 _24331_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06134_));
 sg13g2_mux2_1 _24332_ (.A0(_05592_),
    .A1(_06134_),
    .S(net78),
    .X(_01999_));
 sg13g2_nand2_1 _24333_ (.Y(_06135_),
    .A(\cpu.gpio.r_src_o[5][2] ),
    .B(_06129_));
 sg13g2_o21ai_1 _24334_ (.B1(_06135_),
    .Y(_02000_),
    .A1(net845),
    .A2(net78));
 sg13g2_nand2_1 _24335_ (.Y(_06136_),
    .A(\cpu.gpio.r_src_o[5][3] ),
    .B(_06129_));
 sg13g2_o21ai_1 _24336_ (.B1(_06136_),
    .Y(_02001_),
    .A1(net718),
    .A2(net78));
 sg13g2_nand2_1 _24337_ (.Y(_06137_),
    .A(_04719_),
    .B(_06097_));
 sg13g2_buf_2 _24338_ (.A(_06137_),
    .X(_06138_));
 sg13g2_mux2_1 _24339_ (.A0(net819),
    .A1(_05371_),
    .S(_06138_),
    .X(_02006_));
 sg13g2_buf_1 _24340_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06139_));
 sg13g2_mux2_1 _24341_ (.A0(_05592_),
    .A1(_06139_),
    .S(_06138_),
    .X(_02007_));
 sg13g2_nand2_1 _24342_ (.Y(_06140_),
    .A(\cpu.gpio.r_src_o[7][2] ),
    .B(_06138_));
 sg13g2_o21ai_1 _24343_ (.B1(_06140_),
    .Y(_02008_),
    .A1(net845),
    .A2(_06138_));
 sg13g2_nand2_1 _24344_ (.Y(_06141_),
    .A(\cpu.gpio.r_src_o[7][3] ),
    .B(_06138_));
 sg13g2_o21ai_1 _24345_ (.B1(_06141_),
    .Y(_02009_),
    .A1(_11755_),
    .A2(_06138_));
 sg13g2_buf_1 _24346_ (.A(_12162_),
    .X(_06142_));
 sg13g2_and2_1 _24347_ (.A(net701),
    .B(_08165_),
    .X(_06143_));
 sg13g2_buf_4 _24348_ (.X(_06144_),
    .A(_06143_));
 sg13g2_buf_1 _24349_ (.A(_00253_),
    .X(_06145_));
 sg13g2_nor2_1 _24350_ (.A(\cpu.icache.r_offset[2] ),
    .B(_06145_),
    .Y(_06146_));
 sg13g2_buf_2 _24351_ (.A(_06146_),
    .X(_06147_));
 sg13g2_buf_1 _24352_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06148_));
 sg13g2_buf_1 _24353_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06149_));
 sg13g2_nor2b_1 _24354_ (.A(_06148_),
    .B_N(_06149_),
    .Y(_06150_));
 sg13g2_buf_1 _24355_ (.A(_06150_),
    .X(_06151_));
 sg13g2_and2_1 _24356_ (.A(_06147_),
    .B(_06151_),
    .X(_06152_));
 sg13g2_buf_2 _24357_ (.A(_06152_),
    .X(_06153_));
 sg13g2_nand2_2 _24358_ (.Y(_06154_),
    .A(_06144_),
    .B(_06153_));
 sg13g2_mux2_1 _24359_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06154_),
    .X(_02013_));
 sg13g2_buf_1 _24360_ (.A(net957),
    .X(_06155_));
 sg13g2_inv_1 _24361_ (.Y(_06156_),
    .A(_00254_));
 sg13g2_nand2_1 _24362_ (.Y(_06157_),
    .A(_06148_),
    .B(_06149_));
 sg13g2_buf_2 _24363_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nor3_2 _24364_ (.A(_06145_),
    .B(_06156_),
    .C(_06158_),
    .Y(_06159_));
 sg13g2_nand2_2 _24365_ (.Y(_06160_),
    .A(_06144_),
    .B(_06159_));
 sg13g2_mux2_1 _24366_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06160_),
    .X(_02014_));
 sg13g2_buf_1 _24367_ (.A(_12185_),
    .X(_06161_));
 sg13g2_mux2_1 _24368_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06160_),
    .X(_02015_));
 sg13g2_nor2b_1 _24369_ (.A(_06149_),
    .B_N(_06148_),
    .Y(_06162_));
 sg13g2_buf_1 _24370_ (.A(_06162_),
    .X(_06163_));
 sg13g2_and2_1 _24371_ (.A(_06147_),
    .B(_06163_),
    .X(_06164_));
 sg13g2_buf_2 _24372_ (.A(_06164_),
    .X(_06165_));
 sg13g2_nand2_2 _24373_ (.Y(_06166_),
    .A(_06144_),
    .B(_06165_));
 sg13g2_mux2_1 _24374_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06166_),
    .X(_02016_));
 sg13g2_buf_1 _24375_ (.A(net958),
    .X(_06167_));
 sg13g2_mux2_1 _24376_ (.A0(_06167_),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06166_),
    .X(_02017_));
 sg13g2_mux2_1 _24377_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06166_),
    .X(_02018_));
 sg13g2_mux2_1 _24378_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06166_),
    .X(_02019_));
 sg13g2_nor2_1 _24379_ (.A(_06145_),
    .B(_00254_),
    .Y(_06168_));
 sg13g2_buf_2 _24380_ (.A(_06168_),
    .X(_06169_));
 sg13g2_and2_1 _24381_ (.A(_06151_),
    .B(_06169_),
    .X(_06170_));
 sg13g2_buf_2 _24382_ (.A(_06170_),
    .X(_06171_));
 sg13g2_nand2_2 _24383_ (.Y(_06172_),
    .A(_06144_),
    .B(_06171_));
 sg13g2_mux2_1 _24384_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06172_),
    .X(_02020_));
 sg13g2_mux2_1 _24385_ (.A0(_06167_),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06172_),
    .X(_02021_));
 sg13g2_mux2_1 _24386_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06172_),
    .X(_02022_));
 sg13g2_mux2_1 _24387_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06172_),
    .X(_02023_));
 sg13g2_mux2_1 _24388_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06154_),
    .X(_02024_));
 sg13g2_nor2_2 _24389_ (.A(_06148_),
    .B(_06149_),
    .Y(_06173_));
 sg13g2_and2_1 _24390_ (.A(_06169_),
    .B(_06173_),
    .X(_06174_));
 sg13g2_buf_2 _24391_ (.A(_06174_),
    .X(_06175_));
 sg13g2_nand2_2 _24392_ (.Y(_06176_),
    .A(_06144_),
    .B(_06175_));
 sg13g2_mux2_1 _24393_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06176_),
    .X(_02025_));
 sg13g2_mux2_1 _24394_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06176_),
    .X(_02026_));
 sg13g2_mux2_1 _24395_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06176_),
    .X(_02027_));
 sg13g2_mux2_1 _24396_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06176_),
    .X(_02028_));
 sg13g2_inv_1 _24397_ (.Y(_06177_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_2 _24398_ (.A(_00254_),
    .B(_06177_),
    .C(_06158_),
    .Y(_06178_));
 sg13g2_nand2_1 _24399_ (.Y(_06179_),
    .A(_06144_),
    .B(_06178_));
 sg13g2_buf_1 _24400_ (.A(_06179_),
    .X(_06180_));
 sg13g2_buf_1 _24401_ (.A(_06180_),
    .X(_06181_));
 sg13g2_mux2_1 _24402_ (.A0(_06142_),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(_06181_),
    .X(_02029_));
 sg13g2_mux2_1 _24403_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(_06181_),
    .X(_02030_));
 sg13g2_mux2_1 _24404_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net346),
    .X(_02031_));
 sg13g2_buf_1 _24405_ (.A(_06180_),
    .X(_06182_));
 sg13g2_mux2_1 _24406_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net345),
    .X(_02032_));
 sg13g2_and2_1 _24407_ (.A(_06163_),
    .B(_06169_),
    .X(_06183_));
 sg13g2_buf_2 _24408_ (.A(_06183_),
    .X(_06184_));
 sg13g2_nand2_2 _24409_ (.Y(_06185_),
    .A(_06144_),
    .B(_06184_));
 sg13g2_mux2_1 _24410_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06185_),
    .X(_02033_));
 sg13g2_mux2_1 _24411_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06185_),
    .X(_02034_));
 sg13g2_mux2_1 _24412_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06154_),
    .X(_02035_));
 sg13g2_mux2_1 _24413_ (.A0(_06155_),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06185_),
    .X(_02036_));
 sg13g2_mux2_1 _24414_ (.A0(_06161_),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06185_),
    .X(_02037_));
 sg13g2_mux2_1 _24415_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06154_),
    .X(_02038_));
 sg13g2_and2_1 _24416_ (.A(_06147_),
    .B(_06173_),
    .X(_06186_));
 sg13g2_buf_2 _24417_ (.A(_06186_),
    .X(_06187_));
 sg13g2_nand2_2 _24418_ (.Y(_06188_),
    .A(_06144_),
    .B(_06187_));
 sg13g2_mux2_1 _24419_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06188_),
    .X(_02039_));
 sg13g2_mux2_1 _24420_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06188_),
    .X(_02040_));
 sg13g2_mux2_1 _24421_ (.A0(net797),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06188_),
    .X(_02041_));
 sg13g2_mux2_1 _24422_ (.A0(net796),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06188_),
    .X(_02042_));
 sg13g2_mux2_1 _24423_ (.A0(net798),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06160_),
    .X(_02043_));
 sg13g2_mux2_1 _24424_ (.A0(net795),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06160_),
    .X(_02044_));
 sg13g2_buf_1 _24425_ (.A(_12162_),
    .X(_06189_));
 sg13g2_nand2_1 _24426_ (.Y(_06190_),
    .A(_08093_),
    .B(net694));
 sg13g2_buf_4 _24427_ (.X(_06191_),
    .A(_06190_));
 sg13g2_nand2_2 _24428_ (.Y(_06192_),
    .A(_06147_),
    .B(_06151_));
 sg13g2_nor2_2 _24429_ (.A(_06191_),
    .B(_06192_),
    .Y(_06193_));
 sg13g2_mux2_1 _24430_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net794),
    .S(_06193_),
    .X(_02045_));
 sg13g2_buf_1 _24431_ (.A(net957),
    .X(_06194_));
 sg13g2_or3_1 _24432_ (.A(_06145_),
    .B(_06156_),
    .C(_06158_),
    .X(_06195_));
 sg13g2_buf_2 _24433_ (.A(_06195_),
    .X(_06196_));
 sg13g2_nor2_2 _24434_ (.A(_06191_),
    .B(_06196_),
    .Y(_06197_));
 sg13g2_mux2_1 _24435_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net793),
    .S(_06197_),
    .X(_02046_));
 sg13g2_buf_1 _24436_ (.A(net1057),
    .X(_06198_));
 sg13g2_mux2_1 _24437_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net927),
    .S(_06197_),
    .X(_02047_));
 sg13g2_buf_1 _24438_ (.A(_12162_),
    .X(_06199_));
 sg13g2_nand2_2 _24439_ (.Y(_06200_),
    .A(_06147_),
    .B(_06163_));
 sg13g2_nor2_2 _24440_ (.A(_06191_),
    .B(_06200_),
    .Y(_06201_));
 sg13g2_mux2_1 _24441_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net792),
    .S(_06201_),
    .X(_02048_));
 sg13g2_buf_1 _24442_ (.A(net958),
    .X(_06202_));
 sg13g2_mux2_1 _24443_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net791),
    .S(_06201_),
    .X(_02049_));
 sg13g2_buf_1 _24444_ (.A(net957),
    .X(_06203_));
 sg13g2_mux2_1 _24445_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(_06203_),
    .S(_06201_),
    .X(_02050_));
 sg13g2_buf_1 _24446_ (.A(net1057),
    .X(_06204_));
 sg13g2_mux2_1 _24447_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(_06204_),
    .S(_06201_),
    .X(_02051_));
 sg13g2_nand2_2 _24448_ (.Y(_06205_),
    .A(_06151_),
    .B(_06169_));
 sg13g2_nor2_2 _24449_ (.A(_06191_),
    .B(_06205_),
    .Y(_06206_));
 sg13g2_mux2_1 _24450_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net792),
    .S(_06206_),
    .X(_02052_));
 sg13g2_buf_1 _24451_ (.A(_12469_),
    .X(_06207_));
 sg13g2_mux2_1 _24452_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net789),
    .S(_06206_),
    .X(_02053_));
 sg13g2_mux2_1 _24453_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net790),
    .S(_06206_),
    .X(_02054_));
 sg13g2_mux2_1 _24454_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net926),
    .S(_06206_),
    .X(_02055_));
 sg13g2_mux2_1 _24455_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net789),
    .S(_06193_),
    .X(_02056_));
 sg13g2_nand2_2 _24456_ (.Y(_06208_),
    .A(_06169_),
    .B(_06173_));
 sg13g2_nor2_2 _24457_ (.A(_06191_),
    .B(_06208_),
    .Y(_06209_));
 sg13g2_mux2_1 _24458_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net792),
    .S(_06209_),
    .X(_02057_));
 sg13g2_mux2_1 _24459_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net789),
    .S(_06209_),
    .X(_02058_));
 sg13g2_mux2_1 _24460_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net790),
    .S(_06209_),
    .X(_02059_));
 sg13g2_mux2_1 _24461_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net926),
    .S(_06209_),
    .X(_02060_));
 sg13g2_nand4_1 _24462_ (.B(_06149_),
    .C(_06156_),
    .A(_06148_),
    .Y(_06210_),
    .D(\cpu.i_wstrobe_d ));
 sg13g2_buf_1 _24463_ (.A(_06210_),
    .X(_06211_));
 sg13g2_nor2_1 _24464_ (.A(_06191_),
    .B(_06211_),
    .Y(_06212_));
 sg13g2_buf_2 _24465_ (.A(_06212_),
    .X(_06213_));
 sg13g2_mux2_1 _24466_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net792),
    .S(_06213_),
    .X(_02061_));
 sg13g2_mux2_1 _24467_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net789),
    .S(_06213_),
    .X(_02062_));
 sg13g2_mux2_1 _24468_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(net790),
    .S(_06213_),
    .X(_02063_));
 sg13g2_mux2_1 _24469_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(_06204_),
    .S(_06213_),
    .X(_02064_));
 sg13g2_nand2_2 _24470_ (.Y(_06214_),
    .A(_06163_),
    .B(_06169_));
 sg13g2_nor2_2 _24471_ (.A(_06191_),
    .B(_06214_),
    .Y(_06215_));
 sg13g2_mux2_1 _24472_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net792),
    .S(_06215_),
    .X(_02065_));
 sg13g2_mux2_1 _24473_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net789),
    .S(_06215_),
    .X(_02066_));
 sg13g2_mux2_1 _24474_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net790),
    .S(_06193_),
    .X(_02067_));
 sg13g2_mux2_1 _24475_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(_06203_),
    .S(_06215_),
    .X(_02068_));
 sg13g2_mux2_1 _24476_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net926),
    .S(_06215_),
    .X(_02069_));
 sg13g2_mux2_1 _24477_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net926),
    .S(_06193_),
    .X(_02070_));
 sg13g2_nand2_2 _24478_ (.Y(_06216_),
    .A(_06147_),
    .B(_06173_));
 sg13g2_nor2_2 _24479_ (.A(_06191_),
    .B(_06216_),
    .Y(_06217_));
 sg13g2_mux2_1 _24480_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net792),
    .S(_06217_),
    .X(_02071_));
 sg13g2_mux2_1 _24481_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net789),
    .S(_06217_),
    .X(_02072_));
 sg13g2_mux2_1 _24482_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net790),
    .S(_06217_),
    .X(_02073_));
 sg13g2_mux2_1 _24483_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net926),
    .S(_06217_),
    .X(_02074_));
 sg13g2_mux2_1 _24484_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(_06199_),
    .S(_06197_),
    .X(_02075_));
 sg13g2_mux2_1 _24485_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(net789),
    .S(_06197_),
    .X(_02076_));
 sg13g2_nand2_1 _24486_ (.Y(_06218_),
    .A(_08093_),
    .B(_08117_));
 sg13g2_buf_4 _24487_ (.X(_06219_),
    .A(_06218_));
 sg13g2_nor2_2 _24488_ (.A(_06219_),
    .B(_06192_),
    .Y(_06220_));
 sg13g2_mux2_1 _24489_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(net792),
    .S(_06220_),
    .X(_02077_));
 sg13g2_nor2_2 _24490_ (.A(_06219_),
    .B(_06196_),
    .Y(_06221_));
 sg13g2_mux2_1 _24491_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net790),
    .S(_06221_),
    .X(_02078_));
 sg13g2_mux2_1 _24492_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(net926),
    .S(_06221_),
    .X(_02079_));
 sg13g2_nor2_2 _24493_ (.A(_06219_),
    .B(_06200_),
    .Y(_06222_));
 sg13g2_mux2_1 _24494_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net792),
    .S(_06222_),
    .X(_02080_));
 sg13g2_mux2_1 _24495_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(_06207_),
    .S(_06222_),
    .X(_02081_));
 sg13g2_mux2_1 _24496_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net790),
    .S(_06222_),
    .X(_02082_));
 sg13g2_mux2_1 _24497_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net926),
    .S(_06222_),
    .X(_02083_));
 sg13g2_nor2_2 _24498_ (.A(_06219_),
    .B(_06205_),
    .Y(_06223_));
 sg13g2_mux2_1 _24499_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(_06199_),
    .S(_06223_),
    .X(_02084_));
 sg13g2_mux2_1 _24500_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(_06207_),
    .S(_06223_),
    .X(_02085_));
 sg13g2_mux2_1 _24501_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net790),
    .S(_06223_),
    .X(_02086_));
 sg13g2_mux2_1 _24502_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net926),
    .S(_06223_),
    .X(_02087_));
 sg13g2_mux2_1 _24503_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net789),
    .S(_06220_),
    .X(_02088_));
 sg13g2_buf_1 _24504_ (.A(_12162_),
    .X(_06224_));
 sg13g2_nor2_2 _24505_ (.A(_06219_),
    .B(_06208_),
    .Y(_06225_));
 sg13g2_mux2_1 _24506_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net788),
    .S(_06225_),
    .X(_02089_));
 sg13g2_buf_1 _24507_ (.A(_11743_),
    .X(_06226_));
 sg13g2_mux2_1 _24508_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net925),
    .S(_06225_),
    .X(_02090_));
 sg13g2_buf_1 _24509_ (.A(net957),
    .X(_06227_));
 sg13g2_mux2_1 _24510_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net787),
    .S(_06225_),
    .X(_02091_));
 sg13g2_buf_1 _24511_ (.A(_11833_),
    .X(_06228_));
 sg13g2_mux2_1 _24512_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net924),
    .S(_06225_),
    .X(_02092_));
 sg13g2_nor2_1 _24513_ (.A(_06219_),
    .B(_06211_),
    .Y(_06229_));
 sg13g2_buf_2 _24514_ (.A(_06229_),
    .X(_06230_));
 sg13g2_mux2_1 _24515_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net788),
    .S(_06230_),
    .X(_02093_));
 sg13g2_mux2_1 _24516_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net925),
    .S(_06230_),
    .X(_02094_));
 sg13g2_mux2_1 _24517_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net787),
    .S(_06230_),
    .X(_02095_));
 sg13g2_mux2_1 _24518_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net924),
    .S(_06230_),
    .X(_02096_));
 sg13g2_nor2_2 _24519_ (.A(_06219_),
    .B(_06214_),
    .Y(_06231_));
 sg13g2_mux2_1 _24520_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net788),
    .S(_06231_),
    .X(_02097_));
 sg13g2_mux2_1 _24521_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net925),
    .S(_06231_),
    .X(_02098_));
 sg13g2_mux2_1 _24522_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net787),
    .S(_06220_),
    .X(_02099_));
 sg13g2_mux2_1 _24523_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net787),
    .S(_06231_),
    .X(_02100_));
 sg13g2_mux2_1 _24524_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net924),
    .S(_06231_),
    .X(_02101_));
 sg13g2_mux2_1 _24525_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net924),
    .S(_06220_),
    .X(_02102_));
 sg13g2_nor2_2 _24526_ (.A(_06219_),
    .B(_06216_),
    .Y(_06232_));
 sg13g2_mux2_1 _24527_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(_06224_),
    .S(_06232_),
    .X(_02103_));
 sg13g2_mux2_1 _24528_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net925),
    .S(_06232_),
    .X(_02104_));
 sg13g2_mux2_1 _24529_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net787),
    .S(_06232_),
    .X(_02105_));
 sg13g2_mux2_1 _24530_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net924),
    .S(_06232_),
    .X(_02106_));
 sg13g2_mux2_1 _24531_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net788),
    .S(_06221_),
    .X(_02107_));
 sg13g2_mux2_1 _24532_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net925),
    .S(_06221_),
    .X(_02108_));
 sg13g2_nand2_2 _24533_ (.Y(_06233_),
    .A(net473),
    .B(_06153_));
 sg13g2_mux2_1 _24534_ (.A0(net798),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06233_),
    .X(_02109_));
 sg13g2_and2_1 _24535_ (.A(net473),
    .B(_06159_),
    .X(_06234_));
 sg13g2_buf_1 _24536_ (.A(_06234_),
    .X(_06235_));
 sg13g2_mux2_1 _24537_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net787),
    .S(_06235_),
    .X(_02110_));
 sg13g2_mux2_1 _24538_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net924),
    .S(_06235_),
    .X(_02111_));
 sg13g2_nand2_2 _24539_ (.Y(_06236_),
    .A(net473),
    .B(_06165_));
 sg13g2_mux2_1 _24540_ (.A0(_06142_),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06236_),
    .X(_02112_));
 sg13g2_mux2_1 _24541_ (.A0(net795),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06236_),
    .X(_02113_));
 sg13g2_mux2_1 _24542_ (.A0(net797),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06236_),
    .X(_02114_));
 sg13g2_mux2_1 _24543_ (.A0(_06161_),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06236_),
    .X(_02115_));
 sg13g2_buf_1 _24544_ (.A(_12162_),
    .X(_06237_));
 sg13g2_nand2_2 _24545_ (.Y(_06238_),
    .A(net473),
    .B(_06171_));
 sg13g2_mux2_1 _24546_ (.A0(net786),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06238_),
    .X(_02116_));
 sg13g2_mux2_1 _24547_ (.A0(net795),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06238_),
    .X(_02117_));
 sg13g2_mux2_1 _24548_ (.A0(_06155_),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06238_),
    .X(_02118_));
 sg13g2_mux2_1 _24549_ (.A0(net796),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06238_),
    .X(_02119_));
 sg13g2_buf_1 _24550_ (.A(_12469_),
    .X(_06239_));
 sg13g2_mux2_1 _24551_ (.A0(net785),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06233_),
    .X(_02120_));
 sg13g2_nand2_2 _24552_ (.Y(_06240_),
    .A(_08157_),
    .B(_06175_));
 sg13g2_mux2_1 _24553_ (.A0(net786),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06240_),
    .X(_02121_));
 sg13g2_mux2_1 _24554_ (.A0(net785),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06240_),
    .X(_02122_));
 sg13g2_buf_1 _24555_ (.A(_12473_),
    .X(_06241_));
 sg13g2_mux2_1 _24556_ (.A0(net784),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06240_),
    .X(_02123_));
 sg13g2_buf_1 _24557_ (.A(_12185_),
    .X(_06242_));
 sg13g2_mux2_1 _24558_ (.A0(net783),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06240_),
    .X(_02124_));
 sg13g2_nand2_1 _24559_ (.Y(_06243_),
    .A(net473),
    .B(_06178_));
 sg13g2_buf_1 _24560_ (.A(_06243_),
    .X(_06244_));
 sg13g2_buf_1 _24561_ (.A(_06244_),
    .X(_06245_));
 sg13g2_mux2_1 _24562_ (.A0(net786),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net303),
    .X(_02125_));
 sg13g2_mux2_1 _24563_ (.A0(net785),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net303),
    .X(_02126_));
 sg13g2_mux2_1 _24564_ (.A0(net784),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net303),
    .X(_02127_));
 sg13g2_buf_1 _24565_ (.A(_06244_),
    .X(_06246_));
 sg13g2_mux2_1 _24566_ (.A0(net783),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(_06246_),
    .X(_02128_));
 sg13g2_nand2_2 _24567_ (.Y(_06247_),
    .A(_08157_),
    .B(_06184_));
 sg13g2_mux2_1 _24568_ (.A0(net786),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06247_),
    .X(_02129_));
 sg13g2_mux2_1 _24569_ (.A0(net785),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06247_),
    .X(_02130_));
 sg13g2_mux2_1 _24570_ (.A0(net784),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06233_),
    .X(_02131_));
 sg13g2_mux2_1 _24571_ (.A0(net784),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06247_),
    .X(_02132_));
 sg13g2_mux2_1 _24572_ (.A0(net783),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06247_),
    .X(_02133_));
 sg13g2_mux2_1 _24573_ (.A0(net783),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06233_),
    .X(_02134_));
 sg13g2_nand2_2 _24574_ (.Y(_06248_),
    .A(net473),
    .B(_06187_));
 sg13g2_mux2_1 _24575_ (.A0(net786),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06248_),
    .X(_02135_));
 sg13g2_mux2_1 _24576_ (.A0(net785),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06248_),
    .X(_02136_));
 sg13g2_mux2_1 _24577_ (.A0(net784),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06248_),
    .X(_02137_));
 sg13g2_mux2_1 _24578_ (.A0(net783),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06248_),
    .X(_02138_));
 sg13g2_mux2_1 _24579_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net788),
    .S(_06235_),
    .X(_02139_));
 sg13g2_mux2_1 _24580_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(_06226_),
    .S(_06235_),
    .X(_02140_));
 sg13g2_nand2_2 _24581_ (.Y(_06249_),
    .A(net699),
    .B(_06153_));
 sg13g2_mux2_1 _24582_ (.A0(net786),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06249_),
    .X(_02141_));
 sg13g2_and2_1 _24583_ (.A(net699),
    .B(_06159_),
    .X(_06250_));
 sg13g2_buf_1 _24584_ (.A(_06250_),
    .X(_06251_));
 sg13g2_mux2_1 _24585_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(_06227_),
    .S(_06251_),
    .X(_02142_));
 sg13g2_mux2_1 _24586_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net924),
    .S(_06251_),
    .X(_02143_));
 sg13g2_nand2_2 _24587_ (.Y(_06252_),
    .A(net699),
    .B(_06165_));
 sg13g2_mux2_1 _24588_ (.A0(net786),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06252_),
    .X(_02144_));
 sg13g2_mux2_1 _24589_ (.A0(net785),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06252_),
    .X(_02145_));
 sg13g2_mux2_1 _24590_ (.A0(net784),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06252_),
    .X(_02146_));
 sg13g2_mux2_1 _24591_ (.A0(_06242_),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06252_),
    .X(_02147_));
 sg13g2_nand2_2 _24592_ (.Y(_06253_),
    .A(net699),
    .B(_06171_));
 sg13g2_mux2_1 _24593_ (.A0(_06237_),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06253_),
    .X(_02148_));
 sg13g2_mux2_1 _24594_ (.A0(_06239_),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06253_),
    .X(_02149_));
 sg13g2_mux2_1 _24595_ (.A0(_06241_),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06253_),
    .X(_02150_));
 sg13g2_mux2_1 _24596_ (.A0(_06242_),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06253_),
    .X(_02151_));
 sg13g2_mux2_1 _24597_ (.A0(net785),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06249_),
    .X(_02152_));
 sg13g2_nand2_2 _24598_ (.Y(_06254_),
    .A(net699),
    .B(_06175_));
 sg13g2_mux2_1 _24599_ (.A0(_06237_),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06254_),
    .X(_02153_));
 sg13g2_mux2_1 _24600_ (.A0(_06239_),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06254_),
    .X(_02154_));
 sg13g2_mux2_1 _24601_ (.A0(_06241_),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06254_),
    .X(_02155_));
 sg13g2_mux2_1 _24602_ (.A0(net783),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06254_),
    .X(_02156_));
 sg13g2_and2_1 _24603_ (.A(_08205_),
    .B(_06178_),
    .X(_06255_));
 sg13g2_buf_2 _24604_ (.A(_06255_),
    .X(_06256_));
 sg13g2_mux2_1 _24605_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net788),
    .S(_06256_),
    .X(_02157_));
 sg13g2_mux2_1 _24606_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(_06226_),
    .S(_06256_),
    .X(_02158_));
 sg13g2_mux2_1 _24607_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net787),
    .S(_06256_),
    .X(_02159_));
 sg13g2_mux2_1 _24608_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(_06228_),
    .S(_06256_),
    .X(_02160_));
 sg13g2_nand2_2 _24609_ (.Y(_06257_),
    .A(net699),
    .B(_06184_));
 sg13g2_mux2_1 _24610_ (.A0(net786),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06257_),
    .X(_02161_));
 sg13g2_mux2_1 _24611_ (.A0(net785),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06257_),
    .X(_02162_));
 sg13g2_mux2_1 _24612_ (.A0(net784),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06249_),
    .X(_02163_));
 sg13g2_mux2_1 _24613_ (.A0(net784),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06257_),
    .X(_02164_));
 sg13g2_mux2_1 _24614_ (.A0(net783),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06257_),
    .X(_02165_));
 sg13g2_mux2_1 _24615_ (.A0(net783),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06249_),
    .X(_02166_));
 sg13g2_nand2_2 _24616_ (.Y(_06258_),
    .A(net699),
    .B(_06187_));
 sg13g2_mux2_1 _24617_ (.A0(_06189_),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06258_),
    .X(_02167_));
 sg13g2_mux2_1 _24618_ (.A0(net791),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06258_),
    .X(_02168_));
 sg13g2_mux2_1 _24619_ (.A0(_06194_),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06258_),
    .X(_02169_));
 sg13g2_mux2_1 _24620_ (.A0(net927),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06258_),
    .X(_02170_));
 sg13g2_mux2_1 _24621_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(_06224_),
    .S(_06251_),
    .X(_02171_));
 sg13g2_mux2_1 _24622_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(net925),
    .S(_06251_),
    .X(_02172_));
 sg13g2_nand2_2 _24623_ (.Y(_06259_),
    .A(net595),
    .B(_06153_));
 sg13g2_mux2_1 _24624_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][0] ),
    .S(_06259_),
    .X(_02173_));
 sg13g2_nand2_2 _24625_ (.Y(_06260_),
    .A(_08309_),
    .B(_06159_));
 sg13g2_mux2_1 _24626_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][10] ),
    .S(_06260_),
    .X(_02174_));
 sg13g2_mux2_1 _24627_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][11] ),
    .S(_06260_),
    .X(_02175_));
 sg13g2_nand2_2 _24628_ (.Y(_06261_),
    .A(net595),
    .B(_06165_));
 sg13g2_mux2_1 _24629_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][12] ),
    .S(_06261_),
    .X(_02176_));
 sg13g2_mux2_1 _24630_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][13] ),
    .S(_06261_),
    .X(_02177_));
 sg13g2_mux2_1 _24631_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][14] ),
    .S(_06261_),
    .X(_02178_));
 sg13g2_mux2_1 _24632_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][15] ),
    .S(_06261_),
    .X(_02179_));
 sg13g2_nand2_2 _24633_ (.Y(_06262_),
    .A(net595),
    .B(_06171_));
 sg13g2_mux2_1 _24634_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][16] ),
    .S(_06262_),
    .X(_02180_));
 sg13g2_mux2_1 _24635_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][17] ),
    .S(_06262_),
    .X(_02181_));
 sg13g2_mux2_1 _24636_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][18] ),
    .S(_06262_),
    .X(_02182_));
 sg13g2_mux2_1 _24637_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][19] ),
    .S(_06262_),
    .X(_02183_));
 sg13g2_mux2_1 _24638_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][1] ),
    .S(_06259_),
    .X(_02184_));
 sg13g2_nand2_2 _24639_ (.Y(_06263_),
    .A(net595),
    .B(_06175_));
 sg13g2_mux2_1 _24640_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][20] ),
    .S(_06263_),
    .X(_02185_));
 sg13g2_mux2_1 _24641_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][21] ),
    .S(_06263_),
    .X(_02186_));
 sg13g2_mux2_1 _24642_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][22] ),
    .S(_06263_),
    .X(_02187_));
 sg13g2_mux2_1 _24643_ (.A0(_06198_),
    .A1(\cpu.icache.r_data[5][23] ),
    .S(_06263_),
    .X(_02188_));
 sg13g2_nand2_1 _24644_ (.Y(_06264_),
    .A(net595),
    .B(_06178_));
 sg13g2_buf_2 _24645_ (.A(_06264_),
    .X(_06265_));
 sg13g2_mux2_1 _24646_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][24] ),
    .S(_06265_),
    .X(_02189_));
 sg13g2_mux2_1 _24647_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][25] ),
    .S(_06265_),
    .X(_02190_));
 sg13g2_mux2_1 _24648_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][26] ),
    .S(_06265_),
    .X(_02191_));
 sg13g2_mux2_1 _24649_ (.A0(_06198_),
    .A1(\cpu.icache.r_data[5][27] ),
    .S(_06265_),
    .X(_02192_));
 sg13g2_nand2_2 _24650_ (.Y(_06266_),
    .A(net595),
    .B(_06184_));
 sg13g2_mux2_1 _24651_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][28] ),
    .S(_06266_),
    .X(_02193_));
 sg13g2_mux2_1 _24652_ (.A0(net791),
    .A1(\cpu.icache.r_data[5][29] ),
    .S(_06266_),
    .X(_02194_));
 sg13g2_mux2_1 _24653_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][2] ),
    .S(_06259_),
    .X(_02195_));
 sg13g2_mux2_1 _24654_ (.A0(net793),
    .A1(\cpu.icache.r_data[5][30] ),
    .S(_06266_),
    .X(_02196_));
 sg13g2_mux2_1 _24655_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][31] ),
    .S(_06266_),
    .X(_02197_));
 sg13g2_mux2_1 _24656_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][3] ),
    .S(_06259_),
    .X(_02198_));
 sg13g2_nand2_2 _24657_ (.Y(_06267_),
    .A(_08309_),
    .B(_06187_));
 sg13g2_mux2_1 _24658_ (.A0(_06189_),
    .A1(\cpu.icache.r_data[5][4] ),
    .S(_06267_),
    .X(_02199_));
 sg13g2_mux2_1 _24659_ (.A0(_06202_),
    .A1(\cpu.icache.r_data[5][5] ),
    .S(_06267_),
    .X(_02200_));
 sg13g2_mux2_1 _24660_ (.A0(_06194_),
    .A1(\cpu.icache.r_data[5][6] ),
    .S(_06267_),
    .X(_02201_));
 sg13g2_mux2_1 _24661_ (.A0(net927),
    .A1(\cpu.icache.r_data[5][7] ),
    .S(_06267_),
    .X(_02202_));
 sg13g2_mux2_1 _24662_ (.A0(net794),
    .A1(\cpu.icache.r_data[5][8] ),
    .S(_06260_),
    .X(_02203_));
 sg13g2_mux2_1 _24663_ (.A0(_06202_),
    .A1(\cpu.icache.r_data[5][9] ),
    .S(_06260_),
    .X(_02204_));
 sg13g2_nand2_1 _24664_ (.Y(_06268_),
    .A(_08107_),
    .B(_08117_));
 sg13g2_buf_4 _24665_ (.X(_06269_),
    .A(_06268_));
 sg13g2_nor2_2 _24666_ (.A(_06269_),
    .B(_06192_),
    .Y(_06270_));
 sg13g2_mux2_1 _24667_ (.A0(\cpu.icache.r_data[6][0] ),
    .A1(net788),
    .S(_06270_),
    .X(_02205_));
 sg13g2_nor2_2 _24668_ (.A(_06269_),
    .B(_06196_),
    .Y(_06271_));
 sg13g2_mux2_1 _24669_ (.A0(\cpu.icache.r_data[6][10] ),
    .A1(_06227_),
    .S(_06271_),
    .X(_02206_));
 sg13g2_mux2_1 _24670_ (.A0(\cpu.icache.r_data[6][11] ),
    .A1(net924),
    .S(_06271_),
    .X(_02207_));
 sg13g2_nor2_2 _24671_ (.A(_06269_),
    .B(_06200_),
    .Y(_06272_));
 sg13g2_mux2_1 _24672_ (.A0(\cpu.icache.r_data[6][12] ),
    .A1(net788),
    .S(_06272_),
    .X(_02208_));
 sg13g2_mux2_1 _24673_ (.A0(\cpu.icache.r_data[6][13] ),
    .A1(net925),
    .S(_06272_),
    .X(_02209_));
 sg13g2_mux2_1 _24674_ (.A0(\cpu.icache.r_data[6][14] ),
    .A1(net787),
    .S(_06272_),
    .X(_02210_));
 sg13g2_mux2_1 _24675_ (.A0(\cpu.icache.r_data[6][15] ),
    .A1(_06228_),
    .S(_06272_),
    .X(_02211_));
 sg13g2_buf_1 _24676_ (.A(_12162_),
    .X(_06273_));
 sg13g2_nor2_2 _24677_ (.A(_06269_),
    .B(_06205_),
    .Y(_06274_));
 sg13g2_mux2_1 _24678_ (.A0(\cpu.icache.r_data[6][16] ),
    .A1(net782),
    .S(_06274_),
    .X(_02212_));
 sg13g2_mux2_1 _24679_ (.A0(\cpu.icache.r_data[6][17] ),
    .A1(net925),
    .S(_06274_),
    .X(_02213_));
 sg13g2_buf_2 _24680_ (.A(_11810_),
    .X(_06275_));
 sg13g2_mux2_1 _24681_ (.A0(\cpu.icache.r_data[6][18] ),
    .A1(net923),
    .S(_06274_),
    .X(_02214_));
 sg13g2_buf_1 _24682_ (.A(_11833_),
    .X(_06276_));
 sg13g2_mux2_1 _24683_ (.A0(\cpu.icache.r_data[6][19] ),
    .A1(_06276_),
    .S(_06274_),
    .X(_02215_));
 sg13g2_buf_1 _24684_ (.A(_11743_),
    .X(_06277_));
 sg13g2_mux2_1 _24685_ (.A0(\cpu.icache.r_data[6][1] ),
    .A1(net921),
    .S(_06270_),
    .X(_02216_));
 sg13g2_nor2_2 _24686_ (.A(_06269_),
    .B(_06208_),
    .Y(_06278_));
 sg13g2_mux2_1 _24687_ (.A0(\cpu.icache.r_data[6][20] ),
    .A1(_06273_),
    .S(_06278_),
    .X(_02217_));
 sg13g2_mux2_1 _24688_ (.A0(\cpu.icache.r_data[6][21] ),
    .A1(net921),
    .S(_06278_),
    .X(_02218_));
 sg13g2_mux2_1 _24689_ (.A0(\cpu.icache.r_data[6][22] ),
    .A1(_06275_),
    .S(_06278_),
    .X(_02219_));
 sg13g2_mux2_1 _24690_ (.A0(\cpu.icache.r_data[6][23] ),
    .A1(net922),
    .S(_06278_),
    .X(_02220_));
 sg13g2_nor2_1 _24691_ (.A(_06269_),
    .B(_06211_),
    .Y(_06279_));
 sg13g2_buf_2 _24692_ (.A(_06279_),
    .X(_06280_));
 sg13g2_mux2_1 _24693_ (.A0(\cpu.icache.r_data[6][24] ),
    .A1(net782),
    .S(_06280_),
    .X(_02221_));
 sg13g2_mux2_1 _24694_ (.A0(\cpu.icache.r_data[6][25] ),
    .A1(net921),
    .S(_06280_),
    .X(_02222_));
 sg13g2_mux2_1 _24695_ (.A0(\cpu.icache.r_data[6][26] ),
    .A1(net923),
    .S(_06280_),
    .X(_02223_));
 sg13g2_mux2_1 _24696_ (.A0(\cpu.icache.r_data[6][27] ),
    .A1(net922),
    .S(_06280_),
    .X(_02224_));
 sg13g2_nor2_2 _24697_ (.A(_06269_),
    .B(_06214_),
    .Y(_06281_));
 sg13g2_mux2_1 _24698_ (.A0(\cpu.icache.r_data[6][28] ),
    .A1(net782),
    .S(_06281_),
    .X(_02225_));
 sg13g2_mux2_1 _24699_ (.A0(\cpu.icache.r_data[6][29] ),
    .A1(net921),
    .S(_06281_),
    .X(_02226_));
 sg13g2_mux2_1 _24700_ (.A0(\cpu.icache.r_data[6][2] ),
    .A1(net923),
    .S(_06270_),
    .X(_02227_));
 sg13g2_mux2_1 _24701_ (.A0(\cpu.icache.r_data[6][30] ),
    .A1(net923),
    .S(_06281_),
    .X(_02228_));
 sg13g2_mux2_1 _24702_ (.A0(\cpu.icache.r_data[6][31] ),
    .A1(net922),
    .S(_06281_),
    .X(_02229_));
 sg13g2_mux2_1 _24703_ (.A0(\cpu.icache.r_data[6][3] ),
    .A1(net922),
    .S(_06270_),
    .X(_02230_));
 sg13g2_nor2_2 _24704_ (.A(_06269_),
    .B(_06216_),
    .Y(_06282_));
 sg13g2_mux2_1 _24705_ (.A0(\cpu.icache.r_data[6][4] ),
    .A1(net782),
    .S(_06282_),
    .X(_02231_));
 sg13g2_mux2_1 _24706_ (.A0(\cpu.icache.r_data[6][5] ),
    .A1(_06277_),
    .S(_06282_),
    .X(_02232_));
 sg13g2_mux2_1 _24707_ (.A0(\cpu.icache.r_data[6][6] ),
    .A1(net923),
    .S(_06282_),
    .X(_02233_));
 sg13g2_mux2_1 _24708_ (.A0(\cpu.icache.r_data[6][7] ),
    .A1(net922),
    .S(_06282_),
    .X(_02234_));
 sg13g2_mux2_1 _24709_ (.A0(\cpu.icache.r_data[6][8] ),
    .A1(net782),
    .S(_06271_),
    .X(_02235_));
 sg13g2_mux2_1 _24710_ (.A0(\cpu.icache.r_data[6][9] ),
    .A1(_06277_),
    .S(_06271_),
    .X(_02236_));
 sg13g2_nand2_1 _24711_ (.Y(_06283_),
    .A(net777),
    .B(_08236_));
 sg13g2_buf_4 _24712_ (.X(_06284_),
    .A(_06283_));
 sg13g2_nor2_2 _24713_ (.A(_06284_),
    .B(_06192_),
    .Y(_06285_));
 sg13g2_mux2_1 _24714_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net782),
    .S(_06285_),
    .X(_02237_));
 sg13g2_nor2_2 _24715_ (.A(_06284_),
    .B(_06196_),
    .Y(_06286_));
 sg13g2_mux2_1 _24716_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net923),
    .S(_06286_),
    .X(_02238_));
 sg13g2_mux2_1 _24717_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net922),
    .S(_06286_),
    .X(_02239_));
 sg13g2_nor2_2 _24718_ (.A(_06284_),
    .B(_06200_),
    .Y(_06287_));
 sg13g2_mux2_1 _24719_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(_06273_),
    .S(_06287_),
    .X(_02240_));
 sg13g2_mux2_1 _24720_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net921),
    .S(_06287_),
    .X(_02241_));
 sg13g2_mux2_1 _24721_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(_06275_),
    .S(_06287_),
    .X(_02242_));
 sg13g2_mux2_1 _24722_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net922),
    .S(_06287_),
    .X(_02243_));
 sg13g2_nor2_2 _24723_ (.A(_06284_),
    .B(_06205_),
    .Y(_06288_));
 sg13g2_mux2_1 _24724_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(net782),
    .S(_06288_),
    .X(_02244_));
 sg13g2_mux2_1 _24725_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net921),
    .S(_06288_),
    .X(_02245_));
 sg13g2_mux2_1 _24726_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(net923),
    .S(_06288_),
    .X(_02246_));
 sg13g2_mux2_1 _24727_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(_06276_),
    .S(_06288_),
    .X(_02247_));
 sg13g2_mux2_1 _24728_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net921),
    .S(_06285_),
    .X(_02248_));
 sg13g2_nor2_2 _24729_ (.A(_06284_),
    .B(_06208_),
    .Y(_06289_));
 sg13g2_mux2_1 _24730_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net782),
    .S(_06289_),
    .X(_02249_));
 sg13g2_mux2_1 _24731_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(net921),
    .S(_06289_),
    .X(_02250_));
 sg13g2_mux2_1 _24732_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net923),
    .S(_06289_),
    .X(_02251_));
 sg13g2_mux2_1 _24733_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net922),
    .S(_06289_),
    .X(_02252_));
 sg13g2_nor2_1 _24734_ (.A(_06284_),
    .B(_06211_),
    .Y(_06290_));
 sg13g2_buf_2 _24735_ (.A(_06290_),
    .X(_06291_));
 sg13g2_mux2_1 _24736_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net968),
    .S(_06291_),
    .X(_02253_));
 sg13g2_mux2_1 _24737_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net967),
    .S(_06291_),
    .X(_02254_));
 sg13g2_mux2_1 _24738_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net982),
    .S(_06291_),
    .X(_02255_));
 sg13g2_mux2_1 _24739_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net981),
    .S(_06291_),
    .X(_02256_));
 sg13g2_nor2_2 _24740_ (.A(_06284_),
    .B(_06214_),
    .Y(_06292_));
 sg13g2_mux2_1 _24741_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net968),
    .S(_06292_),
    .X(_02257_));
 sg13g2_mux2_1 _24742_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net967),
    .S(_06292_),
    .X(_02258_));
 sg13g2_mux2_1 _24743_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net982),
    .S(_06285_),
    .X(_02259_));
 sg13g2_mux2_1 _24744_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_11695_),
    .S(_06292_),
    .X(_02260_));
 sg13g2_mux2_1 _24745_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net981),
    .S(_06292_),
    .X(_02261_));
 sg13g2_mux2_1 _24746_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_11712_),
    .S(_06285_),
    .X(_02262_));
 sg13g2_nor2_2 _24747_ (.A(_06284_),
    .B(_06216_),
    .Y(_06293_));
 sg13g2_mux2_1 _24748_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_11866_),
    .S(_06293_),
    .X(_02263_));
 sg13g2_mux2_1 _24749_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_11870_),
    .S(_06293_),
    .X(_02264_));
 sg13g2_mux2_1 _24750_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_11695_),
    .S(_06293_),
    .X(_02265_));
 sg13g2_mux2_1 _24751_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_11712_),
    .S(_06293_),
    .X(_02266_));
 sg13g2_mux2_1 _24752_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_11866_),
    .S(_06286_),
    .X(_02267_));
 sg13g2_mux2_1 _24753_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_11870_),
    .S(_06286_),
    .X(_02268_));
 sg13g2_mux2_1 _24754_ (.A0(net948),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(_06182_),
    .X(_02272_));
 sg13g2_buf_1 _24755_ (.A(_06180_),
    .X(_06294_));
 sg13g2_nand2_1 _24756_ (.Y(_06295_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(_06182_));
 sg13g2_o21ai_1 _24757_ (.B1(_06295_),
    .Y(_02273_),
    .A1(net466),
    .A2(net344));
 sg13g2_nand2_1 _24758_ (.Y(_06296_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net345));
 sg13g2_o21ai_1 _24759_ (.B1(_06296_),
    .Y(_02274_),
    .A1(net470),
    .A2(net344));
 sg13g2_nand2_1 _24760_ (.Y(_06297_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net345));
 sg13g2_o21ai_1 _24761_ (.B1(_06297_),
    .Y(_02275_),
    .A1(net467),
    .A2(net344));
 sg13g2_nand2_1 _24762_ (.Y(_06298_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net345));
 sg13g2_o21ai_1 _24763_ (.B1(_06298_),
    .Y(_02276_),
    .A1(net409),
    .A2(net344));
 sg13g2_nand2_1 _24764_ (.Y(_06299_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(net345));
 sg13g2_o21ai_1 _24765_ (.B1(_06299_),
    .Y(_02277_),
    .A1(net468),
    .A2(net344));
 sg13g2_nand2_1 _24766_ (.Y(_06300_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net345));
 sg13g2_o21ai_1 _24767_ (.B1(_06300_),
    .Y(_02278_),
    .A1(net407),
    .A2(_06294_));
 sg13g2_buf_1 _24768_ (.A(_06180_),
    .X(_06301_));
 sg13g2_nand2_1 _24769_ (.Y(_06302_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net343));
 sg13g2_o21ai_1 _24770_ (.B1(_06302_),
    .Y(_02279_),
    .A1(net408),
    .A2(net344));
 sg13g2_nand2_1 _24771_ (.Y(_06303_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net343));
 sg13g2_o21ai_1 _24772_ (.B1(_06303_),
    .Y(_02280_),
    .A1(net471),
    .A2(net344));
 sg13g2_nand2_1 _24773_ (.Y(_06304_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net343));
 sg13g2_o21ai_1 _24774_ (.B1(_06304_),
    .Y(_02281_),
    .A1(_08327_),
    .A2(net344));
 sg13g2_mux2_1 _24775_ (.A0(net947),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net345),
    .X(_02282_));
 sg13g2_nand2_1 _24776_ (.Y(_06305_),
    .A(\cpu.icache.r_tag[0][7] ),
    .B(net343));
 sg13g2_o21ai_1 _24777_ (.B1(_06305_),
    .Y(_02283_),
    .A1(_08500_),
    .A2(net346));
 sg13g2_nand2_1 _24778_ (.Y(_06306_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(net343));
 sg13g2_o21ai_1 _24779_ (.B1(_06306_),
    .Y(_02284_),
    .A1(net950),
    .A2(net346));
 sg13g2_nand2_1 _24780_ (.Y(_06307_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(net343));
 sg13g2_o21ai_1 _24781_ (.B1(_06307_),
    .Y(_02285_),
    .A1(net888),
    .A2(net346));
 sg13g2_mux2_1 _24782_ (.A0(net946),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net345),
    .X(_02286_));
 sg13g2_nand2_1 _24783_ (.Y(_06308_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(_06301_));
 sg13g2_o21ai_1 _24784_ (.B1(_06308_),
    .Y(_02287_),
    .A1(net1030),
    .A2(net346));
 sg13g2_nand2_1 _24785_ (.Y(_06309_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net343));
 sg13g2_o21ai_1 _24786_ (.B1(_06309_),
    .Y(_02288_),
    .A1(net474),
    .A2(net346));
 sg13g2_nand2_1 _24787_ (.Y(_06310_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(_06301_));
 sg13g2_o21ai_1 _24788_ (.B1(_06310_),
    .Y(_02289_),
    .A1(net478),
    .A2(net346));
 sg13g2_nand2_1 _24789_ (.Y(_06311_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net343));
 sg13g2_o21ai_1 _24790_ (.B1(_06311_),
    .Y(_02290_),
    .A1(_08353_),
    .A2(net346));
 sg13g2_nor2b_1 _24791_ (.A(_06158_),
    .B_N(_06169_),
    .Y(_06312_));
 sg13g2_buf_1 _24792_ (.A(_06312_),
    .X(_06313_));
 sg13g2_nand2_1 _24793_ (.Y(_06314_),
    .A(_08127_),
    .B(_06313_));
 sg13g2_buf_2 _24794_ (.A(_06314_),
    .X(_06315_));
 sg13g2_buf_1 _24795_ (.A(_06315_),
    .X(_06316_));
 sg13g2_mux2_1 _24796_ (.A0(net948),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net377),
    .X(_02291_));
 sg13g2_buf_1 _24797_ (.A(_06315_),
    .X(_06317_));
 sg13g2_nand2_1 _24798_ (.Y(_06318_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net377));
 sg13g2_o21ai_1 _24799_ (.B1(_06318_),
    .Y(_02292_),
    .A1(net466),
    .A2(_06317_));
 sg13g2_buf_1 _24800_ (.A(_06315_),
    .X(_06319_));
 sg13g2_nand2_1 _24801_ (.Y(_06320_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net375));
 sg13g2_o21ai_1 _24802_ (.B1(_06320_),
    .Y(_02293_),
    .A1(net470),
    .A2(net376));
 sg13g2_nand2_1 _24803_ (.Y(_06321_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net375));
 sg13g2_o21ai_1 _24804_ (.B1(_06321_),
    .Y(_02294_),
    .A1(net467),
    .A2(net376));
 sg13g2_nand2_1 _24805_ (.Y(_06322_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net375));
 sg13g2_o21ai_1 _24806_ (.B1(_06322_),
    .Y(_02295_),
    .A1(net409),
    .A2(net376));
 sg13g2_nand2_1 _24807_ (.Y(_06323_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net375));
 sg13g2_o21ai_1 _24808_ (.B1(_06323_),
    .Y(_02296_),
    .A1(net468),
    .A2(net376));
 sg13g2_nand2_1 _24809_ (.Y(_06324_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net375));
 sg13g2_o21ai_1 _24810_ (.B1(_06324_),
    .Y(_02297_),
    .A1(net407),
    .A2(net376));
 sg13g2_nand2_1 _24811_ (.Y(_06325_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net375));
 sg13g2_o21ai_1 _24812_ (.B1(_06325_),
    .Y(_02298_),
    .A1(net408),
    .A2(net376));
 sg13g2_nand2_1 _24813_ (.Y(_06326_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(_06319_));
 sg13g2_o21ai_1 _24814_ (.B1(_06326_),
    .Y(_02299_),
    .A1(net471),
    .A2(_06317_));
 sg13g2_nand2_1 _24815_ (.Y(_06327_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net375));
 sg13g2_o21ai_1 _24816_ (.B1(_06327_),
    .Y(_02300_),
    .A1(net542),
    .A2(net376));
 sg13g2_mux2_1 _24817_ (.A0(net947),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net377),
    .X(_02301_));
 sg13g2_nand2_1 _24818_ (.Y(_06328_),
    .A(\cpu.icache.r_tag[1][7] ),
    .B(net375));
 sg13g2_o21ai_1 _24819_ (.B1(_06328_),
    .Y(_02302_),
    .A1(net1029),
    .A2(net376));
 sg13g2_nand2_1 _24820_ (.Y(_06329_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(_06319_));
 sg13g2_o21ai_1 _24821_ (.B1(_06329_),
    .Y(_02303_),
    .A1(net950),
    .A2(net377));
 sg13g2_nand2_1 _24822_ (.Y(_06330_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(_06315_));
 sg13g2_o21ai_1 _24823_ (.B1(_06330_),
    .Y(_02304_),
    .A1(net888),
    .A2(net377));
 sg13g2_mux2_1 _24824_ (.A0(net946),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net377),
    .X(_02305_));
 sg13g2_nand2_1 _24825_ (.Y(_06331_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(_06315_));
 sg13g2_o21ai_1 _24826_ (.B1(_06331_),
    .Y(_02306_),
    .A1(_08446_),
    .A2(net377));
 sg13g2_nand2_1 _24827_ (.Y(_06332_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06315_));
 sg13g2_o21ai_1 _24828_ (.B1(_06332_),
    .Y(_02307_),
    .A1(net474),
    .A2(_06316_));
 sg13g2_nand2_1 _24829_ (.Y(_06333_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06315_));
 sg13g2_o21ai_1 _24830_ (.B1(_06333_),
    .Y(_02308_),
    .A1(net478),
    .A2(net377));
 sg13g2_nand2_1 _24831_ (.Y(_06334_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06315_));
 sg13g2_o21ai_1 _24832_ (.B1(_06334_),
    .Y(_02309_),
    .A1(net469),
    .A2(_06316_));
 sg13g2_nand2_1 _24833_ (.Y(_06335_),
    .A(net475),
    .B(_06313_));
 sg13g2_buf_2 _24834_ (.A(_06335_),
    .X(_06336_));
 sg13g2_buf_1 _24835_ (.A(_06336_),
    .X(_06337_));
 sg13g2_mux2_1 _24836_ (.A0(net948),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net301),
    .X(_02310_));
 sg13g2_buf_1 _24837_ (.A(_06336_),
    .X(_06338_));
 sg13g2_nand2_1 _24838_ (.Y(_06339_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net301));
 sg13g2_o21ai_1 _24839_ (.B1(_06339_),
    .Y(_02311_),
    .A1(net466),
    .A2(net300));
 sg13g2_buf_1 _24840_ (.A(_06336_),
    .X(_06340_));
 sg13g2_nand2_1 _24841_ (.Y(_06341_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net299));
 sg13g2_o21ai_1 _24842_ (.B1(_06341_),
    .Y(_02312_),
    .A1(net470),
    .A2(net300));
 sg13g2_nand2_1 _24843_ (.Y(_06342_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net299));
 sg13g2_o21ai_1 _24844_ (.B1(_06342_),
    .Y(_02313_),
    .A1(net467),
    .A2(net300));
 sg13g2_nand2_1 _24845_ (.Y(_06343_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net299));
 sg13g2_o21ai_1 _24846_ (.B1(_06343_),
    .Y(_02314_),
    .A1(_08196_),
    .A2(_06338_));
 sg13g2_nand2_1 _24847_ (.Y(_06344_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net299));
 sg13g2_o21ai_1 _24848_ (.B1(_06344_),
    .Y(_02315_),
    .A1(net468),
    .A2(net300));
 sg13g2_nand2_1 _24849_ (.Y(_06345_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net299));
 sg13g2_o21ai_1 _24850_ (.B1(_06345_),
    .Y(_02316_),
    .A1(net407),
    .A2(net300));
 sg13g2_nand2_1 _24851_ (.Y(_06346_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(_06340_));
 sg13g2_o21ai_1 _24852_ (.B1(_06346_),
    .Y(_02317_),
    .A1(net408),
    .A2(_06338_));
 sg13g2_nand2_1 _24853_ (.Y(_06347_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(_06340_));
 sg13g2_o21ai_1 _24854_ (.B1(_06347_),
    .Y(_02318_),
    .A1(net471),
    .A2(net300));
 sg13g2_nand2_1 _24855_ (.Y(_06348_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net299));
 sg13g2_o21ai_1 _24856_ (.B1(_06348_),
    .Y(_02319_),
    .A1(net542),
    .A2(net300));
 sg13g2_mux2_1 _24857_ (.A0(net947),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net301),
    .X(_02320_));
 sg13g2_nand2_1 _24858_ (.Y(_06349_),
    .A(\cpu.icache.r_tag[2][7] ),
    .B(net299));
 sg13g2_o21ai_1 _24859_ (.B1(_06349_),
    .Y(_02321_),
    .A1(net1029),
    .A2(net300));
 sg13g2_nand2_1 _24860_ (.Y(_06350_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(net299));
 sg13g2_o21ai_1 _24861_ (.B1(_06350_),
    .Y(_02322_),
    .A1(net950),
    .A2(net301));
 sg13g2_nand2_1 _24862_ (.Y(_06351_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(_06336_));
 sg13g2_o21ai_1 _24863_ (.B1(_06351_),
    .Y(_02323_),
    .A1(net888),
    .A2(_06337_));
 sg13g2_mux2_1 _24864_ (.A0(net946),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net301),
    .X(_02324_));
 sg13g2_nand2_1 _24865_ (.Y(_06352_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06336_));
 sg13g2_o21ai_1 _24866_ (.B1(_06352_),
    .Y(_02325_),
    .A1(net1030),
    .A2(_06337_));
 sg13g2_nand2_1 _24867_ (.Y(_06353_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06336_));
 sg13g2_o21ai_1 _24868_ (.B1(_06353_),
    .Y(_02326_),
    .A1(net474),
    .A2(net301));
 sg13g2_nand2_1 _24869_ (.Y(_06354_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06336_));
 sg13g2_o21ai_1 _24870_ (.B1(_06354_),
    .Y(_02327_),
    .A1(net478),
    .A2(net301));
 sg13g2_nand2_1 _24871_ (.Y(_06355_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06336_));
 sg13g2_o21ai_1 _24872_ (.B1(_06355_),
    .Y(_02328_),
    .A1(net469),
    .A2(net301));
 sg13g2_mux2_1 _24873_ (.A0(net948),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(_06246_),
    .X(_02329_));
 sg13g2_buf_1 _24874_ (.A(_06244_),
    .X(_06356_));
 sg13g2_nand2_1 _24875_ (.Y(_06357_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net302));
 sg13g2_o21ai_1 _24876_ (.B1(_06357_),
    .Y(_02330_),
    .A1(net466),
    .A2(net298));
 sg13g2_nand2_1 _24877_ (.Y(_06358_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net302));
 sg13g2_o21ai_1 _24878_ (.B1(_06358_),
    .Y(_02331_),
    .A1(net470),
    .A2(net298));
 sg13g2_nand2_1 _24879_ (.Y(_06359_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net302));
 sg13g2_o21ai_1 _24880_ (.B1(_06359_),
    .Y(_02332_),
    .A1(net467),
    .A2(net298));
 sg13g2_nand2_1 _24881_ (.Y(_06360_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net302));
 sg13g2_o21ai_1 _24882_ (.B1(_06360_),
    .Y(_02333_),
    .A1(net409),
    .A2(_06356_));
 sg13g2_nand2_1 _24883_ (.Y(_06361_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net302));
 sg13g2_o21ai_1 _24884_ (.B1(_06361_),
    .Y(_02334_),
    .A1(net468),
    .A2(net298));
 sg13g2_nand2_1 _24885_ (.Y(_06362_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net302));
 sg13g2_o21ai_1 _24886_ (.B1(_06362_),
    .Y(_02335_),
    .A1(net407),
    .A2(net298));
 sg13g2_buf_1 _24887_ (.A(_06244_),
    .X(_06363_));
 sg13g2_nand2_1 _24888_ (.Y(_06364_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(_06363_));
 sg13g2_o21ai_1 _24889_ (.B1(_06364_),
    .Y(_02336_),
    .A1(net408),
    .A2(net298));
 sg13g2_nand2_1 _24890_ (.Y(_06365_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(_06363_));
 sg13g2_o21ai_1 _24891_ (.B1(_06365_),
    .Y(_02337_),
    .A1(net471),
    .A2(net298));
 sg13g2_nand2_1 _24892_ (.Y(_06366_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net297));
 sg13g2_o21ai_1 _24893_ (.B1(_06366_),
    .Y(_02338_),
    .A1(net542),
    .A2(net298));
 sg13g2_mux2_1 _24894_ (.A0(net947),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net302),
    .X(_02339_));
 sg13g2_nand2_1 _24895_ (.Y(_06367_),
    .A(\cpu.icache.r_tag[3][7] ),
    .B(net297));
 sg13g2_o21ai_1 _24896_ (.B1(_06367_),
    .Y(_02340_),
    .A1(net1029),
    .A2(net303));
 sg13g2_nand2_1 _24897_ (.Y(_06368_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net297));
 sg13g2_o21ai_1 _24898_ (.B1(_06368_),
    .Y(_02341_),
    .A1(net950),
    .A2(net303));
 sg13g2_nand2_1 _24899_ (.Y(_06369_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(net297));
 sg13g2_o21ai_1 _24900_ (.B1(_06369_),
    .Y(_02342_),
    .A1(net888),
    .A2(net303));
 sg13g2_mux2_1 _24901_ (.A0(net946),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net302),
    .X(_02343_));
 sg13g2_nand2_1 _24902_ (.Y(_06370_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net297));
 sg13g2_o21ai_1 _24903_ (.B1(_06370_),
    .Y(_02344_),
    .A1(net1030),
    .A2(net303));
 sg13g2_nand2_1 _24904_ (.Y(_06371_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net297));
 sg13g2_o21ai_1 _24905_ (.B1(_06371_),
    .Y(_02345_),
    .A1(net474),
    .A2(_06245_));
 sg13g2_nand2_1 _24906_ (.Y(_06372_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net297));
 sg13g2_o21ai_1 _24907_ (.B1(_06372_),
    .Y(_02346_),
    .A1(net478),
    .A2(_06245_));
 sg13g2_nand2_1 _24908_ (.Y(_06373_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net297));
 sg13g2_o21ai_1 _24909_ (.B1(_06373_),
    .Y(_02347_),
    .A1(net469),
    .A2(net303));
 sg13g2_nand2_1 _24910_ (.Y(_06374_),
    .A(_08205_),
    .B(_06313_));
 sg13g2_buf_2 _24911_ (.A(_06374_),
    .X(_06375_));
 sg13g2_buf_1 _24912_ (.A(_06375_),
    .X(_06376_));
 sg13g2_mux2_1 _24913_ (.A0(net948),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net417),
    .X(_02348_));
 sg13g2_buf_1 _24914_ (.A(_06375_),
    .X(_06377_));
 sg13g2_nand2_1 _24915_ (.Y(_06378_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net417));
 sg13g2_o21ai_1 _24916_ (.B1(_06378_),
    .Y(_02349_),
    .A1(_08425_),
    .A2(_06377_));
 sg13g2_buf_1 _24917_ (.A(_06375_),
    .X(_06379_));
 sg13g2_nand2_1 _24918_ (.Y(_06380_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net415));
 sg13g2_o21ai_1 _24919_ (.B1(_06380_),
    .Y(_02350_),
    .A1(net470),
    .A2(net416));
 sg13g2_nand2_1 _24920_ (.Y(_06381_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net415));
 sg13g2_o21ai_1 _24921_ (.B1(_06381_),
    .Y(_02351_),
    .A1(net467),
    .A2(net416));
 sg13g2_nand2_1 _24922_ (.Y(_06382_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net415));
 sg13g2_o21ai_1 _24923_ (.B1(_06382_),
    .Y(_02352_),
    .A1(net409),
    .A2(net416));
 sg13g2_nand2_1 _24924_ (.Y(_06383_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net415));
 sg13g2_o21ai_1 _24925_ (.B1(_06383_),
    .Y(_02353_),
    .A1(net468),
    .A2(net416));
 sg13g2_nand2_1 _24926_ (.Y(_06384_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(_06379_));
 sg13g2_o21ai_1 _24927_ (.B1(_06384_),
    .Y(_02354_),
    .A1(_08305_),
    .A2(net416));
 sg13g2_nand2_1 _24928_ (.Y(_06385_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net415));
 sg13g2_o21ai_1 _24929_ (.B1(_06385_),
    .Y(_02355_),
    .A1(net408),
    .A2(net416));
 sg13g2_nand2_1 _24930_ (.Y(_06386_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net415));
 sg13g2_o21ai_1 _24931_ (.B1(_06386_),
    .Y(_02356_),
    .A1(net471),
    .A2(net416));
 sg13g2_nand2_1 _24932_ (.Y(_06387_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net415));
 sg13g2_o21ai_1 _24933_ (.B1(_06387_),
    .Y(_02357_),
    .A1(net542),
    .A2(net416));
 sg13g2_mux2_1 _24934_ (.A0(net947),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net417),
    .X(_02358_));
 sg13g2_nand2_1 _24935_ (.Y(_06388_),
    .A(\cpu.icache.r_tag[4][7] ),
    .B(net415));
 sg13g2_o21ai_1 _24936_ (.B1(_06388_),
    .Y(_02359_),
    .A1(net1029),
    .A2(_06377_));
 sg13g2_nand2_1 _24937_ (.Y(_06389_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(_06379_));
 sg13g2_o21ai_1 _24938_ (.B1(_06389_),
    .Y(_02360_),
    .A1(net950),
    .A2(net417));
 sg13g2_nand2_1 _24939_ (.Y(_06390_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(_06375_));
 sg13g2_o21ai_1 _24940_ (.B1(_06390_),
    .Y(_02361_),
    .A1(_08462_),
    .A2(_06376_));
 sg13g2_mux2_1 _24941_ (.A0(net946),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net417),
    .X(_02362_));
 sg13g2_nand2_1 _24942_ (.Y(_06391_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(_06375_));
 sg13g2_o21ai_1 _24943_ (.B1(_06391_),
    .Y(_02363_),
    .A1(net1030),
    .A2(net417));
 sg13g2_nand2_1 _24944_ (.Y(_06392_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06375_));
 sg13g2_o21ai_1 _24945_ (.B1(_06392_),
    .Y(_02364_),
    .A1(net474),
    .A2(_06376_));
 sg13g2_nand2_1 _24946_ (.Y(_06393_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06375_));
 sg13g2_o21ai_1 _24947_ (.B1(_06393_),
    .Y(_02365_),
    .A1(net478),
    .A2(net417));
 sg13g2_nand2_1 _24948_ (.Y(_06394_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06375_));
 sg13g2_o21ai_1 _24949_ (.B1(_06394_),
    .Y(_02366_),
    .A1(net469),
    .A2(net417));
 sg13g2_nand2_1 _24950_ (.Y(_06395_),
    .A(net595),
    .B(_06313_));
 sg13g2_buf_2 _24951_ (.A(_06395_),
    .X(_06396_));
 sg13g2_buf_1 _24952_ (.A(_06396_),
    .X(_06397_));
 sg13g2_mux2_1 _24953_ (.A0(net948),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net374),
    .X(_02367_));
 sg13g2_buf_1 _24954_ (.A(_06396_),
    .X(_06398_));
 sg13g2_nand2_1 _24955_ (.Y(_06399_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net374));
 sg13g2_o21ai_1 _24956_ (.B1(_06399_),
    .Y(_02368_),
    .A1(net466),
    .A2(net373));
 sg13g2_buf_1 _24957_ (.A(_06396_),
    .X(_06400_));
 sg13g2_nand2_1 _24958_ (.Y(_06401_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net372));
 sg13g2_o21ai_1 _24959_ (.B1(_06401_),
    .Y(_02369_),
    .A1(net470),
    .A2(net373));
 sg13g2_nand2_1 _24960_ (.Y(_06402_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net372));
 sg13g2_o21ai_1 _24961_ (.B1(_06402_),
    .Y(_02370_),
    .A1(net467),
    .A2(net373));
 sg13g2_nand2_1 _24962_ (.Y(_06403_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net372));
 sg13g2_o21ai_1 _24963_ (.B1(_06403_),
    .Y(_02371_),
    .A1(net409),
    .A2(_06398_));
 sg13g2_nand2_1 _24964_ (.Y(_06404_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net372));
 sg13g2_o21ai_1 _24965_ (.B1(_06404_),
    .Y(_02372_),
    .A1(net468),
    .A2(net373));
 sg13g2_nand2_1 _24966_ (.Y(_06405_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net372));
 sg13g2_o21ai_1 _24967_ (.B1(_06405_),
    .Y(_02373_),
    .A1(net407),
    .A2(net373));
 sg13g2_nand2_1 _24968_ (.Y(_06406_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(_06400_));
 sg13g2_o21ai_1 _24969_ (.B1(_06406_),
    .Y(_02374_),
    .A1(net408),
    .A2(net373));
 sg13g2_nand2_1 _24970_ (.Y(_06407_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(_06400_));
 sg13g2_o21ai_1 _24971_ (.B1(_06407_),
    .Y(_02375_),
    .A1(_08253_),
    .A2(_06398_));
 sg13g2_nand2_1 _24972_ (.Y(_06408_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net372));
 sg13g2_o21ai_1 _24973_ (.B1(_06408_),
    .Y(_02376_),
    .A1(net542),
    .A2(net373));
 sg13g2_mux2_1 _24974_ (.A0(net947),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(net374),
    .X(_02377_));
 sg13g2_nand2_1 _24975_ (.Y(_06409_),
    .A(\cpu.icache.r_tag[5][7] ),
    .B(net372));
 sg13g2_o21ai_1 _24976_ (.B1(_06409_),
    .Y(_02378_),
    .A1(net1029),
    .A2(net373));
 sg13g2_nand2_1 _24977_ (.Y(_06410_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net372));
 sg13g2_o21ai_1 _24978_ (.B1(_06410_),
    .Y(_02379_),
    .A1(net950),
    .A2(net374));
 sg13g2_nand2_1 _24979_ (.Y(_06411_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(_06396_));
 sg13g2_o21ai_1 _24980_ (.B1(_06411_),
    .Y(_02380_),
    .A1(net888),
    .A2(net374));
 sg13g2_mux2_1 _24981_ (.A0(net946),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net374),
    .X(_02381_));
 sg13g2_nand2_1 _24982_ (.Y(_06412_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(_06396_));
 sg13g2_o21ai_1 _24983_ (.B1(_06412_),
    .Y(_02382_),
    .A1(net1030),
    .A2(net374));
 sg13g2_nand2_1 _24984_ (.Y(_06413_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06396_));
 sg13g2_o21ai_1 _24985_ (.B1(_06413_),
    .Y(_02383_),
    .A1(net474),
    .A2(net374));
 sg13g2_nand2_1 _24986_ (.Y(_06414_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06396_));
 sg13g2_o21ai_1 _24987_ (.B1(_06414_),
    .Y(_02384_),
    .A1(_08087_),
    .A2(_06397_));
 sg13g2_nand2_1 _24988_ (.Y(_06415_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06396_));
 sg13g2_o21ai_1 _24989_ (.B1(_06415_),
    .Y(_02385_),
    .A1(net469),
    .A2(_06397_));
 sg13g2_nand2_1 _24990_ (.Y(_06416_),
    .A(_08155_),
    .B(_06313_));
 sg13g2_buf_2 _24991_ (.A(_06416_),
    .X(_06417_));
 sg13g2_buf_1 _24992_ (.A(_06417_),
    .X(_06418_));
 sg13g2_mux2_1 _24993_ (.A0(_04412_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net342),
    .X(_02386_));
 sg13g2_buf_1 _24994_ (.A(_06417_),
    .X(_06419_));
 sg13g2_nand2_1 _24995_ (.Y(_06420_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net342));
 sg13g2_o21ai_1 _24996_ (.B1(_06420_),
    .Y(_02387_),
    .A1(net466),
    .A2(_06419_));
 sg13g2_buf_1 _24997_ (.A(_06417_),
    .X(_06421_));
 sg13g2_nand2_1 _24998_ (.Y(_06422_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net340));
 sg13g2_o21ai_1 _24999_ (.B1(_06422_),
    .Y(_02388_),
    .A1(net470),
    .A2(net341));
 sg13g2_nand2_1 _25000_ (.Y(_06423_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net340));
 sg13g2_o21ai_1 _25001_ (.B1(_06423_),
    .Y(_02389_),
    .A1(net467),
    .A2(net341));
 sg13g2_nand2_1 _25002_ (.Y(_06424_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net340));
 sg13g2_o21ai_1 _25003_ (.B1(_06424_),
    .Y(_02390_),
    .A1(net409),
    .A2(net341));
 sg13g2_nand2_1 _25004_ (.Y(_06425_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net340));
 sg13g2_o21ai_1 _25005_ (.B1(_06425_),
    .Y(_02391_),
    .A1(net468),
    .A2(net341));
 sg13g2_nand2_1 _25006_ (.Y(_06426_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(_06421_));
 sg13g2_o21ai_1 _25007_ (.B1(_06426_),
    .Y(_02392_),
    .A1(net407),
    .A2(net341));
 sg13g2_nand2_1 _25008_ (.Y(_06427_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net340));
 sg13g2_o21ai_1 _25009_ (.B1(_06427_),
    .Y(_02393_),
    .A1(net408),
    .A2(net341));
 sg13g2_nand2_1 _25010_ (.Y(_06428_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(_06421_));
 sg13g2_o21ai_1 _25011_ (.B1(_06428_),
    .Y(_02394_),
    .A1(net471),
    .A2(net341));
 sg13g2_nand2_1 _25012_ (.Y(_06429_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net340));
 sg13g2_o21ai_1 _25013_ (.B1(_06429_),
    .Y(_02395_),
    .A1(net542),
    .A2(net341));
 sg13g2_mux2_1 _25014_ (.A0(_04447_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net342),
    .X(_02396_));
 sg13g2_nand2_1 _25015_ (.Y(_06430_),
    .A(\cpu.icache.r_tag[6][7] ),
    .B(net340));
 sg13g2_o21ai_1 _25016_ (.B1(_06430_),
    .Y(_02397_),
    .A1(net1029),
    .A2(_06419_));
 sg13g2_nand2_1 _25017_ (.Y(_06431_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(net340));
 sg13g2_o21ai_1 _25018_ (.B1(_06431_),
    .Y(_02398_),
    .A1(_04096_),
    .A2(net342));
 sg13g2_nand2_1 _25019_ (.Y(_06432_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(_06417_));
 sg13g2_o21ai_1 _25020_ (.B1(_06432_),
    .Y(_02399_),
    .A1(net888),
    .A2(_06418_));
 sg13g2_mux2_1 _25021_ (.A0(_04570_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(_06418_),
    .X(_02400_));
 sg13g2_nand2_1 _25022_ (.Y(_06433_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06417_));
 sg13g2_o21ai_1 _25023_ (.B1(_06433_),
    .Y(_02401_),
    .A1(net1030),
    .A2(net342));
 sg13g2_nand2_1 _25024_ (.Y(_06434_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06417_));
 sg13g2_o21ai_1 _25025_ (.B1(_06434_),
    .Y(_02402_),
    .A1(_08152_),
    .A2(net342));
 sg13g2_nand2_1 _25026_ (.Y(_06435_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06417_));
 sg13g2_o21ai_1 _25027_ (.B1(_06435_),
    .Y(_02403_),
    .A1(net478),
    .A2(net342));
 sg13g2_nand2_1 _25028_ (.Y(_06436_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06417_));
 sg13g2_o21ai_1 _25029_ (.B1(_06436_),
    .Y(_02404_),
    .A1(net469),
    .A2(net342));
 sg13g2_nand2_1 _25030_ (.Y(_06437_),
    .A(net697),
    .B(_06313_));
 sg13g2_buf_2 _25031_ (.A(_06437_),
    .X(_06438_));
 sg13g2_buf_1 _25032_ (.A(_06438_),
    .X(_06439_));
 sg13g2_mux2_1 _25033_ (.A0(_04412_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net414),
    .X(_02405_));
 sg13g2_buf_1 _25034_ (.A(_06438_),
    .X(_06440_));
 sg13g2_nand2_1 _25035_ (.Y(_06441_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net414));
 sg13g2_o21ai_1 _25036_ (.B1(_06441_),
    .Y(_02406_),
    .A1(net466),
    .A2(net413));
 sg13g2_buf_1 _25037_ (.A(_06438_),
    .X(_06442_));
 sg13g2_nand2_1 _25038_ (.Y(_06443_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net412));
 sg13g2_o21ai_1 _25039_ (.B1(_06443_),
    .Y(_02407_),
    .A1(net470),
    .A2(net413));
 sg13g2_nand2_1 _25040_ (.Y(_06444_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net412));
 sg13g2_o21ai_1 _25041_ (.B1(_06444_),
    .Y(_02408_),
    .A1(_08403_),
    .A2(net413));
 sg13g2_nand2_1 _25042_ (.Y(_06445_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(_06442_));
 sg13g2_o21ai_1 _25043_ (.B1(_06445_),
    .Y(_02409_),
    .A1(net409),
    .A2(_06440_));
 sg13g2_nand2_1 _25044_ (.Y(_06446_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net412));
 sg13g2_o21ai_1 _25045_ (.B1(_06446_),
    .Y(_02410_),
    .A1(_08380_),
    .A2(net413));
 sg13g2_nand2_1 _25046_ (.Y(_06447_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net412));
 sg13g2_o21ai_1 _25047_ (.B1(_06447_),
    .Y(_02411_),
    .A1(net407),
    .A2(net413));
 sg13g2_nand2_1 _25048_ (.Y(_06448_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(_06442_));
 sg13g2_o21ai_1 _25049_ (.B1(_06448_),
    .Y(_02412_),
    .A1(_08228_),
    .A2(_06440_));
 sg13g2_nand2_1 _25050_ (.Y(_06449_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net412));
 sg13g2_o21ai_1 _25051_ (.B1(_06449_),
    .Y(_02413_),
    .A1(net471),
    .A2(net413));
 sg13g2_nand2_1 _25052_ (.Y(_06450_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net412));
 sg13g2_o21ai_1 _25053_ (.B1(_06450_),
    .Y(_02414_),
    .A1(net542),
    .A2(net413));
 sg13g2_mux2_1 _25054_ (.A0(_04447_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net414),
    .X(_02415_));
 sg13g2_nand2_1 _25055_ (.Y(_06451_),
    .A(\cpu.icache.r_tag[7][7] ),
    .B(net412));
 sg13g2_o21ai_1 _25056_ (.B1(_06451_),
    .Y(_02416_),
    .A1(net1029),
    .A2(net413));
 sg13g2_nand2_1 _25057_ (.Y(_06452_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net412));
 sg13g2_o21ai_1 _25058_ (.B1(_06452_),
    .Y(_02417_),
    .A1(_04096_),
    .A2(net414));
 sg13g2_nand2_1 _25059_ (.Y(_06453_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(_06438_));
 sg13g2_o21ai_1 _25060_ (.B1(_06453_),
    .Y(_02418_),
    .A1(net888),
    .A2(net414));
 sg13g2_mux2_1 _25061_ (.A0(_04570_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(_06439_),
    .X(_02419_));
 sg13g2_nand2_1 _25062_ (.Y(_06454_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06438_));
 sg13g2_o21ai_1 _25063_ (.B1(_06454_),
    .Y(_02420_),
    .A1(net1030),
    .A2(net414));
 sg13g2_nand2_1 _25064_ (.Y(_06455_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06438_));
 sg13g2_o21ai_1 _25065_ (.B1(_06455_),
    .Y(_02421_),
    .A1(net474),
    .A2(net414));
 sg13g2_nand2_1 _25066_ (.Y(_06456_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06438_));
 sg13g2_o21ai_1 _25067_ (.B1(_06456_),
    .Y(_02422_),
    .A1(net478),
    .A2(_06439_));
 sg13g2_nand2_1 _25068_ (.Y(_06457_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06438_));
 sg13g2_o21ai_1 _25069_ (.B1(_06457_),
    .Y(_02423_),
    .A1(net469),
    .A2(net414));
 sg13g2_nand2_1 _25070_ (.Y(_06458_),
    .A(net183),
    .B(net554));
 sg13g2_buf_1 _25071_ (.A(_06458_),
    .X(_06459_));
 sg13g2_buf_1 _25072_ (.A(_06459_),
    .X(_06460_));
 sg13g2_buf_1 _25073_ (.A(_06459_),
    .X(_06461_));
 sg13g2_nand2_1 _25074_ (.Y(_06462_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(net98));
 sg13g2_o21ai_1 _25075_ (.B1(_06462_),
    .Y(_02433_),
    .A1(net872),
    .A2(net99));
 sg13g2_nand2_1 _25076_ (.Y(_06463_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(net98));
 sg13g2_o21ai_1 _25077_ (.B1(_06463_),
    .Y(_02434_),
    .A1(_11702_),
    .A2(net99));
 sg13g2_mux2_1 _25078_ (.A0(_09937_),
    .A1(\cpu.intr.r_clock_cmp[11] ),
    .S(net99),
    .X(_02435_));
 sg13g2_mux2_1 _25079_ (.A0(_09942_),
    .A1(\cpu.intr.r_clock_cmp[12] ),
    .S(net99),
    .X(_02436_));
 sg13g2_nand2_1 _25080_ (.Y(_06464_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(net98));
 sg13g2_o21ai_1 _25081_ (.B1(_06464_),
    .Y(_02437_),
    .A1(_11737_),
    .A2(net99));
 sg13g2_nand2_1 _25082_ (.Y(_06465_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(net98));
 sg13g2_o21ai_1 _25083_ (.B1(_06465_),
    .Y(_02438_),
    .A1(_11747_),
    .A2(net99));
 sg13g2_mux2_1 _25084_ (.A0(_09958_),
    .A1(\cpu.intr.r_clock_cmp[15] ),
    .S(_06461_),
    .X(_02439_));
 sg13g2_nand2_1 _25085_ (.Y(_06466_),
    .A(net183),
    .B(net553));
 sg13g2_buf_1 _25086_ (.A(_06466_),
    .X(_06467_));
 sg13g2_buf_1 _25087_ (.A(_06467_),
    .X(_06468_));
 sg13g2_buf_1 _25088_ (.A(_06467_),
    .X(_06469_));
 sg13g2_nand2_1 _25089_ (.Y(_06470_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(net96));
 sg13g2_o21ai_1 _25090_ (.B1(_06470_),
    .Y(_02440_),
    .A1(net872),
    .A2(net97));
 sg13g2_mux2_1 _25091_ (.A0(net871),
    .A1(\cpu.intr.r_clock_cmp[17] ),
    .S(_06468_),
    .X(_02441_));
 sg13g2_mux2_1 _25092_ (.A0(net870),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(net97),
    .X(_02442_));
 sg13g2_nand2_1 _25093_ (.Y(_06471_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(net96));
 sg13g2_o21ai_1 _25094_ (.B1(_06471_),
    .Y(_02443_),
    .A1(net849),
    .A2(net97));
 sg13g2_mux2_1 _25095_ (.A0(net871),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .S(net98),
    .X(_02444_));
 sg13g2_mux2_1 _25096_ (.A0(net819),
    .A1(\cpu.intr.r_clock_cmp[20] ),
    .S(_06469_),
    .X(_02445_));
 sg13g2_mux2_1 _25097_ (.A0(net818),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .S(_06469_),
    .X(_02446_));
 sg13g2_nand2_1 _25098_ (.Y(_06472_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(net96));
 sg13g2_o21ai_1 _25099_ (.B1(_06472_),
    .Y(_02447_),
    .A1(net845),
    .A2(net97));
 sg13g2_nand2_1 _25100_ (.Y(_06473_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(net96));
 sg13g2_o21ai_1 _25101_ (.B1(_06473_),
    .Y(_02448_),
    .A1(net848),
    .A2(_06468_));
 sg13g2_inv_1 _25102_ (.Y(_06474_),
    .A(_09921_));
 sg13g2_nand2_1 _25103_ (.Y(_06475_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_06467_));
 sg13g2_o21ai_1 _25104_ (.B1(_06475_),
    .Y(_02449_),
    .A1(_06474_),
    .A2(net97));
 sg13g2_mux2_1 _25105_ (.A0(_09926_),
    .A1(\cpu.intr.r_clock_cmp[25] ),
    .S(net96),
    .X(_02450_));
 sg13g2_nand2_1 _25106_ (.Y(_06476_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_06467_));
 sg13g2_o21ai_1 _25107_ (.B1(_06476_),
    .Y(_02451_),
    .A1(_11702_),
    .A2(net97));
 sg13g2_mux2_1 _25108_ (.A0(_09937_),
    .A1(\cpu.intr.r_clock_cmp[27] ),
    .S(net96),
    .X(_02452_));
 sg13g2_mux2_1 _25109_ (.A0(_09942_),
    .A1(\cpu.intr.r_clock_cmp[28] ),
    .S(net96),
    .X(_02453_));
 sg13g2_nand2_1 _25110_ (.Y(_06477_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_06467_));
 sg13g2_o21ai_1 _25111_ (.B1(_06477_),
    .Y(_02454_),
    .A1(_11737_),
    .A2(net97));
 sg13g2_mux2_1 _25112_ (.A0(net870),
    .A1(\cpu.intr.r_clock_cmp[2] ),
    .S(net98),
    .X(_02455_));
 sg13g2_nand2_1 _25113_ (.Y(_06478_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_06467_));
 sg13g2_o21ai_1 _25114_ (.B1(_06478_),
    .Y(_02456_),
    .A1(_11747_),
    .A2(net97));
 sg13g2_mux2_1 _25115_ (.A0(_09958_),
    .A1(\cpu.intr.r_clock_cmp[31] ),
    .S(net96),
    .X(_02457_));
 sg13g2_nand2_1 _25116_ (.Y(_06479_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_06459_));
 sg13g2_o21ai_1 _25117_ (.B1(_06479_),
    .Y(_02458_),
    .A1(net849),
    .A2(net99));
 sg13g2_mux2_1 _25118_ (.A0(net819),
    .A1(\cpu.intr.r_clock_cmp[4] ),
    .S(_06461_),
    .X(_02459_));
 sg13g2_mux2_1 _25119_ (.A0(net818),
    .A1(\cpu.intr.r_clock_cmp[5] ),
    .S(net98),
    .X(_02460_));
 sg13g2_nand2_1 _25120_ (.Y(_06480_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_06459_));
 sg13g2_o21ai_1 _25121_ (.B1(_06480_),
    .Y(_02461_),
    .A1(net845),
    .A2(_06460_));
 sg13g2_nand2_1 _25122_ (.Y(_06481_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_06459_));
 sg13g2_o21ai_1 _25123_ (.B1(_06481_),
    .Y(_02462_),
    .A1(net848),
    .A2(net99));
 sg13g2_nand2_1 _25124_ (.Y(_06482_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_06459_));
 sg13g2_o21ai_1 _25125_ (.B1(_06482_),
    .Y(_02463_),
    .A1(_06474_),
    .A2(_06460_));
 sg13g2_mux2_1 _25126_ (.A0(_09926_),
    .A1(\cpu.intr.r_clock_cmp[9] ),
    .S(net98),
    .X(_02464_));
 sg13g2_nand2_1 _25127_ (.Y(_06483_),
    .A(net183),
    .B(_04928_));
 sg13g2_buf_1 _25128_ (.A(_06483_),
    .X(_06484_));
 sg13g2_buf_1 _25129_ (.A(_06484_),
    .X(_06485_));
 sg13g2_buf_1 _25130_ (.A(_06484_),
    .X(_06486_));
 sg13g2_nand2_1 _25131_ (.Y(_06487_),
    .A(\cpu.intr.r_timer_reload[0] ),
    .B(net94));
 sg13g2_o21ai_1 _25132_ (.B1(_06487_),
    .Y(_02488_),
    .A1(net872),
    .A2(net95));
 sg13g2_nand2_1 _25133_ (.Y(_06488_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net94));
 sg13g2_o21ai_1 _25134_ (.B1(_06488_),
    .Y(_02489_),
    .A1(_11702_),
    .A2(net95));
 sg13g2_mux2_1 _25135_ (.A0(_09937_),
    .A1(\cpu.intr.r_timer_reload[11] ),
    .S(net95),
    .X(_02490_));
 sg13g2_mux2_1 _25136_ (.A0(_09942_),
    .A1(\cpu.intr.r_timer_reload[12] ),
    .S(net95),
    .X(_02491_));
 sg13g2_nand2_1 _25137_ (.Y(_06489_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net94));
 sg13g2_o21ai_1 _25138_ (.B1(_06489_),
    .Y(_02492_),
    .A1(_11737_),
    .A2(net95));
 sg13g2_nand2_1 _25139_ (.Y(_06490_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net94));
 sg13g2_o21ai_1 _25140_ (.B1(_06490_),
    .Y(_02493_),
    .A1(_11747_),
    .A2(net95));
 sg13g2_mux2_1 _25141_ (.A0(_09958_),
    .A1(\cpu.intr.r_timer_reload[15] ),
    .S(net94),
    .X(_02494_));
 sg13g2_mux2_1 _25142_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net821),
    .S(_09813_),
    .X(_02495_));
 sg13g2_mux2_1 _25143_ (.A0(\cpu.intr.r_timer_reload[17] ),
    .A1(net847),
    .S(net153),
    .X(_02496_));
 sg13g2_mux2_1 _25144_ (.A0(\cpu.intr.r_timer_reload[18] ),
    .A1(net846),
    .S(net153),
    .X(_02497_));
 sg13g2_inv_1 _25145_ (.Y(_06491_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25146_ (.B1(_09834_),
    .Y(_02498_),
    .A1(_06491_),
    .A2(net154));
 sg13g2_mux2_1 _25147_ (.A0(net871),
    .A1(\cpu.intr.r_timer_reload[1] ),
    .S(net94),
    .X(_02499_));
 sg13g2_o21ai_1 _25148_ (.B1(_09841_),
    .Y(_02500_),
    .A1(_09835_),
    .A2(net154));
 sg13g2_inv_1 _25149_ (.Y(_06492_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25150_ (.B1(_09847_),
    .Y(_02501_),
    .A1(_06492_),
    .A2(net154));
 sg13g2_inv_1 _25151_ (.Y(_06493_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25152_ (.B1(_09852_),
    .Y(_02502_),
    .A1(_06493_),
    .A2(_09812_));
 sg13g2_mux2_1 _25153_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net1005),
    .S(net153),
    .X(_02503_));
 sg13g2_mux2_1 _25154_ (.A0(net870),
    .A1(\cpu.intr.r_timer_reload[2] ),
    .S(net94),
    .X(_02504_));
 sg13g2_nand2_1 _25155_ (.Y(_06494_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(_06484_));
 sg13g2_o21ai_1 _25156_ (.B1(_06494_),
    .Y(_02505_),
    .A1(net849),
    .A2(net95));
 sg13g2_mux2_1 _25157_ (.A0(net819),
    .A1(\cpu.intr.r_timer_reload[4] ),
    .S(_06486_),
    .X(_02506_));
 sg13g2_mux2_1 _25158_ (.A0(net818),
    .A1(\cpu.intr.r_timer_reload[5] ),
    .S(_06486_),
    .X(_02507_));
 sg13g2_nand2_1 _25159_ (.Y(_06495_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(_06484_));
 sg13g2_o21ai_1 _25160_ (.B1(_06495_),
    .Y(_02508_),
    .A1(net845),
    .A2(_06485_));
 sg13g2_nand2_1 _25161_ (.Y(_06496_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_06484_));
 sg13g2_o21ai_1 _25162_ (.B1(_06496_),
    .Y(_02509_),
    .A1(net848),
    .A2(_06485_));
 sg13g2_nand2_1 _25163_ (.Y(_06497_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(_06484_));
 sg13g2_o21ai_1 _25164_ (.B1(_06497_),
    .Y(_02510_),
    .A1(_06474_),
    .A2(net95));
 sg13g2_mux2_1 _25165_ (.A0(_09926_),
    .A1(\cpu.intr.r_timer_reload[9] ),
    .S(net94),
    .X(_02511_));
 sg13g2_inv_1 _25166_ (.Y(_06498_),
    .A(_09580_));
 sg13g2_nor2_1 _25167_ (.A(_09589_),
    .B(_09577_),
    .Y(_06499_));
 sg13g2_nor4_2 _25168_ (.A(_11549_),
    .B(_11569_),
    .C(_09601_),
    .Y(_06500_),
    .D(\cpu.qspi.r_state[11] ));
 sg13g2_nor3_1 _25169_ (.A(_11570_),
    .B(_11551_),
    .C(_11571_),
    .Y(_06501_));
 sg13g2_nand4_1 _25170_ (.B(_06499_),
    .C(_06500_),
    .A(_09576_),
    .Y(_06502_),
    .D(_06501_));
 sg13g2_a21oi_1 _25171_ (.A1(_09129_),
    .A2(_09623_),
    .Y(_06503_),
    .B1(_06502_));
 sg13g2_buf_1 _25172_ (.A(_06503_),
    .X(_06504_));
 sg13g2_and2_1 _25173_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_09615_),
    .X(_06505_));
 sg13g2_a221oi_1 _25174_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06505_),
    .B1(_09619_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06506_),
    .A2(_09617_));
 sg13g2_nor2_1 _25175_ (.A(_09588_),
    .B(net1082),
    .Y(_06507_));
 sg13g2_nor2_1 _25176_ (.A(_09600_),
    .B(_09593_),
    .Y(_06508_));
 sg13g2_nand2_1 _25177_ (.Y(_06509_),
    .A(_06507_),
    .B(_06508_));
 sg13g2_a221oi_1 _25178_ (.B2(_06509_),
    .C1(_09598_),
    .B1(_00183_),
    .A1(_09627_),
    .Y(_06510_),
    .A2(_06498_));
 sg13g2_o21ai_1 _25179_ (.B1(_06510_),
    .Y(_06511_),
    .A1(_09670_),
    .A2(_06506_));
 sg13g2_nand2_1 _25180_ (.Y(_06512_),
    .A(_06504_),
    .B(_06511_));
 sg13g2_o21ai_1 _25181_ (.B1(_06512_),
    .Y(_02512_),
    .A1(_06498_),
    .A2(_06504_));
 sg13g2_inv_1 _25182_ (.Y(_06513_),
    .A(_09581_));
 sg13g2_and2_1 _25183_ (.A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_09615_),
    .X(_06514_));
 sg13g2_a221oi_1 _25184_ (.B2(\cpu.qspi.r_read_delay[0][1] ),
    .C1(_06514_),
    .B1(_09619_),
    .A1(\cpu.qspi.r_read_delay[2][1] ),
    .Y(_06515_),
    .A2(_09617_));
 sg13g2_nor2_1 _25185_ (.A(_09627_),
    .B(_06509_),
    .Y(_06516_));
 sg13g2_xor2_1 _25186_ (.B(_09581_),
    .A(_09580_),
    .X(_06517_));
 sg13g2_nor2_1 _25187_ (.A(_06516_),
    .B(_06517_),
    .Y(_06518_));
 sg13g2_a21oi_1 _25188_ (.A1(_09670_),
    .A2(_06516_),
    .Y(_06519_),
    .B1(_06518_));
 sg13g2_o21ai_1 _25189_ (.B1(_06519_),
    .Y(_06520_),
    .A1(_09670_),
    .A2(_06515_));
 sg13g2_o21ai_1 _25190_ (.B1(net27),
    .Y(_06521_),
    .A1(_09598_),
    .A2(_06520_));
 sg13g2_o21ai_1 _25191_ (.B1(_06521_),
    .Y(_02513_),
    .A1(_06513_),
    .A2(net27));
 sg13g2_nor2_1 _25192_ (.A(_09580_),
    .B(_09581_),
    .Y(_06522_));
 sg13g2_xor2_1 _25193_ (.B(_06522_),
    .A(_00184_),
    .X(_06523_));
 sg13g2_and2_1 _25194_ (.A(_06507_),
    .B(_06508_),
    .X(_06524_));
 sg13g2_buf_1 _25195_ (.A(_06524_),
    .X(_06525_));
 sg13g2_o21ai_1 _25196_ (.B1(_09671_),
    .Y(_06526_),
    .A1(_09627_),
    .A2(_06525_));
 sg13g2_a22oi_1 _25197_ (.Y(_06527_),
    .B1(_06523_),
    .B2(_06526_),
    .A2(_06516_),
    .A1(_09669_));
 sg13g2_a22oi_1 _25198_ (.Y(_06528_),
    .B1(_09615_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09617_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25199_ (.Y(_06529_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09619_));
 sg13g2_a21oi_1 _25200_ (.A1(_06528_),
    .A2(_06529_),
    .Y(_06530_),
    .B1(_09670_));
 sg13g2_nor3_1 _25201_ (.A(_09598_),
    .B(_06527_),
    .C(_06530_),
    .Y(_06531_));
 sg13g2_nor2_1 _25202_ (.A(_09582_),
    .B(net27),
    .Y(_06532_));
 sg13g2_a21oi_1 _25203_ (.A1(net27),
    .A2(_06531_),
    .Y(_02514_),
    .B1(_06532_));
 sg13g2_a21oi_1 _25204_ (.A1(_09671_),
    .A2(_06525_),
    .Y(_06533_),
    .B1(_09583_));
 sg13g2_nand2b_1 _25205_ (.Y(_06534_),
    .B(net27),
    .A_N(_06533_));
 sg13g2_nand2_1 _25206_ (.Y(_06535_),
    .A(_09671_),
    .B(_06525_));
 sg13g2_a22oi_1 _25207_ (.Y(_06536_),
    .B1(_09615_),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(_09617_),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_nand2_1 _25208_ (.Y(_06537_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_09619_));
 sg13g2_nand2_1 _25209_ (.Y(_06538_),
    .A(_06536_),
    .B(_06537_));
 sg13g2_a22oi_1 _25210_ (.Y(_06539_),
    .B1(_06538_),
    .B2(_09669_),
    .A2(_06535_),
    .A1(_09585_));
 sg13g2_nor2b_1 _25211_ (.A(_06539_),
    .B_N(net27),
    .Y(_06540_));
 sg13g2_a21o_1 _25212_ (.A2(_06534_),
    .A1(\cpu.qspi.r_count[3] ),
    .B1(_06540_),
    .X(_02515_));
 sg13g2_and2_1 _25213_ (.A(_09585_),
    .B(_06509_),
    .X(_06541_));
 sg13g2_nor3_1 _25214_ (.A(_09579_),
    .B(_09585_),
    .C(_06516_),
    .Y(_06542_));
 sg13g2_a21oi_1 _25215_ (.A1(_09579_),
    .A2(_06541_),
    .Y(_06543_),
    .B1(_06542_));
 sg13g2_nor2_1 _25216_ (.A(\cpu.qspi.r_count[4] ),
    .B(net27),
    .Y(_06544_));
 sg13g2_a21oi_1 _25217_ (.A1(net27),
    .A2(_06543_),
    .Y(_02516_),
    .B1(_06544_));
 sg13g2_nand2_1 _25218_ (.Y(_06545_),
    .A(_09734_),
    .B(_06093_));
 sg13g2_buf_1 _25219_ (.A(_06545_),
    .X(_06546_));
 sg13g2_nor2_1 _25220_ (.A(_04693_),
    .B(net137),
    .Y(_06547_));
 sg13g2_buf_1 _25221_ (.A(_06547_),
    .X(_06548_));
 sg13g2_nand2_1 _25222_ (.Y(_06549_),
    .A(net821),
    .B(_06548_));
 sg13g2_nand3_1 _25223_ (.B(_09734_),
    .C(_06093_),
    .A(_08966_),
    .Y(_06550_));
 sg13g2_buf_1 _25224_ (.A(_06550_),
    .X(_06551_));
 sg13g2_nand2_1 _25225_ (.Y(_06552_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06551_));
 sg13g2_a21oi_1 _25226_ (.A1(_06549_),
    .A2(_06552_),
    .Y(_02527_),
    .B1(net688));
 sg13g2_nand2_1 _25227_ (.Y(_06553_),
    .A(net959),
    .B(_06548_));
 sg13g2_nand2_1 _25228_ (.Y(_06554_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06551_));
 sg13g2_a21oi_1 _25229_ (.A1(_06553_),
    .A2(_06554_),
    .Y(_02528_),
    .B1(net688));
 sg13g2_nand2_1 _25230_ (.Y(_06555_),
    .A(net844),
    .B(_06548_));
 sg13g2_nand2_1 _25231_ (.Y(_06556_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06551_));
 sg13g2_nand3_1 _25232_ (.B(_06555_),
    .C(_06556_),
    .A(net622),
    .Y(_02529_));
 sg13g2_nand2_1 _25233_ (.Y(_06557_),
    .A(_06116_),
    .B(_06548_));
 sg13g2_nand2_1 _25234_ (.Y(_06558_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06551_));
 sg13g2_a21oi_1 _25235_ (.A1(_06557_),
    .A2(_06558_),
    .Y(_02530_),
    .B1(net688));
 sg13g2_nor2_1 _25236_ (.A(net557),
    .B(net137),
    .Y(_06559_));
 sg13g2_nand2_1 _25237_ (.Y(_06560_),
    .A(net821),
    .B(_06559_));
 sg13g2_or2_1 _25238_ (.X(_06561_),
    .B(net137),
    .A(_04737_));
 sg13g2_buf_1 _25239_ (.A(_06561_),
    .X(_06562_));
 sg13g2_nand2_1 _25240_ (.Y(_06563_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06562_));
 sg13g2_a21oi_1 _25241_ (.A1(_06560_),
    .A2(_06563_),
    .Y(_02531_),
    .B1(net688));
 sg13g2_nand2_1 _25242_ (.Y(_06564_),
    .A(_12263_),
    .B(_06559_));
 sg13g2_nand2_1 _25243_ (.Y(_06565_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06562_));
 sg13g2_a21oi_1 _25244_ (.A1(_06564_),
    .A2(_06565_),
    .Y(_02532_),
    .B1(net688));
 sg13g2_nand2_1 _25245_ (.Y(_06566_),
    .A(_12292_),
    .B(_06559_));
 sg13g2_nand2_1 _25246_ (.Y(_06567_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06562_));
 sg13g2_nand3_1 _25247_ (.B(_06566_),
    .C(_06567_),
    .A(net622),
    .Y(_02533_));
 sg13g2_nand2_1 _25248_ (.Y(_06568_),
    .A(net928),
    .B(_06559_));
 sg13g2_nand2_1 _25249_ (.Y(_06569_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06562_));
 sg13g2_buf_1 _25250_ (.A(_09103_),
    .X(_06570_));
 sg13g2_a21oi_1 _25251_ (.A1(_06568_),
    .A2(_06569_),
    .Y(_02534_),
    .B1(net615));
 sg13g2_nor2_1 _25252_ (.A(net558),
    .B(net137),
    .Y(_06571_));
 sg13g2_buf_2 _25253_ (.A(_06571_),
    .X(_06572_));
 sg13g2_nand2_1 _25254_ (.Y(_06573_),
    .A(_05565_),
    .B(_06572_));
 sg13g2_or2_1 _25255_ (.X(_06574_),
    .B(net137),
    .A(net558));
 sg13g2_buf_1 _25256_ (.A(_06574_),
    .X(_06575_));
 sg13g2_nand2_1 _25257_ (.Y(_06576_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06575_));
 sg13g2_a21oi_1 _25258_ (.A1(_06573_),
    .A2(_06576_),
    .Y(_02535_),
    .B1(_06570_));
 sg13g2_nand2_1 _25259_ (.Y(_06577_),
    .A(_12263_),
    .B(_06572_));
 sg13g2_nand2_1 _25260_ (.Y(_06578_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06575_));
 sg13g2_a21oi_1 _25261_ (.A1(_06577_),
    .A2(_06578_),
    .Y(_02536_),
    .B1(net615));
 sg13g2_nand2_1 _25262_ (.Y(_06579_),
    .A(_12292_),
    .B(_06572_));
 sg13g2_nand2_1 _25263_ (.Y(_06580_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06575_));
 sg13g2_nand3_1 _25264_ (.B(_06579_),
    .C(_06580_),
    .A(net622),
    .Y(_02537_));
 sg13g2_nand2_1 _25265_ (.Y(_06581_),
    .A(_06116_),
    .B(_06572_));
 sg13g2_nand2_1 _25266_ (.Y(_06582_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06575_));
 sg13g2_a21oi_1 _25267_ (.A1(_06581_),
    .A2(_06582_),
    .Y(_02538_),
    .B1(net615));
 sg13g2_nand2_1 _25268_ (.Y(_06583_),
    .A(_06498_),
    .B(_09581_));
 sg13g2_mux2_1 _25269_ (.A0(_06583_),
    .A1(_09581_),
    .S(net128),
    .X(_06584_));
 sg13g2_nand2_1 _25270_ (.Y(_06585_),
    .A(net1082),
    .B(_09578_));
 sg13g2_a21o_1 _25271_ (.A2(_06585_),
    .A1(_00183_),
    .B1(_09581_),
    .X(_06586_));
 sg13g2_o21ai_1 _25272_ (.B1(_06586_),
    .Y(_06587_),
    .A1(net1082),
    .A2(_06584_));
 sg13g2_nand2b_1 _25273_ (.Y(_06588_),
    .B(net128),
    .A_N(_09581_));
 sg13g2_a21oi_1 _25274_ (.A1(_06583_),
    .A2(_06588_),
    .Y(_06589_),
    .B1(_09604_));
 sg13g2_nand3_1 _25275_ (.B(_09580_),
    .C(_09578_),
    .A(net1082),
    .Y(_06590_));
 sg13g2_o21ai_1 _25276_ (.B1(_06590_),
    .Y(_06591_),
    .A1(_09578_),
    .A2(_06583_));
 sg13g2_nor3_1 _25277_ (.A(_09582_),
    .B(_06589_),
    .C(_06591_),
    .Y(_06592_));
 sg13g2_a21o_1 _25278_ (.A2(_06587_),
    .A1(_09582_),
    .B1(_06592_),
    .X(_06593_));
 sg13g2_o21ai_1 _25279_ (.B1(_06593_),
    .Y(_06594_),
    .A1(_09600_),
    .A2(net1082));
 sg13g2_buf_1 _25280_ (.A(net1015),
    .X(_06595_));
 sg13g2_buf_1 _25281_ (.A(net129),
    .X(_06596_));
 sg13g2_mux2_1 _25282_ (.A0(_09497_),
    .A1(_09503_),
    .S(_06596_),
    .X(_06597_));
 sg13g2_nand2_1 _25283_ (.Y(_06598_),
    .A(net1015),
    .B(_10681_));
 sg13g2_o21ai_1 _25284_ (.B1(_06598_),
    .Y(_06599_),
    .A1(net781),
    .A2(_06597_));
 sg13g2_nand2_1 _25285_ (.Y(_06600_),
    .A(_11569_),
    .B(_06599_));
 sg13g2_nor2b_1 _25286_ (.A(net128),
    .B_N(_09601_),
    .Y(_06601_));
 sg13g2_nor2b_1 _25287_ (.A(_11794_),
    .B_N(_11677_),
    .Y(_06602_));
 sg13g2_nor2_1 _25288_ (.A(_11767_),
    .B(_06602_),
    .Y(_06603_));
 sg13g2_and2_1 _25289_ (.A(_11767_),
    .B(_11680_),
    .X(_06604_));
 sg13g2_mux2_1 _25290_ (.A0(_05020_),
    .A1(_04664_),
    .S(_11655_),
    .X(_06605_));
 sg13g2_nor2_1 _25291_ (.A(_11655_),
    .B(_05013_),
    .Y(_06606_));
 sg13g2_a21oi_1 _25292_ (.A1(_11655_),
    .A2(_04635_),
    .Y(_06607_),
    .B1(_06606_));
 sg13g2_a22oi_1 _25293_ (.Y(_06608_),
    .B1(_06607_),
    .B2(_11652_),
    .A2(_06605_),
    .A1(_11677_));
 sg13g2_and2_1 _25294_ (.A(_11655_),
    .B(_11677_),
    .X(_06609_));
 sg13g2_nor2b_1 _25295_ (.A(_11729_),
    .B_N(_11652_),
    .Y(_06610_));
 sg13g2_a221oi_1 _25296_ (.B2(_05330_),
    .C1(net979),
    .B1(_06610_),
    .A1(_04656_),
    .Y(_06611_),
    .A2(_06609_));
 sg13g2_a21oi_1 _25297_ (.A1(net979),
    .A2(_06608_),
    .Y(_06612_),
    .B1(_06611_));
 sg13g2_a221oi_1 _25298_ (.B2(_04644_),
    .C1(_06612_),
    .B1(_06604_),
    .A1(_05323_),
    .Y(_06613_),
    .A2(_06603_));
 sg13g2_buf_1 _25299_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06614_));
 sg13g2_nand2_1 _25300_ (.Y(_06615_),
    .A(net1038),
    .B(_09130_));
 sg13g2_o21ai_1 _25301_ (.B1(_06615_),
    .Y(_06616_),
    .A1(_09130_),
    .A2(_11607_));
 sg13g2_a221oi_1 _25302_ (.B2(_11571_),
    .C1(_11549_),
    .B1(_06616_),
    .A1(_09629_),
    .Y(_06617_),
    .A2(_06614_));
 sg13g2_o21ai_1 _25303_ (.B1(_06617_),
    .Y(_06618_),
    .A1(_11552_),
    .A2(_06613_));
 sg13g2_nor2_1 _25304_ (.A(_06601_),
    .B(_06618_),
    .Y(_06619_));
 sg13g2_mux2_1 _25305_ (.A0(_09235_),
    .A1(_09215_),
    .S(net129),
    .X(_06620_));
 sg13g2_nor2_1 _25306_ (.A(net1015),
    .B(_06620_),
    .Y(_06621_));
 sg13g2_a21oi_1 _25307_ (.A1(net781),
    .A2(_08152_),
    .Y(_06622_),
    .B1(_06621_));
 sg13g2_buf_1 _25308_ (.A(_09609_),
    .X(_06623_));
 sg13g2_mux2_1 _25309_ (.A0(_09285_),
    .A1(_09291_),
    .S(net129),
    .X(_06624_));
 sg13g2_nand2_1 _25310_ (.Y(_06625_),
    .A(_09609_),
    .B(_06624_));
 sg13g2_o21ai_1 _25311_ (.B1(_06625_),
    .Y(_06626_),
    .A1(net780),
    .A2(_08276_));
 sg13g2_a22oi_1 _25312_ (.Y(_06627_),
    .B1(_06626_),
    .B2(_11570_),
    .A2(_06622_),
    .A1(_11551_));
 sg13g2_nand4_1 _25313_ (.B(_06600_),
    .C(_06619_),
    .A(_06594_),
    .Y(_06628_),
    .D(_06627_));
 sg13g2_xor2_1 _25314_ (.B(_09622_),
    .A(net128),
    .X(_06629_));
 sg13g2_nand2_1 _25315_ (.Y(_06630_),
    .A(_06501_),
    .B(_06508_));
 sg13g2_nor2_1 _25316_ (.A(_09598_),
    .B(_06630_),
    .Y(_06631_));
 sg13g2_nor2b_1 _25317_ (.A(net1082),
    .B_N(_06500_),
    .Y(_06632_));
 sg13g2_and3_1 _25318_ (.X(_06633_),
    .A(_09603_),
    .B(_06631_),
    .C(_06632_));
 sg13g2_buf_1 _25319_ (.A(_06633_),
    .X(_06634_));
 sg13g2_mux2_1 _25320_ (.A0(_06628_),
    .A1(_06629_),
    .S(_06634_),
    .X(_06635_));
 sg13g2_and2_1 _25321_ (.A(\cpu.qspi.r_mask[1] ),
    .B(_09615_),
    .X(_06636_));
 sg13g2_a221oi_1 _25322_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06636_),
    .B1(_09619_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06637_),
    .A2(_09617_));
 sg13g2_nor3_2 _25323_ (.A(_09588_),
    .B(_09589_),
    .C(_09577_),
    .Y(_06638_));
 sg13g2_nor2_1 _25324_ (.A(_09669_),
    .B(_09627_),
    .Y(_06639_));
 sg13g2_nand3_1 _25325_ (.B(_06638_),
    .C(_06639_),
    .A(_09576_),
    .Y(_06640_));
 sg13g2_a21oi_1 _25326_ (.A1(_11549_),
    .A2(_06637_),
    .Y(_06641_),
    .B1(_06640_));
 sg13g2_buf_2 _25327_ (.A(_06641_),
    .X(_06642_));
 sg13g2_mux2_1 _25328_ (.A0(net11),
    .A1(_06635_),
    .S(_06642_),
    .X(_02543_));
 sg13g2_or2_1 _25329_ (.X(_06643_),
    .B(_06634_),
    .A(_11549_));
 sg13g2_buf_1 _25330_ (.A(_06643_),
    .X(_06644_));
 sg13g2_mux2_1 _25331_ (.A0(_05044_),
    .A1(_05128_),
    .S(net980),
    .X(_06645_));
 sg13g2_a22oi_1 _25332_ (.Y(_06646_),
    .B1(_06645_),
    .B2(net979),
    .A2(_05111_),
    .A1(_11680_));
 sg13g2_nand2b_1 _25333_ (.Y(_06647_),
    .B(net984),
    .A_N(_06646_));
 sg13g2_mux4_1 _25334_ (.S0(net980),
    .A0(_05402_),
    .A1(_05118_),
    .A2(_05038_),
    .A3(_05134_),
    .S1(net979),
    .X(_06648_));
 sg13g2_a22oi_1 _25335_ (.Y(_06649_),
    .B1(_06648_),
    .B2(net976),
    .A2(_06603_),
    .A1(_05395_));
 sg13g2_a21oi_1 _25336_ (.A1(_06647_),
    .A2(_06649_),
    .Y(_06650_),
    .B1(_11552_));
 sg13g2_nor3_1 _25337_ (.A(_06601_),
    .B(_06644_),
    .C(_06650_),
    .Y(_06651_));
 sg13g2_nor2_1 _25338_ (.A(_00237_),
    .B(_09571_),
    .Y(_06652_));
 sg13g2_a21o_1 _25339_ (.A2(net93),
    .A1(_09450_),
    .B1(_06652_),
    .X(_06653_));
 sg13g2_mux2_1 _25340_ (.A0(_10718_),
    .A1(_06653_),
    .S(_09609_),
    .X(_06654_));
 sg13g2_mux2_1 _25341_ (.A0(_09350_),
    .A1(_09356_),
    .S(net129),
    .X(_06655_));
 sg13g2_nand2_1 _25342_ (.Y(_06656_),
    .A(net780),
    .B(_06655_));
 sg13g2_o21ai_1 _25343_ (.B1(_06656_),
    .Y(_06657_),
    .A1(_06623_),
    .A2(_08403_));
 sg13g2_a22oi_1 _25344_ (.Y(_06658_),
    .B1(_06657_),
    .B2(_11570_),
    .A2(_06654_),
    .A1(_11569_));
 sg13g2_mux2_1 _25345_ (.A0(_09206_),
    .A1(_09180_),
    .S(net129),
    .X(_06659_));
 sg13g2_nor2_1 _25346_ (.A(net1015),
    .B(_06659_),
    .Y(_06660_));
 sg13g2_a21oi_1 _25347_ (.A1(net781),
    .A2(_08087_),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_buf_1 _25348_ (.A(net1015),
    .X(_06662_));
 sg13g2_mux2_1 _25349_ (.A0(_05363_),
    .A1(_09485_),
    .S(net93),
    .X(_06663_));
 sg13g2_nand2_1 _25350_ (.Y(_06664_),
    .A(net1015),
    .B(_10929_));
 sg13g2_o21ai_1 _25351_ (.B1(_06664_),
    .Y(_06665_),
    .A1(net779),
    .A2(_06663_));
 sg13g2_a22oi_1 _25352_ (.Y(_06666_),
    .B1(_06665_),
    .B2(_11571_),
    .A2(_06661_),
    .A1(_11551_));
 sg13g2_and2_1 _25353_ (.A(_06658_),
    .B(_06666_),
    .X(_06667_));
 sg13g2_a22oi_1 _25354_ (.Y(_06668_),
    .B1(_06651_),
    .B2(_06667_),
    .A2(_06634_),
    .A1(_09622_));
 sg13g2_mux2_1 _25355_ (.A0(net12),
    .A1(_06668_),
    .S(_06642_),
    .X(_02544_));
 sg13g2_inv_1 _25356_ (.Y(_06669_),
    .A(net13));
 sg13g2_inv_1 _25357_ (.Y(_06670_),
    .A(_00185_));
 sg13g2_nand2_1 _25358_ (.Y(_06671_),
    .A(net770),
    .B(net781));
 sg13g2_o21ai_1 _25359_ (.B1(_06671_),
    .Y(_06672_),
    .A1(net779),
    .A2(net632));
 sg13g2_a21oi_1 _25360_ (.A1(_06670_),
    .A2(_06672_),
    .Y(_06673_),
    .B1(_06644_));
 sg13g2_nand2_1 _25361_ (.Y(_06674_),
    .A(net984),
    .B(_05070_));
 sg13g2_a22oi_1 _25362_ (.Y(_06675_),
    .B1(_04950_),
    .B2(_11678_),
    .A2(_04943_),
    .A1(_11652_));
 sg13g2_nand2b_1 _25363_ (.Y(_06676_),
    .B(net980),
    .A_N(_06675_));
 sg13g2_o21ai_1 _25364_ (.B1(_06676_),
    .Y(_06677_),
    .A1(net980),
    .A2(_06674_));
 sg13g2_mux2_1 _25365_ (.A0(_05505_),
    .A1(_05196_),
    .S(net980),
    .X(_06678_));
 sg13g2_nand2b_1 _25366_ (.Y(_06679_),
    .B(_06678_),
    .A_N(net979));
 sg13g2_nand2b_1 _25367_ (.Y(_06680_),
    .B(_11731_),
    .A_N(_05064_));
 sg13g2_nand2_1 _25368_ (.Y(_06681_),
    .A(_06679_),
    .B(_06680_));
 sg13g2_inv_1 _25369_ (.Y(_06682_),
    .A(_06603_));
 sg13g2_nand3_1 _25370_ (.B(_11680_),
    .C(_05190_),
    .A(net984),
    .Y(_06683_));
 sg13g2_o21ai_1 _25371_ (.B1(_06683_),
    .Y(_06684_),
    .A1(_05514_),
    .A2(_06682_));
 sg13g2_a221oi_1 _25372_ (.B2(net976),
    .C1(_06684_),
    .B1(_06681_),
    .A1(net979),
    .Y(_06685_),
    .A2(_06677_));
 sg13g2_nand2b_1 _25373_ (.Y(_06686_),
    .B(_09593_),
    .A_N(_06685_));
 sg13g2_mux2_1 _25374_ (.A0(_09527_),
    .A1(_09533_),
    .S(net129),
    .X(_06687_));
 sg13g2_nand2_1 _25375_ (.Y(_06688_),
    .A(net780),
    .B(_06687_));
 sg13g2_o21ai_1 _25376_ (.B1(_06688_),
    .Y(_06689_),
    .A1(net780),
    .A2(_08196_));
 sg13g2_mux2_1 _25377_ (.A0(net366),
    .A1(_09413_),
    .S(net93),
    .X(_06690_));
 sg13g2_nor2_1 _25378_ (.A(net781),
    .B(_06690_),
    .Y(_06691_));
 sg13g2_a21oi_1 _25379_ (.A1(net779),
    .A2(_08353_),
    .Y(_06692_),
    .B1(_06691_));
 sg13g2_a22oi_1 _25380_ (.Y(_06693_),
    .B1(_06692_),
    .B2(_11551_),
    .A2(_06689_),
    .A1(_11570_));
 sg13g2_mux2_1 _25381_ (.A0(_00239_),
    .A1(_09495_),
    .S(net93),
    .X(_06694_));
 sg13g2_nand2_1 _25382_ (.Y(_06695_),
    .A(net781),
    .B(_10527_));
 sg13g2_o21ai_1 _25383_ (.B1(_06695_),
    .Y(_06696_),
    .A1(net779),
    .A2(_06694_));
 sg13g2_mux2_1 _25384_ (.A0(_00231_),
    .A1(_09510_),
    .S(net93),
    .X(_06697_));
 sg13g2_nand2_1 _25385_ (.Y(_06698_),
    .A(net781),
    .B(_10982_));
 sg13g2_o21ai_1 _25386_ (.B1(_06698_),
    .Y(_06699_),
    .A1(net779),
    .A2(_06697_));
 sg13g2_a22oi_1 _25387_ (.Y(_06700_),
    .B1(_06699_),
    .B2(_11571_),
    .A2(_06696_),
    .A1(_11569_));
 sg13g2_nand4_1 _25388_ (.B(_06686_),
    .C(_06693_),
    .A(_06673_),
    .Y(_06701_),
    .D(_06700_));
 sg13g2_o21ai_1 _25389_ (.B1(_06634_),
    .Y(_06702_),
    .A1(_09597_),
    .A2(_09622_));
 sg13g2_nand3_1 _25390_ (.B(_06701_),
    .C(_06702_),
    .A(_06642_),
    .Y(_06703_));
 sg13g2_o21ai_1 _25391_ (.B1(_06703_),
    .Y(_02545_),
    .A1(_06669_),
    .A2(_06642_));
 sg13g2_inv_1 _25392_ (.Y(_06704_),
    .A(net14));
 sg13g2_mux2_1 _25393_ (.A0(_09554_),
    .A1(_09540_),
    .S(net129),
    .X(_06705_));
 sg13g2_nor2_1 _25394_ (.A(_06595_),
    .B(_06705_),
    .Y(_06706_));
 sg13g2_a21oi_1 _25395_ (.A1(_06662_),
    .A2(_08425_),
    .Y(_06707_),
    .B1(_06706_));
 sg13g2_nand2_1 _25396_ (.Y(_06708_),
    .A(_09335_),
    .B(net93));
 sg13g2_o21ai_1 _25397_ (.B1(_06708_),
    .Y(_06709_),
    .A1(_02861_),
    .A2(net93));
 sg13g2_nand2_1 _25398_ (.Y(_06710_),
    .A(net780),
    .B(_06709_));
 sg13g2_o21ai_1 _25399_ (.B1(_06710_),
    .Y(_06711_),
    .A1(net780),
    .A2(_08327_));
 sg13g2_nor3_1 _25400_ (.A(_09608_),
    .B(_09606_),
    .C(_11547_),
    .Y(_06712_));
 sg13g2_a22oi_1 _25401_ (.Y(_06713_),
    .B1(_06711_),
    .B2(_06712_),
    .A2(_06707_),
    .A1(_11551_));
 sg13g2_nand2_1 _25402_ (.Y(_06714_),
    .A(net703),
    .B(net1015));
 sg13g2_nand2_1 _25403_ (.Y(_06715_),
    .A(_09609_),
    .B(_08947_));
 sg13g2_a21oi_1 _25404_ (.A1(_06714_),
    .A2(_06715_),
    .Y(_06716_),
    .B1(_00185_));
 sg13g2_mux2_1 _25405_ (.A0(_04908_),
    .A1(_04994_),
    .S(net980),
    .X(_06717_));
 sg13g2_nand3_1 _25406_ (.B(_11678_),
    .C(_06717_),
    .A(net979),
    .Y(_06718_));
 sg13g2_mux4_1 _25407_ (.S0(net980),
    .A0(_04899_),
    .A1(_05267_),
    .A2(_04914_),
    .A3(_04986_),
    .S1(net979),
    .X(_06719_));
 sg13g2_nor2_1 _25408_ (.A(_11729_),
    .B(_11652_),
    .Y(_06720_));
 sg13g2_a21oi_1 _25409_ (.A1(_05260_),
    .A2(_06609_),
    .Y(_06721_),
    .B1(_06720_));
 sg13g2_or2_1 _25410_ (.X(_06722_),
    .B(_11677_),
    .A(_11652_));
 sg13g2_o21ai_1 _25411_ (.B1(_06722_),
    .Y(_06723_),
    .A1(_11730_),
    .A2(_06721_));
 sg13g2_a21oi_1 _25412_ (.A1(net976),
    .A2(_06719_),
    .Y(_06724_),
    .B1(_06723_));
 sg13g2_a221oi_1 _25413_ (.B2(_06724_),
    .C1(_11552_),
    .B1(_06718_),
    .A1(_04891_),
    .Y(_06725_),
    .A2(_06603_));
 sg13g2_nor4_1 _25414_ (.A(_09601_),
    .B(_06644_),
    .C(_06716_),
    .D(_06725_),
    .Y(_06726_));
 sg13g2_mux2_1 _25415_ (.A0(_00233_),
    .A1(_09464_),
    .S(_06596_),
    .X(_06727_));
 sg13g2_nand2_1 _25416_ (.Y(_06728_),
    .A(net781),
    .B(_10945_));
 sg13g2_o21ai_1 _25417_ (.B1(_06728_),
    .Y(_06729_),
    .A1(net779),
    .A2(_06727_));
 sg13g2_nand2_1 _25418_ (.Y(_06730_),
    .A(_11571_),
    .B(_06729_));
 sg13g2_mux2_1 _25419_ (.A0(_09306_),
    .A1(_09312_),
    .S(net129),
    .X(_06731_));
 sg13g2_nand2_1 _25420_ (.Y(_06732_),
    .A(net780),
    .B(_06731_));
 sg13g2_o21ai_1 _25421_ (.B1(_06732_),
    .Y(_06733_),
    .A1(net780),
    .A2(_08380_));
 sg13g2_mux2_1 _25422_ (.A0(_00241_),
    .A1(_09474_),
    .S(net93),
    .X(_06734_));
 sg13g2_nand2_1 _25423_ (.Y(_06735_),
    .A(_06595_),
    .B(_03465_));
 sg13g2_o21ai_1 _25424_ (.B1(_06735_),
    .Y(_06736_),
    .A1(net779),
    .A2(_06734_));
 sg13g2_a22oi_1 _25425_ (.Y(_06737_),
    .B1(_06736_),
    .B2(_11569_),
    .A2(_06733_),
    .A1(_11570_));
 sg13g2_nand4_1 _25426_ (.B(_06726_),
    .C(_06730_),
    .A(_06713_),
    .Y(_06738_),
    .D(_06737_));
 sg13g2_nand3_1 _25427_ (.B(_06702_),
    .C(_06738_),
    .A(_06642_),
    .Y(_06739_));
 sg13g2_o21ai_1 _25428_ (.B1(_06739_),
    .Y(_02546_),
    .A1(_06704_),
    .A2(_06642_));
 sg13g2_mux4_1 _25429_ (.S0(_05360_),
    .A0(_08974_),
    .A1(_08981_),
    .A2(_08969_),
    .A3(_08976_),
    .S1(_06111_),
    .X(_06740_));
 sg13g2_mux4_1 _25430_ (.S0(_05360_),
    .A0(_08980_),
    .A1(_08973_),
    .A2(_08984_),
    .A3(_08988_),
    .S1(_06111_),
    .X(_06741_));
 sg13g2_nor2b_1 _25431_ (.A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B_N(_06741_),
    .Y(_06742_));
 sg13g2_a21oi_1 _25432_ (.A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .A2(_06740_),
    .Y(_06743_),
    .B1(_06742_));
 sg13g2_mux4_1 _25433_ (.S0(_05360_),
    .A0(_08978_),
    .A1(_08986_),
    .A2(_08989_),
    .A3(_08971_),
    .S1(_06111_),
    .X(_06744_));
 sg13g2_nand3b_1 _25434_ (.B(\cpu.gpio.r_spi_miso_src[1][3] ),
    .C(_06744_),
    .Y(_06745_),
    .A_N(_00150_));
 sg13g2_o21ai_1 _25435_ (.B1(_06745_),
    .Y(_06746_),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .A2(_06743_));
 sg13g2_mux4_1 _25436_ (.S0(_04722_),
    .A0(_08974_),
    .A1(_08981_),
    .A2(_08969_),
    .A3(_08976_),
    .S1(_06109_),
    .X(_06747_));
 sg13g2_mux4_1 _25437_ (.S0(_04722_),
    .A0(_08980_),
    .A1(_08973_),
    .A2(_08984_),
    .A3(_08988_),
    .S1(_06109_),
    .X(_06748_));
 sg13g2_nor2b_1 _25438_ (.A(\cpu.gpio.r_spi_miso_src[0][2] ),
    .B_N(_06748_),
    .Y(_06749_));
 sg13g2_a21oi_1 _25439_ (.A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .A2(_06747_),
    .Y(_06750_),
    .B1(_06749_));
 sg13g2_mux4_1 _25440_ (.S0(_04722_),
    .A0(_08978_),
    .A1(_08986_),
    .A2(_08989_),
    .A3(_08971_),
    .S1(_06109_),
    .X(_06751_));
 sg13g2_nand3b_1 _25441_ (.B(\cpu.gpio.r_spi_miso_src[0][3] ),
    .C(_06751_),
    .Y(_06752_),
    .A_N(_00110_));
 sg13g2_o21ai_1 _25442_ (.B1(_06752_),
    .Y(_06753_),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .A2(_06750_));
 sg13g2_mux2_1 _25443_ (.A0(_06746_),
    .A1(_06753_),
    .S(_11591_),
    .X(_06754_));
 sg13g2_nor2_1 _25444_ (.A(net1083),
    .B(_11637_),
    .Y(_06755_));
 sg13g2_nor2b_1 _25445_ (.A(net1017),
    .B_N(net1083),
    .Y(_06756_));
 sg13g2_a22oi_1 _25446_ (.Y(_06757_),
    .B1(_06756_),
    .B2(net520),
    .A2(_06755_),
    .A1(net1017));
 sg13g2_nor3_1 _25447_ (.A(net877),
    .B(net406),
    .C(_06757_),
    .Y(_06758_));
 sg13g2_buf_4 _25448_ (.X(_06759_),
    .A(_06758_));
 sg13g2_mux2_1 _25449_ (.A0(_09072_),
    .A1(_06754_),
    .S(_06759_),
    .X(_02586_));
 sg13g2_mux2_1 _25450_ (.A0(_09071_),
    .A1(_09072_),
    .S(_06759_),
    .X(_02587_));
 sg13g2_mux2_1 _25451_ (.A0(_09075_),
    .A1(_09071_),
    .S(_06759_),
    .X(_02588_));
 sg13g2_mux2_1 _25452_ (.A0(_09069_),
    .A1(_09075_),
    .S(_06759_),
    .X(_02589_));
 sg13g2_mux2_1 _25453_ (.A0(_09077_),
    .A1(_09069_),
    .S(_06759_),
    .X(_02590_));
 sg13g2_mux2_1 _25454_ (.A0(_09076_),
    .A1(_09077_),
    .S(_06759_),
    .X(_02591_));
 sg13g2_mux2_1 _25455_ (.A0(_09070_),
    .A1(_09076_),
    .S(_06759_),
    .X(_02592_));
 sg13g2_mux2_1 _25456_ (.A0(\cpu.spi.r_in[7] ),
    .A1(_09070_),
    .S(_06759_),
    .X(_02593_));
 sg13g2_nor2_1 _25457_ (.A(_09019_),
    .B(net850),
    .Y(_06760_));
 sg13g2_buf_2 _25458_ (.A(_06760_),
    .X(_06761_));
 sg13g2_a22oi_1 _25459_ (.Y(_06762_),
    .B1(_06761_),
    .B2(_09032_),
    .A2(_11641_),
    .A1(_09088_));
 sg13g2_nand4_1 _25460_ (.B(_09044_),
    .C(_11645_),
    .A(_09034_),
    .Y(_06763_),
    .D(_06762_));
 sg13g2_buf_1 _25461_ (.A(_06763_),
    .X(_06764_));
 sg13g2_buf_1 _25462_ (.A(_00225_),
    .X(_06765_));
 sg13g2_nor2b_1 _25463_ (.A(net520),
    .B_N(_00223_),
    .Y(_06766_));
 sg13g2_o21ai_1 _25464_ (.B1(_09084_),
    .Y(_06767_),
    .A1(_06765_),
    .A2(_06766_));
 sg13g2_o21ai_1 _25465_ (.B1(_06767_),
    .Y(_06768_),
    .A1(_09084_),
    .A2(net942));
 sg13g2_a21oi_1 _25466_ (.A1(_11578_),
    .A2(_06768_),
    .Y(_06769_),
    .B1(net72));
 sg13g2_a21o_1 _25467_ (.A2(net72),
    .A1(\cpu.spi.r_out[0] ),
    .B1(_06769_),
    .X(_02601_));
 sg13g2_buf_1 _25468_ (.A(_09020_),
    .X(_06770_));
 sg13g2_mux2_1 _25469_ (.A0(_00178_),
    .A1(_00223_),
    .S(net520),
    .X(_06771_));
 sg13g2_a22oi_1 _25470_ (.Y(_06772_),
    .B1(_06761_),
    .B2(_09818_),
    .A2(net850),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _25471_ (.B1(_06772_),
    .Y(_06773_),
    .A1(net778),
    .A2(_06771_));
 sg13g2_mux2_1 _25472_ (.A0(_06773_),
    .A1(\cpu.spi.r_out[1] ),
    .S(net72),
    .X(_02602_));
 sg13g2_mux2_1 _25473_ (.A0(_00179_),
    .A1(_00178_),
    .S(net520),
    .X(_06774_));
 sg13g2_a22oi_1 _25474_ (.Y(_06775_),
    .B1(_06761_),
    .B2(_09826_),
    .A2(net850),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _25475_ (.B1(_06775_),
    .Y(_06776_),
    .A1(net778),
    .A2(_06774_));
 sg13g2_mux2_1 _25476_ (.A0(_06776_),
    .A1(\cpu.spi.r_out[2] ),
    .S(net72),
    .X(_02603_));
 sg13g2_mux2_1 _25477_ (.A0(_00287_),
    .A1(_00179_),
    .S(net520),
    .X(_06777_));
 sg13g2_a22oi_1 _25478_ (.Y(_06778_),
    .B1(_06761_),
    .B2(_09833_),
    .A2(net850),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _25479_ (.B1(_06778_),
    .Y(_06779_),
    .A1(net778),
    .A2(_06777_));
 sg13g2_mux2_1 _25480_ (.A0(_06779_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net72),
    .X(_02604_));
 sg13g2_mux2_1 _25481_ (.A0(_00180_),
    .A1(_00287_),
    .S(net520),
    .X(_06780_));
 sg13g2_a22oi_1 _25482_ (.Y(_06781_),
    .B1(_06761_),
    .B2(_09839_),
    .A2(net850),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _25483_ (.B1(_06781_),
    .Y(_06782_),
    .A1(net778),
    .A2(_06780_));
 sg13g2_mux2_1 _25484_ (.A0(_06782_),
    .A1(\cpu.spi.r_out[4] ),
    .S(net72),
    .X(_02605_));
 sg13g2_mux2_1 _25485_ (.A0(_00181_),
    .A1(_00180_),
    .S(net520),
    .X(_06783_));
 sg13g2_a22oi_1 _25486_ (.Y(_06784_),
    .B1(_06761_),
    .B2(_09845_),
    .A2(net850),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _25487_ (.B1(_06784_),
    .Y(_06785_),
    .A1(net778),
    .A2(_06783_));
 sg13g2_mux2_1 _25488_ (.A0(_06785_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net72),
    .X(_02606_));
 sg13g2_buf_1 _25489_ (.A(_00182_),
    .X(_06786_));
 sg13g2_mux2_1 _25490_ (.A0(_06786_),
    .A1(_00181_),
    .S(_11638_),
    .X(_06787_));
 sg13g2_a22oi_1 _25491_ (.Y(_06788_),
    .B1(_06761_),
    .B2(_09851_),
    .A2(net850),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _25492_ (.B1(_06788_),
    .Y(_06789_),
    .A1(_06770_),
    .A2(_06787_));
 sg13g2_mux2_1 _25493_ (.A0(_06789_),
    .A1(\cpu.spi.r_out[6] ),
    .S(_06764_),
    .X(_02607_));
 sg13g2_buf_1 _25494_ (.A(_00281_),
    .X(_06790_));
 sg13g2_mux2_1 _25495_ (.A0(_06790_),
    .A1(_06786_),
    .S(_11638_),
    .X(_06791_));
 sg13g2_a22oi_1 _25496_ (.Y(_06792_),
    .B1(_06761_),
    .B2(_09856_),
    .A2(_11627_),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _25497_ (.B1(_06792_),
    .Y(_06793_),
    .A1(_06770_),
    .A2(_06791_));
 sg13g2_mux2_1 _25498_ (.A0(_06793_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net72),
    .X(_02608_));
 sg13g2_or2_1 _25499_ (.X(_06794_),
    .B(_09098_),
    .A(net877));
 sg13g2_buf_1 _25500_ (.A(_06794_),
    .X(_06795_));
 sg13g2_nand2_1 _25501_ (.Y(_06796_),
    .A(net853),
    .B(_06795_));
 sg13g2_o21ai_1 _25502_ (.B1(_06796_),
    .Y(_02611_),
    .A1(_03612_),
    .A2(_06795_));
 sg13g2_nand2_1 _25503_ (.Y(_06797_),
    .A(_11580_),
    .B(_06795_));
 sg13g2_o21ai_1 _25504_ (.B1(_06797_),
    .Y(_02612_),
    .A1(net716),
    .A2(_06795_));
 sg13g2_nand2b_1 _25505_ (.Y(_06798_),
    .B(_04873_),
    .A_N(_09024_));
 sg13g2_buf_1 _25506_ (.A(_06798_),
    .X(_06799_));
 sg13g2_buf_1 _25507_ (.A(_06799_),
    .X(_06800_));
 sg13g2_nand2_1 _25508_ (.Y(_06801_),
    .A(\cpu.spi.r_timeout[0] ),
    .B(net92));
 sg13g2_o21ai_1 _25509_ (.B1(_06801_),
    .Y(_02616_),
    .A1(net872),
    .A2(net92));
 sg13g2_mux2_1 _25510_ (.A0(net871),
    .A1(\cpu.spi.r_timeout[1] ),
    .S(net92),
    .X(_02617_));
 sg13g2_mux2_1 _25511_ (.A0(net870),
    .A1(\cpu.spi.r_timeout[2] ),
    .S(net92),
    .X(_02618_));
 sg13g2_nand2_1 _25512_ (.Y(_06802_),
    .A(\cpu.spi.r_timeout[3] ),
    .B(net92));
 sg13g2_o21ai_1 _25513_ (.B1(_06802_),
    .Y(_02619_),
    .A1(net849),
    .A2(net92));
 sg13g2_mux2_1 _25514_ (.A0(_05591_),
    .A1(\cpu.spi.r_timeout[4] ),
    .S(net92),
    .X(_02620_));
 sg13g2_mux2_1 _25515_ (.A0(net818),
    .A1(\cpu.spi.r_timeout[5] ),
    .S(_06800_),
    .X(_02621_));
 sg13g2_nand2_1 _25516_ (.Y(_06803_),
    .A(\cpu.spi.r_timeout[6] ),
    .B(_06799_));
 sg13g2_o21ai_1 _25517_ (.B1(_06803_),
    .Y(_02622_),
    .A1(_11808_),
    .A2(_06800_));
 sg13g2_nand2_1 _25518_ (.Y(_06804_),
    .A(\cpu.spi.r_timeout[7] ),
    .B(_06799_));
 sg13g2_o21ai_1 _25519_ (.B1(_06804_),
    .Y(_02623_),
    .A1(net848),
    .A2(net92));
 sg13g2_nand2_1 _25520_ (.Y(_06805_),
    .A(net1084),
    .B(_09026_));
 sg13g2_nand2_1 _25521_ (.Y(_06806_),
    .A(_09020_),
    .B(_09045_));
 sg13g2_o21ai_1 _25522_ (.B1(_09045_),
    .Y(_06807_),
    .A1(net406),
    .A2(_09081_));
 sg13g2_or4_1 _25523_ (.A(_00226_),
    .B(_08939_),
    .C(_09052_),
    .D(_09081_),
    .X(_06808_));
 sg13g2_nand3_1 _25524_ (.B(_06807_),
    .C(_06808_),
    .A(net1018),
    .Y(_06809_));
 sg13g2_a21o_1 _25525_ (.A2(_06806_),
    .A1(_06805_),
    .B1(_06809_),
    .X(_06810_));
 sg13g2_buf_2 _25526_ (.A(_06810_),
    .X(_06811_));
 sg13g2_buf_1 _25527_ (.A(_06811_),
    .X(_06812_));
 sg13g2_and2_1 _25528_ (.A(net878),
    .B(\cpu.spi.r_timeout[0] ),
    .X(_06813_));
 sg13g2_a21oi_1 _25529_ (.A1(net778),
    .A2(_00284_),
    .Y(_06814_),
    .B1(_06813_));
 sg13g2_nand2_1 _25530_ (.Y(_06815_),
    .A(_09054_),
    .B(net71));
 sg13g2_o21ai_1 _25531_ (.B1(_06815_),
    .Y(_02624_),
    .A1(net71),
    .A2(_06814_));
 sg13g2_nor3_1 _25532_ (.A(_09054_),
    .B(_09055_),
    .C(_06811_),
    .Y(_06816_));
 sg13g2_a21oi_1 _25533_ (.A1(_09054_),
    .A2(_09055_),
    .Y(_06817_),
    .B1(_06816_));
 sg13g2_nor2_1 _25534_ (.A(net778),
    .B(_06811_),
    .Y(_06818_));
 sg13g2_buf_2 _25535_ (.A(_06818_),
    .X(_06819_));
 sg13g2_a22oi_1 _25536_ (.Y(_06820_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[1] ),
    .A2(net71),
    .A1(_09055_));
 sg13g2_o21ai_1 _25537_ (.B1(_06820_),
    .Y(_02625_),
    .A1(net878),
    .A2(_06817_));
 sg13g2_a22oi_1 _25538_ (.Y(_06821_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[2] ),
    .A2(net71),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_o21ai_1 _25539_ (.B1(\cpu.spi.r_timeout_count[2] ),
    .Y(_06822_),
    .A1(_09054_),
    .A2(_09055_));
 sg13g2_o21ai_1 _25540_ (.B1(_06822_),
    .Y(_06823_),
    .A1(_09057_),
    .A2(net71));
 sg13g2_nand2_1 _25541_ (.Y(_06824_),
    .A(net778),
    .B(_06823_));
 sg13g2_nand2_1 _25542_ (.Y(_02626_),
    .A(_06821_),
    .B(_06824_));
 sg13g2_nor2_1 _25543_ (.A(_09059_),
    .B(_06811_),
    .Y(_06825_));
 sg13g2_a21oi_1 _25544_ (.A1(\cpu.spi.r_timeout_count[3] ),
    .A2(_09057_),
    .Y(_06826_),
    .B1(_06825_));
 sg13g2_a22oi_1 _25545_ (.Y(_06827_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[3] ),
    .A2(net71),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_o21ai_1 _25546_ (.B1(_06827_),
    .Y(_02627_),
    .A1(net878),
    .A2(_06826_));
 sg13g2_nor2_1 _25547_ (.A(_09061_),
    .B(_06811_),
    .Y(_06828_));
 sg13g2_a21oi_1 _25548_ (.A1(\cpu.spi.r_timeout_count[4] ),
    .A2(_09059_),
    .Y(_06829_),
    .B1(_06828_));
 sg13g2_a22oi_1 _25549_ (.Y(_06830_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[4] ),
    .A2(net71),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_o21ai_1 _25550_ (.B1(_06830_),
    .Y(_02628_),
    .A1(net878),
    .A2(_06829_));
 sg13g2_nor2_1 _25551_ (.A(_09063_),
    .B(_06811_),
    .Y(_06831_));
 sg13g2_a21oi_1 _25552_ (.A1(\cpu.spi.r_timeout_count[5] ),
    .A2(_09061_),
    .Y(_06832_),
    .B1(_06831_));
 sg13g2_a22oi_1 _25553_ (.Y(_06833_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[5] ),
    .A2(net71),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_o21ai_1 _25554_ (.B1(_06833_),
    .Y(_02629_),
    .A1(net878),
    .A2(_06832_));
 sg13g2_nor2_1 _25555_ (.A(_09065_),
    .B(_06811_),
    .Y(_06834_));
 sg13g2_a21oi_1 _25556_ (.A1(\cpu.spi.r_timeout_count[6] ),
    .A2(_09063_),
    .Y(_06835_),
    .B1(_06834_));
 sg13g2_a22oi_1 _25557_ (.Y(_06836_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[6] ),
    .A2(_06812_),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_o21ai_1 _25558_ (.B1(_06836_),
    .Y(_02630_),
    .A1(net878),
    .A2(_06835_));
 sg13g2_nor3_1 _25559_ (.A(_09053_),
    .B(_09065_),
    .C(_06811_),
    .Y(_06837_));
 sg13g2_a21oi_1 _25560_ (.A1(_09053_),
    .A2(_09065_),
    .Y(_06838_),
    .B1(_06837_));
 sg13g2_a22oi_1 _25561_ (.Y(_06839_),
    .B1(_06819_),
    .B2(\cpu.spi.r_timeout[7] ),
    .A2(_06812_),
    .A1(_09053_));
 sg13g2_o21ai_1 _25562_ (.B1(_06839_),
    .Y(_02631_),
    .A1(net878),
    .A2(_06838_));
 sg13g2_buf_1 _25563_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_06840_));
 sg13g2_nor2_1 _25564_ (.A(_06840_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_06841_));
 sg13g2_nand2_1 _25565_ (.Y(_06842_),
    .A(net337),
    .B(_06841_));
 sg13g2_nor2_1 _25566_ (.A(net1019),
    .B(_06842_),
    .Y(_06843_));
 sg13g2_buf_1 _25567_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_06844_));
 sg13g2_buf_1 _25568_ (.A(net1051),
    .X(_06845_));
 sg13g2_buf_1 _25569_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_06846_));
 sg13g2_buf_1 _25570_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_06847_));
 sg13g2_buf_1 _25571_ (.A(_06847_),
    .X(_06848_));
 sg13g2_nor2_2 _25572_ (.A(net1050),
    .B(_06848_),
    .Y(_06849_));
 sg13g2_buf_2 _25573_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_06850_));
 sg13g2_inv_1 _25574_ (.Y(_06851_),
    .A(_06850_));
 sg13g2_nand3_1 _25575_ (.B(net920),
    .C(_06849_),
    .A(_06851_),
    .Y(_06852_));
 sg13g2_o21ai_1 _25576_ (.B1(_06852_),
    .Y(_06853_),
    .A1(net920),
    .A2(_06849_));
 sg13g2_and2_1 _25577_ (.A(_06843_),
    .B(_06853_),
    .X(_06854_));
 sg13g2_buf_2 _25578_ (.A(_06854_),
    .X(_06855_));
 sg13g2_mux2_1 _25579_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_06855_),
    .X(_02644_));
 sg13g2_mux2_1 _25580_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_06855_),
    .X(_02645_));
 sg13g2_mux2_1 _25581_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_06855_),
    .X(_02646_));
 sg13g2_mux2_1 _25582_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_06855_),
    .X(_02647_));
 sg13g2_mux2_1 _25583_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_06855_),
    .X(_02648_));
 sg13g2_mux2_1 _25584_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_06855_),
    .X(_02649_));
 sg13g2_xor2_1 _25585_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_06856_));
 sg13g2_mux2_1 _25586_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_06856_),
    .S(_06855_),
    .X(_02650_));
 sg13g2_and4_1 _25587_ (.A(_06850_),
    .B(net920),
    .C(_06843_),
    .D(_06849_),
    .X(_06857_));
 sg13g2_buf_1 _25588_ (.A(_06857_),
    .X(_06858_));
 sg13g2_mux2_1 _25589_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net163),
    .X(_02651_));
 sg13g2_mux2_1 _25590_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net163),
    .X(_02652_));
 sg13g2_mux2_1 _25591_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net163),
    .X(_02653_));
 sg13g2_mux2_1 _25592_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net163),
    .X(_02654_));
 sg13g2_mux2_1 _25593_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net163),
    .X(_02655_));
 sg13g2_mux2_1 _25594_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net163),
    .X(_02656_));
 sg13g2_mux2_1 _25595_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net163),
    .X(_02657_));
 sg13g2_mux2_1 _25596_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_06856_),
    .S(_06858_),
    .X(_02658_));
 sg13g2_buf_1 _25597_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_06859_));
 sg13g2_buf_1 _25598_ (.A(_06859_),
    .X(_06860_));
 sg13g2_buf_1 _25599_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_06861_));
 sg13g2_inv_2 _25600_ (.Y(_06862_),
    .A(net1049));
 sg13g2_buf_1 _25601_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_06863_));
 sg13g2_buf_1 _25602_ (.A(_06863_),
    .X(_06864_));
 sg13g2_inv_1 _25603_ (.Y(_06865_),
    .A(_06864_));
 sg13g2_nor2_1 _25604_ (.A(net1085),
    .B(net956),
    .Y(_06866_));
 sg13g2_nand3_1 _25605_ (.B(_06866_),
    .C(_06093_),
    .A(net1010),
    .Y(_06867_));
 sg13g2_buf_1 _25606_ (.A(_06867_),
    .X(_06868_));
 sg13g2_nor3_1 _25607_ (.A(net627),
    .B(net557),
    .C(_06868_),
    .Y(_06869_));
 sg13g2_buf_2 _25608_ (.A(_06869_),
    .X(_06870_));
 sg13g2_buf_2 _25609_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_06871_));
 sg13g2_a21oi_1 _25610_ (.A1(_06865_),
    .A2(_06870_),
    .Y(_06872_),
    .B1(_06871_));
 sg13g2_nand2_1 _25611_ (.Y(_06873_),
    .A(_06871_),
    .B(_06863_));
 sg13g2_nor3_1 _25612_ (.A(_06862_),
    .B(_06870_),
    .C(_06873_),
    .Y(_06874_));
 sg13g2_a21oi_1 _25613_ (.A1(_06862_),
    .A2(_06872_),
    .Y(_06875_),
    .B1(_06874_));
 sg13g2_nor2_1 _25614_ (.A(_06860_),
    .B(_06875_),
    .Y(_06876_));
 sg13g2_buf_1 _25615_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_06877_));
 sg13g2_nor2_1 _25616_ (.A(_06877_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_06878_));
 sg13g2_and2_1 _25617_ (.A(net337),
    .B(_06878_),
    .X(_06879_));
 sg13g2_buf_2 _25618_ (.A(_06879_),
    .X(_06880_));
 sg13g2_inv_2 _25619_ (.Y(_06881_),
    .A(_06871_));
 sg13g2_nor2_1 _25620_ (.A(_06862_),
    .B(_06880_),
    .Y(_06882_));
 sg13g2_a21oi_1 _25621_ (.A1(_06863_),
    .A2(\cpu.uart.r_xstate[3] ),
    .Y(_06883_),
    .B1(_06881_));
 sg13g2_a21oi_1 _25622_ (.A1(_06881_),
    .A2(_06882_),
    .Y(_06884_),
    .B1(_06883_));
 sg13g2_inv_2 _25623_ (.Y(_06885_),
    .A(_06859_));
 sg13g2_a22oi_1 _25624_ (.Y(_06886_),
    .B1(_06884_),
    .B2(_06885_),
    .A2(_06880_),
    .A1(_06862_));
 sg13g2_nor3_1 _25625_ (.A(net1019),
    .B(_06876_),
    .C(_06886_),
    .Y(_06887_));
 sg13g2_buf_2 _25626_ (.A(_06887_),
    .X(_06888_));
 sg13g2_buf_1 _25627_ (.A(_06888_),
    .X(_06889_));
 sg13g2_nor2_1 _25628_ (.A(_06871_),
    .B(_06859_),
    .Y(_06890_));
 sg13g2_xnor2_1 _25629_ (.Y(_06891_),
    .A(net1049),
    .B(_06890_));
 sg13g2_buf_1 _25630_ (.A(_06891_),
    .X(_06892_));
 sg13g2_buf_1 _25631_ (.A(_06892_),
    .X(_06893_));
 sg13g2_nor2_1 _25632_ (.A(_09809_),
    .B(net614),
    .Y(_06894_));
 sg13g2_a21oi_1 _25633_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net614),
    .Y(_06895_),
    .B1(_06894_));
 sg13g2_nor2_1 _25634_ (.A(\cpu.uart.r_out[0] ),
    .B(net29),
    .Y(_06896_));
 sg13g2_a21oi_1 _25635_ (.A1(net29),
    .A2(_06895_),
    .Y(_02659_),
    .B1(_06896_));
 sg13g2_nor2b_1 _25636_ (.A(_06892_),
    .B_N(_09818_),
    .Y(_06897_));
 sg13g2_a21oi_1 _25637_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net614),
    .Y(_06898_),
    .B1(_06897_));
 sg13g2_nor2_1 _25638_ (.A(\cpu.uart.r_out[1] ),
    .B(_06889_),
    .Y(_06899_));
 sg13g2_a21oi_1 _25639_ (.A1(net29),
    .A2(_06898_),
    .Y(_02660_),
    .B1(_06899_));
 sg13g2_nor2b_1 _25640_ (.A(_06892_),
    .B_N(_09825_),
    .Y(_06900_));
 sg13g2_a21oi_1 _25641_ (.A1(\cpu.uart.r_out[3] ),
    .A2(_06893_),
    .Y(_06901_),
    .B1(_06900_));
 sg13g2_nor2_1 _25642_ (.A(\cpu.uart.r_out[2] ),
    .B(_06888_),
    .Y(_06902_));
 sg13g2_a21oi_1 _25643_ (.A1(net29),
    .A2(_06901_),
    .Y(_02661_),
    .B1(_06902_));
 sg13g2_nor2_1 _25644_ (.A(net849),
    .B(net614),
    .Y(_06903_));
 sg13g2_a21oi_1 _25645_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net614),
    .Y(_06904_),
    .B1(_06903_));
 sg13g2_nor2_1 _25646_ (.A(\cpu.uart.r_out[3] ),
    .B(_06888_),
    .Y(_06905_));
 sg13g2_a21oi_1 _25647_ (.A1(net29),
    .A2(_06904_),
    .Y(_02662_),
    .B1(_06905_));
 sg13g2_nor2b_1 _25648_ (.A(_06892_),
    .B_N(_09839_),
    .Y(_06906_));
 sg13g2_a21oi_1 _25649_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net614),
    .Y(_06907_),
    .B1(_06906_));
 sg13g2_nor2_1 _25650_ (.A(\cpu.uart.r_out[4] ),
    .B(_06888_),
    .Y(_06908_));
 sg13g2_a21oi_1 _25651_ (.A1(net29),
    .A2(_06907_),
    .Y(_02663_),
    .B1(_06908_));
 sg13g2_nor2b_1 _25652_ (.A(_06892_),
    .B_N(_09845_),
    .Y(_06909_));
 sg13g2_a21oi_1 _25653_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net614),
    .Y(_06910_),
    .B1(_06909_));
 sg13g2_nor2_1 _25654_ (.A(\cpu.uart.r_out[5] ),
    .B(_06888_),
    .Y(_06911_));
 sg13g2_a21oi_1 _25655_ (.A1(net29),
    .A2(_06910_),
    .Y(_02664_),
    .B1(_06911_));
 sg13g2_nor2_1 _25656_ (.A(_11746_),
    .B(_06892_),
    .Y(_06912_));
 sg13g2_a21oi_1 _25657_ (.A1(\cpu.uart.r_out[7] ),
    .A2(_06893_),
    .Y(_06913_),
    .B1(_06912_));
 sg13g2_nor2_1 _25658_ (.A(\cpu.uart.r_out[6] ),
    .B(_06888_),
    .Y(_06914_));
 sg13g2_a21oi_1 _25659_ (.A1(net29),
    .A2(_06913_),
    .Y(_02665_),
    .B1(_06914_));
 sg13g2_nor2_1 _25660_ (.A(_06790_),
    .B(net614),
    .Y(_06915_));
 sg13g2_mux2_1 _25661_ (.A0(\cpu.uart.r_out[7] ),
    .A1(_06915_),
    .S(_06889_),
    .X(_02666_));
 sg13g2_nand2b_1 _25662_ (.Y(_06916_),
    .B(_09723_),
    .A_N(_09684_));
 sg13g2_nor3_1 _25663_ (.A(net1050),
    .B(_06847_),
    .C(net1051),
    .Y(_06917_));
 sg13g2_a22oi_1 _25664_ (.Y(_06918_),
    .B1(_06916_),
    .B2(_06917_),
    .A2(net1051),
    .A1(net1050));
 sg13g2_nor4_1 _25665_ (.A(_06850_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_06847_),
    .D(_06844_),
    .Y(_06919_));
 sg13g2_a21o_1 _25666_ (.A2(_06916_),
    .A1(net1050),
    .B1(_06847_),
    .X(_06920_));
 sg13g2_a22oi_1 _25667_ (.Y(_06921_),
    .B1(_06920_),
    .B2(net1051),
    .A2(_06919_),
    .A1(_06856_));
 sg13g2_o21ai_1 _25668_ (.B1(_06921_),
    .Y(_06922_),
    .A1(_06851_),
    .A2(_06918_));
 sg13g2_nor2_1 _25669_ (.A(_06851_),
    .B(net1050),
    .Y(_06923_));
 sg13g2_nor2b_1 _25670_ (.A(net1051),
    .B_N(_06856_),
    .Y(_06924_));
 sg13g2_nand2_1 _25671_ (.Y(_06925_),
    .A(_06846_),
    .B(net1051));
 sg13g2_nor2_1 _25672_ (.A(_06850_),
    .B(_06925_),
    .Y(_06926_));
 sg13g2_a21oi_1 _25673_ (.A1(_06923_),
    .A2(_06924_),
    .Y(_06927_),
    .B1(_06926_));
 sg13g2_nor3_1 _25674_ (.A(net919),
    .B(_06842_),
    .C(_06927_),
    .Y(_06928_));
 sg13g2_xor2_1 _25675_ (.B(_06849_),
    .A(net920),
    .X(_06929_));
 sg13g2_o21ai_1 _25676_ (.B1(net1018),
    .Y(_06930_),
    .A1(_09695_),
    .A2(_06929_));
 sg13g2_nor3_1 _25677_ (.A(_06922_),
    .B(_06928_),
    .C(_06930_),
    .Y(_06931_));
 sg13g2_and2_1 _25678_ (.A(_06850_),
    .B(net1050),
    .X(_06932_));
 sg13g2_buf_1 _25679_ (.A(_06932_),
    .X(_06933_));
 sg13g2_o21ai_1 _25680_ (.B1(net920),
    .Y(_06934_),
    .A1(net919),
    .A2(_06933_));
 sg13g2_nor2b_1 _25681_ (.A(_06919_),
    .B_N(_06934_),
    .Y(_06935_));
 sg13g2_and2_1 _25682_ (.A(_06931_),
    .B(_06935_),
    .X(_06936_));
 sg13g2_nor2_1 _25683_ (.A(_06840_),
    .B(_06931_),
    .Y(_06937_));
 sg13g2_a21oi_1 _25684_ (.A1(_06840_),
    .A2(_06936_),
    .Y(_02669_),
    .B1(_06937_));
 sg13g2_nand2_1 _25685_ (.Y(_06938_),
    .A(_06840_),
    .B(_06935_));
 sg13g2_inv_1 _25686_ (.Y(_06939_),
    .A(\cpu.uart.r_rcnt[1] ));
 sg13g2_a21oi_1 _25687_ (.A1(_06931_),
    .A2(_06938_),
    .Y(_06940_),
    .B1(_06939_));
 sg13g2_a21o_1 _25688_ (.A2(_06936_),
    .A1(_06841_),
    .B1(_06940_),
    .X(_02670_));
 sg13g2_nor3_2 _25689_ (.A(_06881_),
    .B(_06862_),
    .C(_06860_),
    .Y(_06941_));
 sg13g2_nor2_1 _25690_ (.A(_06862_),
    .B(net918),
    .Y(_06942_));
 sg13g2_nor2_1 _25691_ (.A(_06861_),
    .B(_06885_),
    .Y(_06943_));
 sg13g2_or2_1 _25692_ (.X(_06944_),
    .B(_06863_),
    .A(_06871_));
 sg13g2_buf_1 _25693_ (.A(_06944_),
    .X(_06945_));
 sg13g2_nor3_1 _25694_ (.A(_06942_),
    .B(_06943_),
    .C(_06945_),
    .Y(_06946_));
 sg13g2_nor3_1 _25695_ (.A(net877),
    .B(_06941_),
    .C(_06946_),
    .Y(_06947_));
 sg13g2_nand2_1 _25696_ (.Y(_06948_),
    .A(\cpu.uart.r_out[0] ),
    .B(_06892_));
 sg13g2_xor2_1 _25697_ (.B(_06948_),
    .A(\cpu.uart.r_x_invert ),
    .X(_06949_));
 sg13g2_nor2_1 _25698_ (.A(_00280_),
    .B(_06947_),
    .Y(_06950_));
 sg13g2_a21oi_1 _25699_ (.A1(_06947_),
    .A2(_06949_),
    .Y(_06951_),
    .B1(_06950_));
 sg13g2_buf_1 _25700_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_06952_));
 sg13g2_nand3_1 _25701_ (.B(_06870_),
    .C(_06941_),
    .A(net917),
    .Y(_06953_));
 sg13g2_buf_1 _25702_ (.A(_06953_),
    .X(_06954_));
 sg13g2_nand2_1 _25703_ (.Y(_06955_),
    .A(net1049),
    .B(net918));
 sg13g2_o21ai_1 _25704_ (.B1(_06955_),
    .Y(_06956_),
    .A1(net1049),
    .A2(net337));
 sg13g2_nand2b_1 _25705_ (.Y(_06957_),
    .B(_06890_),
    .A_N(_06880_));
 sg13g2_o21ai_1 _25706_ (.B1(_06957_),
    .Y(_06958_),
    .A1(_06881_),
    .A2(_06885_));
 sg13g2_nor2_1 _25707_ (.A(_06883_),
    .B(_06943_),
    .Y(_06959_));
 sg13g2_nor2_1 _25708_ (.A(_06880_),
    .B(_06959_),
    .Y(_06960_));
 sg13g2_a221oi_1 _25709_ (.B2(net1049),
    .C1(_06960_),
    .B1(_06958_),
    .A1(_06863_),
    .Y(_06961_),
    .A2(_06956_));
 sg13g2_a21oi_1 _25710_ (.A1(_06954_),
    .A2(_06961_),
    .Y(_06962_),
    .B1(net877));
 sg13g2_mux2_1 _25711_ (.A0(_06951_),
    .A1(_06952_),
    .S(_06962_),
    .X(_02675_));
 sg13g2_a21oi_1 _25712_ (.A1(net917),
    .A2(_06878_),
    .Y(_06963_),
    .B1(net918));
 sg13g2_o21ai_1 _25713_ (.B1(net918),
    .Y(_06964_),
    .A1(net917),
    .A2(_06878_));
 sg13g2_o21ai_1 _25714_ (.B1(_06964_),
    .Y(_06965_),
    .A1(_06881_),
    .A2(_06963_));
 sg13g2_nand2_1 _25715_ (.Y(_06966_),
    .A(_06861_),
    .B(_06965_));
 sg13g2_nor3_1 _25716_ (.A(_06871_),
    .B(net1049),
    .C(net918),
    .Y(_06967_));
 sg13g2_nand2b_1 _25717_ (.Y(_06968_),
    .B(_06967_),
    .A_N(_06863_));
 sg13g2_nand4_1 _25718_ (.B(net337),
    .C(_06966_),
    .A(net879),
    .Y(_06969_),
    .D(_06968_));
 sg13g2_nor2b_1 _25719_ (.A(_06969_),
    .B_N(_06954_),
    .Y(_06970_));
 sg13g2_nor2_1 _25720_ (.A(_06862_),
    .B(_06885_),
    .Y(_06971_));
 sg13g2_a21oi_1 _25721_ (.A1(_06971_),
    .A2(_06945_),
    .Y(_06972_),
    .B1(_06967_));
 sg13g2_nand2_1 _25722_ (.Y(_06973_),
    .A(_06970_),
    .B(_06972_));
 sg13g2_nor2b_1 _25723_ (.A(_06877_),
    .B_N(_06970_),
    .Y(_06974_));
 sg13g2_a21oi_1 _25724_ (.A1(_06877_),
    .A2(_06973_),
    .Y(_06975_),
    .B1(_06974_));
 sg13g2_inv_1 _25725_ (.Y(_02678_),
    .A(_06975_));
 sg13g2_nand2_1 _25726_ (.Y(_06976_),
    .A(_06877_),
    .B(_06972_));
 sg13g2_nand2_1 _25727_ (.Y(_06977_),
    .A(_06970_),
    .B(_06976_));
 sg13g2_o21ai_1 _25728_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_06978_),
    .A1(_06877_),
    .A2(_06973_));
 sg13g2_o21ai_1 _25729_ (.B1(_06978_),
    .Y(_02679_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_06977_));
 sg13g2_nor2_1 _25730_ (.A(net529),
    .B(net125),
    .Y(_06979_));
 sg13g2_buf_1 _25731_ (.A(_06979_),
    .X(_06980_));
 sg13g2_nand4_1 _25732_ (.B(_09950_),
    .C(_09955_),
    .A(_09944_),
    .Y(_06981_),
    .D(_04741_));
 sg13g2_nor3_2 _25733_ (.A(_09917_),
    .B(_09946_),
    .C(_06981_),
    .Y(_06982_));
 sg13g2_nand4_1 _25734_ (.B(_09950_),
    .C(_09955_),
    .A(_09944_),
    .Y(_06983_),
    .D(_09951_));
 sg13g2_nand2_1 _25735_ (.Y(_06984_),
    .A(net530),
    .B(_09873_));
 sg13g2_buf_2 _25736_ (.A(_06984_),
    .X(_06985_));
 sg13g2_o21ai_1 _25737_ (.B1(_06985_),
    .Y(_06986_),
    .A1(_09873_),
    .A2(_06983_));
 sg13g2_nor2_1 _25738_ (.A(_04741_),
    .B(_06986_),
    .Y(_06987_));
 sg13g2_a221oi_1 _25739_ (.B2(net107),
    .C1(_06987_),
    .B1(_06982_),
    .A1(net872),
    .Y(_02465_),
    .A2(net83));
 sg13g2_inv_1 _25740_ (.Y(_06988_),
    .A(_05169_));
 sg13g2_nand2_1 _25741_ (.Y(_06989_),
    .A(net529),
    .B(_09873_));
 sg13g2_buf_1 _25742_ (.A(_06989_),
    .X(_06990_));
 sg13g2_o21ai_1 _25743_ (.B1(net116),
    .Y(_06991_),
    .A1(net152),
    .A2(_06982_));
 sg13g2_nand3_1 _25744_ (.B(net107),
    .C(_06982_),
    .A(_05169_),
    .Y(_06992_));
 sg13g2_o21ai_1 _25745_ (.B1(_06992_),
    .Y(_06993_),
    .A1(net1009),
    .A2(_06985_));
 sg13g2_a21oi_1 _25746_ (.A1(_06988_),
    .A2(_06991_),
    .Y(_02466_),
    .B1(_06993_));
 sg13g2_a21o_1 _25747_ (.A2(_06982_),
    .A1(_05169_),
    .B1(_09873_),
    .X(_06994_));
 sg13g2_a21oi_1 _25748_ (.A1(net116),
    .A2(_06994_),
    .Y(_06995_),
    .B1(_05233_));
 sg13g2_nor2_1 _25749_ (.A(net1008),
    .B(_06985_),
    .Y(_06996_));
 sg13g2_nand3_1 _25750_ (.B(_05233_),
    .C(_06982_),
    .A(_05169_),
    .Y(_06997_));
 sg13g2_buf_1 _25751_ (.A(_06997_),
    .X(_06998_));
 sg13g2_nor2_1 _25752_ (.A(_09873_),
    .B(_06998_),
    .Y(_06999_));
 sg13g2_nor3_1 _25753_ (.A(_06995_),
    .B(_06996_),
    .C(_06999_),
    .Y(_02467_));
 sg13g2_inv_1 _25754_ (.Y(_07000_),
    .A(_05295_));
 sg13g2_inv_1 _25755_ (.Y(_07001_),
    .A(_06981_));
 sg13g2_nand4_1 _25756_ (.B(_05233_),
    .C(_09947_),
    .A(_05169_),
    .Y(_07002_),
    .D(_07001_));
 sg13g2_buf_1 _25757_ (.A(_07002_),
    .X(_07003_));
 sg13g2_nor2_1 _25758_ (.A(net530),
    .B(net125),
    .Y(_07004_));
 sg13g2_a21oi_1 _25759_ (.A1(net107),
    .A2(_07003_),
    .Y(_07005_),
    .B1(_07004_));
 sg13g2_nor2_1 _25760_ (.A(_09873_),
    .B(_07003_),
    .Y(_07006_));
 sg13g2_a22oi_1 _25761_ (.Y(_07007_),
    .B1(_07006_),
    .B2(_07000_),
    .A2(net83),
    .A1(net1078));
 sg13g2_o21ai_1 _25762_ (.B1(_07007_),
    .Y(_02468_),
    .A1(_07000_),
    .A2(_07005_));
 sg13g2_o21ai_1 _25763_ (.B1(_09865_),
    .Y(_07008_),
    .A1(_07000_),
    .A2(_06998_));
 sg13g2_a21oi_1 _25764_ (.A1(net116),
    .A2(_07008_),
    .Y(_07009_),
    .B1(_05343_));
 sg13g2_nand3_1 _25765_ (.B(_05343_),
    .C(_06999_),
    .A(_05295_),
    .Y(_07010_));
 sg13g2_o21ai_1 _25766_ (.B1(_07010_),
    .Y(_07011_),
    .A1(net1007),
    .A2(_06985_));
 sg13g2_nor2_1 _25767_ (.A(_07009_),
    .B(_07011_),
    .Y(_02469_));
 sg13g2_nand2_1 _25768_ (.Y(_07012_),
    .A(_05295_),
    .B(_05343_));
 sg13g2_o21ai_1 _25769_ (.B1(_09865_),
    .Y(_07013_),
    .A1(_07003_),
    .A2(_07012_));
 sg13g2_a21oi_1 _25770_ (.A1(net116),
    .A2(_07013_),
    .Y(_07014_),
    .B1(_05442_));
 sg13g2_nand4_1 _25771_ (.B(_05343_),
    .C(_05442_),
    .A(_05295_),
    .Y(_07015_),
    .D(_07006_));
 sg13g2_o21ai_1 _25772_ (.B1(_07015_),
    .Y(_07016_),
    .A1(net1006),
    .A2(_06985_));
 sg13g2_nor2_1 _25773_ (.A(_07014_),
    .B(_07016_),
    .Y(_02470_));
 sg13g2_inv_1 _25774_ (.Y(_07017_),
    .A(_05470_));
 sg13g2_nand3_1 _25775_ (.B(_05343_),
    .C(_05442_),
    .A(_05295_),
    .Y(_07018_));
 sg13g2_nor2_1 _25776_ (.A(_07017_),
    .B(_07018_),
    .Y(_07019_));
 sg13g2_o21ai_1 _25777_ (.B1(net125),
    .Y(_07020_),
    .A1(_06998_),
    .A2(_07018_));
 sg13g2_a21oi_1 _25778_ (.A1(_06990_),
    .A2(_07020_),
    .Y(_07021_),
    .B1(_05470_));
 sg13g2_a221oi_1 _25779_ (.B2(_07019_),
    .C1(_07021_),
    .B1(_06999_),
    .A1(net845),
    .Y(_02471_),
    .A2(_06980_));
 sg13g2_nand2_2 _25780_ (.Y(_07022_),
    .A(_04859_),
    .B(_07019_));
 sg13g2_inv_1 _25781_ (.Y(_07023_),
    .A(_07022_));
 sg13g2_inv_1 _25782_ (.Y(_07024_),
    .A(_07019_));
 sg13g2_o21ai_1 _25783_ (.B1(_09864_),
    .Y(_07025_),
    .A1(_07003_),
    .A2(_07024_));
 sg13g2_a21oi_1 _25784_ (.A1(_06990_),
    .A2(_07025_),
    .Y(_07026_),
    .B1(_04859_));
 sg13g2_a221oi_1 _25785_ (.B2(_07023_),
    .C1(_07026_),
    .B1(_07006_),
    .A1(net848),
    .Y(_02472_),
    .A2(_06980_));
 sg13g2_inv_1 _25786_ (.Y(_07027_),
    .A(_05531_));
 sg13g2_nor3_1 _25787_ (.A(_07027_),
    .B(_06998_),
    .C(_07022_),
    .Y(_07028_));
 sg13g2_o21ai_1 _25788_ (.B1(net125),
    .Y(_07029_),
    .A1(_06998_),
    .A2(_07022_));
 sg13g2_a21oi_1 _25789_ (.A1(net116),
    .A2(_07029_),
    .Y(_07030_),
    .B1(_05531_));
 sg13g2_a221oi_1 _25790_ (.B2(net107),
    .C1(_07030_),
    .B1(_07028_),
    .A1(_06474_),
    .Y(_02473_),
    .A2(net83));
 sg13g2_and2_1 _25791_ (.A(_05546_),
    .B(_07028_),
    .X(_07031_));
 sg13g2_buf_1 _25792_ (.A(_07031_),
    .X(_07032_));
 sg13g2_o21ai_1 _25793_ (.B1(net116),
    .Y(_07033_),
    .A1(net152),
    .A2(_07028_));
 sg13g2_inv_1 _25794_ (.Y(_07034_),
    .A(_05546_));
 sg13g2_nor2_1 _25795_ (.A(_09926_),
    .B(_06985_),
    .Y(_07035_));
 sg13g2_a221oi_1 _25796_ (.B2(_07034_),
    .C1(_07035_),
    .B1(_07033_),
    .A1(net107),
    .Y(_02474_),
    .A2(_07032_));
 sg13g2_o21ai_1 _25797_ (.B1(_06989_),
    .Y(_07036_),
    .A1(net152),
    .A2(_07032_));
 sg13g2_inv_1 _25798_ (.Y(_07037_),
    .A(_04930_));
 sg13g2_nand2_1 _25799_ (.Y(_07038_),
    .A(_04930_),
    .B(_07032_));
 sg13g2_nor2_1 _25800_ (.A(_09873_),
    .B(_07038_),
    .Y(_07039_));
 sg13g2_a221oi_1 _25801_ (.B2(_07037_),
    .C1(_07039_),
    .B1(_07036_),
    .A1(_11702_),
    .Y(_02475_),
    .A2(net83));
 sg13g2_nand3_1 _25802_ (.B(_05546_),
    .C(_04930_),
    .A(_05531_),
    .Y(_07040_));
 sg13g2_nor3_2 _25803_ (.A(_07003_),
    .B(_07022_),
    .C(_07040_),
    .Y(_07041_));
 sg13g2_o21ai_1 _25804_ (.B1(_06989_),
    .Y(_07042_),
    .A1(_09874_),
    .A2(_07041_));
 sg13g2_nand2_1 _25805_ (.Y(_07043_),
    .A(_04978_),
    .B(_07042_));
 sg13g2_nor2b_1 _25806_ (.A(_09874_),
    .B_N(_07041_),
    .Y(_07044_));
 sg13g2_inv_1 _25807_ (.Y(_07045_),
    .A(_04978_));
 sg13g2_a22oi_1 _25808_ (.Y(_07046_),
    .B1(_07044_),
    .B2(_07045_),
    .A2(net83),
    .A1(_09937_));
 sg13g2_nand2_1 _25809_ (.Y(_02476_),
    .A(_07043_),
    .B(_07046_));
 sg13g2_o21ai_1 _25810_ (.B1(net125),
    .Y(_07047_),
    .A1(_07045_),
    .A2(_07038_));
 sg13g2_a21oi_1 _25811_ (.A1(net116),
    .A2(_07047_),
    .Y(_07048_),
    .B1(_05005_));
 sg13g2_nand3_1 _25812_ (.B(_05005_),
    .C(_07039_),
    .A(_04978_),
    .Y(_07049_));
 sg13g2_o21ai_1 _25813_ (.B1(_07049_),
    .Y(_07050_),
    .A1(_09942_),
    .A2(_06985_));
 sg13g2_nor2_1 _25814_ (.A(_07048_),
    .B(_07050_),
    .Y(_02477_));
 sg13g2_and3_1 _25815_ (.X(_07051_),
    .A(_04978_),
    .B(_05005_),
    .C(_05030_));
 sg13g2_buf_1 _25816_ (.A(_07051_),
    .X(_07052_));
 sg13g2_nand3_1 _25817_ (.B(_05005_),
    .C(_07041_),
    .A(_04978_),
    .Y(_07053_));
 sg13g2_nand2_1 _25818_ (.Y(_07054_),
    .A(net125),
    .B(_07053_));
 sg13g2_a21oi_1 _25819_ (.A1(net116),
    .A2(_07054_),
    .Y(_07055_),
    .B1(_05030_));
 sg13g2_a221oi_1 _25820_ (.B2(_07052_),
    .C1(_07055_),
    .B1(_07044_),
    .A1(_11737_),
    .Y(_02478_),
    .A2(net83));
 sg13g2_nand3_1 _25821_ (.B(_07032_),
    .C(_07052_),
    .A(_04930_),
    .Y(_07056_));
 sg13g2_a21oi_1 _25822_ (.A1(net107),
    .A2(_07056_),
    .Y(_07057_),
    .B1(_07004_));
 sg13g2_nand2b_1 _25823_ (.Y(_07058_),
    .B(_07057_),
    .A_N(_05051_));
 sg13g2_o21ai_1 _25824_ (.B1(_05051_),
    .Y(_07059_),
    .A1(net152),
    .A2(_07056_));
 sg13g2_a22oi_1 _25825_ (.Y(_02479_),
    .B1(_07058_),
    .B2(_07059_),
    .A2(net83),
    .A1(_11747_));
 sg13g2_nand3_1 _25826_ (.B(_07041_),
    .C(_07052_),
    .A(_05051_),
    .Y(_07060_));
 sg13g2_a21o_1 _25827_ (.A2(_07060_),
    .A1(net125),
    .B1(_07004_),
    .X(_07061_));
 sg13g2_nor3_1 _25828_ (.A(_05085_),
    .B(net152),
    .C(_07060_),
    .Y(_07062_));
 sg13g2_a221oi_1 _25829_ (.B2(_05085_),
    .C1(_07062_),
    .B1(_07061_),
    .A1(_09958_),
    .Y(_07063_),
    .A2(net83));
 sg13g2_inv_1 _25830_ (.Y(_02480_),
    .A(_07063_));
 sg13g2_nor2_1 _25831_ (.A(\cpu.r_clk_invert ),
    .B(net747),
    .Y(_07064_));
 sg13g2_a21oi_1 _25832_ (.A1(_08976_),
    .A2(net690),
    .Y(_02547_),
    .B1(_07064_));
 sg13g2_nand2b_1 _25833_ (.Y(_07065_),
    .B(net879),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _25834_ (.A(_07065_),
    .X(_07066_));
 sg13g2_nor2b_1 _25835_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net459),
    .Y(_07067_));
 sg13g2_nand4_1 _25836_ (.B(_02838_),
    .C(net976),
    .A(_09131_),
    .Y(_07068_),
    .D(_11657_));
 sg13g2_buf_2 _25837_ (.A(_07068_),
    .X(_07069_));
 sg13g2_nor2_1 _25838_ (.A(net570),
    .B(_07069_),
    .Y(_07070_));
 sg13g2_nor3_1 _25839_ (.A(_07066_),
    .B(_07067_),
    .C(_07070_),
    .Y(_00741_));
 sg13g2_nor2_1 _25840_ (.A(\cpu.dcache.r_valid[1] ),
    .B(_02883_),
    .Y(_07071_));
 sg13g2_nor2_1 _25841_ (.A(net568),
    .B(_07069_),
    .Y(_07072_));
 sg13g2_nor3_1 _25842_ (.A(_07066_),
    .B(_07071_),
    .C(_07072_),
    .Y(_00742_));
 sg13g2_nor2_1 _25843_ (.A(\cpu.dcache.r_valid[2] ),
    .B(_12065_),
    .Y(_07073_));
 sg13g2_nor2_1 _25844_ (.A(net641),
    .B(_07069_),
    .Y(_07074_));
 sg13g2_nor3_1 _25845_ (.A(_07066_),
    .B(_07073_),
    .C(_07074_),
    .Y(_00743_));
 sg13g2_nor2_1 _25846_ (.A(\cpu.dcache.r_valid[3] ),
    .B(_02893_),
    .Y(_07075_));
 sg13g2_nor2_1 _25847_ (.A(net640),
    .B(_07069_),
    .Y(_07076_));
 sg13g2_nor3_1 _25848_ (.A(_07066_),
    .B(_07075_),
    .C(_07076_),
    .Y(_00744_));
 sg13g2_inv_1 _25849_ (.Y(_07077_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _25850_ (.Y(_07078_),
    .A(_07069_));
 sg13g2_a221oi_1 _25851_ (.B2(_09860_),
    .C1(_07066_),
    .B1(_07078_),
    .A1(_07077_),
    .Y(_00745_),
    .A2(_02894_));
 sg13g2_nor2_1 _25852_ (.A(\cpu.dcache.r_valid[5] ),
    .B(_12386_),
    .Y(_07079_));
 sg13g2_nor2_1 _25853_ (.A(net638),
    .B(_07069_),
    .Y(_07080_));
 sg13g2_nor3_1 _25854_ (.A(_07066_),
    .B(_07079_),
    .C(_07080_),
    .Y(_00746_));
 sg13g2_nor2_1 _25855_ (.A(\cpu.dcache.r_valid[6] ),
    .B(net453),
    .Y(_07081_));
 sg13g2_nor2_1 _25856_ (.A(_12431_),
    .B(_07069_),
    .Y(_07082_));
 sg13g2_nor3_1 _25857_ (.A(_07066_),
    .B(_07081_),
    .C(_07082_),
    .Y(_00747_));
 sg13g2_nor2_1 _25858_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net385),
    .Y(_07083_));
 sg13g2_nor2_1 _25859_ (.A(net567),
    .B(_07069_),
    .Y(_07084_));
 sg13g2_nor3_1 _25860_ (.A(_07066_),
    .B(_07083_),
    .C(_07084_),
    .Y(_00748_));
 sg13g2_nand3_1 _25861_ (.B(_09986_),
    .C(_04584_),
    .A(_09969_),
    .Y(_07085_));
 sg13g2_buf_2 _25862_ (.A(_07085_),
    .X(_07086_));
 sg13g2_nand2_1 _25863_ (.Y(_07087_),
    .A(_08516_),
    .B(_07086_));
 sg13g2_o21ai_1 _25864_ (.B1(_07087_),
    .Y(_07088_),
    .A1(net708),
    .A2(_07086_));
 sg13g2_and3_1 _25865_ (.X(_00797_),
    .A(net186),
    .B(_09093_),
    .C(_07088_));
 sg13g2_and4_1 _25866_ (.A(net710),
    .B(_11021_),
    .C(\cpu.dec.do_flush_all ),
    .D(net646),
    .X(_00930_));
 sg13g2_and4_1 _25867_ (.A(net710),
    .B(_11048_),
    .C(\cpu.dec.do_flush_all ),
    .D(_11385_),
    .X(_00948_));
 sg13g2_nand4_1 _25868_ (.B(_03907_),
    .C(_11385_),
    .A(net710),
    .Y(_07089_),
    .D(_10888_));
 sg13g2_mux2_1 _25869_ (.A0(_10796_),
    .A1(_09007_),
    .S(_07089_),
    .X(_07090_));
 sg13g2_mux2_1 _25870_ (.A0(net831),
    .A1(_07090_),
    .S(_07086_),
    .X(_07091_));
 sg13g2_nand3_1 _25871_ (.B(_11207_),
    .C(_07091_),
    .A(net759),
    .Y(_07092_));
 sg13g2_a21oi_1 _25872_ (.A1(_04013_),
    .A2(_05098_),
    .Y(_00949_),
    .B1(_07092_));
 sg13g2_nand2b_1 _25873_ (.Y(_07093_),
    .B(_04832_),
    .A_N(_04809_));
 sg13g2_nor4_2 _25874_ (.A(_00310_),
    .B(_08561_),
    .C(_09095_),
    .Y(_07094_),
    .D(_09108_));
 sg13g2_o21ai_1 _25875_ (.B1(_07094_),
    .Y(_07095_),
    .A1(_00298_),
    .A2(_07093_));
 sg13g2_a22oi_1 _25876_ (.Y(_07096_),
    .B1(_11659_),
    .B2(_09036_),
    .A2(_09564_),
    .A1(_09131_));
 sg13g2_nand3_1 _25877_ (.B(_11228_),
    .C(_07096_),
    .A(_11227_),
    .Y(_07097_));
 sg13g2_nand2_1 _25878_ (.Y(_07098_),
    .A(_08561_),
    .B(_07097_));
 sg13g2_nand2_1 _25879_ (.Y(_07099_),
    .A(net761),
    .B(_07098_));
 sg13g2_a21oi_1 _25880_ (.A1(_08560_),
    .A2(_07095_),
    .Y(_01068_),
    .B1(_07099_));
 sg13g2_o21ai_1 _25881_ (.B1(_07094_),
    .Y(_07100_),
    .A1(_11553_),
    .A2(_04833_));
 sg13g2_a21oi_1 _25882_ (.A1(_08559_),
    .A2(_07100_),
    .Y(_01069_),
    .B1(_07099_));
 sg13g2_inv_1 _25883_ (.Y(_07101_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _25884_ (.Y(_07102_),
    .B(net879),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _25885_ (.A(_07102_),
    .X(_07103_));
 sg13g2_a21oi_1 _25886_ (.A1(_07101_),
    .A2(_06294_),
    .Y(_02424_),
    .B1(_07103_));
 sg13g2_nor2_1 _25887_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06213_),
    .Y(_07104_));
 sg13g2_nor2_1 _25888_ (.A(_07103_),
    .B(_07104_),
    .Y(_02425_));
 sg13g2_nor2_1 _25889_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06230_),
    .Y(_07105_));
 sg13g2_nor2_1 _25890_ (.A(_07103_),
    .B(_07105_),
    .Y(_02426_));
 sg13g2_inv_1 _25891_ (.Y(_07106_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _25892_ (.A1(_07106_),
    .A2(_06356_),
    .Y(_02427_),
    .B1(_07103_));
 sg13g2_nor2_1 _25893_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06256_),
    .Y(_07107_));
 sg13g2_nor2_1 _25894_ (.A(_07103_),
    .B(_07107_),
    .Y(_02428_));
 sg13g2_inv_1 _25895_ (.Y(_07108_),
    .A(\cpu.icache.r_valid[5] ));
 sg13g2_a21oi_1 _25896_ (.A1(_07108_),
    .A2(_06265_),
    .Y(_02429_),
    .B1(_07103_));
 sg13g2_nor2_1 _25897_ (.A(\cpu.icache.r_valid[6] ),
    .B(_06280_),
    .Y(_07109_));
 sg13g2_nor2_1 _25898_ (.A(_07103_),
    .B(_07109_),
    .Y(_02430_));
 sg13g2_nor2_1 _25899_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06291_),
    .Y(_07110_));
 sg13g2_nor2_1 _25900_ (.A(_07103_),
    .B(_07110_),
    .Y(_02431_));
 sg13g2_nand3_1 _25901_ (.B(net183),
    .C(_04766_),
    .A(net1078),
    .Y(_07111_));
 sg13g2_nor3_2 _25902_ (.A(_09022_),
    .B(net583),
    .C(_04697_),
    .Y(_07112_));
 sg13g2_a22oi_1 _25903_ (.Y(_07113_),
    .B1(_07112_),
    .B2(net928),
    .A2(_07111_),
    .A1(_08995_));
 sg13g2_nor2_1 _25904_ (.A(net667),
    .B(_07113_),
    .Y(_00317_));
 sg13g2_nor2_1 _25905_ (.A(_02838_),
    .B(net985),
    .Y(_07114_));
 sg13g2_nor2b_1 _25906_ (.A(_07114_),
    .B_N(_00315_),
    .Y(_00586_));
 sg13g2_nor2_1 _25907_ (.A(_11680_),
    .B(_11731_),
    .Y(_07115_));
 sg13g2_nor2_1 _25908_ (.A(_07114_),
    .B(_07115_),
    .Y(_00587_));
 sg13g2_xnor2_1 _25909_ (.Y(_07116_),
    .A(net984),
    .B(_11657_));
 sg13g2_nor2b_1 _25910_ (.A(_07114_),
    .B_N(_07116_),
    .Y(_00588_));
 sg13g2_nor2_1 _25911_ (.A(_09041_),
    .B(_07086_),
    .Y(_07117_));
 sg13g2_a21oi_1 _25912_ (.A1(net1042),
    .A2(_07086_),
    .Y(_07118_),
    .B1(_07117_));
 sg13g2_nor2_1 _25913_ (.A(net667),
    .B(_07118_),
    .Y(_00798_));
 sg13g2_nand2_1 _25914_ (.Y(_07119_),
    .A(_08589_),
    .B(net646));
 sg13g2_o21ai_1 _25915_ (.B1(_11207_),
    .Y(_07120_),
    .A1(_03911_),
    .A2(_07119_));
 sg13g2_buf_1 _25916_ (.A(_07120_),
    .X(_07121_));
 sg13g2_nand2_1 _25917_ (.Y(_07122_),
    .A(net710),
    .B(_07121_));
 sg13g2_nor2_1 _25918_ (.A(_10659_),
    .B(_09108_),
    .Y(_07123_));
 sg13g2_nand3_1 _25919_ (.B(_10888_),
    .C(_07123_),
    .A(_03907_),
    .Y(_07124_));
 sg13g2_a21oi_1 _25920_ (.A1(net710),
    .A2(_07124_),
    .Y(_07125_),
    .B1(_09030_));
 sg13g2_nor2_1 _25921_ (.A(_03594_),
    .B(_07125_),
    .Y(_07126_));
 sg13g2_mux2_1 _25922_ (.A0(_10659_),
    .A1(_03339_),
    .S(_07126_),
    .X(_07127_));
 sg13g2_nand2b_1 _25923_ (.Y(_07128_),
    .B(_07127_),
    .A_N(_07121_));
 sg13g2_nand3_1 _25924_ (.B(_07122_),
    .C(_07128_),
    .A(_05644_),
    .Y(_00799_));
 sg13g2_mux2_1 _25925_ (.A0(net956),
    .A1(_10388_),
    .S(_07086_),
    .X(_07129_));
 sg13g2_and2_1 _25926_ (.A(_09039_),
    .B(_07129_),
    .X(_00800_));
 sg13g2_nor3_1 _25927_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11205_),
    .C(_03294_),
    .Y(_07130_));
 sg13g2_nand3_1 _25928_ (.B(net646),
    .C(_07130_),
    .A(_08536_),
    .Y(_07131_));
 sg13g2_nand3_1 _25929_ (.B(_07098_),
    .C(_07131_),
    .A(_11199_),
    .Y(_07132_));
 sg13g2_and3_1 _25930_ (.X(_07133_),
    .A(_08589_),
    .B(_11210_),
    .C(_07132_));
 sg13g2_nor3_1 _25931_ (.A(_06662_),
    .B(_04626_),
    .C(_07133_),
    .Y(_07134_));
 sg13g2_nor2_1 _25932_ (.A(_06623_),
    .B(net104),
    .Y(_07135_));
 sg13g2_o21ai_1 _25933_ (.B1(_05631_),
    .Y(_00946_),
    .A1(_07134_),
    .A2(_07135_));
 sg13g2_nand2_1 _25934_ (.Y(_07136_),
    .A(_09131_),
    .B(_09108_));
 sg13g2_nand3_1 _25935_ (.B(\cpu.dec.do_flush_write ),
    .C(_04013_),
    .A(net710),
    .Y(_07137_));
 sg13g2_a21oi_1 _25936_ (.A1(_07136_),
    .A2(_07137_),
    .Y(_00947_),
    .B1(net615));
 sg13g2_nand2_1 _25937_ (.Y(_07138_),
    .A(\cpu.dec.io ),
    .B(_04013_));
 sg13g2_nand2_1 _25938_ (.Y(_07139_),
    .A(_04627_),
    .B(_09108_));
 sg13g2_a21oi_1 _25939_ (.A1(_07138_),
    .A2(_07139_),
    .Y(_00950_),
    .B1(net615));
 sg13g2_and2_1 _25940_ (.A(_09008_),
    .B(_07121_),
    .X(_07140_));
 sg13g2_nand2_1 _25941_ (.Y(_07141_),
    .A(_10796_),
    .B(_07086_));
 sg13g2_o21ai_1 _25942_ (.B1(_07141_),
    .Y(_07142_),
    .A1(_09881_),
    .A2(_07086_));
 sg13g2_nor2_1 _25943_ (.A(_07121_),
    .B(_07142_),
    .Y(_07143_));
 sg13g2_nor3_1 _25944_ (.A(_09591_),
    .B(_07140_),
    .C(_07143_),
    .Y(_00997_));
 sg13g2_a22oi_1 _25945_ (.Y(_07144_),
    .B1(_03392_),
    .B2(net1091),
    .A2(_04013_),
    .A1(_11205_));
 sg13g2_nor2_1 _25946_ (.A(net667),
    .B(_07144_),
    .Y(_00998_));
 sg13g2_nor2b_1 _25947_ (.A(net951),
    .B_N(_05611_),
    .Y(_07145_));
 sg13g2_buf_2 _25948_ (.A(_07145_),
    .X(_07146_));
 sg13g2_nand2_1 _25949_ (.Y(_07147_),
    .A(net538),
    .B(_07146_));
 sg13g2_o21ai_1 _25950_ (.B1(_07147_),
    .Y(_07148_),
    .A1(_11095_),
    .A2(_07146_));
 sg13g2_nand2_1 _25951_ (.Y(_07149_),
    .A(net186),
    .B(_07148_));
 sg13g2_a21oi_1 _25952_ (.A1(_11207_),
    .A2(_07149_),
    .Y(_01074_),
    .B1(_06570_));
 sg13g2_nand2_1 _25953_ (.Y(_07150_),
    .A(net565),
    .B(_07146_));
 sg13g2_o21ai_1 _25954_ (.B1(_07150_),
    .Y(_07151_),
    .A1(_05670_),
    .A2(_07146_));
 sg13g2_nor2_1 _25955_ (.A(_09181_),
    .B(_05602_),
    .Y(_07152_));
 sg13g2_a21oi_1 _25956_ (.A1(_05602_),
    .A2(_07151_),
    .Y(_07153_),
    .B1(_07152_));
 sg13g2_nor2_1 _25957_ (.A(net667),
    .B(_07153_),
    .Y(_01075_));
 sg13g2_mux2_1 _25958_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_09869_),
    .S(_07146_),
    .X(_07154_));
 sg13g2_a21oi_1 _25959_ (.A1(_10653_),
    .A2(_07154_),
    .Y(_07155_),
    .B1(_08617_));
 sg13g2_nor2_1 _25960_ (.A(net667),
    .B(_07155_),
    .Y(_01076_));
 sg13g2_nor2_2 _25961_ (.A(net1072),
    .B(net1073),
    .Y(_07156_));
 sg13g2_nand2_1 _25962_ (.Y(_07157_),
    .A(_00288_),
    .B(_07156_));
 sg13g2_nor4_2 _25963_ (.A(_10576_),
    .B(_10317_),
    .C(_10220_),
    .Y(_07158_),
    .D(_07157_));
 sg13g2_inv_1 _25964_ (.Y(_07159_),
    .A(_00255_));
 sg13g2_nor2b_1 _25965_ (.A(_00257_),
    .B_N(_05609_),
    .Y(_07160_));
 sg13g2_nand2_1 _25966_ (.Y(_07161_),
    .A(_05608_),
    .B(_07160_));
 sg13g2_a21oi_1 _25967_ (.A1(net951),
    .A2(_07159_),
    .Y(_07162_),
    .B1(_07161_));
 sg13g2_nand2_1 _25968_ (.Y(_07163_),
    .A(_08619_),
    .B(_07162_));
 sg13g2_buf_1 _25969_ (.A(_07163_),
    .X(_07164_));
 sg13g2_a21oi_1 _25970_ (.A1(_03171_),
    .A2(_11021_),
    .Y(_07165_),
    .B1(_07162_));
 sg13g2_nor2b_1 _25971_ (.A(_07165_),
    .B_N(net253),
    .Y(_07166_));
 sg13g2_buf_2 _25972_ (.A(_07166_),
    .X(_07167_));
 sg13g2_o21ai_1 _25973_ (.B1(_07167_),
    .Y(_07168_),
    .A1(_07158_),
    .A2(net185));
 sg13g2_nor2_1 _25974_ (.A(_09880_),
    .B(_07163_),
    .Y(_07169_));
 sg13g2_buf_2 _25975_ (.A(_07169_),
    .X(_07170_));
 sg13g2_buf_1 _25976_ (.A(_07170_),
    .X(_07171_));
 sg13g2_a22oi_1 _25977_ (.Y(_07172_),
    .B1(net136),
    .B2(_07158_),
    .A2(_07168_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _25978_ (.A(_09592_),
    .B(_07172_),
    .Y(_01077_));
 sg13g2_nor3_1 _25979_ (.A(net940),
    .B(_04628_),
    .C(net706),
    .Y(_07173_));
 sg13g2_buf_2 _25980_ (.A(_07173_),
    .X(_07174_));
 sg13g2_nor2_1 _25981_ (.A(_10220_),
    .B(_07157_),
    .Y(_07175_));
 sg13g2_a21oi_1 _25982_ (.A1(net1052),
    .A2(_07156_),
    .Y(_07176_),
    .B1(_10892_));
 sg13g2_a21oi_1 _25983_ (.A1(net941),
    .A2(_07175_),
    .Y(_07177_),
    .B1(_07176_));
 sg13g2_nand2_1 _25984_ (.Y(_07178_),
    .A(_05717_),
    .B(_07175_));
 sg13g2_o21ai_1 _25985_ (.B1(_07178_),
    .Y(_07179_),
    .A1(net938),
    .A2(_07177_));
 sg13g2_buf_2 _25986_ (.A(_07179_),
    .X(_07180_));
 sg13g2_nor2b_2 _25987_ (.A(net185),
    .B_N(_07180_),
    .Y(_07181_));
 sg13g2_buf_1 _25988_ (.A(net185),
    .X(_07182_));
 sg13g2_buf_1 _25989_ (.A(_07167_),
    .X(_07183_));
 sg13g2_o21ai_1 _25990_ (.B1(_07183_),
    .Y(_07184_),
    .A1(_05673_),
    .A2(net162));
 sg13g2_a22oi_1 _25991_ (.Y(_07185_),
    .B1(_07184_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07181_),
    .A1(_07174_));
 sg13g2_nor2_1 _25992_ (.A(_09592_),
    .B(_07185_),
    .Y(_01078_));
 sg13g2_buf_1 _25993_ (.A(net747),
    .X(_07186_));
 sg13g2_o21ai_1 _25994_ (.B1(_07183_),
    .Y(_07187_),
    .A1(_05678_),
    .A2(net162));
 sg13g2_a22oi_1 _25995_ (.Y(_07188_),
    .B1(_07187_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07170_),
    .A1(_05678_));
 sg13g2_nor2_1 _25996_ (.A(net613),
    .B(_07188_),
    .Y(_01079_));
 sg13g2_nand2_1 _25997_ (.Y(_07189_),
    .A(net940),
    .B(_11688_));
 sg13g2_nor3_1 _25998_ (.A(net941),
    .B(net1072),
    .C(_07189_),
    .Y(_07190_));
 sg13g2_buf_2 _25999_ (.A(_07190_),
    .X(_07191_));
 sg13g2_buf_1 _26000_ (.A(net185),
    .X(_07192_));
 sg13g2_nor2_1 _26001_ (.A(net1073),
    .B(net816),
    .Y(_07193_));
 sg13g2_nor3_1 _26002_ (.A(net941),
    .B(net1072),
    .C(_05632_),
    .Y(_07194_));
 sg13g2_o21ai_1 _26003_ (.B1(_05612_),
    .Y(_07195_),
    .A1(_07193_),
    .A2(_07194_));
 sg13g2_buf_1 _26004_ (.A(_07195_),
    .X(_07196_));
 sg13g2_nor2b_1 _26005_ (.A(_07196_),
    .B_N(_07180_),
    .Y(_07197_));
 sg13g2_o21ai_1 _26006_ (.B1(net135),
    .Y(_07198_),
    .A1(net161),
    .A2(_07197_));
 sg13g2_a22oi_1 _26007_ (.Y(_07199_),
    .B1(_07198_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07191_),
    .A1(_07181_));
 sg13g2_nor2_1 _26008_ (.A(net613),
    .B(_07199_),
    .Y(_01080_));
 sg13g2_nor2_1 _26009_ (.A(net817),
    .B(_05689_),
    .Y(_07200_));
 sg13g2_and2_1 _26010_ (.A(_07180_),
    .B(_07200_),
    .X(_07201_));
 sg13g2_buf_1 _26011_ (.A(_07201_),
    .X(_07202_));
 sg13g2_o21ai_1 _26012_ (.B1(net135),
    .Y(_07203_),
    .A1(net161),
    .A2(_07202_));
 sg13g2_a22oi_1 _26013_ (.Y(_07204_),
    .B1(_07203_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07202_),
    .A1(net136));
 sg13g2_nor2_1 _26014_ (.A(net613),
    .B(_07204_),
    .Y(_01081_));
 sg13g2_nor2_1 _26015_ (.A(net706),
    .B(_07189_),
    .Y(_07205_));
 sg13g2_buf_2 _26016_ (.A(_07205_),
    .X(_07206_));
 sg13g2_and2_1 _26017_ (.A(_05809_),
    .B(_07180_),
    .X(_07207_));
 sg13g2_o21ai_1 _26018_ (.B1(net135),
    .Y(_07208_),
    .A1(net161),
    .A2(_07207_));
 sg13g2_a22oi_1 _26019_ (.Y(_07209_),
    .B1(_07208_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07206_),
    .A1(_07181_));
 sg13g2_nor2_1 _26020_ (.A(net613),
    .B(_07209_),
    .Y(_01082_));
 sg13g2_and2_1 _26021_ (.A(_05637_),
    .B(_07180_),
    .X(_07210_));
 sg13g2_buf_1 _26022_ (.A(_07210_),
    .X(_07211_));
 sg13g2_o21ai_1 _26023_ (.B1(net135),
    .Y(_07212_),
    .A1(net161),
    .A2(_07211_));
 sg13g2_a22oi_1 _26024_ (.Y(_07213_),
    .B1(_07212_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07211_),
    .A1(net136));
 sg13g2_nor2_1 _26025_ (.A(net613),
    .B(_07213_),
    .Y(_01083_));
 sg13g2_a21oi_1 _26026_ (.A1(net1052),
    .A2(_05656_),
    .Y(_07214_),
    .B1(_04628_));
 sg13g2_and2_1 _26027_ (.A(_05888_),
    .B(_07214_),
    .X(_07215_));
 sg13g2_buf_2 _26028_ (.A(_07215_),
    .X(_07216_));
 sg13g2_nand2_1 _26029_ (.Y(_07217_),
    .A(net1073),
    .B(_05624_));
 sg13g2_o21ai_1 _26030_ (.B1(_07217_),
    .Y(_07218_),
    .A1(_05656_),
    .A2(_05707_));
 sg13g2_nand2_1 _26031_ (.Y(_07219_),
    .A(_05612_),
    .B(_07218_));
 sg13g2_nor2b_1 _26032_ (.A(_07219_),
    .B_N(_07180_),
    .Y(_07220_));
 sg13g2_a21oi_1 _26033_ (.A1(_03171_),
    .A2(_11078_),
    .Y(_07221_),
    .B1(_07162_));
 sg13g2_nor2b_1 _26034_ (.A(_07221_),
    .B_N(net253),
    .Y(_07222_));
 sg13g2_buf_2 _26035_ (.A(_07222_),
    .X(_07223_));
 sg13g2_buf_1 _26036_ (.A(_07223_),
    .X(_07224_));
 sg13g2_o21ai_1 _26037_ (.B1(net134),
    .Y(_07225_),
    .A1(_07192_),
    .A2(_07220_));
 sg13g2_a22oi_1 _26038_ (.Y(_07226_),
    .B1(_07225_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07216_),
    .A1(_07181_));
 sg13g2_nor2_1 _26039_ (.A(net613),
    .B(_07226_),
    .Y(_01084_));
 sg13g2_nor4_1 _26040_ (.A(net938),
    .B(net941),
    .C(net939),
    .D(net1052),
    .Y(_07227_));
 sg13g2_nand3_1 _26041_ (.B(net939),
    .C(net1052),
    .A(net938),
    .Y(_07228_));
 sg13g2_nand2b_1 _26042_ (.Y(_07229_),
    .B(_07228_),
    .A_N(_07227_));
 sg13g2_nand2b_1 _26043_ (.Y(_07230_),
    .B(net941),
    .A_N(net1052));
 sg13g2_a21oi_1 _26044_ (.A1(_07156_),
    .A2(_07230_),
    .Y(_07231_),
    .B1(net939));
 sg13g2_a22oi_1 _26045_ (.Y(_07232_),
    .B1(_07231_),
    .B2(_05704_),
    .A2(_07229_),
    .A1(_07156_));
 sg13g2_buf_2 _26046_ (.A(_07232_),
    .X(_07233_));
 sg13g2_nor2_1 _26047_ (.A(net940),
    .B(_05689_),
    .Y(_07234_));
 sg13g2_nor2b_2 _26048_ (.A(_07233_),
    .B_N(_07234_),
    .Y(_07235_));
 sg13g2_o21ai_1 _26049_ (.B1(_07224_),
    .Y(_07236_),
    .A1(net161),
    .A2(_07235_));
 sg13g2_a22oi_1 _26050_ (.Y(_07237_),
    .B1(_07236_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07235_),
    .A1(net136));
 sg13g2_nor2_1 _26051_ (.A(net613),
    .B(_07237_),
    .Y(_01085_));
 sg13g2_nor2_1 _26052_ (.A(_07164_),
    .B(_07233_),
    .Y(_07238_));
 sg13g2_o21ai_1 _26053_ (.B1(net134),
    .Y(_07239_),
    .A1(_05719_),
    .A2(net162));
 sg13g2_a22oi_1 _26054_ (.Y(_07240_),
    .B1(_07239_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07238_),
    .A1(_07174_));
 sg13g2_nor2_1 _26055_ (.A(_07186_),
    .B(_07240_),
    .Y(_01086_));
 sg13g2_o21ai_1 _26056_ (.B1(_07224_),
    .Y(_07241_),
    .A1(_05728_),
    .A2(net162));
 sg13g2_a22oi_1 _26057_ (.Y(_07242_),
    .B1(_07241_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07170_),
    .A1(_05728_));
 sg13g2_nor2_1 _26058_ (.A(_07186_),
    .B(_07242_),
    .Y(_01087_));
 sg13g2_nor2_1 _26059_ (.A(_05647_),
    .B(net1052),
    .Y(_07243_));
 sg13g2_a22oi_1 _26060_ (.Y(_07244_),
    .B1(_05717_),
    .B2(_07243_),
    .A2(_05683_),
    .A1(net1052));
 sg13g2_nor2b_1 _26061_ (.A(_07244_),
    .B_N(_07156_),
    .Y(_07245_));
 sg13g2_a21oi_1 _26062_ (.A1(_05670_),
    .A2(_07231_),
    .Y(_07246_),
    .B1(_07245_));
 sg13g2_buf_2 _26063_ (.A(_07246_),
    .X(_07247_));
 sg13g2_nor2b_2 _26064_ (.A(_07247_),
    .B_N(_07234_),
    .Y(_07248_));
 sg13g2_o21ai_1 _26065_ (.B1(net135),
    .Y(_07249_),
    .A1(net161),
    .A2(_07248_));
 sg13g2_a22oi_1 _26066_ (.Y(_07250_),
    .B1(_07249_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07248_),
    .A1(net136));
 sg13g2_nor2_1 _26067_ (.A(net613),
    .B(_07250_),
    .Y(_01088_));
 sg13g2_buf_1 _26068_ (.A(net747),
    .X(_07251_));
 sg13g2_nor2_1 _26069_ (.A(_07196_),
    .B(_07233_),
    .Y(_07252_));
 sg13g2_o21ai_1 _26070_ (.B1(net134),
    .Y(_07253_),
    .A1(net161),
    .A2(_07252_));
 sg13g2_a22oi_1 _26071_ (.Y(_07254_),
    .B1(_07253_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07238_),
    .A1(_07191_));
 sg13g2_nor2_1 _26072_ (.A(net612),
    .B(_07254_),
    .Y(_01089_));
 sg13g2_nor2b_2 _26073_ (.A(_07233_),
    .B_N(_07200_),
    .Y(_07255_));
 sg13g2_o21ai_1 _26074_ (.B1(net134),
    .Y(_07256_),
    .A1(_07192_),
    .A2(_07255_));
 sg13g2_a22oi_1 _26075_ (.Y(_07257_),
    .B1(_07256_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07255_),
    .A1(net136));
 sg13g2_nor2_1 _26076_ (.A(net612),
    .B(_07257_),
    .Y(_01090_));
 sg13g2_nor2b_1 _26077_ (.A(_07233_),
    .B_N(_05809_),
    .Y(_07258_));
 sg13g2_o21ai_1 _26078_ (.B1(net134),
    .Y(_07259_),
    .A1(net161),
    .A2(_07258_));
 sg13g2_a22oi_1 _26079_ (.Y(_07260_),
    .B1(_07259_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07238_),
    .A1(_07206_));
 sg13g2_nor2_1 _26080_ (.A(_07251_),
    .B(_07260_),
    .Y(_01091_));
 sg13g2_nor2_2 _26081_ (.A(_07217_),
    .B(_05706_),
    .Y(_07261_));
 sg13g2_buf_1 _26082_ (.A(net185),
    .X(_07262_));
 sg13g2_o21ai_1 _26083_ (.B1(net134),
    .Y(_07263_),
    .A1(_07262_),
    .A2(_07261_));
 sg13g2_a22oi_1 _26084_ (.Y(_07264_),
    .B1(_07263_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07261_),
    .A1(net136));
 sg13g2_nor2_1 _26085_ (.A(_07251_),
    .B(_07264_),
    .Y(_01092_));
 sg13g2_nor2_1 _26086_ (.A(_07219_),
    .B(_07233_),
    .Y(_07265_));
 sg13g2_o21ai_1 _26087_ (.B1(net134),
    .Y(_07266_),
    .A1(_07262_),
    .A2(_07265_));
 sg13g2_a22oi_1 _26088_ (.Y(_07267_),
    .B1(_07266_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07238_),
    .A1(_07216_));
 sg13g2_nor2_1 _26089_ (.A(net612),
    .B(_07267_),
    .Y(_01093_));
 sg13g2_nor2_1 _26090_ (.A(_05670_),
    .B(_07177_),
    .Y(_07268_));
 sg13g2_or2_1 _26091_ (.X(_07269_),
    .B(_07268_),
    .A(_07158_));
 sg13g2_buf_1 _26092_ (.A(_07269_),
    .X(_07270_));
 sg13g2_and2_1 _26093_ (.A(_07234_),
    .B(_07270_),
    .X(_07271_));
 sg13g2_buf_1 _26094_ (.A(_07271_),
    .X(_07272_));
 sg13g2_o21ai_1 _26095_ (.B1(net134),
    .Y(_07273_),
    .A1(net160),
    .A2(_07272_));
 sg13g2_a22oi_1 _26096_ (.Y(_07274_),
    .B1(_07273_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07272_),
    .A1(_07171_));
 sg13g2_nor2_1 _26097_ (.A(net612),
    .B(_07274_),
    .Y(_01094_));
 sg13g2_nor2b_1 _26098_ (.A(_07164_),
    .B_N(_07270_),
    .Y(_07275_));
 sg13g2_o21ai_1 _26099_ (.B1(_07223_),
    .Y(_07276_),
    .A1(_05763_),
    .A2(_07182_));
 sg13g2_a22oi_1 _26100_ (.Y(_07277_),
    .B1(_07276_),
    .B2(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A2(_07275_),
    .A1(_07174_));
 sg13g2_nor2_1 _26101_ (.A(net612),
    .B(_07277_),
    .Y(_01095_));
 sg13g2_o21ai_1 _26102_ (.B1(_07223_),
    .Y(_07278_),
    .A1(_05769_),
    .A2(_07182_));
 sg13g2_a22oi_1 _26103_ (.Y(_07279_),
    .B1(_07278_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07170_),
    .A1(_05769_));
 sg13g2_nor2_1 _26104_ (.A(net612),
    .B(_07279_),
    .Y(_01096_));
 sg13g2_nor2b_1 _26105_ (.A(_07196_),
    .B_N(_07270_),
    .Y(_07280_));
 sg13g2_o21ai_1 _26106_ (.B1(_07223_),
    .Y(_07281_),
    .A1(net160),
    .A2(_07280_));
 sg13g2_a22oi_1 _26107_ (.Y(_07282_),
    .B1(_07281_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07275_),
    .A1(_07191_));
 sg13g2_nor2_1 _26108_ (.A(net612),
    .B(_07282_),
    .Y(_01097_));
 sg13g2_and2_1 _26109_ (.A(_07200_),
    .B(_07270_),
    .X(_07283_));
 sg13g2_buf_1 _26110_ (.A(_07283_),
    .X(_07284_));
 sg13g2_o21ai_1 _26111_ (.B1(_07223_),
    .Y(_07285_),
    .A1(net160),
    .A2(_07284_));
 sg13g2_a22oi_1 _26112_ (.Y(_07286_),
    .B1(_07285_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07284_),
    .A1(_07171_));
 sg13g2_nor2_1 _26113_ (.A(net612),
    .B(_07286_),
    .Y(_01098_));
 sg13g2_buf_1 _26114_ (.A(net747),
    .X(_07287_));
 sg13g2_nor3_1 _26115_ (.A(net940),
    .B(net706),
    .C(_07247_),
    .Y(_07288_));
 sg13g2_o21ai_1 _26116_ (.B1(_07167_),
    .Y(_07289_),
    .A1(net185),
    .A2(_07288_));
 sg13g2_and2_1 _26117_ (.A(_11688_),
    .B(_07288_),
    .X(_07290_));
 sg13g2_inv_1 _26118_ (.Y(_07291_),
    .A(net162));
 sg13g2_a22oi_1 _26119_ (.Y(_07292_),
    .B1(_07290_),
    .B2(_07291_),
    .A2(_07289_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26120_ (.A(net611),
    .B(_07292_),
    .Y(_01099_));
 sg13g2_and2_1 _26121_ (.A(_05809_),
    .B(_07270_),
    .X(_07293_));
 sg13g2_o21ai_1 _26122_ (.B1(_07223_),
    .Y(_07294_),
    .A1(net160),
    .A2(_07293_));
 sg13g2_a22oi_1 _26123_ (.Y(_07295_),
    .B1(_07294_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07275_),
    .A1(_07206_));
 sg13g2_nor2_1 _26124_ (.A(_07287_),
    .B(_07295_),
    .Y(_01100_));
 sg13g2_and2_1 _26125_ (.A(_05637_),
    .B(_07270_),
    .X(_07296_));
 sg13g2_buf_1 _26126_ (.A(_07296_),
    .X(_07297_));
 sg13g2_o21ai_1 _26127_ (.B1(_07223_),
    .Y(_07298_),
    .A1(net160),
    .A2(_07297_));
 sg13g2_a22oi_1 _26128_ (.Y(_07299_),
    .B1(_07298_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07297_),
    .A1(net136));
 sg13g2_nor2_1 _26129_ (.A(_07287_),
    .B(_07299_),
    .Y(_01101_));
 sg13g2_nor2b_2 _26130_ (.A(_07247_),
    .B_N(_07193_),
    .Y(_07300_));
 sg13g2_o21ai_1 _26131_ (.B1(net135),
    .Y(_07301_),
    .A1(net160),
    .A2(_07300_));
 sg13g2_a22oi_1 _26132_ (.Y(_07302_),
    .B1(_07301_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07300_),
    .A1(_07170_));
 sg13g2_nor2_1 _26133_ (.A(net611),
    .B(_07302_),
    .Y(_01102_));
 sg13g2_nor2_1 _26134_ (.A(net185),
    .B(_07247_),
    .Y(_07303_));
 sg13g2_nor2_1 _26135_ (.A(_07196_),
    .B(_07247_),
    .Y(_07304_));
 sg13g2_o21ai_1 _26136_ (.B1(net135),
    .Y(_07305_),
    .A1(net160),
    .A2(_07304_));
 sg13g2_a22oi_1 _26137_ (.Y(_07306_),
    .B1(_07305_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07303_),
    .A1(_07191_));
 sg13g2_nor2_1 _26138_ (.A(net611),
    .B(_07306_),
    .Y(_01103_));
 sg13g2_o21ai_1 _26139_ (.B1(net135),
    .Y(_07307_),
    .A1(_05805_),
    .A2(net162));
 sg13g2_a22oi_1 _26140_ (.Y(_07308_),
    .B1(_07307_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07170_),
    .A1(_05805_));
 sg13g2_nor2_1 _26141_ (.A(net611),
    .B(_07308_),
    .Y(_01104_));
 sg13g2_o21ai_1 _26142_ (.B1(_07167_),
    .Y(_07309_),
    .A1(_05811_),
    .A2(net162));
 sg13g2_a22oi_1 _26143_ (.Y(_07310_),
    .B1(_07309_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07303_),
    .A1(_07206_));
 sg13g2_nor2_1 _26144_ (.A(net611),
    .B(_07310_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26145_ (.B1(_07167_),
    .Y(_07311_),
    .A1(_05816_),
    .A2(net162));
 sg13g2_a22oi_1 _26146_ (.Y(_07312_),
    .B1(_07311_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07170_),
    .A1(_05816_));
 sg13g2_nor2_1 _26147_ (.A(net611),
    .B(_07312_),
    .Y(_01106_));
 sg13g2_nor2_1 _26148_ (.A(_07219_),
    .B(_07247_),
    .Y(_07313_));
 sg13g2_o21ai_1 _26149_ (.B1(_07167_),
    .Y(_07314_),
    .A1(net160),
    .A2(_07313_));
 sg13g2_a22oi_1 _26150_ (.Y(_07315_),
    .B1(_07314_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07303_),
    .A1(_07216_));
 sg13g2_nor2_1 _26151_ (.A(net611),
    .B(_07315_),
    .Y(_01107_));
 sg13g2_and2_1 _26152_ (.A(_07180_),
    .B(_07234_),
    .X(_07316_));
 sg13g2_buf_1 _26153_ (.A(_07316_),
    .X(_07317_));
 sg13g2_o21ai_1 _26154_ (.B1(_07167_),
    .Y(_07318_),
    .A1(net185),
    .A2(_07317_));
 sg13g2_a22oi_1 _26155_ (.Y(_07319_),
    .B1(_07318_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07317_),
    .A1(_07170_));
 sg13g2_nor2_1 _26156_ (.A(net611),
    .B(_07319_),
    .Y(_01108_));
 sg13g2_buf_1 _26157_ (.A(net747),
    .X(_07320_));
 sg13g2_a21oi_1 _26158_ (.A1(net951),
    .A2(_00255_),
    .Y(_07321_),
    .B1(_07161_));
 sg13g2_nand2_1 _26159_ (.Y(_07322_),
    .A(_08619_),
    .B(_07321_));
 sg13g2_buf_1 _26160_ (.A(_07322_),
    .X(_07323_));
 sg13g2_a22oi_1 _26161_ (.Y(_07324_),
    .B1(_05607_),
    .B2(_03171_),
    .A2(_00255_),
    .A1(net951));
 sg13g2_a22oi_1 _26162_ (.Y(_07325_),
    .B1(_07160_),
    .B2(_07324_),
    .A2(_11048_),
    .A1(_03171_));
 sg13g2_nor3_1 _26163_ (.A(_08557_),
    .B(_08617_),
    .C(_07325_),
    .Y(_07326_));
 sg13g2_buf_2 _26164_ (.A(_07326_),
    .X(_07327_));
 sg13g2_o21ai_1 _26165_ (.B1(_07327_),
    .Y(_07328_),
    .A1(_07158_),
    .A2(net184));
 sg13g2_nor2_1 _26166_ (.A(_09880_),
    .B(_07322_),
    .Y(_07329_));
 sg13g2_buf_2 _26167_ (.A(_07329_),
    .X(_07330_));
 sg13g2_buf_1 _26168_ (.A(_07330_),
    .X(_07331_));
 sg13g2_a22oi_1 _26169_ (.Y(_07332_),
    .B1(net133),
    .B2(_07158_),
    .A2(_07328_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26170_ (.A(net610),
    .B(_07332_),
    .Y(_01109_));
 sg13g2_nor2b_1 _26171_ (.A(net184),
    .B_N(_07180_),
    .Y(_07333_));
 sg13g2_buf_1 _26172_ (.A(net184),
    .X(_07334_));
 sg13g2_buf_1 _26173_ (.A(_07327_),
    .X(_07335_));
 sg13g2_o21ai_1 _26174_ (.B1(net215),
    .Y(_07336_),
    .A1(_05673_),
    .A2(net159));
 sg13g2_a22oi_1 _26175_ (.Y(_07337_),
    .B1(_07336_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07333_),
    .A1(_07174_));
 sg13g2_nor2_1 _26176_ (.A(net610),
    .B(_07337_),
    .Y(_01110_));
 sg13g2_o21ai_1 _26177_ (.B1(net215),
    .Y(_07338_),
    .A1(_05678_),
    .A2(net159));
 sg13g2_a22oi_1 _26178_ (.Y(_07339_),
    .B1(_07338_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(net133),
    .A1(_05678_));
 sg13g2_nor2_1 _26179_ (.A(net610),
    .B(_07339_),
    .Y(_01111_));
 sg13g2_o21ai_1 _26180_ (.B1(net215),
    .Y(_07340_),
    .A1(_07197_),
    .A2(net159));
 sg13g2_a22oi_1 _26181_ (.Y(_07341_),
    .B1(_07340_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07333_),
    .A1(_07191_));
 sg13g2_nor2_1 _26182_ (.A(net610),
    .B(_07341_),
    .Y(_01112_));
 sg13g2_o21ai_1 _26183_ (.B1(net215),
    .Y(_07342_),
    .A1(_07202_),
    .A2(net159));
 sg13g2_a22oi_1 _26184_ (.Y(_07343_),
    .B1(_07342_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net133),
    .A1(_07202_));
 sg13g2_nor2_1 _26185_ (.A(net610),
    .B(_07343_),
    .Y(_01113_));
 sg13g2_o21ai_1 _26186_ (.B1(_07335_),
    .Y(_07344_),
    .A1(_07207_),
    .A2(net159));
 sg13g2_a22oi_1 _26187_ (.Y(_07345_),
    .B1(_07344_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07333_),
    .A1(_07206_));
 sg13g2_nor2_1 _26188_ (.A(net610),
    .B(_07345_),
    .Y(_01114_));
 sg13g2_o21ai_1 _26189_ (.B1(_07335_),
    .Y(_07346_),
    .A1(_07211_),
    .A2(net159));
 sg13g2_a22oi_1 _26190_ (.Y(_07347_),
    .B1(_07346_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net133),
    .A1(_07211_));
 sg13g2_nor2_1 _26191_ (.A(net610),
    .B(_07347_),
    .Y(_01115_));
 sg13g2_a21oi_1 _26192_ (.A1(_03171_),
    .A2(_11112_),
    .Y(_07348_),
    .B1(_07321_));
 sg13g2_nor2b_1 _26193_ (.A(_07348_),
    .B_N(_08619_),
    .Y(_07349_));
 sg13g2_buf_2 _26194_ (.A(_07349_),
    .X(_07350_));
 sg13g2_buf_1 _26195_ (.A(_07350_),
    .X(_07351_));
 sg13g2_o21ai_1 _26196_ (.B1(net158),
    .Y(_07352_),
    .A1(_07220_),
    .A2(net159));
 sg13g2_a22oi_1 _26197_ (.Y(_07353_),
    .B1(_07352_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07333_),
    .A1(_07216_));
 sg13g2_nor2_1 _26198_ (.A(_07320_),
    .B(_07353_),
    .Y(_01116_));
 sg13g2_o21ai_1 _26199_ (.B1(_07351_),
    .Y(_07354_),
    .A1(_07235_),
    .A2(_07334_));
 sg13g2_a22oi_1 _26200_ (.Y(_07355_),
    .B1(_07354_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net133),
    .A1(_07235_));
 sg13g2_nor2_1 _26201_ (.A(_07320_),
    .B(_07355_),
    .Y(_01117_));
 sg13g2_nor2_1 _26202_ (.A(_07233_),
    .B(net184),
    .Y(_07356_));
 sg13g2_o21ai_1 _26203_ (.B1(net158),
    .Y(_07357_),
    .A1(_05719_),
    .A2(_07334_));
 sg13g2_a22oi_1 _26204_ (.Y(_07358_),
    .B1(_07357_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07356_),
    .A1(_07174_));
 sg13g2_nor2_1 _26205_ (.A(net610),
    .B(_07358_),
    .Y(_01118_));
 sg13g2_buf_1 _26206_ (.A(_09103_),
    .X(_07359_));
 sg13g2_buf_1 _26207_ (.A(_07323_),
    .X(_07360_));
 sg13g2_o21ai_1 _26208_ (.B1(net158),
    .Y(_07361_),
    .A1(_05728_),
    .A2(net157));
 sg13g2_a22oi_1 _26209_ (.Y(_07362_),
    .B1(_07361_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net133),
    .A1(_05728_));
 sg13g2_nor2_1 _26210_ (.A(net609),
    .B(_07362_),
    .Y(_01119_));
 sg13g2_o21ai_1 _26211_ (.B1(net215),
    .Y(_07363_),
    .A1(_07248_),
    .A2(net157));
 sg13g2_a22oi_1 _26212_ (.Y(_07364_),
    .B1(_07363_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net133),
    .A1(_07248_));
 sg13g2_nor2_1 _26213_ (.A(net609),
    .B(_07364_),
    .Y(_01120_));
 sg13g2_o21ai_1 _26214_ (.B1(net158),
    .Y(_07365_),
    .A1(_07252_),
    .A2(net157));
 sg13g2_a22oi_1 _26215_ (.Y(_07366_),
    .B1(_07365_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07356_),
    .A1(_07191_));
 sg13g2_nor2_1 _26216_ (.A(net609),
    .B(_07366_),
    .Y(_01121_));
 sg13g2_o21ai_1 _26217_ (.B1(net158),
    .Y(_07367_),
    .A1(_07255_),
    .A2(net157));
 sg13g2_a22oi_1 _26218_ (.Y(_07368_),
    .B1(_07367_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net133),
    .A1(_07255_));
 sg13g2_nor2_1 _26219_ (.A(net609),
    .B(_07368_),
    .Y(_01122_));
 sg13g2_o21ai_1 _26220_ (.B1(net158),
    .Y(_07369_),
    .A1(_07258_),
    .A2(net157));
 sg13g2_a22oi_1 _26221_ (.Y(_07370_),
    .B1(_07369_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07356_),
    .A1(_07206_));
 sg13g2_nor2_1 _26222_ (.A(net609),
    .B(_07370_),
    .Y(_01123_));
 sg13g2_o21ai_1 _26223_ (.B1(net158),
    .Y(_07371_),
    .A1(_07261_),
    .A2(_07360_));
 sg13g2_a22oi_1 _26224_ (.Y(_07372_),
    .B1(_07371_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(_07331_),
    .A1(_07261_));
 sg13g2_nor2_1 _26225_ (.A(_07359_),
    .B(_07372_),
    .Y(_01124_));
 sg13g2_o21ai_1 _26226_ (.B1(_07351_),
    .Y(_07373_),
    .A1(_07265_),
    .A2(_07360_));
 sg13g2_a22oi_1 _26227_ (.Y(_07374_),
    .B1(_07373_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07356_),
    .A1(_07216_));
 sg13g2_nor2_1 _26228_ (.A(net609),
    .B(_07374_),
    .Y(_01125_));
 sg13g2_o21ai_1 _26229_ (.B1(net158),
    .Y(_07375_),
    .A1(_07272_),
    .A2(net157));
 sg13g2_a22oi_1 _26230_ (.Y(_07376_),
    .B1(_07375_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(_07331_),
    .A1(_07272_));
 sg13g2_nor2_1 _26231_ (.A(_07359_),
    .B(_07376_),
    .Y(_01126_));
 sg13g2_nor2b_1 _26232_ (.A(_07323_),
    .B_N(_07270_),
    .Y(_07377_));
 sg13g2_o21ai_1 _26233_ (.B1(_07350_),
    .Y(_07378_),
    .A1(_05763_),
    .A2(net157));
 sg13g2_a22oi_1 _26234_ (.Y(_07379_),
    .B1(_07378_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07377_),
    .A1(_07174_));
 sg13g2_nor2_1 _26235_ (.A(net609),
    .B(_07379_),
    .Y(_01127_));
 sg13g2_o21ai_1 _26236_ (.B1(_07350_),
    .Y(_07380_),
    .A1(_05769_),
    .A2(net157));
 sg13g2_a22oi_1 _26237_ (.Y(_07381_),
    .B1(_07380_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07330_),
    .A1(_05769_));
 sg13g2_nor2_1 _26238_ (.A(net609),
    .B(_07381_),
    .Y(_01128_));
 sg13g2_buf_1 _26239_ (.A(_09103_),
    .X(_07382_));
 sg13g2_buf_1 _26240_ (.A(net184),
    .X(_07383_));
 sg13g2_o21ai_1 _26241_ (.B1(_07350_),
    .Y(_07384_),
    .A1(_07280_),
    .A2(net156));
 sg13g2_a22oi_1 _26242_ (.Y(_07385_),
    .B1(_07384_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07377_),
    .A1(_07191_));
 sg13g2_nor2_1 _26243_ (.A(net608),
    .B(_07385_),
    .Y(_01129_));
 sg13g2_o21ai_1 _26244_ (.B1(_07350_),
    .Y(_07386_),
    .A1(_07284_),
    .A2(net156));
 sg13g2_a22oi_1 _26245_ (.Y(_07387_),
    .B1(_07386_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07330_),
    .A1(_07284_));
 sg13g2_nor2_1 _26246_ (.A(_07382_),
    .B(_07387_),
    .Y(_01130_));
 sg13g2_inv_1 _26247_ (.Y(_07388_),
    .A(net159));
 sg13g2_o21ai_1 _26248_ (.B1(net215),
    .Y(_07389_),
    .A1(_07288_),
    .A2(net156));
 sg13g2_a22oi_1 _26249_ (.Y(_07390_),
    .B1(_07389_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07388_),
    .A1(_07290_));
 sg13g2_nor2_1 _26250_ (.A(net608),
    .B(_07390_),
    .Y(_01131_));
 sg13g2_o21ai_1 _26251_ (.B1(_07350_),
    .Y(_07391_),
    .A1(_07293_),
    .A2(_07383_));
 sg13g2_a22oi_1 _26252_ (.Y(_07392_),
    .B1(_07391_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07377_),
    .A1(_07206_));
 sg13g2_nor2_1 _26253_ (.A(net608),
    .B(_07392_),
    .Y(_01132_));
 sg13g2_o21ai_1 _26254_ (.B1(_07350_),
    .Y(_07393_),
    .A1(_07297_),
    .A2(_07383_));
 sg13g2_a22oi_1 _26255_ (.Y(_07394_),
    .B1(_07393_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07330_),
    .A1(_07297_));
 sg13g2_nor2_1 _26256_ (.A(_07382_),
    .B(_07394_),
    .Y(_01133_));
 sg13g2_o21ai_1 _26257_ (.B1(net215),
    .Y(_07395_),
    .A1(_07300_),
    .A2(net156));
 sg13g2_a22oi_1 _26258_ (.Y(_07396_),
    .B1(_07395_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07330_),
    .A1(_07300_));
 sg13g2_nor2_1 _26259_ (.A(net608),
    .B(_07396_),
    .Y(_01134_));
 sg13g2_nor2_1 _26260_ (.A(_07247_),
    .B(net184),
    .Y(_07397_));
 sg13g2_o21ai_1 _26261_ (.B1(net215),
    .Y(_07398_),
    .A1(_07304_),
    .A2(net156));
 sg13g2_a22oi_1 _26262_ (.Y(_07399_),
    .B1(_07398_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07397_),
    .A1(_07191_));
 sg13g2_nor2_1 _26263_ (.A(net608),
    .B(_07399_),
    .Y(_01135_));
 sg13g2_o21ai_1 _26264_ (.B1(_07327_),
    .Y(_07400_),
    .A1(_05805_),
    .A2(net156));
 sg13g2_a22oi_1 _26265_ (.Y(_07401_),
    .B1(_07400_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07330_),
    .A1(_05805_));
 sg13g2_nor2_1 _26266_ (.A(net608),
    .B(_07401_),
    .Y(_01136_));
 sg13g2_o21ai_1 _26267_ (.B1(_07327_),
    .Y(_07402_),
    .A1(_05811_),
    .A2(net156));
 sg13g2_a22oi_1 _26268_ (.Y(_07403_),
    .B1(_07402_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07397_),
    .A1(_07206_));
 sg13g2_nor2_1 _26269_ (.A(net608),
    .B(_07403_),
    .Y(_01137_));
 sg13g2_o21ai_1 _26270_ (.B1(_07327_),
    .Y(_07404_),
    .A1(_05816_),
    .A2(net156));
 sg13g2_a22oi_1 _26271_ (.Y(_07405_),
    .B1(_07404_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07330_),
    .A1(_05816_));
 sg13g2_nor2_1 _26272_ (.A(net608),
    .B(_07405_),
    .Y(_01138_));
 sg13g2_buf_1 _26273_ (.A(_09103_),
    .X(_07406_));
 sg13g2_o21ai_1 _26274_ (.B1(_07327_),
    .Y(_07407_),
    .A1(_07313_),
    .A2(net184));
 sg13g2_a22oi_1 _26275_ (.Y(_07408_),
    .B1(_07407_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07397_),
    .A1(_07216_));
 sg13g2_nor2_1 _26276_ (.A(_07406_),
    .B(_07408_),
    .Y(_01139_));
 sg13g2_o21ai_1 _26277_ (.B1(_07327_),
    .Y(_07409_),
    .A1(_07317_),
    .A2(net184));
 sg13g2_a22oi_1 _26278_ (.Y(_07410_),
    .B1(_07409_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07330_),
    .A1(_07317_));
 sg13g2_nor2_1 _26279_ (.A(_07406_),
    .B(_07410_),
    .Y(_01140_));
 sg13g2_nor3_1 _26280_ (.A(_11612_),
    .B(_04697_),
    .C(net138),
    .Y(_07411_));
 sg13g2_buf_2 _26281_ (.A(_07411_),
    .X(_07412_));
 sg13g2_nand2_1 _26282_ (.Y(_07413_),
    .A(_05565_),
    .B(_07412_));
 sg13g2_nand4_1 _26283_ (.B(_09497_),
    .C(_04699_),
    .A(net956),
    .Y(_07414_),
    .D(_06093_));
 sg13g2_buf_2 _26284_ (.A(_07414_),
    .X(_07415_));
 sg13g2_nand2_1 _26285_ (.Y(_07416_),
    .A(\cpu.gpio.r_enable_in[0] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26286_ (.A1(_07413_),
    .A2(_07416_),
    .Y(_01941_),
    .B1(net615));
 sg13g2_nand2_1 _26287_ (.Y(_07417_),
    .A(net1004),
    .B(_07412_));
 sg13g2_nand2_1 _26288_ (.Y(_07418_),
    .A(\cpu.gpio.r_enable_in[1] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26289_ (.A1(_07417_),
    .A2(_07418_),
    .Y(_01942_),
    .B1(net615));
 sg13g2_nand2_1 _26290_ (.Y(_07419_),
    .A(net869),
    .B(_07412_));
 sg13g2_nand2_1 _26291_ (.Y(_07420_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26292_ (.A1(_07419_),
    .A2(_07420_),
    .Y(_01943_),
    .B1(net615));
 sg13g2_nand2_1 _26293_ (.Y(_07421_),
    .A(net928),
    .B(_07412_));
 sg13g2_nand2_1 _26294_ (.Y(_07422_),
    .A(\cpu.gpio.r_enable_in[3] ),
    .B(_07415_));
 sg13g2_buf_1 _26295_ (.A(_09103_),
    .X(_07423_));
 sg13g2_a21oi_1 _26296_ (.A1(_07421_),
    .A2(_07422_),
    .Y(_01944_),
    .B1(net606));
 sg13g2_nand2_1 _26297_ (.Y(_07424_),
    .A(net964),
    .B(_07412_));
 sg13g2_nand2_1 _26298_ (.Y(_07425_),
    .A(\cpu.gpio.r_enable_in[4] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26299_ (.A1(_07424_),
    .A2(_07425_),
    .Y(_01945_),
    .B1(_07423_));
 sg13g2_nand2_1 _26300_ (.Y(_07426_),
    .A(_11988_),
    .B(_07412_));
 sg13g2_nand2_1 _26301_ (.Y(_07427_),
    .A(\cpu.gpio.r_enable_in[5] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26302_ (.A1(_07426_),
    .A2(_07427_),
    .Y(_01946_),
    .B1(_07423_));
 sg13g2_nand2_1 _26303_ (.Y(_07428_),
    .A(_06100_),
    .B(_07412_));
 sg13g2_nand2_1 _26304_ (.Y(_07429_),
    .A(_08968_),
    .B(_07415_));
 sg13g2_a21oi_1 _26305_ (.A1(_07428_),
    .A2(_07429_),
    .Y(_01947_),
    .B1(net606));
 sg13g2_nand2_1 _26306_ (.Y(_07430_),
    .A(net1005),
    .B(_07412_));
 sg13g2_nand2_1 _26307_ (.Y(_07431_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_07415_));
 sg13g2_a21oi_1 _26308_ (.A1(_07430_),
    .A2(_07431_),
    .Y(_01948_),
    .B1(net606));
 sg13g2_nor2_1 _26309_ (.A(net381),
    .B(net138),
    .Y(_07432_));
 sg13g2_nand2_1 _26310_ (.Y(_07433_),
    .A(net1007),
    .B(_07432_));
 sg13g2_buf_1 _26311_ (.A(net138),
    .X(_07434_));
 sg13g2_o21ai_1 _26312_ (.B1(_08977_),
    .Y(_07435_),
    .A1(net381),
    .A2(net115));
 sg13g2_a21oi_1 _26313_ (.A1(_07433_),
    .A2(_07435_),
    .Y(_01949_),
    .B1(net606));
 sg13g2_nand2_1 _26314_ (.Y(_07436_),
    .A(net1006),
    .B(_07432_));
 sg13g2_o21ai_1 _26315_ (.B1(_08985_),
    .Y(_07437_),
    .A1(net381),
    .A2(net115));
 sg13g2_a21oi_1 _26316_ (.A1(_07436_),
    .A2(_07437_),
    .Y(_01950_),
    .B1(net606));
 sg13g2_nand2_1 _26317_ (.Y(_07438_),
    .A(net929),
    .B(_07432_));
 sg13g2_o21ai_1 _26318_ (.B1(\cpu.gpio.r_enable_io[6] ),
    .Y(_07439_),
    .A1(net381),
    .A2(net115));
 sg13g2_a21oi_1 _26319_ (.A1(_07438_),
    .A2(_07439_),
    .Y(_01951_),
    .B1(net606));
 sg13g2_nand2_1 _26320_ (.Y(_07440_),
    .A(net1005),
    .B(_07432_));
 sg13g2_o21ai_1 _26321_ (.B1(_08970_),
    .Y(_07441_),
    .A1(net381),
    .A2(net115));
 sg13g2_a21oi_1 _26322_ (.A1(_07440_),
    .A2(_07441_),
    .Y(_01952_),
    .B1(net606));
 sg13g2_nand2_2 _26323_ (.Y(_07442_),
    .A(net822),
    .B(_04973_));
 sg13g2_nor2_1 _26324_ (.A(net138),
    .B(_07442_),
    .Y(_07443_));
 sg13g2_nand2_1 _26325_ (.Y(_07444_),
    .A(_09840_),
    .B(_07443_));
 sg13g2_o21ai_1 _26326_ (.B1(net7),
    .Y(_07445_),
    .A1(net115),
    .A2(_07442_));
 sg13g2_a21oi_1 _26327_ (.A1(_07444_),
    .A2(_07445_),
    .Y(_01953_),
    .B1(net606));
 sg13g2_nand2_1 _26328_ (.Y(_07446_),
    .A(_09846_),
    .B(_07443_));
 sg13g2_o21ai_1 _26329_ (.B1(net8),
    .Y(_07447_),
    .A1(net115),
    .A2(_07442_));
 sg13g2_buf_1 _26330_ (.A(_09103_),
    .X(_07448_));
 sg13g2_a21oi_1 _26331_ (.A1(_07446_),
    .A2(_07447_),
    .Y(_01954_),
    .B1(net605));
 sg13g2_nand2_1 _26332_ (.Y(_07449_),
    .A(net929),
    .B(_07443_));
 sg13g2_o21ai_1 _26333_ (.B1(net9),
    .Y(_07450_),
    .A1(net138),
    .A2(_07442_));
 sg13g2_a21oi_1 _26334_ (.A1(_07449_),
    .A2(_07450_),
    .Y(_01955_),
    .B1(net605));
 sg13g2_nand2_1 _26335_ (.Y(_07451_),
    .A(net1005),
    .B(_07443_));
 sg13g2_o21ai_1 _26336_ (.B1(net10),
    .Y(_07452_),
    .A1(net138),
    .A2(_07442_));
 sg13g2_a21oi_1 _26337_ (.A1(_07451_),
    .A2(_07452_),
    .Y(_01956_),
    .B1(net605));
 sg13g2_nor3_1 _26338_ (.A(net942),
    .B(net352),
    .C(net115),
    .Y(_07453_));
 sg13g2_nor2_1 _26339_ (.A(net352),
    .B(_06095_),
    .Y(_07454_));
 sg13g2_nor2_1 _26340_ (.A(_04720_),
    .B(_07454_),
    .Y(_07455_));
 sg13g2_o21ai_1 _26341_ (.B1(net623),
    .Y(_02002_),
    .A1(_07453_),
    .A2(_07455_));
 sg13g2_nand2_1 _26342_ (.Y(_07456_),
    .A(_09883_),
    .B(_07454_));
 sg13g2_buf_1 _26343_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07457_));
 sg13g2_o21ai_1 _26344_ (.B1(_07457_),
    .Y(_07458_),
    .A1(net352),
    .A2(_07434_));
 sg13g2_a21oi_1 _26345_ (.A1(_07456_),
    .A2(_07458_),
    .Y(_02003_),
    .B1(net605));
 sg13g2_nand2_1 _26346_ (.Y(_07459_),
    .A(_09889_),
    .B(_07454_));
 sg13g2_o21ai_1 _26347_ (.B1(\cpu.gpio.r_src_o[6][2] ),
    .Y(_07460_),
    .A1(net352),
    .A2(_07434_));
 sg13g2_a21oi_1 _26348_ (.A1(_07459_),
    .A2(_07460_),
    .Y(_02004_),
    .B1(net605));
 sg13g2_nand2_1 _26349_ (.Y(_07461_),
    .A(net928),
    .B(_07454_));
 sg13g2_o21ai_1 _26350_ (.B1(\cpu.gpio.r_src_o[6][3] ),
    .Y(_07462_),
    .A1(net352),
    .A2(net115));
 sg13g2_a21oi_1 _26351_ (.A1(_07461_),
    .A2(_07462_),
    .Y(_02005_),
    .B1(net605));
 sg13g2_nor4_2 _26352_ (.A(net643),
    .B(net530),
    .C(net717),
    .Y(_07463_),
    .D(net138));
 sg13g2_mux2_1 _26353_ (.A0(_04725_),
    .A1(_05564_),
    .S(_07463_),
    .X(_07464_));
 sg13g2_and2_1 _26354_ (.A(net691),
    .B(_07464_),
    .X(_02010_));
 sg13g2_nand2_1 _26355_ (.Y(_07465_),
    .A(_09883_),
    .B(_07463_));
 sg13g2_nand2b_1 _26356_ (.Y(_07466_),
    .B(\cpu.gpio.r_uart_rx_src[1] ),
    .A_N(_07463_));
 sg13g2_a21oi_1 _26357_ (.A1(_07465_),
    .A2(_07466_),
    .Y(_02011_),
    .B1(_07448_));
 sg13g2_nand2_1 _26358_ (.Y(_07467_),
    .A(net869),
    .B(_07463_));
 sg13g2_nand2b_1 _26359_ (.Y(_07468_),
    .B(\cpu.gpio.r_uart_rx_src[2] ),
    .A_N(_07463_));
 sg13g2_a21oi_1 _26360_ (.A1(_07467_),
    .A2(_07468_),
    .Y(_02012_),
    .B1(_07448_));
 sg13g2_and2_1 _26361_ (.A(\cpu.i_wstrobe_d ),
    .B(_00316_),
    .X(_02269_));
 sg13g2_nor2_1 _26362_ (.A(_06151_),
    .B(_06163_),
    .Y(_07469_));
 sg13g2_nor2_1 _26363_ (.A(_06177_),
    .B(_07469_),
    .Y(_02270_));
 sg13g2_xor2_1 _26364_ (.B(_06158_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_07470_));
 sg13g2_nor2_1 _26365_ (.A(_06177_),
    .B(_07470_),
    .Y(_02271_));
 sg13g2_xnor2_1 _26366_ (.Y(_07471_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_04978_));
 sg13g2_xnor2_1 _26367_ (.Y(_07472_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_09911_));
 sg13g2_xnor2_1 _26368_ (.Y(_07473_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05546_));
 sg13g2_xnor2_1 _26369_ (.Y(_07474_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_09916_));
 sg13g2_nand4_1 _26370_ (.B(_07472_),
    .C(_07473_),
    .A(_07471_),
    .Y(_07475_),
    .D(_07474_));
 sg13g2_xnor2_1 _26371_ (.Y(_07476_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05531_));
 sg13g2_xnor2_1 _26372_ (.Y(_07477_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05233_));
 sg13g2_xnor2_1 _26373_ (.Y(_07478_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05442_));
 sg13g2_xnor2_1 _26374_ (.Y(_07479_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_09939_));
 sg13g2_nand4_1 _26375_ (.B(_07477_),
    .C(_07478_),
    .A(_07476_),
    .Y(_07480_),
    .D(_07479_));
 sg13g2_xnor2_1 _26376_ (.Y(_07481_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_09923_));
 sg13g2_xnor2_1 _26377_ (.Y(_07482_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_09928_));
 sg13g2_xnor2_1 _26378_ (.Y(_07483_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_09906_));
 sg13g2_xnor2_1 _26379_ (.Y(_07484_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_09955_));
 sg13g2_nand4_1 _26380_ (.B(_07482_),
    .C(_07483_),
    .A(_07481_),
    .Y(_07485_),
    .D(_07484_));
 sg13g2_xnor2_1 _26381_ (.Y(_07486_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_09944_));
 sg13g2_xnor2_1 _26382_ (.Y(_07487_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_09950_));
 sg13g2_xnor2_1 _26383_ (.Y(_07488_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_04859_));
 sg13g2_xnor2_1 _26384_ (.Y(_07489_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_09891_));
 sg13g2_nand4_1 _26385_ (.B(_07487_),
    .C(_07488_),
    .A(_07486_),
    .Y(_07490_),
    .D(_07489_));
 sg13g2_nor4_1 _26386_ (.A(_07475_),
    .B(_07480_),
    .C(_07485_),
    .D(_07490_),
    .Y(_07491_));
 sg13g2_xnor2_1 _26387_ (.Y(_07492_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05295_));
 sg13g2_xnor2_1 _26388_ (.Y(_07493_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05085_));
 sg13g2_xnor2_1 _26389_ (.Y(_07494_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_09896_));
 sg13g2_xnor2_1 _26390_ (.Y(_07495_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_09877_));
 sg13g2_nand4_1 _26391_ (.B(_07493_),
    .C(_07494_),
    .A(_07492_),
    .Y(_07496_),
    .D(_07495_));
 sg13g2_xnor2_1 _26392_ (.Y(_07497_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05169_));
 sg13g2_xnor2_1 _26393_ (.Y(_07498_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_09901_));
 sg13g2_xnor2_1 _26394_ (.Y(_07499_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05051_));
 sg13g2_xnor2_1 _26395_ (.Y(_07500_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05030_));
 sg13g2_nand4_1 _26396_ (.B(_07498_),
    .C(_07499_),
    .A(_07497_),
    .Y(_07501_),
    .D(_07500_));
 sg13g2_xnor2_1 _26397_ (.Y(_07502_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05470_));
 sg13g2_xnor2_1 _26398_ (.Y(_07503_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05005_));
 sg13g2_xnor2_1 _26399_ (.Y(_07504_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_09932_));
 sg13g2_xnor2_1 _26400_ (.Y(_07505_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_09886_));
 sg13g2_nand4_1 _26401_ (.B(_07503_),
    .C(_07504_),
    .A(_07502_),
    .Y(_07506_),
    .D(_07505_));
 sg13g2_xnor2_1 _26402_ (.Y(_07507_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04741_));
 sg13g2_xnor2_1 _26403_ (.Y(_07508_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_09876_));
 sg13g2_xnor2_1 _26404_ (.Y(_07509_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_04930_));
 sg13g2_xnor2_1 _26405_ (.Y(_07510_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05343_));
 sg13g2_nand4_1 _26406_ (.B(_07508_),
    .C(_07509_),
    .A(_07507_),
    .Y(_07511_),
    .D(_07510_));
 sg13g2_nor4_1 _26407_ (.A(_07496_),
    .B(_07501_),
    .C(_07506_),
    .D(_07511_),
    .Y(_07512_));
 sg13g2_a22oi_1 _26408_ (.Y(_07513_),
    .B1(_07491_),
    .B2(_07512_),
    .A2(_07112_),
    .A1(net1009));
 sg13g2_nand3_1 _26409_ (.B(net183),
    .C(_04766_),
    .A(net1009),
    .Y(_07514_));
 sg13g2_nand2_1 _26410_ (.Y(_07515_),
    .A(\cpu.intr.r_clock ),
    .B(_07514_));
 sg13g2_a21oi_1 _26411_ (.A1(_07513_),
    .A2(_07515_),
    .Y(_02432_),
    .B1(net605));
 sg13g2_and2_1 _26412_ (.A(net183),
    .B(net431),
    .X(_07516_));
 sg13g2_buf_1 _26413_ (.A(_07516_),
    .X(_07517_));
 sg13g2_nand2_1 _26414_ (.Y(_07518_),
    .A(net821),
    .B(_07517_));
 sg13g2_nand2_1 _26415_ (.Y(_07519_),
    .A(net183),
    .B(_04735_));
 sg13g2_buf_1 _26416_ (.A(_07519_),
    .X(_07520_));
 sg13g2_nand2_1 _26417_ (.Y(_07521_),
    .A(_09003_),
    .B(_07520_));
 sg13g2_a21oi_1 _26418_ (.A1(_07518_),
    .A2(_07521_),
    .Y(_02481_),
    .B1(net605));
 sg13g2_nand2_1 _26419_ (.Y(_07522_),
    .A(net1004),
    .B(_07517_));
 sg13g2_nand2_1 _26420_ (.Y(_07523_),
    .A(_08997_),
    .B(_07520_));
 sg13g2_buf_1 _26421_ (.A(_09096_),
    .X(_07524_));
 sg13g2_a21oi_1 _26422_ (.A1(_07522_),
    .A2(_07523_),
    .Y(_02482_),
    .B1(net604));
 sg13g2_nand2_1 _26423_ (.Y(_07525_),
    .A(net869),
    .B(_07517_));
 sg13g2_nand2_1 _26424_ (.Y(_07526_),
    .A(\cpu.intr.r_enable[2] ),
    .B(_07520_));
 sg13g2_a21oi_1 _26425_ (.A1(_07525_),
    .A2(_07526_),
    .Y(_02483_),
    .B1(net604));
 sg13g2_nand2_1 _26426_ (.Y(_07527_),
    .A(net928),
    .B(_07517_));
 sg13g2_nand2_1 _26427_ (.Y(_07528_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07520_));
 sg13g2_a21oi_1 _26428_ (.A1(_07527_),
    .A2(_07528_),
    .Y(_02484_),
    .B1(net604));
 sg13g2_nand2_1 _26429_ (.Y(_07529_),
    .A(net1007),
    .B(_07517_));
 sg13g2_nand2_1 _26430_ (.Y(_07530_),
    .A(_08992_),
    .B(_07520_));
 sg13g2_a21oi_1 _26431_ (.A1(_07529_),
    .A2(_07530_),
    .Y(_02485_),
    .B1(net604));
 sg13g2_nand2_1 _26432_ (.Y(_07531_),
    .A(net1006),
    .B(_07517_));
 sg13g2_nand2_1 _26433_ (.Y(_07532_),
    .A(_08999_),
    .B(_07520_));
 sg13g2_a21oi_1 _26434_ (.A1(_07531_),
    .A2(_07532_),
    .Y(_02486_),
    .B1(net604));
 sg13g2_nand3_1 _26435_ (.B(net183),
    .C(_04766_),
    .A(_09825_),
    .Y(_07533_));
 sg13g2_inv_1 _26436_ (.Y(_07534_),
    .A(_09769_));
 sg13g2_a221oi_1 _26437_ (.B2(_08994_),
    .C1(_07534_),
    .B1(_07533_),
    .A1(net1008),
    .Y(_07535_),
    .A2(_07112_));
 sg13g2_nor2_1 _26438_ (.A(net607),
    .B(_07535_),
    .Y(_02487_));
 sg13g2_and2_1 _26439_ (.A(_09576_),
    .B(_06631_),
    .X(_07536_));
 sg13g2_nand4_1 _26440_ (.B(_06639_),
    .C(_06632_),
    .A(_09626_),
    .Y(_07537_),
    .D(_07536_));
 sg13g2_buf_1 _26441_ (.A(_07537_),
    .X(_07538_));
 sg13g2_o21ai_1 _26442_ (.B1(net761),
    .Y(_07539_),
    .A1(_06638_),
    .A2(_07538_));
 sg13g2_nor2b_1 _26443_ (.A(_09619_),
    .B_N(_09603_),
    .Y(_07540_));
 sg13g2_o21ai_1 _26444_ (.B1(net19),
    .Y(_07541_),
    .A1(_07538_),
    .A2(_07540_));
 sg13g2_nand2b_1 _26445_ (.Y(_02517_),
    .B(_07541_),
    .A_N(_07539_));
 sg13g2_nand3b_1 _26446_ (.B(_06614_),
    .C(_09578_),
    .Y(_07542_),
    .A_N(_09603_));
 sg13g2_a21o_1 _26447_ (.A2(_07542_),
    .A1(_06638_),
    .B1(_07538_),
    .X(_07543_));
 sg13g2_nand2_1 _26448_ (.Y(_07544_),
    .A(_09603_),
    .B(_06638_));
 sg13g2_nor2_1 _26449_ (.A(_09615_),
    .B(_07544_),
    .Y(_07545_));
 sg13g2_o21ai_1 _26450_ (.B1(net20),
    .Y(_07546_),
    .A1(_07538_),
    .A2(_07545_));
 sg13g2_nand3_1 _26451_ (.B(_07543_),
    .C(_07546_),
    .A(net622),
    .Y(_02518_));
 sg13g2_nor2b_1 _26452_ (.A(_09617_),
    .B_N(_09603_),
    .Y(_07547_));
 sg13g2_buf_1 _26453_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07548_));
 sg13g2_o21ai_1 _26454_ (.B1(_07548_),
    .Y(_07549_),
    .A1(_07538_),
    .A2(_07547_));
 sg13g2_nand2b_1 _26455_ (.Y(_02519_),
    .B(_07549_),
    .A_N(_07539_));
 sg13g2_nor3_1 _26456_ (.A(_09129_),
    .B(_09589_),
    .C(_06614_),
    .Y(_07550_));
 sg13g2_nand3_1 _26457_ (.B(_06507_),
    .C(_07550_),
    .A(_06500_),
    .Y(_07551_));
 sg13g2_nor3_1 _26458_ (.A(_09598_),
    .B(_06630_),
    .C(_07551_),
    .Y(_07552_));
 sg13g2_a21oi_1 _26459_ (.A1(_06639_),
    .A2(_07552_),
    .Y(_07553_),
    .B1(_09578_));
 sg13g2_nor2_1 _26460_ (.A(net607),
    .B(_07553_),
    .Y(_02520_));
 sg13g2_nand2_1 _26461_ (.Y(_07554_),
    .A(_09857_),
    .B(_06548_));
 sg13g2_nand2_1 _26462_ (.Y(_07555_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06551_));
 sg13g2_a21oi_1 _26463_ (.A1(_07554_),
    .A2(_07555_),
    .Y(_02521_),
    .B1(_07524_));
 sg13g2_nor4_1 _26464_ (.A(net945),
    .B(_06790_),
    .C(_04749_),
    .D(net137),
    .Y(_07556_));
 sg13g2_a21oi_1 _26465_ (.A1(\cpu.qspi.r_mask[1] ),
    .A2(_06562_),
    .Y(_07557_),
    .B1(_07556_));
 sg13g2_nand2_1 _26466_ (.Y(_02522_),
    .A(net623),
    .B(_07557_));
 sg13g2_nand2_1 _26467_ (.Y(_07558_),
    .A(_06790_),
    .B(_06572_));
 sg13g2_o21ai_1 _26468_ (.B1(_07558_),
    .Y(_07559_),
    .A1(\cpu.qspi.r_mask[2] ),
    .A2(_06572_));
 sg13g2_nor2_1 _26469_ (.A(net607),
    .B(_07559_),
    .Y(_02523_));
 sg13g2_nand2_1 _26470_ (.Y(_07560_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06551_));
 sg13g2_nand2_1 _26471_ (.Y(_07561_),
    .A(_06100_),
    .B(_06548_));
 sg13g2_nand3_1 _26472_ (.B(_07560_),
    .C(_07561_),
    .A(net622),
    .Y(_02524_));
 sg13g2_nor4_1 _26473_ (.A(net945),
    .B(_06786_),
    .C(_04749_),
    .D(net137),
    .Y(_07562_));
 sg13g2_a21oi_1 _26474_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06562_),
    .Y(_07563_),
    .B1(_07562_));
 sg13g2_nor2_1 _26475_ (.A(net607),
    .B(_07563_),
    .Y(_02525_));
 sg13g2_nand2_1 _26476_ (.Y(_07564_),
    .A(_06786_),
    .B(_06572_));
 sg13g2_o21ai_1 _26477_ (.B1(_07564_),
    .Y(_07565_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06572_));
 sg13g2_nand2_1 _26478_ (.Y(_02526_),
    .A(net623),
    .B(_07565_));
 sg13g2_nor2_1 _26479_ (.A(_04714_),
    .B(_06546_),
    .Y(_07566_));
 sg13g2_nand2_1 _26480_ (.Y(_07567_),
    .A(net821),
    .B(_07566_));
 sg13g2_o21ai_1 _26481_ (.B1(_09607_),
    .Y(_07568_),
    .A1(_04714_),
    .A2(net137));
 sg13g2_nand3_1 _26482_ (.B(_07567_),
    .C(_07568_),
    .A(net622),
    .Y(_02539_));
 sg13g2_nor3_1 _26483_ (.A(_09819_),
    .B(_04714_),
    .C(_06546_),
    .Y(_07569_));
 sg13g2_nor2_1 _26484_ (.A(_09606_),
    .B(_07566_),
    .Y(_07570_));
 sg13g2_o21ai_1 _26485_ (.B1(net623),
    .Y(_02540_),
    .A1(_07569_),
    .A2(_07570_));
 sg13g2_inv_1 _26486_ (.Y(_07571_),
    .A(_06614_));
 sg13g2_nor4_1 _26487_ (.A(_11549_),
    .B(_09627_),
    .C(\cpu.qspi.r_state[11] ),
    .D(_06614_),
    .Y(_07572_));
 sg13g2_nand2_1 _26488_ (.Y(_07573_),
    .A(_06499_),
    .B(_07572_));
 sg13g2_nand3_1 _26489_ (.B(_07571_),
    .C(_07573_),
    .A(_11547_),
    .Y(_07574_));
 sg13g2_nand2b_1 _26490_ (.Y(_07575_),
    .B(_11549_),
    .A_N(_06637_));
 sg13g2_nor3_1 _26491_ (.A(_11569_),
    .B(_09669_),
    .C(_09601_),
    .Y(_07576_));
 sg13g2_and4_1 _26492_ (.A(_06507_),
    .B(_07536_),
    .C(_07575_),
    .D(_07576_),
    .X(_07577_));
 sg13g2_buf_1 _26493_ (.A(_07577_),
    .X(_07578_));
 sg13g2_mux2_1 _26494_ (.A0(net3),
    .A1(_07574_),
    .S(_07578_),
    .X(_07579_));
 sg13g2_and2_1 _26495_ (.A(net691),
    .B(_07579_),
    .X(_02541_));
 sg13g2_nand2b_1 _26496_ (.Y(_07580_),
    .B(net6),
    .A_N(_07578_));
 sg13g2_o21ai_1 _26497_ (.B1(_11547_),
    .Y(_07581_),
    .A1(_09622_),
    .A2(_07573_));
 sg13g2_nand2_1 _26498_ (.Y(_07582_),
    .A(_07578_),
    .B(_07581_));
 sg13g2_a21oi_1 _26499_ (.A1(_07580_),
    .A2(_07582_),
    .Y(_02542_),
    .B1(_07524_));
 sg13g2_nor3_1 _26500_ (.A(_09031_),
    .B(net1084),
    .C(_09045_),
    .Y(_07583_));
 sg13g2_a221oi_1 _26501_ (.B2(net1017),
    .C1(_07583_),
    .B1(net406),
    .A1(net1084),
    .Y(_07584_),
    .A2(net130));
 sg13g2_buf_1 _26502_ (.A(_07584_),
    .X(_07585_));
 sg13g2_nand3_1 _26503_ (.B(net1017),
    .C(_07585_),
    .A(_09050_),
    .Y(_07586_));
 sg13g2_o21ai_1 _26504_ (.B1(_07586_),
    .Y(_07587_),
    .A1(_09050_),
    .A2(_07585_));
 sg13g2_nand2_1 _26505_ (.Y(_02548_),
    .A(net623),
    .B(_07587_));
 sg13g2_nand2_1 _26506_ (.Y(_07588_),
    .A(_09050_),
    .B(_11577_));
 sg13g2_a21oi_1 _26507_ (.A1(_07585_),
    .A2(_07588_),
    .Y(_07589_),
    .B1(_09051_));
 sg13g2_inv_1 _26508_ (.Y(_07590_),
    .A(_09050_));
 sg13g2_and4_1 _26509_ (.A(_07590_),
    .B(_09051_),
    .C(_11577_),
    .D(_07585_),
    .X(_07591_));
 sg13g2_o21ai_1 _26510_ (.B1(net623),
    .Y(_02549_),
    .A1(_07589_),
    .A2(_07591_));
 sg13g2_nor2_1 _26511_ (.A(_09050_),
    .B(_09051_),
    .Y(_07592_));
 sg13g2_or2_1 _26512_ (.X(_07593_),
    .B(_07592_),
    .A(_00226_));
 sg13g2_a21oi_1 _26513_ (.A1(_07585_),
    .A2(_07593_),
    .Y(_07594_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _26514_ (.A(\cpu.spi.r_bits[2] ),
    .B(_11577_),
    .C(_07592_),
    .D(_07585_),
    .X(_07595_));
 sg13g2_o21ai_1 _26515_ (.B1(net623),
    .Y(_02550_),
    .A1(_07594_),
    .A2(_07595_));
 sg13g2_nor3_1 _26516_ (.A(net852),
    .B(_04778_),
    .C(_09024_),
    .Y(_07596_));
 sg13g2_buf_2 _26517_ (.A(_07596_),
    .X(_07597_));
 sg13g2_and2_1 _26518_ (.A(_04783_),
    .B(_07597_),
    .X(_07598_));
 sg13g2_buf_2 _26519_ (.A(_07598_),
    .X(_07599_));
 sg13g2_nand2_1 _26520_ (.Y(_07600_),
    .A(net942),
    .B(_07599_));
 sg13g2_nand2_1 _26521_ (.Y(_07601_),
    .A(_04783_),
    .B(_07597_));
 sg13g2_buf_2 _26522_ (.A(_07601_),
    .X(_07602_));
 sg13g2_nand2_1 _26523_ (.Y(_07603_),
    .A(\cpu.spi.r_clk_count[0][0] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26524_ (.A1(_07600_),
    .A2(_07603_),
    .Y(_02551_),
    .B1(net604));
 sg13g2_nand2_1 _26525_ (.Y(_07604_),
    .A(net1004),
    .B(_07599_));
 sg13g2_nand2_1 _26526_ (.Y(_07605_),
    .A(\cpu.spi.r_clk_count[0][1] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26527_ (.A1(_07604_),
    .A2(_07605_),
    .Y(_02552_),
    .B1(net604));
 sg13g2_nand2_1 _26528_ (.Y(_07606_),
    .A(net869),
    .B(_07599_));
 sg13g2_nand2_1 _26529_ (.Y(_07607_),
    .A(\cpu.spi.r_clk_count[0][2] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26530_ (.A1(_07606_),
    .A2(_07607_),
    .Y(_02553_),
    .B1(net604));
 sg13g2_nand2_1 _26531_ (.Y(_07608_),
    .A(net928),
    .B(_07599_));
 sg13g2_nand2_1 _26532_ (.Y(_07609_),
    .A(\cpu.spi.r_clk_count[0][3] ),
    .B(_07602_));
 sg13g2_buf_1 _26533_ (.A(_09096_),
    .X(_07610_));
 sg13g2_a21oi_1 _26534_ (.A1(_07608_),
    .A2(_07609_),
    .Y(_02554_),
    .B1(_07610_));
 sg13g2_nand2_1 _26535_ (.Y(_07611_),
    .A(net1007),
    .B(_07599_));
 sg13g2_nand2_1 _26536_ (.Y(_07612_),
    .A(\cpu.spi.r_clk_count[0][4] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26537_ (.A1(_07611_),
    .A2(_07612_),
    .Y(_02555_),
    .B1(net603));
 sg13g2_nand2_1 _26538_ (.Y(_07613_),
    .A(net1006),
    .B(_07599_));
 sg13g2_nand2_1 _26539_ (.Y(_07614_),
    .A(\cpu.spi.r_clk_count[0][5] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26540_ (.A1(_07613_),
    .A2(_07614_),
    .Y(_02556_),
    .B1(net603));
 sg13g2_nand2_1 _26541_ (.Y(_07615_),
    .A(net929),
    .B(_07599_));
 sg13g2_nand2_1 _26542_ (.Y(_07616_),
    .A(\cpu.spi.r_clk_count[0][6] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26543_ (.A1(_07615_),
    .A2(_07616_),
    .Y(_02557_),
    .B1(net603));
 sg13g2_nand2_1 _26544_ (.Y(_07617_),
    .A(_09856_),
    .B(_07599_));
 sg13g2_nand2_1 _26545_ (.Y(_07618_),
    .A(\cpu.spi.r_clk_count[0][7] ),
    .B(_07602_));
 sg13g2_a21oi_1 _26546_ (.A1(_07617_),
    .A2(_07618_),
    .Y(_02558_),
    .B1(_07610_));
 sg13g2_nand2_1 _26547_ (.Y(_07619_),
    .A(net573),
    .B(_07597_));
 sg13g2_or2_1 _26548_ (.X(_07620_),
    .B(_07619_),
    .A(net557));
 sg13g2_buf_2 _26549_ (.A(_07620_),
    .X(_07621_));
 sg13g2_nand2_1 _26550_ (.Y(_07622_),
    .A(\cpu.spi.r_clk_count[1][0] ),
    .B(_07621_));
 sg13g2_nor2_1 _26551_ (.A(net557),
    .B(_07619_),
    .Y(_07623_));
 sg13g2_buf_2 _26552_ (.A(_07623_),
    .X(_07624_));
 sg13g2_nand2_1 _26553_ (.Y(_07625_),
    .A(net942),
    .B(_07624_));
 sg13g2_a21oi_1 _26554_ (.A1(_07622_),
    .A2(_07625_),
    .Y(_02559_),
    .B1(net603));
 sg13g2_nand2_1 _26555_ (.Y(_07626_),
    .A(\cpu.spi.r_clk_count[1][1] ),
    .B(_07621_));
 sg13g2_nand2_1 _26556_ (.Y(_07627_),
    .A(net1004),
    .B(_07624_));
 sg13g2_a21oi_1 _26557_ (.A1(_07626_),
    .A2(_07627_),
    .Y(_02560_),
    .B1(net603));
 sg13g2_nand2_1 _26558_ (.Y(_07628_),
    .A(\cpu.spi.r_clk_count[1][2] ),
    .B(_07621_));
 sg13g2_nand2_1 _26559_ (.Y(_07629_),
    .A(net869),
    .B(_07624_));
 sg13g2_a21oi_1 _26560_ (.A1(_07628_),
    .A2(_07629_),
    .Y(_02561_),
    .B1(net603));
 sg13g2_nand2_1 _26561_ (.Y(_07630_),
    .A(\cpu.spi.r_clk_count[1][3] ),
    .B(_07621_));
 sg13g2_nand2_1 _26562_ (.Y(_07631_),
    .A(net1078),
    .B(_07624_));
 sg13g2_a21oi_1 _26563_ (.A1(_07630_),
    .A2(_07631_),
    .Y(_02562_),
    .B1(net603));
 sg13g2_nand2_1 _26564_ (.Y(_07632_),
    .A(\cpu.spi.r_clk_count[1][4] ),
    .B(_07621_));
 sg13g2_nand2_1 _26565_ (.Y(_07633_),
    .A(_09840_),
    .B(_07624_));
 sg13g2_a21oi_1 _26566_ (.A1(_07632_),
    .A2(_07633_),
    .Y(_02563_),
    .B1(net603));
 sg13g2_nand2_1 _26567_ (.Y(_07634_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(_07621_));
 sg13g2_nand2_1 _26568_ (.Y(_07635_),
    .A(net1006),
    .B(_07624_));
 sg13g2_buf_1 _26569_ (.A(_09096_),
    .X(_07636_));
 sg13g2_a21oi_1 _26570_ (.A1(_07634_),
    .A2(_07635_),
    .Y(_02564_),
    .B1(net602));
 sg13g2_nand2_1 _26571_ (.Y(_07637_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_07621_));
 sg13g2_nand2_1 _26572_ (.Y(_07638_),
    .A(net929),
    .B(_07624_));
 sg13g2_a21oi_1 _26573_ (.A1(_07637_),
    .A2(_07638_),
    .Y(_02565_),
    .B1(net602));
 sg13g2_nand2_1 _26574_ (.Y(_07639_),
    .A(\cpu.spi.r_clk_count[1][7] ),
    .B(_07621_));
 sg13g2_nand2_1 _26575_ (.Y(_07640_),
    .A(_09856_),
    .B(_07624_));
 sg13g2_a21oi_1 _26576_ (.A1(_07639_),
    .A2(_07640_),
    .Y(_02566_),
    .B1(net602));
 sg13g2_nor2_1 _26577_ (.A(_04778_),
    .B(_09024_),
    .Y(_07641_));
 sg13g2_nand3_1 _26578_ (.B(_04783_),
    .C(_07641_),
    .A(_11611_),
    .Y(_07642_));
 sg13g2_buf_1 _26579_ (.A(_07642_),
    .X(_07643_));
 sg13g2_buf_1 _26580_ (.A(_07643_),
    .X(_07644_));
 sg13g2_or2_1 _26581_ (.X(_07645_),
    .B(_07644_),
    .A(_09810_));
 sg13g2_nand2_1 _26582_ (.Y(_07646_),
    .A(_04794_),
    .B(net82));
 sg13g2_a21oi_1 _26583_ (.A1(_07645_),
    .A2(_07646_),
    .Y(_02567_),
    .B1(net602));
 sg13g2_mux2_1 _26584_ (.A0(net1009),
    .A1(_05141_),
    .S(net82),
    .X(_07647_));
 sg13g2_and2_1 _26585_ (.A(net691),
    .B(_07647_),
    .X(_02568_));
 sg13g2_mux2_1 _26586_ (.A0(net1008),
    .A1(_05207_),
    .S(_07644_),
    .X(_07648_));
 sg13g2_and2_1 _26587_ (.A(net691),
    .B(_07648_),
    .X(_02569_));
 sg13g2_nand2_1 _26588_ (.Y(_07649_),
    .A(_05286_),
    .B(net82));
 sg13g2_o21ai_1 _26589_ (.B1(_07649_),
    .Y(_07650_),
    .A1(net849),
    .A2(net82));
 sg13g2_and2_1 _26590_ (.A(net691),
    .B(_07650_),
    .X(_02570_));
 sg13g2_mux2_1 _26591_ (.A0(_09839_),
    .A1(_05336_),
    .S(net82),
    .X(_07651_));
 sg13g2_and2_1 _26592_ (.A(net691),
    .B(_07651_),
    .X(_02571_));
 sg13g2_mux2_1 _26593_ (.A0(_09845_),
    .A1(_05431_),
    .S(net82),
    .X(_07652_));
 sg13g2_and2_1 _26594_ (.A(net691),
    .B(_07652_),
    .X(_02572_));
 sg13g2_nand2_1 _26595_ (.Y(_07653_),
    .A(_05463_),
    .B(_07643_));
 sg13g2_o21ai_1 _26596_ (.B1(_07653_),
    .Y(_07654_),
    .A1(_11808_),
    .A2(net82));
 sg13g2_and2_1 _26597_ (.A(net645),
    .B(_07654_),
    .X(_02573_));
 sg13g2_nand2_1 _26598_ (.Y(_07655_),
    .A(_04871_),
    .B(_07643_));
 sg13g2_o21ai_1 _26599_ (.B1(_07655_),
    .Y(_07656_),
    .A1(net848),
    .A2(net82));
 sg13g2_and2_1 _26600_ (.A(net645),
    .B(_07656_),
    .X(_02574_));
 sg13g2_o21ai_1 _26601_ (.B1(_09027_),
    .Y(_07657_),
    .A1(_09048_),
    .A2(_09018_));
 sg13g2_nor2_1 _26602_ (.A(\cpu.spi.r_state[3] ),
    .B(\cpu.spi.r_state[5] ),
    .Y(_07658_));
 sg13g2_and2_1 _26603_ (.A(_11572_),
    .B(_07658_),
    .X(_07659_));
 sg13g2_buf_1 _26604_ (.A(_07659_),
    .X(_07660_));
 sg13g2_nand2_1 _26605_ (.Y(_07661_),
    .A(_06765_),
    .B(_07660_));
 sg13g2_buf_1 _26606_ (.A(_07661_),
    .X(_07662_));
 sg13g2_nor2_1 _26607_ (.A(_09031_),
    .B(_07662_),
    .Y(_07663_));
 sg13g2_nor3_1 _26608_ (.A(_06765_),
    .B(net130),
    .C(_09047_),
    .Y(_07664_));
 sg13g2_nor3_1 _26609_ (.A(_09033_),
    .B(_07663_),
    .C(_07664_),
    .Y(_07665_));
 sg13g2_nand2_1 _26610_ (.Y(_07666_),
    .A(_07657_),
    .B(_07665_));
 sg13g2_buf_1 _26611_ (.A(_07666_),
    .X(_07667_));
 sg13g2_buf_1 _26612_ (.A(_07667_),
    .X(_07668_));
 sg13g2_buf_1 _26613_ (.A(_07662_),
    .X(_07669_));
 sg13g2_nand2b_1 _26614_ (.Y(_07670_),
    .B(net572),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _26615_ (.B1(_07670_),
    .Y(_07671_),
    .A1(net572),
    .A2(_04794_));
 sg13g2_mux2_1 _26616_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net571),
    .X(_07672_));
 sg13g2_nor2_1 _26617_ (.A(net643),
    .B(_07672_),
    .Y(_07673_));
 sg13g2_a21oi_1 _26618_ (.A1(net635),
    .A2(_07671_),
    .Y(_07674_),
    .B1(_07673_));
 sg13g2_buf_1 _26619_ (.A(_11583_),
    .X(_07675_));
 sg13g2_nor2_1 _26620_ (.A(net916),
    .B(_04794_),
    .Y(_07676_));
 sg13g2_a21oi_1 _26621_ (.A1(net916),
    .A2(_00314_),
    .Y(_07677_),
    .B1(_07676_));
 sg13g2_buf_1 _26622_ (.A(_11579_),
    .X(_07678_));
 sg13g2_mux2_1 _26623_ (.A0(_00314_),
    .A1(_00313_),
    .S(_11586_),
    .X(_07679_));
 sg13g2_nor2_1 _26624_ (.A(net915),
    .B(_07679_),
    .Y(_07680_));
 sg13g2_a21oi_1 _26625_ (.A1(net988),
    .A2(_07677_),
    .Y(_07681_),
    .B1(_07680_));
 sg13g2_nand2_1 _26626_ (.Y(_07682_),
    .A(net371),
    .B(_07681_));
 sg13g2_buf_1 _26627_ (.A(_07660_),
    .X(_07683_));
 sg13g2_nor2_1 _26628_ (.A(_08931_),
    .B(net601),
    .Y(_07684_));
 sg13g2_nand2b_1 _26629_ (.Y(_07685_),
    .B(net110),
    .A_N(_07681_));
 sg13g2_o21ai_1 _26630_ (.B1(_07685_),
    .Y(_07686_),
    .A1(_08931_),
    .A2(net110));
 sg13g2_a22oi_1 _26631_ (.Y(_07687_),
    .B1(_07686_),
    .B2(net1016),
    .A2(_07684_),
    .A1(_07682_));
 sg13g2_nand2_1 _26632_ (.Y(_07688_),
    .A(net479),
    .B(_07687_));
 sg13g2_o21ai_1 _26633_ (.B1(_07688_),
    .Y(_07689_),
    .A1(net479),
    .A2(_07674_));
 sg13g2_nor2_1 _26634_ (.A(_07668_),
    .B(_07689_),
    .Y(_07690_));
 sg13g2_a21oi_1 _26635_ (.A1(_08931_),
    .A2(_07668_),
    .Y(_07691_),
    .B1(_07690_));
 sg13g2_nor2_1 _26636_ (.A(net607),
    .B(_07691_),
    .Y(_02575_));
 sg13g2_mux2_1 _26637_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net644),
    .X(_07692_));
 sg13g2_nand2_1 _26638_ (.Y(_07693_),
    .A(net851),
    .B(_05141_));
 sg13g2_nand2_1 _26639_ (.Y(_07694_),
    .A(net644),
    .B(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_nand3_1 _26640_ (.B(_07693_),
    .C(_07694_),
    .A(_11611_),
    .Y(_07695_));
 sg13g2_o21ai_1 _26641_ (.B1(_07695_),
    .Y(_07696_),
    .A1(net725),
    .A2(_07692_));
 sg13g2_nand2b_1 _26642_ (.Y(_07697_),
    .B(_07696_),
    .A_N(_07662_));
 sg13g2_nand3_1 _26643_ (.B(_09027_),
    .C(_07697_),
    .A(_08931_),
    .Y(_07698_));
 sg13g2_nand2b_1 _26644_ (.Y(_07699_),
    .B(_07698_),
    .A_N(_07667_));
 sg13g2_nor2_1 _26645_ (.A(net853),
    .B(_05141_),
    .Y(_07700_));
 sg13g2_a21oi_1 _26646_ (.A1(net853),
    .A2(_00095_),
    .Y(_07701_),
    .B1(_07700_));
 sg13g2_mux2_1 _26647_ (.A0(_00095_),
    .A1(_00094_),
    .S(net853),
    .X(_07702_));
 sg13g2_nor2_1 _26648_ (.A(net988),
    .B(_07702_),
    .Y(_07703_));
 sg13g2_a21oi_1 _26649_ (.A1(net988),
    .A2(_07701_),
    .Y(_07704_),
    .B1(_07703_));
 sg13g2_nand2_1 _26650_ (.Y(_07705_),
    .A(net130),
    .B(_08933_));
 sg13g2_o21ai_1 _26651_ (.B1(_07705_),
    .Y(_07706_),
    .A1(net130),
    .A2(_07704_));
 sg13g2_nand2_1 _26652_ (.Y(_07707_),
    .A(_08931_),
    .B(_08932_));
 sg13g2_or2_1 _26653_ (.X(_07708_),
    .B(_08932_),
    .A(_08931_));
 sg13g2_a221oi_1 _26654_ (.B2(_07708_),
    .C1(net601),
    .B1(_07707_),
    .A1(net371),
    .Y(_07709_),
    .A2(_07704_));
 sg13g2_a221oi_1 _26655_ (.B2(net1016),
    .C1(_07709_),
    .B1(_07706_),
    .A1(_06765_),
    .Y(_07710_),
    .A2(net601));
 sg13g2_nor2_1 _26656_ (.A(_07667_),
    .B(_07710_),
    .Y(_07711_));
 sg13g2_a22oi_1 _26657_ (.Y(_07712_),
    .B1(_07711_),
    .B2(_07697_),
    .A2(_07699_),
    .A1(_08932_));
 sg13g2_nor2_1 _26658_ (.A(net607),
    .B(_07712_),
    .Y(_02576_));
 sg13g2_nand2b_1 _26659_ (.Y(_07713_),
    .B(_11617_),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _26660_ (.B1(_07713_),
    .Y(_07714_),
    .A1(net572),
    .A2(_05207_));
 sg13g2_mux2_1 _26661_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net571),
    .X(_07715_));
 sg13g2_nor2_1 _26662_ (.A(net725),
    .B(_07715_),
    .Y(_07716_));
 sg13g2_a21oi_1 _26663_ (.A1(net635),
    .A2(_07714_),
    .Y(_07717_),
    .B1(_07716_));
 sg13g2_nor2_1 _26664_ (.A(_07675_),
    .B(_05207_),
    .Y(_07718_));
 sg13g2_a21oi_1 _26665_ (.A1(net853),
    .A2(_00105_),
    .Y(_07719_),
    .B1(_07718_));
 sg13g2_mux2_1 _26666_ (.A0(_00105_),
    .A1(_00104_),
    .S(_07675_),
    .X(_07720_));
 sg13g2_nor2_1 _26667_ (.A(_07678_),
    .B(_07720_),
    .Y(_07721_));
 sg13g2_a21oi_1 _26668_ (.A1(net988),
    .A2(_07719_),
    .Y(_07722_),
    .B1(_07721_));
 sg13g2_nand2_1 _26669_ (.Y(_07723_),
    .A(\cpu.spi.r_count[2] ),
    .B(_07708_));
 sg13g2_a21o_1 _26670_ (.A2(_07723_),
    .A1(_08935_),
    .B1(net131),
    .X(_07724_));
 sg13g2_o21ai_1 _26671_ (.B1(_07724_),
    .Y(_07725_),
    .A1(net130),
    .A2(_07722_));
 sg13g2_a221oi_1 _26672_ (.B2(_08935_),
    .C1(_07683_),
    .B1(_07723_),
    .A1(net405),
    .Y(_07726_),
    .A2(_07722_));
 sg13g2_a21oi_1 _26673_ (.A1(net1084),
    .A2(_07725_),
    .Y(_07727_),
    .B1(_07726_));
 sg13g2_nand2_1 _26674_ (.Y(_07728_),
    .A(net479),
    .B(_07727_));
 sg13g2_o21ai_1 _26675_ (.B1(_07728_),
    .Y(_07729_),
    .A1(_07669_),
    .A2(_07717_));
 sg13g2_nor2_1 _26676_ (.A(net34),
    .B(_07729_),
    .Y(_07730_));
 sg13g2_a21oi_1 _26677_ (.A1(\cpu.spi.r_count[2] ),
    .A2(net34),
    .Y(_07731_),
    .B1(_07730_));
 sg13g2_nor2_1 _26678_ (.A(net607),
    .B(_07731_),
    .Y(_02577_));
 sg13g2_nand2b_1 _26679_ (.Y(_07732_),
    .B(net571),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _26680_ (.B1(_07732_),
    .Y(_07733_),
    .A1(net572),
    .A2(_05286_));
 sg13g2_mux2_1 _26681_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net571),
    .X(_07734_));
 sg13g2_nor2_1 _26682_ (.A(net725),
    .B(_07734_),
    .Y(_07735_));
 sg13g2_a21oi_1 _26683_ (.A1(net635),
    .A2(_07733_),
    .Y(_07736_),
    .B1(_07735_));
 sg13g2_xor2_1 _26684_ (.B(_08935_),
    .A(_08930_),
    .X(_07737_));
 sg13g2_nor2_1 _26685_ (.A(net601),
    .B(_07737_),
    .Y(_07738_));
 sg13g2_nor2_1 _26686_ (.A(net916),
    .B(_05286_),
    .Y(_07739_));
 sg13g2_a21oi_1 _26687_ (.A1(net916),
    .A2(_00115_),
    .Y(_07740_),
    .B1(_07739_));
 sg13g2_mux2_1 _26688_ (.A0(_00115_),
    .A1(_00114_),
    .S(net987),
    .X(_07741_));
 sg13g2_nor2_1 _26689_ (.A(net915),
    .B(_07741_),
    .Y(_07742_));
 sg13g2_a21oi_1 _26690_ (.A1(net988),
    .A2(_07740_),
    .Y(_07743_),
    .B1(_07742_));
 sg13g2_nand2_1 _26691_ (.Y(_07744_),
    .A(net405),
    .B(_07743_));
 sg13g2_nand2b_1 _26692_ (.Y(_07745_),
    .B(net110),
    .A_N(_07743_));
 sg13g2_o21ai_1 _26693_ (.B1(_07745_),
    .Y(_07746_),
    .A1(net110),
    .A2(_07737_));
 sg13g2_a22oi_1 _26694_ (.Y(_07747_),
    .B1(_07746_),
    .B2(net1016),
    .A2(_07744_),
    .A1(_07738_));
 sg13g2_nand2_1 _26695_ (.Y(_07748_),
    .A(_07662_),
    .B(_07747_));
 sg13g2_o21ai_1 _26696_ (.B1(_07748_),
    .Y(_07749_),
    .A1(net479),
    .A2(_07736_));
 sg13g2_nor2_1 _26697_ (.A(net34),
    .B(_07749_),
    .Y(_07750_));
 sg13g2_a21oi_1 _26698_ (.A1(_08930_),
    .A2(net34),
    .Y(_07751_),
    .B1(_07750_));
 sg13g2_nor2_1 _26699_ (.A(net607),
    .B(_07751_),
    .Y(_02578_));
 sg13g2_nand2b_1 _26700_ (.Y(_07752_),
    .B(net571),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _26701_ (.B1(_07752_),
    .Y(_07753_),
    .A1(net572),
    .A2(_05336_));
 sg13g2_mux2_1 _26702_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net571),
    .X(_07754_));
 sg13g2_nor2_1 _26703_ (.A(net725),
    .B(_07754_),
    .Y(_07755_));
 sg13g2_a21oi_1 _26704_ (.A1(net643),
    .A2(_07753_),
    .Y(_07756_),
    .B1(_07755_));
 sg13g2_nor2_1 _26705_ (.A(_08930_),
    .B(_08935_),
    .Y(_07757_));
 sg13g2_xnor2_1 _26706_ (.Y(_07758_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07757_));
 sg13g2_nor2_1 _26707_ (.A(net601),
    .B(_07758_),
    .Y(_07759_));
 sg13g2_nor2_1 _26708_ (.A(net987),
    .B(_05336_),
    .Y(_07760_));
 sg13g2_a21oi_1 _26709_ (.A1(net916),
    .A2(_00126_),
    .Y(_07761_),
    .B1(_07760_));
 sg13g2_mux2_1 _26710_ (.A0(_00126_),
    .A1(_00125_),
    .S(net987),
    .X(_07762_));
 sg13g2_nor2_1 _26711_ (.A(net915),
    .B(_07762_),
    .Y(_07763_));
 sg13g2_a21oi_1 _26712_ (.A1(net988),
    .A2(_07761_),
    .Y(_07764_),
    .B1(_07763_));
 sg13g2_nand2_1 _26713_ (.Y(_07765_),
    .A(net405),
    .B(_07764_));
 sg13g2_nand2b_1 _26714_ (.Y(_07766_),
    .B(net131),
    .A_N(_07764_));
 sg13g2_o21ai_1 _26715_ (.B1(_07766_),
    .Y(_07767_),
    .A1(net110),
    .A2(_07758_));
 sg13g2_a22oi_1 _26716_ (.Y(_07768_),
    .B1(_07767_),
    .B2(net1016),
    .A2(_07765_),
    .A1(_07759_));
 sg13g2_nand2_1 _26717_ (.Y(_07769_),
    .A(_07662_),
    .B(_07768_));
 sg13g2_o21ai_1 _26718_ (.B1(_07769_),
    .Y(_07770_),
    .A1(net479),
    .A2(_07756_));
 sg13g2_nor2_1 _26719_ (.A(net34),
    .B(_07770_),
    .Y(_07771_));
 sg13g2_a21oi_1 _26720_ (.A1(\cpu.spi.r_count[4] ),
    .A2(net34),
    .Y(_07772_),
    .B1(_07771_));
 sg13g2_nor2_1 _26721_ (.A(net689),
    .B(_07772_),
    .Y(_02579_));
 sg13g2_nand2b_1 _26722_ (.Y(_07773_),
    .B(net571),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _26723_ (.B1(_07773_),
    .Y(_07774_),
    .A1(net572),
    .A2(_05431_));
 sg13g2_mux2_1 _26724_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net644),
    .X(_07775_));
 sg13g2_nor2_1 _26725_ (.A(net725),
    .B(_07775_),
    .Y(_07776_));
 sg13g2_a21oi_1 _26726_ (.A1(net643),
    .A2(_07774_),
    .Y(_07777_),
    .B1(_07776_));
 sg13g2_nor2_1 _26727_ (.A(net987),
    .B(_05431_),
    .Y(_07778_));
 sg13g2_a21oi_1 _26728_ (.A1(net916),
    .A2(_00133_),
    .Y(_07779_),
    .B1(_07778_));
 sg13g2_mux2_1 _26729_ (.A0(_00133_),
    .A1(_00132_),
    .S(net987),
    .X(_07780_));
 sg13g2_nor2_1 _26730_ (.A(net915),
    .B(_07780_),
    .Y(_07781_));
 sg13g2_a21oi_1 _26731_ (.A1(net915),
    .A2(_07779_),
    .Y(_07782_),
    .B1(_07781_));
 sg13g2_nand2_1 _26732_ (.Y(_07783_),
    .A(net371),
    .B(_07782_));
 sg13g2_xnor2_1 _26733_ (.Y(_07784_),
    .A(\cpu.spi.r_count[5] ),
    .B(_08936_));
 sg13g2_nor2_1 _26734_ (.A(net601),
    .B(_07784_),
    .Y(_07785_));
 sg13g2_nand2b_1 _26735_ (.Y(_07786_),
    .B(net131),
    .A_N(_07782_));
 sg13g2_o21ai_1 _26736_ (.B1(_07786_),
    .Y(_07787_),
    .A1(net110),
    .A2(_07784_));
 sg13g2_a22oi_1 _26737_ (.Y(_07788_),
    .B1(_07787_),
    .B2(net1016),
    .A2(_07785_),
    .A1(_07783_));
 sg13g2_nand2_1 _26738_ (.Y(_07789_),
    .A(_07662_),
    .B(_07788_));
 sg13g2_o21ai_1 _26739_ (.B1(_07789_),
    .Y(_07790_),
    .A1(net479),
    .A2(_07777_));
 sg13g2_nor2_1 _26740_ (.A(_07667_),
    .B(_07790_),
    .Y(_07791_));
 sg13g2_a21oi_1 _26741_ (.A1(\cpu.spi.r_count[5] ),
    .A2(net34),
    .Y(_07792_),
    .B1(_07791_));
 sg13g2_nor2_1 _26742_ (.A(net689),
    .B(_07792_),
    .Y(_02580_));
 sg13g2_nand2b_1 _26743_ (.Y(_07793_),
    .B(net571),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _26744_ (.B1(_07793_),
    .Y(_07794_),
    .A1(net572),
    .A2(_05463_));
 sg13g2_mux2_1 _26745_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(_11604_),
    .X(_07795_));
 sg13g2_nor2_1 _26746_ (.A(net725),
    .B(_07795_),
    .Y(_07796_));
 sg13g2_a21oi_1 _26747_ (.A1(net643),
    .A2(_07794_),
    .Y(_07797_),
    .B1(_07796_));
 sg13g2_nor2_1 _26748_ (.A(net987),
    .B(_05463_),
    .Y(_07798_));
 sg13g2_a21oi_1 _26749_ (.A1(net916),
    .A2(_00145_),
    .Y(_07799_),
    .B1(_07798_));
 sg13g2_mux2_1 _26750_ (.A0(_00145_),
    .A1(_00144_),
    .S(net987),
    .X(_07800_));
 sg13g2_nor2_1 _26751_ (.A(net915),
    .B(_07800_),
    .Y(_07801_));
 sg13g2_a21oi_1 _26752_ (.A1(net915),
    .A2(_07799_),
    .Y(_07802_),
    .B1(_07801_));
 sg13g2_nand2_1 _26753_ (.Y(_07803_),
    .A(net405),
    .B(_07802_));
 sg13g2_xnor2_1 _26754_ (.Y(_07804_),
    .A(\cpu.spi.r_count[6] ),
    .B(_08937_));
 sg13g2_nor2_1 _26755_ (.A(net601),
    .B(_07804_),
    .Y(_07805_));
 sg13g2_nand2b_1 _26756_ (.Y(_07806_),
    .B(net131),
    .A_N(_07802_));
 sg13g2_o21ai_1 _26757_ (.B1(_07806_),
    .Y(_07807_),
    .A1(net110),
    .A2(_07804_));
 sg13g2_a22oi_1 _26758_ (.Y(_07808_),
    .B1(_07807_),
    .B2(net1016),
    .A2(_07805_),
    .A1(_07803_));
 sg13g2_nand2_1 _26759_ (.Y(_07809_),
    .A(_07662_),
    .B(_07808_));
 sg13g2_o21ai_1 _26760_ (.B1(_07809_),
    .Y(_07810_),
    .A1(net479),
    .A2(_07797_));
 sg13g2_nor2_1 _26761_ (.A(_07667_),
    .B(_07810_),
    .Y(_07811_));
 sg13g2_a21oi_1 _26762_ (.A1(\cpu.spi.r_count[6] ),
    .A2(net34),
    .Y(_07812_),
    .B1(_07811_));
 sg13g2_nor2_1 _26763_ (.A(net689),
    .B(_07812_),
    .Y(_02581_));
 sg13g2_mux2_1 _26764_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(_11614_),
    .X(_07813_));
 sg13g2_nand2_1 _26765_ (.Y(_07814_),
    .A(net851),
    .B(_04871_));
 sg13g2_nand2_1 _26766_ (.Y(_07815_),
    .A(_11614_),
    .B(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_nand3_1 _26767_ (.B(_07814_),
    .C(_07815_),
    .A(net643),
    .Y(_07816_));
 sg13g2_o21ai_1 _26768_ (.B1(_07816_),
    .Y(_07817_),
    .A1(net635),
    .A2(_07813_));
 sg13g2_nand2b_1 _26769_ (.Y(_07818_),
    .B(_08929_),
    .A_N(_08938_));
 sg13g2_a21oi_1 _26770_ (.A1(_09044_),
    .A2(net601),
    .Y(_07819_),
    .B1(_07818_));
 sg13g2_nor2_1 _26771_ (.A(_11586_),
    .B(_04871_),
    .Y(_07820_));
 sg13g2_a21oi_1 _26772_ (.A1(net916),
    .A2(_00157_),
    .Y(_07821_),
    .B1(_07820_));
 sg13g2_mux2_1 _26773_ (.A0(_00157_),
    .A1(_00156_),
    .S(_11583_),
    .X(_07822_));
 sg13g2_nor2_1 _26774_ (.A(_07678_),
    .B(_07822_),
    .Y(_07823_));
 sg13g2_a21oi_1 _26775_ (.A1(net915),
    .A2(_07821_),
    .Y(_07824_),
    .B1(_07823_));
 sg13g2_nor2_1 _26776_ (.A(_07683_),
    .B(_07824_),
    .Y(_07825_));
 sg13g2_o21ai_1 _26777_ (.B1(net405),
    .Y(_07826_),
    .A1(_09027_),
    .A2(_07825_));
 sg13g2_o21ai_1 _26778_ (.B1(_07826_),
    .Y(_07827_),
    .A1(_06805_),
    .A2(_07824_));
 sg13g2_o21ai_1 _26779_ (.B1(net479),
    .Y(_07828_),
    .A1(_07819_),
    .A2(_07827_));
 sg13g2_o21ai_1 _26780_ (.B1(_07828_),
    .Y(_07829_),
    .A1(_07669_),
    .A2(_07817_));
 sg13g2_mux2_1 _26781_ (.A0(_07829_),
    .A1(_08929_),
    .S(_07667_),
    .X(_07830_));
 sg13g2_and2_1 _26782_ (.A(_11550_),
    .B(_07830_),
    .X(_02582_));
 sg13g2_inv_1 _26783_ (.Y(_07831_),
    .A(\cpu.spi.r_state[3] ));
 sg13g2_nand2_1 _26784_ (.Y(_07832_),
    .A(_07831_),
    .B(_09020_));
 sg13g2_nor3_1 _26785_ (.A(_09088_),
    .B(net405),
    .C(_07832_),
    .Y(_07833_));
 sg13g2_a21oi_1 _26786_ (.A1(net988),
    .A2(_11587_),
    .Y(_07834_),
    .B1(_08940_));
 sg13g2_nor3_1 _26787_ (.A(_00278_),
    .B(_07833_),
    .C(_07834_),
    .Y(_07835_));
 sg13g2_inv_1 _26788_ (.Y(_07836_),
    .A(_00278_));
 sg13g2_a21oi_1 _26789_ (.A1(_09049_),
    .A2(_07832_),
    .Y(_07837_),
    .B1(_07836_));
 sg13g2_a21oi_1 _26790_ (.A1(_09043_),
    .A2(_09018_),
    .Y(_07838_),
    .B1(_06765_));
 sg13g2_nor3_1 _26791_ (.A(_07835_),
    .B(_07837_),
    .C(_07838_),
    .Y(_07839_));
 sg13g2_a21oi_1 _26792_ (.A1(_07832_),
    .A2(_07839_),
    .Y(_07840_),
    .B1(net747));
 sg13g2_nand2_1 _26793_ (.Y(_07841_),
    .A(_11594_),
    .B(_07839_));
 sg13g2_buf_1 _26794_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_07842_));
 sg13g2_o21ai_1 _26795_ (.B1(net1046),
    .Y(_07843_),
    .A1(_11587_),
    .A2(_07841_));
 sg13g2_nand2_1 _26796_ (.Y(_02583_),
    .A(_07840_),
    .B(_07843_));
 sg13g2_buf_1 _26797_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_07844_));
 sg13g2_o21ai_1 _26798_ (.B1(net1045),
    .Y(_07845_),
    .A1(_11584_),
    .A2(_07841_));
 sg13g2_nand2_1 _26799_ (.Y(_02584_),
    .A(_07840_),
    .B(_07845_));
 sg13g2_buf_1 _26800_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_07846_));
 sg13g2_nand2_1 _26801_ (.Y(_07847_),
    .A(_11598_),
    .B(_07839_));
 sg13g2_nand2_1 _26802_ (.Y(_07848_),
    .A(net1044),
    .B(_07847_));
 sg13g2_nand2_1 _26803_ (.Y(_02585_),
    .A(_07840_),
    .B(_07848_));
 sg13g2_nand2_1 _26804_ (.Y(_07849_),
    .A(_09048_),
    .B(_09081_));
 sg13g2_a21o_1 _26805_ (.A2(_07849_),
    .A1(net1017),
    .B1(_07583_),
    .X(_07850_));
 sg13g2_buf_1 _26806_ (.A(_07850_),
    .X(_07851_));
 sg13g2_nor3_1 _26807_ (.A(_06765_),
    .B(net131),
    .C(_09018_),
    .Y(_07852_));
 sg13g2_or2_1 _26808_ (.X(_07853_),
    .B(_07852_),
    .A(_09033_));
 sg13g2_buf_1 _26809_ (.A(_07853_),
    .X(_07854_));
 sg13g2_or3_1 _26810_ (.A(_09089_),
    .B(_07851_),
    .C(_07854_),
    .X(_07855_));
 sg13g2_o21ai_1 _26811_ (.B1(_08998_),
    .Y(_07856_),
    .A1(_07851_),
    .A2(_07854_));
 sg13g2_a21oi_1 _26812_ (.A1(_07855_),
    .A2(_07856_),
    .Y(_02594_),
    .B1(net602));
 sg13g2_nand3_1 _26813_ (.B(_04695_),
    .C(_07597_),
    .A(_05564_),
    .Y(_07857_));
 sg13g2_nand2_1 _26814_ (.Y(_07858_),
    .A(_04695_),
    .B(_07597_));
 sg13g2_nand2_1 _26815_ (.Y(_07859_),
    .A(\cpu.spi.r_mode[0][0] ),
    .B(_07858_));
 sg13g2_a21oi_1 _26816_ (.A1(_07857_),
    .A2(_07859_),
    .Y(_02595_),
    .B1(net602));
 sg13g2_nand3_1 _26817_ (.B(_04695_),
    .C(_07597_),
    .A(_09819_),
    .Y(_07860_));
 sg13g2_nand2_1 _26818_ (.Y(_07861_),
    .A(_11595_),
    .B(_07858_));
 sg13g2_a21oi_1 _26819_ (.A1(_07860_),
    .A2(_07861_),
    .Y(_02596_),
    .B1(_07636_));
 sg13g2_nand3_1 _26820_ (.B(_08966_),
    .C(_07597_),
    .A(net573),
    .Y(_07862_));
 sg13g2_buf_1 _26821_ (.A(_07862_),
    .X(_07863_));
 sg13g2_nand2_1 _26822_ (.Y(_07864_),
    .A(\cpu.spi.r_mode[1][0] ),
    .B(_07863_));
 sg13g2_o21ai_1 _26823_ (.B1(_07864_),
    .Y(_07865_),
    .A1(net872),
    .A2(_07863_));
 sg13g2_and2_1 _26824_ (.A(net645),
    .B(_07865_),
    .X(_02597_));
 sg13g2_mux2_1 _26825_ (.A0(net1009),
    .A1(_11596_),
    .S(_07863_),
    .X(_07866_));
 sg13g2_and2_1 _26826_ (.A(net645),
    .B(_07866_),
    .X(_02598_));
 sg13g2_nand3_1 _26827_ (.B(_04695_),
    .C(_07641_),
    .A(_11612_),
    .Y(_07867_));
 sg13g2_buf_1 _26828_ (.A(_07867_),
    .X(_07868_));
 sg13g2_or2_1 _26829_ (.X(_07869_),
    .B(_07868_),
    .A(_09809_));
 sg13g2_nand2_1 _26830_ (.Y(_07870_),
    .A(\cpu.spi.r_mode[2][0] ),
    .B(_07868_));
 sg13g2_a21oi_1 _26831_ (.A1(_07869_),
    .A2(_07870_),
    .Y(_02599_),
    .B1(net602));
 sg13g2_mux2_1 _26832_ (.A0(net1009),
    .A1(_11599_),
    .S(_07868_),
    .X(_07871_));
 sg13g2_and2_1 _26833_ (.A(net645),
    .B(_07871_),
    .X(_02600_));
 sg13g2_a221oi_1 _26834_ (.B2(_07831_),
    .C1(_07854_),
    .B1(_07583_),
    .A1(net1017),
    .Y(_07872_),
    .A2(_07849_));
 sg13g2_nand3_1 _26835_ (.B(_09044_),
    .C(_07872_),
    .A(_07831_),
    .Y(_07873_));
 sg13g2_o21ai_1 _26836_ (.B1(_07873_),
    .Y(_07874_),
    .A1(\cpu.spi.r_ready ),
    .A2(_09049_));
 sg13g2_nand2_1 _26837_ (.Y(_07875_),
    .A(_09089_),
    .B(_07874_));
 sg13g2_o21ai_1 _26838_ (.B1(_07875_),
    .Y(_07876_),
    .A1(\cpu.spi.r_ready ),
    .A2(_07872_));
 sg13g2_nand2_1 _26839_ (.Y(_02609_),
    .A(net623),
    .B(_07876_));
 sg13g2_nor3_1 _26840_ (.A(_08966_),
    .B(net130),
    .C(_07851_),
    .Y(_07877_));
 sg13g2_a21o_1 _26841_ (.A2(net130),
    .A1(_09066_),
    .B1(_07877_),
    .X(_07878_));
 sg13g2_a22oi_1 _26842_ (.Y(_07879_),
    .B1(_07878_),
    .B2(_09085_),
    .A2(_07851_),
    .A1(_09066_));
 sg13g2_nor2_1 _26843_ (.A(_09100_),
    .B(_07879_),
    .Y(_02610_));
 sg13g2_nand3_1 _26844_ (.B(_04695_),
    .C(_07597_),
    .A(_09889_),
    .Y(_07880_));
 sg13g2_nand2_1 _26845_ (.Y(_07881_),
    .A(\cpu.spi.r_src[0] ),
    .B(_07858_));
 sg13g2_a21oi_1 _26846_ (.A1(_07880_),
    .A2(_07881_),
    .Y(_02613_),
    .B1(_07636_));
 sg13g2_mux2_1 _26847_ (.A0(net1008),
    .A1(\cpu.spi.r_src[1] ),
    .S(_07863_),
    .X(_07882_));
 sg13g2_and2_1 _26848_ (.A(net645),
    .B(_07882_),
    .X(_02614_));
 sg13g2_mux2_1 _26849_ (.A0(net1008),
    .A1(_11582_),
    .S(_07868_),
    .X(_07883_));
 sg13g2_and2_1 _26850_ (.A(net645),
    .B(_07883_),
    .X(_02615_));
 sg13g2_buf_1 _26851_ (.A(_06868_),
    .X(_07884_));
 sg13g2_nor2_1 _26852_ (.A(_04697_),
    .B(net114),
    .Y(_07885_));
 sg13g2_buf_2 _26853_ (.A(_07885_),
    .X(_07886_));
 sg13g2_nand2_1 _26854_ (.Y(_07887_),
    .A(net821),
    .B(_07886_));
 sg13g2_inv_1 _26855_ (.Y(_07888_),
    .A(net114));
 sg13g2_nand2_1 _26856_ (.Y(_07889_),
    .A(net429),
    .B(_07888_));
 sg13g2_buf_2 _26857_ (.A(_07889_),
    .X(_07890_));
 sg13g2_nand2_1 _26858_ (.Y(_07891_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_07890_));
 sg13g2_nand3_1 _26859_ (.B(_07887_),
    .C(_07891_),
    .A(net622),
    .Y(_02632_));
 sg13g2_nor2_1 _26860_ (.A(net428),
    .B(_07884_),
    .Y(_07892_));
 sg13g2_nand2_1 _26861_ (.Y(_07893_),
    .A(net869),
    .B(_07892_));
 sg13g2_o21ai_1 _26862_ (.B1(_09717_),
    .Y(_07894_),
    .A1(net428),
    .A2(_07884_));
 sg13g2_a21oi_1 _26863_ (.A1(_07893_),
    .A2(_07894_),
    .Y(_02633_),
    .B1(net602));
 sg13g2_nand2_1 _26864_ (.Y(_07895_),
    .A(net928),
    .B(_07892_));
 sg13g2_o21ai_1 _26865_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_07896_),
    .A1(net428),
    .A2(net114));
 sg13g2_buf_1 _26866_ (.A(_09096_),
    .X(_07897_));
 sg13g2_a21oi_1 _26867_ (.A1(_07895_),
    .A2(_07896_),
    .Y(_02634_),
    .B1(net600));
 sg13g2_nand2_1 _26868_ (.Y(_07898_),
    .A(net1004),
    .B(_07886_));
 sg13g2_nand2_1 _26869_ (.Y(_07899_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26870_ (.A1(_07898_),
    .A2(_07899_),
    .Y(_02635_),
    .B1(net600));
 sg13g2_nand2_1 _26871_ (.Y(_07900_),
    .A(net869),
    .B(_07886_));
 sg13g2_nand2_1 _26872_ (.Y(_07901_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26873_ (.A1(_07900_),
    .A2(_07901_),
    .Y(_02636_),
    .B1(net600));
 sg13g2_nand2_1 _26874_ (.Y(_07902_),
    .A(net1078),
    .B(_07886_));
 sg13g2_nand2_1 _26875_ (.Y(_07903_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26876_ (.A1(_07902_),
    .A2(_07903_),
    .Y(_02637_),
    .B1(net600));
 sg13g2_nand2_1 _26877_ (.Y(_07904_),
    .A(net1007),
    .B(_07886_));
 sg13g2_nand2_1 _26878_ (.Y(_07905_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26879_ (.A1(_07904_),
    .A2(_07905_),
    .Y(_02638_),
    .B1(net600));
 sg13g2_nand2_1 _26880_ (.Y(_07906_),
    .A(_09846_),
    .B(_07886_));
 sg13g2_nand2_1 _26881_ (.Y(_07907_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26882_ (.A1(_07906_),
    .A2(_07907_),
    .Y(_02639_),
    .B1(net600));
 sg13g2_nand2_1 _26883_ (.Y(_07908_),
    .A(net929),
    .B(_07886_));
 sg13g2_nand2_1 _26884_ (.Y(_07909_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26885_ (.A1(_07908_),
    .A2(_07909_),
    .Y(_02640_),
    .B1(_07897_));
 sg13g2_nand2_1 _26886_ (.Y(_07910_),
    .A(_09856_),
    .B(_07886_));
 sg13g2_nand2_1 _26887_ (.Y(_07911_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_07890_));
 sg13g2_a21oi_1 _26888_ (.A1(_07910_),
    .A2(_07911_),
    .Y(_02641_),
    .B1(net600));
 sg13g2_nand2_1 _26889_ (.Y(_07912_),
    .A(net942),
    .B(_07892_));
 sg13g2_o21ai_1 _26890_ (.B1(\cpu.uart.r_div_value[8] ),
    .Y(_07913_),
    .A1(net428),
    .A2(net114));
 sg13g2_a21oi_1 _26891_ (.A1(_07912_),
    .A2(_07913_),
    .Y(_02642_),
    .B1(_07897_));
 sg13g2_nand2_1 _26892_ (.Y(_07914_),
    .A(net1004),
    .B(_07892_));
 sg13g2_o21ai_1 _26893_ (.B1(\cpu.uart.r_div_value[9] ),
    .Y(_07915_),
    .A1(net428),
    .A2(net114));
 sg13g2_a21oi_1 _26894_ (.A1(_07914_),
    .A2(_07915_),
    .Y(_02643_),
    .B1(net600));
 sg13g2_nand3_1 _26895_ (.B(net431),
    .C(_07888_),
    .A(_09818_),
    .Y(_07916_));
 sg13g2_nand3_1 _26896_ (.B(_08590_),
    .C(_06866_),
    .A(net635),
    .Y(_07917_));
 sg13g2_or4_1 _26897_ (.A(net1022),
    .B(_09012_),
    .C(net627),
    .D(_07917_),
    .X(_07918_));
 sg13g2_nand4_1 _26898_ (.B(net761),
    .C(_07916_),
    .A(_09002_),
    .Y(_07919_),
    .D(_07918_));
 sg13g2_nand2b_1 _26899_ (.Y(_02667_),
    .B(_07919_),
    .A_N(net163));
 sg13g2_nor2_1 _26900_ (.A(_05420_),
    .B(net114),
    .Y(_07920_));
 sg13g2_nand2_1 _26901_ (.Y(_07921_),
    .A(net1004),
    .B(_07920_));
 sg13g2_o21ai_1 _26902_ (.B1(\cpu.uart.r_r_invert ),
    .Y(_07922_),
    .A1(_05420_),
    .A2(net114));
 sg13g2_a21oi_1 _26903_ (.A1(_07921_),
    .A2(_07922_),
    .Y(_02668_),
    .B1(net690));
 sg13g2_a21oi_1 _26904_ (.A1(_06850_),
    .A2(net337),
    .Y(_07923_),
    .B1(net1051));
 sg13g2_a21oi_1 _26905_ (.A1(_06851_),
    .A2(net337),
    .Y(_07924_),
    .B1(_06925_));
 sg13g2_a221oi_1 _26906_ (.B2(_07923_),
    .C1(_07924_),
    .B1(_06849_),
    .A1(net919),
    .Y(_07925_),
    .A2(net1051));
 sg13g2_a21oi_1 _26907_ (.A1(_06842_),
    .A2(_07925_),
    .Y(_07926_),
    .B1(_06922_));
 sg13g2_buf_2 _26908_ (.A(_07926_),
    .X(_07927_));
 sg13g2_o21ai_1 _26909_ (.B1(_07927_),
    .Y(_07928_),
    .A1(net919),
    .A2(_06925_));
 sg13g2_xnor2_1 _26910_ (.Y(_07929_),
    .A(_06851_),
    .B(_07928_));
 sg13g2_nor2_1 _26911_ (.A(net689),
    .B(_07929_),
    .Y(_02671_));
 sg13g2_o21ai_1 _26912_ (.B1(_07927_),
    .Y(_07930_),
    .A1(_06850_),
    .A2(net920));
 sg13g2_nand2_1 _26913_ (.Y(_07931_),
    .A(_06846_),
    .B(_07930_));
 sg13g2_nand2b_1 _26914_ (.Y(_07932_),
    .B(_06848_),
    .A_N(net920));
 sg13g2_o21ai_1 _26915_ (.B1(_07932_),
    .Y(_07933_),
    .A1(net919),
    .A2(_06924_));
 sg13g2_nand3_1 _26916_ (.B(_07927_),
    .C(_07933_),
    .A(_06923_),
    .Y(_07934_));
 sg13g2_a21oi_1 _26917_ (.A1(_07931_),
    .A2(_07934_),
    .Y(_02672_),
    .B1(net690));
 sg13g2_nand2_1 _26918_ (.Y(_07935_),
    .A(_06850_),
    .B(net1050));
 sg13g2_nor3_1 _26919_ (.A(net919),
    .B(net920),
    .C(_07935_),
    .Y(_07936_));
 sg13g2_o21ai_1 _26920_ (.B1(_07927_),
    .Y(_07937_),
    .A1(_06845_),
    .A2(_06933_));
 sg13g2_a22oi_1 _26921_ (.Y(_07938_),
    .B1(_07937_),
    .B2(net919),
    .A2(_07936_),
    .A1(_07927_));
 sg13g2_nor2_1 _26922_ (.A(net689),
    .B(_07938_),
    .Y(_02673_));
 sg13g2_a21oi_1 _26923_ (.A1(_06933_),
    .A2(_07927_),
    .Y(_07939_),
    .B1(_06845_));
 sg13g2_nor2b_1 _26924_ (.A(net919),
    .B_N(net1050),
    .Y(_07940_));
 sg13g2_a21oi_1 _26925_ (.A1(_07927_),
    .A2(_07940_),
    .Y(_07941_),
    .B1(_09103_));
 sg13g2_nor2b_1 _26926_ (.A(_07939_),
    .B_N(_07941_),
    .Y(_02674_));
 sg13g2_nor2b_1 _26927_ (.A(net917),
    .B_N(_06941_),
    .Y(_07942_));
 sg13g2_o21ai_1 _26928_ (.B1(_07942_),
    .Y(_07943_),
    .A1(_09001_),
    .A2(_06880_));
 sg13g2_o21ai_1 _26929_ (.B1(net557),
    .Y(_07944_),
    .A1(_00223_),
    .A2(net558));
 sg13g2_nor2b_1 _26930_ (.A(_06968_),
    .B_N(_07944_),
    .Y(_07945_));
 sg13g2_a21o_1 _26931_ (.A2(net431),
    .A1(net942),
    .B1(net382),
    .X(_07946_));
 sg13g2_a22oi_1 _26932_ (.Y(_07947_),
    .B1(_07946_),
    .B2(_06941_),
    .A2(_07945_),
    .A1(_09454_));
 sg13g2_o21ai_1 _26933_ (.B1(_09001_),
    .Y(_07948_),
    .A1(net114),
    .A2(_07947_));
 sg13g2_a21oi_1 _26934_ (.A1(_07943_),
    .A2(_07948_),
    .Y(_02676_),
    .B1(net690));
 sg13g2_mux2_1 _26935_ (.A0(\cpu.uart.r_x_invert ),
    .A1(net942),
    .S(_07920_),
    .X(_07949_));
 sg13g2_and2_1 _26936_ (.A(net645),
    .B(_07949_),
    .X(_02677_));
 sg13g2_o21ai_1 _26937_ (.B1(_06961_),
    .Y(_07950_),
    .A1(_06870_),
    .A2(_06968_));
 sg13g2_nor2_1 _26938_ (.A(_06885_),
    .B(_06945_),
    .Y(_07951_));
 sg13g2_nor3_1 _26939_ (.A(net918),
    .B(_06870_),
    .C(_06873_),
    .Y(_07952_));
 sg13g2_o21ai_1 _26940_ (.B1(_06882_),
    .Y(_07953_),
    .A1(_07951_),
    .A2(_07952_));
 sg13g2_nor2b_1 _26941_ (.A(_07950_),
    .B_N(_07953_),
    .Y(_07954_));
 sg13g2_buf_2 _26942_ (.A(_07954_),
    .X(_07955_));
 sg13g2_nand4_1 _26943_ (.B(_06870_),
    .C(_06880_),
    .A(_06864_),
    .Y(_07956_),
    .D(_06941_));
 sg13g2_nand4_1 _26944_ (.B(_06955_),
    .C(_07955_),
    .A(net917),
    .Y(_07957_),
    .D(_07956_));
 sg13g2_o21ai_1 _26945_ (.B1(_07957_),
    .Y(_07958_),
    .A1(net917),
    .A2(_07955_));
 sg13g2_nor2_1 _26946_ (.A(net689),
    .B(_07958_),
    .Y(_02680_));
 sg13g2_o21ai_1 _26947_ (.B1(_07955_),
    .Y(_07959_),
    .A1(net917),
    .A2(_06971_));
 sg13g2_nand2_1 _26948_ (.Y(_07960_),
    .A(_06871_),
    .B(_07959_));
 sg13g2_nand4_1 _26949_ (.B(net917),
    .C(_06955_),
    .A(_06881_),
    .Y(_07961_),
    .D(_07955_));
 sg13g2_a21oi_1 _26950_ (.A1(_07960_),
    .A2(_07961_),
    .Y(_02681_),
    .B1(net690));
 sg13g2_inv_1 _26951_ (.Y(_07962_),
    .A(_06873_));
 sg13g2_nand3_1 _26952_ (.B(_07962_),
    .C(_07955_),
    .A(_06885_),
    .Y(_07963_));
 sg13g2_nand2_1 _26953_ (.Y(_07964_),
    .A(net918),
    .B(_06873_));
 sg13g2_a21oi_1 _26954_ (.A1(_07963_),
    .A2(_07964_),
    .Y(_07965_),
    .B1(net1049));
 sg13g2_nor2_1 _26955_ (.A(_06880_),
    .B(_06954_),
    .Y(_07966_));
 sg13g2_nor2_1 _26956_ (.A(_06885_),
    .B(_07955_),
    .Y(_07967_));
 sg13g2_nor3_1 _26957_ (.A(_07965_),
    .B(_07966_),
    .C(_07967_),
    .Y(_07968_));
 sg13g2_nor2_1 _26958_ (.A(net689),
    .B(_07968_),
    .Y(_02682_));
 sg13g2_o21ai_1 _26959_ (.B1(_07955_),
    .Y(_07969_),
    .A1(net918),
    .A2(_07962_));
 sg13g2_a21o_1 _26960_ (.A2(_06943_),
    .A1(_07962_),
    .B1(_07966_),
    .X(_07970_));
 sg13g2_a22oi_1 _26961_ (.Y(_07971_),
    .B1(_07970_),
    .B2(_07955_),
    .A2(_07969_),
    .A1(net1049));
 sg13g2_nor2_1 _26962_ (.A(net689),
    .B(_07971_),
    .Y(_02683_));
 sg13g2_nand2b_1 _26963_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07125_),
    .A_N(_07121_));
 sg13g2_nor4_1 _26964_ (.A(_09669_),
    .B(_09577_),
    .C(_06630_),
    .D(_07551_),
    .Y(_07972_));
 sg13g2_nor2b_1 _26965_ (.A(_09627_),
    .B_N(_07972_),
    .Y(_07973_));
 sg13g2_a22oi_1 _26966_ (.Y(_07974_),
    .B1(net128),
    .B2(_07973_),
    .A2(net584),
    .A1(_09593_));
 sg13g2_inv_1 _26967_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_07974_));
 sg13g2_nor2_1 _26968_ (.A(_09598_),
    .B(net584),
    .Y(_07975_));
 sg13g2_a22oi_1 _26969_ (.Y(_07976_),
    .B1(_07972_),
    .B2(_07975_),
    .A2(net584),
    .A1(_09588_));
 sg13g2_nor2_1 _26970_ (.A(net779),
    .B(_07976_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _26971_ (.A(_00189_),
    .B(_07976_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _26972_ (.S0(_04725_),
    .A0(_08980_),
    .A1(_08973_),
    .A2(_08984_),
    .A3(_08988_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_07977_));
 sg13g2_mux4_1 _26973_ (.S0(_04725_),
    .A0(_08974_),
    .A1(_08981_),
    .A2(_08969_),
    .A3(_08976_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_07978_));
 sg13g2_mux2_1 _26974_ (.A0(_07977_),
    .A1(_07978_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _26975_ (.S0(_04710_),
    .A0(_11630_),
    .A1(net1069),
    .A2(net1046),
    .A3(net1045),
    .S1(_05151_),
    .X(_07979_));
 sg13g2_mux4_1 _26976_ (.S0(_04710_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1048),
    .A2(_11648_),
    .A3(_11632_),
    .S1(_05151_),
    .X(_07980_));
 sg13g2_nor2b_1 _26977_ (.A(_05217_),
    .B_N(_07980_),
    .Y(_07981_));
 sg13g2_a21oi_1 _26978_ (.A1(_05217_),
    .A2(_07979_),
    .Y(_07982_),
    .B1(_07981_));
 sg13g2_nand2b_1 _26979_ (.Y(_07983_),
    .B(net1044),
    .A_N(_04710_));
 sg13g2_nand3_1 _26980_ (.B(_05151_),
    .C(net1047),
    .A(_04710_),
    .Y(_07984_));
 sg13g2_o21ai_1 _26981_ (.B1(_07984_),
    .Y(_07985_),
    .A1(_05151_),
    .A2(_07983_));
 sg13g2_nand3_1 _26982_ (.B(_00187_),
    .C(_07985_),
    .A(_05279_),
    .Y(_07986_));
 sg13g2_o21ai_1 _26983_ (.B1(_07986_),
    .Y(net15),
    .A1(_05279_),
    .A2(_07982_));
 sg13g2_mux4_1 _26984_ (.S0(_05368_),
    .A0(net1068),
    .A1(net1069),
    .A2(net1046),
    .A3(net1045),
    .S1(_05425_),
    .X(_07987_));
 sg13g2_mux4_1 _26985_ (.S0(_05368_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_05425_),
    .X(_07988_));
 sg13g2_nor2b_1 _26986_ (.A(_05484_),
    .B_N(_07988_),
    .Y(_07989_));
 sg13g2_a21oi_1 _26987_ (.A1(_05484_),
    .A2(_07987_),
    .Y(_07990_),
    .B1(_07989_));
 sg13g2_nand2b_1 _26988_ (.Y(_07991_),
    .B(net1044),
    .A_N(_05368_));
 sg13g2_nand3_1 _26989_ (.B(_05425_),
    .C(_07548_),
    .A(_05368_),
    .Y(_07992_));
 sg13g2_o21ai_1 _26990_ (.B1(_07992_),
    .Y(_07993_),
    .A1(_05425_),
    .A2(_07991_));
 sg13g2_nand3_1 _26991_ (.B(_00186_),
    .C(_07993_),
    .A(_04849_),
    .Y(_07994_));
 sg13g2_o21ai_1 _26992_ (.B1(_07994_),
    .Y(net16),
    .A1(_04849_),
    .A2(_07990_));
 sg13g2_mux4_1 _26993_ (.S0(_04711_),
    .A0(net1068),
    .A1(net1069),
    .A2(net1046),
    .A3(net1045),
    .S1(_06121_),
    .X(_07995_));
 sg13g2_mux4_1 _26994_ (.S0(_04711_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_06121_),
    .X(_07996_));
 sg13g2_nor2b_1 _26995_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_07996_),
    .Y(_07997_));
 sg13g2_a21oi_1 _26996_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_07995_),
    .Y(_07998_),
    .B1(_07997_));
 sg13g2_nand2b_1 _26997_ (.Y(_07999_),
    .B(_07846_),
    .A_N(_04711_));
 sg13g2_nand3_1 _26998_ (.B(net1047),
    .C(_06121_),
    .A(_04711_),
    .Y(_08000_));
 sg13g2_o21ai_1 _26999_ (.B1(_08000_),
    .Y(_08001_),
    .A1(_06121_),
    .A2(_07999_));
 sg13g2_nand3_1 _27000_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08001_),
    .A(_00106_),
    .Y(_08002_));
 sg13g2_o21ai_1 _27001_ (.B1(_08002_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_07998_));
 sg13g2_mux4_1 _27002_ (.S0(_05369_),
    .A0(net1068),
    .A1(net1069),
    .A2(net1046),
    .A3(net1045),
    .S1(_06123_),
    .X(_08003_));
 sg13g2_mux4_1 _27003_ (.S0(_05369_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_06123_),
    .X(_08004_));
 sg13g2_nor2b_1 _27004_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08004_),
    .Y(_08005_));
 sg13g2_a21oi_1 _27005_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08003_),
    .Y(_08006_),
    .B1(_08005_));
 sg13g2_nand2b_1 _27006_ (.Y(_08007_),
    .B(net1044),
    .A_N(_05369_));
 sg13g2_nand3_1 _27007_ (.B(net1047),
    .C(_06123_),
    .A(_05369_),
    .Y(_08008_));
 sg13g2_o21ai_1 _27008_ (.B1(_08008_),
    .Y(_08009_),
    .A1(_06123_),
    .A2(_08007_));
 sg13g2_nand3_1 _27009_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08009_),
    .A(_00146_),
    .Y(_08010_));
 sg13g2_o21ai_1 _27010_ (.B1(_08010_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08006_));
 sg13g2_xor2_1 _27011_ (.B(clknet_leaf_68_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27012_ (.S0(_05372_),
    .A0(net1068),
    .A1(net1069),
    .A2(_07842_),
    .A3(net1045),
    .S1(_06128_),
    .X(_08011_));
 sg13g2_mux4_1 _27013_ (.S0(_05372_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_06128_),
    .X(_08012_));
 sg13g2_nor2b_1 _27014_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08012_),
    .Y(_08013_));
 sg13g2_a21oi_1 _27015_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08011_),
    .Y(_08014_),
    .B1(_08013_));
 sg13g2_nand2b_1 _27016_ (.Y(_08015_),
    .B(net1044),
    .A_N(_05372_));
 sg13g2_nand3_1 _27017_ (.B(net1047),
    .C(_06128_),
    .A(_05372_),
    .Y(_08016_));
 sg13g2_o21ai_1 _27018_ (.B1(_08016_),
    .Y(_08017_),
    .A1(_06128_),
    .A2(_08015_));
 sg13g2_nand3_1 _27019_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08017_),
    .A(_00149_),
    .Y(_08018_));
 sg13g2_o21ai_1 _27020_ (.B1(_08018_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08014_));
 sg13g2_mux4_1 _27021_ (.S0(_04706_),
    .A0(net1068),
    .A1(_11623_),
    .A2(net1046),
    .A3(net1045),
    .S1(_06132_),
    .X(_08019_));
 sg13g2_mux4_1 _27022_ (.S0(_04706_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(_06952_),
    .A2(net1066),
    .A3(net1067),
    .S1(_06132_),
    .X(_08020_));
 sg13g2_nor2b_1 _27023_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08020_),
    .Y(_08021_));
 sg13g2_a21oi_1 _27024_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08019_),
    .Y(_08022_),
    .B1(_08021_));
 sg13g2_nand2b_1 _27025_ (.Y(_08023_),
    .B(net1044),
    .A_N(_04706_));
 sg13g2_nand3_1 _27026_ (.B(net1047),
    .C(_06132_),
    .A(_04706_),
    .Y(_08024_));
 sg13g2_o21ai_1 _27027_ (.B1(_08024_),
    .Y(_08025_),
    .A1(_06132_),
    .A2(_08023_));
 sg13g2_nand3_1 _27028_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08025_),
    .A(_00108_),
    .Y(_08026_));
 sg13g2_o21ai_1 _27029_ (.B1(_08026_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08022_));
 sg13g2_mux4_1 _27030_ (.S0(_05366_),
    .A0(net1068),
    .A1(net1069),
    .A2(net1046),
    .A3(net1045),
    .S1(_06134_),
    .X(_08027_));
 sg13g2_mux4_1 _27031_ (.S0(_05366_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_06134_),
    .X(_08028_));
 sg13g2_nor2b_1 _27032_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08028_),
    .Y(_08029_));
 sg13g2_a21oi_1 _27033_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08027_),
    .Y(_08030_),
    .B1(_08029_));
 sg13g2_nand2b_1 _27034_ (.Y(_08031_),
    .B(net1044),
    .A_N(_05366_));
 sg13g2_nand3_1 _27035_ (.B(net1047),
    .C(_06134_),
    .A(_05366_),
    .Y(_08032_));
 sg13g2_o21ai_1 _27036_ (.B1(_08032_),
    .Y(_08033_),
    .A1(_06134_),
    .A2(_08031_));
 sg13g2_nand3_1 _27037_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08033_),
    .A(_00148_),
    .Y(_08034_));
 sg13g2_o21ai_1 _27038_ (.B1(_08034_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08030_));
 sg13g2_mux4_1 _27039_ (.S0(_04720_),
    .A0(net1068),
    .A1(net1069),
    .A2(net1046),
    .A3(_07844_),
    .S1(_07457_),
    .X(_08035_));
 sg13g2_mux4_1 _27040_ (.S0(_04720_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_07457_),
    .X(_08036_));
 sg13g2_nor2b_1 _27041_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08036_),
    .Y(_08037_));
 sg13g2_a21oi_1 _27042_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08035_),
    .Y(_08038_),
    .B1(_08037_));
 sg13g2_nand2b_1 _27043_ (.Y(_08039_),
    .B(net1044),
    .A_N(_04720_));
 sg13g2_nand3_1 _27044_ (.B(net1047),
    .C(_07457_),
    .A(_04720_),
    .Y(_08040_));
 sg13g2_o21ai_1 _27045_ (.B1(_08040_),
    .Y(_08041_),
    .A1(_07457_),
    .A2(_08039_));
 sg13g2_nand3_1 _27046_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08041_),
    .A(_00107_),
    .Y(_08042_));
 sg13g2_o21ai_1 _27047_ (.B1(_08042_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08038_));
 sg13g2_mux4_1 _27048_ (.S0(_05371_),
    .A0(_11630_),
    .A1(net1069),
    .A2(_07842_),
    .A3(_07844_),
    .S1(_06139_),
    .X(_08043_));
 sg13g2_mux4_1 _27049_ (.S0(_05371_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1048),
    .A2(net1066),
    .A3(net1067),
    .S1(_06139_),
    .X(_08044_));
 sg13g2_nor2b_1 _27050_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08044_),
    .Y(_08045_));
 sg13g2_a21oi_1 _27051_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08043_),
    .Y(_08046_),
    .B1(_08045_));
 sg13g2_nand2b_1 _27052_ (.Y(_08047_),
    .B(_07846_),
    .A_N(_05371_));
 sg13g2_nand3_1 _27053_ (.B(net1047),
    .C(_06139_),
    .A(_05371_),
    .Y(_08048_));
 sg13g2_o21ai_1 _27054_ (.B1(_08048_),
    .Y(_08049_),
    .A1(_06139_),
    .A2(_08047_));
 sg13g2_nand3_1 _27055_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08049_),
    .A(_00147_),
    .Y(_08050_));
 sg13g2_o21ai_1 _27056_ (.B1(_08050_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08046_));
 sg13g2_dfrbp_1 _27057_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1097),
    .D(_00317_),
    .Q_N(_14653_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27058_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1098),
    .D(_00318_),
    .Q_N(_14652_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27059_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1099),
    .D(_00319_),
    .Q_N(_14651_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27060_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1100),
    .D(_00320_),
    .Q_N(_14650_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27061_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1101),
    .D(_00321_),
    .Q_N(_14649_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27063_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27064_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1102),
    .D(_00322_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1103),
    .D(_00323_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1104),
    .D(_00324_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1105),
    .D(_00325_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1106),
    .D(_00326_),
    .Q_N(_00131_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1107),
    .D(_00327_),
    .Q_N(_00143_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1108),
    .D(_00328_),
    .Q_N(_00155_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1109),
    .D(_00329_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1110),
    .D(_00330_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1111),
    .D(_00331_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1112),
    .D(_00332_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1113),
    .D(_00333_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1114),
    .D(_00334_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1115),
    .D(_00335_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1116),
    .D(_00336_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1117),
    .D(_00337_),
    .Q_N(_00153_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1118),
    .D(_00338_),
    .Q_N(_00311_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1119),
    .D(_00339_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1120),
    .D(_00340_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1121),
    .D(_00341_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1122),
    .D(_00342_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1123),
    .D(_00343_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1124),
    .D(_00344_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1125),
    .D(_00345_),
    .Q_N(_00142_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1126),
    .D(_00346_),
    .Q_N(_00154_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1127),
    .D(_00347_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1128),
    .D(_00348_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1129),
    .D(_00349_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1130),
    .D(_00350_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1131),
    .D(_00351_),
    .Q_N(_00152_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1132),
    .D(_00352_),
    .Q_N(_00312_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1133),
    .D(_00353_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1134),
    .D(_00354_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1135),
    .D(_00355_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1136),
    .D(_00356_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1137),
    .D(_00357_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1138),
    .D(_00358_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1139),
    .D(_00359_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1140),
    .D(_00360_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1141),
    .D(_00361_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1142),
    .D(_00362_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1143),
    .D(_00363_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1144),
    .D(_00364_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1145),
    .D(_00365_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1146),
    .D(_00366_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1147),
    .D(_00367_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1148),
    .D(_00368_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1149),
    .D(_00369_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1150),
    .D(_00370_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1151),
    .D(_00371_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1152),
    .D(_00372_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1153),
    .D(_00373_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1154),
    .D(_00374_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1155),
    .D(_00375_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1156),
    .D(_00376_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1157),
    .D(_00377_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1158),
    .D(_00378_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1159),
    .D(_00379_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1160),
    .D(_00380_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1161),
    .D(_00381_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1162),
    .D(_00382_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1163),
    .D(_00383_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1164),
    .D(_00384_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1165),
    .D(_00385_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1166),
    .D(_00386_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1167),
    .D(_00387_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1168),
    .D(_00388_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1169),
    .D(_00389_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1170),
    .D(_00390_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1171),
    .D(_00391_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1172),
    .D(_00392_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1173),
    .D(_00393_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1174),
    .D(_00394_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1175),
    .D(_00395_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1176),
    .D(_00396_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1177),
    .D(_00397_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1178),
    .D(_00398_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1179),
    .D(_00399_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1180),
    .D(_00400_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1181),
    .D(_00401_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1182),
    .D(_00402_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1183),
    .D(_00403_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1184),
    .D(_00404_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1185),
    .D(_00405_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1186),
    .D(_00406_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1187),
    .D(_00407_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1188),
    .D(_00408_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1189),
    .D(_00409_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1190),
    .D(_00410_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1191),
    .D(_00411_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1192),
    .D(_00412_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1193),
    .D(_00413_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1194),
    .D(_00414_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1195),
    .D(_00415_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1196),
    .D(_00416_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1197),
    .D(_00417_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1198),
    .D(_00418_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1199),
    .D(_00419_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1200),
    .D(_00420_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1201),
    .D(_00421_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1202),
    .D(_00422_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1203),
    .D(_00423_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1204),
    .D(_00424_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1205),
    .D(_00425_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1206),
    .D(_00426_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1207),
    .D(_00427_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1208),
    .D(_00428_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1209),
    .D(_00429_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1210),
    .D(_00430_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1211),
    .D(_00431_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1212),
    .D(_00432_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1213),
    .D(_00433_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1214),
    .D(_00434_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1215),
    .D(_00435_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1216),
    .D(_00436_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1217),
    .D(_00437_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1218),
    .D(_00438_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1219),
    .D(_00439_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1220),
    .D(_00440_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1221),
    .D(_00441_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1222),
    .D(_00442_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1223),
    .D(_00443_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1224),
    .D(_00444_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1225),
    .D(_00445_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1226),
    .D(_00446_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1227),
    .D(_00447_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1228),
    .D(_00448_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1229),
    .D(_00449_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1230),
    .D(_00450_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1231),
    .D(_00451_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1232),
    .D(_00452_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1233),
    .D(_00453_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1234),
    .D(_00454_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1235),
    .D(_00455_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1236),
    .D(_00456_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1237),
    .D(_00457_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1238),
    .D(_00458_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1239),
    .D(_00459_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1240),
    .D(_00460_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1241),
    .D(_00461_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1242),
    .D(_00462_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1243),
    .D(_00463_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1244),
    .D(_00464_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1245),
    .D(_00465_),
    .Q_N(_14532_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1246),
    .D(_00466_),
    .Q_N(_14531_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1247),
    .D(_00467_),
    .Q_N(_14530_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1248),
    .D(_00468_),
    .Q_N(_14529_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1249),
    .D(_00469_),
    .Q_N(_14528_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1250),
    .D(_00470_),
    .Q_N(_14527_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1251),
    .D(_00471_),
    .Q_N(_14526_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1252),
    .D(_00472_),
    .Q_N(_14525_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1253),
    .D(_00473_),
    .Q_N(_14524_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1254),
    .D(_00474_),
    .Q_N(_14523_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1255),
    .D(_00475_),
    .Q_N(_14522_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1256),
    .D(_00476_),
    .Q_N(_14521_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1257),
    .D(_00477_),
    .Q_N(_14520_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1258),
    .D(_00478_),
    .Q_N(_14519_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1259),
    .D(_00479_),
    .Q_N(_14518_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1260),
    .D(_00480_),
    .Q_N(_14517_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1261),
    .D(_00481_),
    .Q_N(_14516_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1262),
    .D(_00482_),
    .Q_N(_14515_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1263),
    .D(_00483_),
    .Q_N(_14514_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1264),
    .D(_00484_),
    .Q_N(_14513_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1265),
    .D(_00485_),
    .Q_N(_14512_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1266),
    .D(_00486_),
    .Q_N(_14511_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1267),
    .D(_00487_),
    .Q_N(_14510_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1268),
    .D(_00488_),
    .Q_N(_14509_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1269),
    .D(_00489_),
    .Q_N(_14508_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1270),
    .D(_00490_),
    .Q_N(_14507_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1271),
    .D(_00491_),
    .Q_N(_14506_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1272),
    .D(_00492_),
    .Q_N(_14505_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1273),
    .D(_00493_),
    .Q_N(_14504_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1274),
    .D(_00494_),
    .Q_N(_14503_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1275),
    .D(_00495_),
    .Q_N(_14502_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1276),
    .D(_00496_),
    .Q_N(_14501_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1277),
    .D(_00497_),
    .Q_N(_14500_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1278),
    .D(_00498_),
    .Q_N(_14499_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1279),
    .D(_00499_),
    .Q_N(_14498_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1280),
    .D(_00500_),
    .Q_N(_14497_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1281),
    .D(_00501_),
    .Q_N(_14496_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1282),
    .D(_00502_),
    .Q_N(_14495_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1283),
    .D(_00503_),
    .Q_N(_14494_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1284),
    .D(_00504_),
    .Q_N(_14493_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1285),
    .D(_00505_),
    .Q_N(_14492_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1286),
    .D(_00506_),
    .Q_N(_14491_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1287),
    .D(_00507_),
    .Q_N(_14490_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1288),
    .D(_00508_),
    .Q_N(_14489_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1289),
    .D(_00509_),
    .Q_N(_14488_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1290),
    .D(_00510_),
    .Q_N(_14487_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1291),
    .D(_00511_),
    .Q_N(_14486_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1292),
    .D(_00512_),
    .Q_N(_14485_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1293),
    .D(_00513_),
    .Q_N(_14484_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1294),
    .D(_00514_),
    .Q_N(_14483_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1295),
    .D(_00515_),
    .Q_N(_14482_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1296),
    .D(_00516_),
    .Q_N(_14481_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1297),
    .D(_00517_),
    .Q_N(_14480_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1298),
    .D(_00518_),
    .Q_N(_14479_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1299),
    .D(_00519_),
    .Q_N(_14478_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1300),
    .D(_00520_),
    .Q_N(_14477_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1301),
    .D(_00521_),
    .Q_N(_14476_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1302),
    .D(_00522_),
    .Q_N(_14475_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1303),
    .D(_00523_),
    .Q_N(_14474_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1304),
    .D(_00524_),
    .Q_N(_14473_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1305),
    .D(_00525_),
    .Q_N(_14472_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1306),
    .D(_00526_),
    .Q_N(_14471_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1307),
    .D(_00527_),
    .Q_N(_14470_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1308),
    .D(_00528_),
    .Q_N(_14469_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1309),
    .D(_00529_),
    .Q_N(_14468_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1310),
    .D(_00530_),
    .Q_N(_14467_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1311),
    .D(_00531_),
    .Q_N(_14466_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1312),
    .D(_00532_),
    .Q_N(_14465_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1313),
    .D(_00533_),
    .Q_N(_14464_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1314),
    .D(_00534_),
    .Q_N(_14463_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1315),
    .D(_00535_),
    .Q_N(_14462_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1316),
    .D(_00536_),
    .Q_N(_14461_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1317),
    .D(_00537_),
    .Q_N(_14460_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1318),
    .D(_00538_),
    .Q_N(_14459_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1319),
    .D(_00539_),
    .Q_N(_14458_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1320),
    .D(_00540_),
    .Q_N(_14457_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1321),
    .D(_00541_),
    .Q_N(_14456_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1322),
    .D(_00542_),
    .Q_N(_14455_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1323),
    .D(_00543_),
    .Q_N(_14454_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1324),
    .D(_00544_),
    .Q_N(_14453_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1325),
    .D(_00545_),
    .Q_N(_14452_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1326),
    .D(_00546_),
    .Q_N(_14451_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1327),
    .D(_00547_),
    .Q_N(_14450_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1328),
    .D(_00548_),
    .Q_N(_14449_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1329),
    .D(_00549_),
    .Q_N(_14448_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1330),
    .D(_00550_),
    .Q_N(_14447_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1331),
    .D(_00551_),
    .Q_N(_14446_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1332),
    .D(_00552_),
    .Q_N(_14445_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1333),
    .D(_00553_),
    .Q_N(_14444_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1334),
    .D(_00554_),
    .Q_N(_14443_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1335),
    .D(_00555_),
    .Q_N(_14442_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1336),
    .D(_00556_),
    .Q_N(_14441_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1337),
    .D(_00557_),
    .Q_N(_14440_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1338),
    .D(_00558_),
    .Q_N(_14439_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1339),
    .D(_00559_),
    .Q_N(_14438_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1340),
    .D(_00560_),
    .Q_N(_14437_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1341),
    .D(_00561_),
    .Q_N(_14436_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1342),
    .D(_00562_),
    .Q_N(_14435_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1343),
    .D(_00563_),
    .Q_N(_14434_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1344),
    .D(_00564_),
    .Q_N(_14433_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1345),
    .D(_00565_),
    .Q_N(_14432_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1346),
    .D(_00566_),
    .Q_N(_14431_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1347),
    .D(_00567_),
    .Q_N(_14430_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1348),
    .D(_00568_),
    .Q_N(_14429_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1349),
    .D(_00569_),
    .Q_N(_14428_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1350),
    .D(_00570_),
    .Q_N(_14427_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1351),
    .D(_00571_),
    .Q_N(_14426_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1352),
    .D(_00572_),
    .Q_N(_14425_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1353),
    .D(_00573_),
    .Q_N(_14424_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1354),
    .D(_00574_),
    .Q_N(_14423_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1355),
    .D(_00575_),
    .Q_N(_14422_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1356),
    .D(_00576_),
    .Q_N(_14421_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1357),
    .D(_00577_),
    .Q_N(_14420_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1358),
    .D(_00578_),
    .Q_N(_14419_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1359),
    .D(_00579_),
    .Q_N(_14418_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1360),
    .D(_00580_),
    .Q_N(_14417_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1361),
    .D(_00581_),
    .Q_N(_14416_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1362),
    .D(_00582_),
    .Q_N(_14415_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1363),
    .D(_00583_),
    .Q_N(_14414_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1364),
    .D(_00584_),
    .Q_N(_14413_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1365),
    .D(_00585_),
    .Q_N(_14412_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1366),
    .D(_00586_),
    .Q_N(_00315_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1367),
    .D(_00587_),
    .Q_N(_14411_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1368),
    .D(_00588_),
    .Q_N(_00276_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1369),
    .D(_00589_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1370),
    .D(_00590_),
    .Q_N(_00246_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1371),
    .D(_00591_),
    .Q_N(_00247_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1372),
    .D(_00592_),
    .Q_N(_00248_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1373),
    .D(_00593_),
    .Q_N(_00249_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1374),
    .D(_00594_),
    .Q_N(_00250_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1375),
    .D(_00595_),
    .Q_N(_14410_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1376),
    .D(_00596_),
    .Q_N(_14409_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1377),
    .D(_00597_),
    .Q_N(_14408_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1378),
    .D(_00598_),
    .Q_N(_00251_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1379),
    .D(_00599_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1380),
    .D(_00600_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1381),
    .D(_00601_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1382),
    .D(_00602_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1383),
    .D(_00603_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1384),
    .D(_00604_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1385),
    .D(_00605_),
    .Q_N(_00243_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1386),
    .D(_00606_),
    .Q_N(_00244_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1387),
    .D(_00607_),
    .Q_N(_00245_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1388),
    .D(_00608_),
    .Q_N(_14407_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1389),
    .D(_00609_),
    .Q_N(_14406_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1390),
    .D(_00610_),
    .Q_N(_14405_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1391),
    .D(_00611_),
    .Q_N(_14404_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1392),
    .D(_00612_),
    .Q_N(_14403_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1393),
    .D(_00613_),
    .Q_N(_14402_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1394),
    .D(_00614_),
    .Q_N(_14401_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1395),
    .D(_00615_),
    .Q_N(_14400_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1396),
    .D(_00616_),
    .Q_N(_14399_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1397),
    .D(_00617_),
    .Q_N(_14398_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1398),
    .D(_00618_),
    .Q_N(_14397_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1399),
    .D(_00619_),
    .Q_N(_14396_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1400),
    .D(_00620_),
    .Q_N(_14395_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1401),
    .D(_00621_),
    .Q_N(_14394_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1402),
    .D(_00622_),
    .Q_N(_14393_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1403),
    .D(_00623_),
    .Q_N(_14392_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1404),
    .D(_00624_),
    .Q_N(_14391_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1405),
    .D(_00625_),
    .Q_N(_14390_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1406),
    .D(_00626_),
    .Q_N(_14389_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1407),
    .D(_00627_),
    .Q_N(_14388_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1408),
    .D(_00628_),
    .Q_N(_14387_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1409),
    .D(_00629_),
    .Q_N(_14386_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1410),
    .D(_00630_),
    .Q_N(_14385_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1411),
    .D(_00631_),
    .Q_N(_14384_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1412),
    .D(_00632_),
    .Q_N(_14383_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1413),
    .D(_00633_),
    .Q_N(_14382_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1414),
    .D(_00634_),
    .Q_N(_14381_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1415),
    .D(_00635_),
    .Q_N(_14380_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1416),
    .D(_00636_),
    .Q_N(_14379_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1417),
    .D(_00637_),
    .Q_N(_14378_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1418),
    .D(_00638_),
    .Q_N(_14377_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1419),
    .D(_00639_),
    .Q_N(_14376_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1420),
    .D(_00640_),
    .Q_N(_14375_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1421),
    .D(_00641_),
    .Q_N(_14374_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1422),
    .D(_00642_),
    .Q_N(_14373_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1423),
    .D(_00643_),
    .Q_N(_14372_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1424),
    .D(_00644_),
    .Q_N(_14371_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1425),
    .D(_00645_),
    .Q_N(_14370_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1426),
    .D(_00646_),
    .Q_N(_14369_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1427),
    .D(_00647_),
    .Q_N(_14368_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1428),
    .D(_00648_),
    .Q_N(_14367_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1429),
    .D(_00649_),
    .Q_N(_14366_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1430),
    .D(_00650_),
    .Q_N(_14365_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1431),
    .D(_00651_),
    .Q_N(_14364_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1432),
    .D(_00652_),
    .Q_N(_14363_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1433),
    .D(_00653_),
    .Q_N(_14362_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1434),
    .D(_00654_),
    .Q_N(_14361_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1435),
    .D(_00655_),
    .Q_N(_14360_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1436),
    .D(_00656_),
    .Q_N(_14359_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1437),
    .D(_00657_),
    .Q_N(_14358_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1438),
    .D(_00658_),
    .Q_N(_14357_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1439),
    .D(_00659_),
    .Q_N(_14356_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1440),
    .D(_00660_),
    .Q_N(_14355_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1441),
    .D(_00661_),
    .Q_N(_14354_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1442),
    .D(_00662_),
    .Q_N(_14353_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1443),
    .D(_00663_),
    .Q_N(_14352_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1444),
    .D(_00664_),
    .Q_N(_14351_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1445),
    .D(_00665_),
    .Q_N(_14350_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1446),
    .D(_00666_),
    .Q_N(_14349_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1447),
    .D(_00667_),
    .Q_N(_14348_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1448),
    .D(_00668_),
    .Q_N(_14347_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1449),
    .D(_00669_),
    .Q_N(_14346_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1450),
    .D(_00670_),
    .Q_N(_14345_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1451),
    .D(_00671_),
    .Q_N(_14344_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1452),
    .D(_00672_),
    .Q_N(_14343_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1453),
    .D(_00673_),
    .Q_N(_14342_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1454),
    .D(_00674_),
    .Q_N(_14341_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1455),
    .D(_00675_),
    .Q_N(_14340_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1456),
    .D(_00676_),
    .Q_N(_14339_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1457),
    .D(_00677_),
    .Q_N(_14338_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1458),
    .D(_00678_),
    .Q_N(_14337_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1459),
    .D(_00679_),
    .Q_N(_14336_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1460),
    .D(_00680_),
    .Q_N(_14335_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1461),
    .D(_00681_),
    .Q_N(_14334_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1462),
    .D(_00682_),
    .Q_N(_14333_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1463),
    .D(_00683_),
    .Q_N(_14332_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1464),
    .D(_00684_),
    .Q_N(_14331_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1465),
    .D(_00685_),
    .Q_N(_14330_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1466),
    .D(_00686_),
    .Q_N(_14329_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1467),
    .D(_00687_),
    .Q_N(_14328_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1468),
    .D(_00688_),
    .Q_N(_14327_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1469),
    .D(_00689_),
    .Q_N(_14326_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1470),
    .D(_00690_),
    .Q_N(_14325_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1471),
    .D(_00691_),
    .Q_N(_14324_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1472),
    .D(_00692_),
    .Q_N(_14323_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1473),
    .D(_00693_),
    .Q_N(_14322_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1474),
    .D(_00694_),
    .Q_N(_14321_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1475),
    .D(_00695_),
    .Q_N(_14320_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1476),
    .D(_00696_),
    .Q_N(_14319_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1477),
    .D(_00697_),
    .Q_N(_14318_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1478),
    .D(_00698_),
    .Q_N(_14317_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1479),
    .D(_00699_),
    .Q_N(_14316_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1480),
    .D(_00700_),
    .Q_N(_14315_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1481),
    .D(_00701_),
    .Q_N(_14314_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1482),
    .D(_00702_),
    .Q_N(_14313_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1483),
    .D(_00703_),
    .Q_N(_14312_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1484),
    .D(_00704_),
    .Q_N(_14311_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1485),
    .D(_00705_),
    .Q_N(_14310_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1486),
    .D(_00706_),
    .Q_N(_14309_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1487),
    .D(_00707_),
    .Q_N(_14308_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1488),
    .D(_00708_),
    .Q_N(_14307_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1489),
    .D(_00709_),
    .Q_N(_14306_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1490),
    .D(_00710_),
    .Q_N(_14305_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1491),
    .D(_00711_),
    .Q_N(_14304_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1492),
    .D(_00712_),
    .Q_N(_14303_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1493),
    .D(_00713_),
    .Q_N(_14302_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1494),
    .D(_00714_),
    .Q_N(_14301_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1495),
    .D(_00715_),
    .Q_N(_14300_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1496),
    .D(_00716_),
    .Q_N(_14299_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1497),
    .D(_00717_),
    .Q_N(_14298_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1498),
    .D(_00718_),
    .Q_N(_14297_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1499),
    .D(_00719_),
    .Q_N(_14296_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1500),
    .D(_00720_),
    .Q_N(_14295_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1501),
    .D(_00721_),
    .Q_N(_14294_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1502),
    .D(_00722_),
    .Q_N(_14293_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1503),
    .D(_00723_),
    .Q_N(_14292_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1504),
    .D(_00724_),
    .Q_N(_14291_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1505),
    .D(_00725_),
    .Q_N(_14290_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1506),
    .D(_00726_),
    .Q_N(_14289_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1507),
    .D(_00727_),
    .Q_N(_14288_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1508),
    .D(_00728_),
    .Q_N(_14287_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1509),
    .D(_00729_),
    .Q_N(_14286_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1510),
    .D(_00730_),
    .Q_N(_14285_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1511),
    .D(_00731_),
    .Q_N(_14284_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1512),
    .D(_00732_),
    .Q_N(_14283_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1513),
    .D(_00733_),
    .Q_N(_14282_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1514),
    .D(_00734_),
    .Q_N(_14281_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1515),
    .D(_00735_),
    .Q_N(_14280_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1516),
    .D(_00736_),
    .Q_N(_14279_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1517),
    .D(_00737_),
    .Q_N(_14278_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1518),
    .D(_00738_),
    .Q_N(_14277_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1519),
    .D(_00739_),
    .Q_N(_14276_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1520),
    .D(_00740_),
    .Q_N(_14275_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1521),
    .D(_00741_),
    .Q_N(_14274_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1522),
    .D(_00742_),
    .Q_N(_14273_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1523),
    .D(_00743_),
    .Q_N(_14272_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1524),
    .D(_00744_),
    .Q_N(_14271_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1525),
    .D(_00745_),
    .Q_N(_14270_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1526),
    .D(_00746_),
    .Q_N(_14269_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1527),
    .D(_00747_),
    .Q_N(_14268_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1528),
    .D(_00748_),
    .Q_N(_14267_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1529),
    .D(_00749_),
    .Q_N(_14266_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1530),
    .D(_00750_),
    .Q_N(_00298_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1531),
    .D(_00751_),
    .Q_N(_14265_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1532),
    .D(_00752_),
    .Q_N(_00273_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1533),
    .D(_00753_),
    .Q_N(_14264_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1534),
    .D(_00754_),
    .Q_N(_14263_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1535),
    .D(_00755_),
    .Q_N(_14262_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1536),
    .D(_00756_),
    .Q_N(_14261_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1537),
    .D(_00757_),
    .Q_N(_14260_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1538),
    .D(_00758_),
    .Q_N(_14259_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1539),
    .D(_00759_),
    .Q_N(_14258_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1540),
    .D(_00760_),
    .Q_N(_14257_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1541),
    .D(_00761_),
    .Q_N(_14256_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1542),
    .D(_00762_),
    .Q_N(_14255_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1543),
    .D(_00763_),
    .Q_N(_14254_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1544),
    .D(_00764_),
    .Q_N(_14253_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1545),
    .D(_00765_),
    .Q_N(_14252_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1546),
    .D(_00766_),
    .Q_N(_14251_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1547),
    .D(_00767_),
    .Q_N(_14250_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1548),
    .D(_00768_),
    .Q_N(_14249_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1549),
    .D(_00769_),
    .Q_N(_14248_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1550),
    .D(_00770_),
    .Q_N(_14247_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1551),
    .D(_00771_),
    .Q_N(_14246_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1552),
    .D(_00772_),
    .Q_N(_14245_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1553),
    .D(_00773_),
    .Q_N(_14244_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1554),
    .D(_00774_),
    .Q_N(_00258_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1555),
    .D(_00775_),
    .Q_N(_14243_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1556),
    .D(_00776_),
    .Q_N(_14242_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1557),
    .D(_00777_),
    .Q_N(_14654_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1558),
    .D(_00011_),
    .Q_N(_14655_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1559),
    .D(_00012_),
    .Q_N(_14656_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1560),
    .D(_00013_),
    .Q_N(_14657_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1561),
    .D(_00014_),
    .Q_N(_14658_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1562),
    .D(_00015_),
    .Q_N(_14659_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1563),
    .D(_00016_),
    .Q_N(_14660_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1564),
    .D(_00017_),
    .Q_N(_14661_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1565),
    .D(_00018_),
    .Q_N(_14662_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1566),
    .D(_00019_),
    .Q_N(_14663_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1567),
    .D(_00020_),
    .Q_N(_14241_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1568),
    .D(_00778_),
    .Q_N(_14240_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1569),
    .D(_00779_),
    .Q_N(_14239_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1570),
    .D(_00780_),
    .Q_N(_14238_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1571),
    .D(_00781_),
    .Q_N(_14664_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1572),
    .D(_00052_),
    .Q_N(_14237_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1573),
    .D(_00782_),
    .Q_N(_14236_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1574),
    .D(_00783_),
    .Q_N(_14235_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1575),
    .D(_00784_),
    .Q_N(_14234_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1576),
    .D(_00785_),
    .Q_N(_14233_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1577),
    .D(_00786_),
    .Q_N(_14232_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1578),
    .D(_00787_),
    .Q_N(_14231_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1579),
    .D(_00788_),
    .Q_N(_14230_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1580),
    .D(_00789_),
    .Q_N(_14229_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_inv$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1581),
    .D(_00790_),
    .Q_N(_14228_),
    .Q(\cpu.dec.r_rs2_inv ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1582),
    .D(_00791_),
    .Q_N(_14227_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1583),
    .D(_00792_),
    .Q_N(_14226_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1584),
    .D(_00793_),
    .Q_N(_00310_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1585),
    .D(_00794_),
    .Q_N(_14225_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1586),
    .D(_00795_),
    .Q_N(_00274_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1587),
    .D(_00796_),
    .Q_N(_14224_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1588),
    .D(_00797_),
    .Q_N(_14223_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1589),
    .D(_00798_),
    .Q_N(_00192_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1590),
    .D(_00799_),
    .Q_N(_14665_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1591),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00193_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1592),
    .D(_00800_),
    .Q_N(_14222_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1593),
    .D(_00801_),
    .Q_N(_14221_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1594),
    .D(_00802_),
    .Q_N(_14220_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1595),
    .D(_00803_),
    .Q_N(_14219_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1596),
    .D(_00804_),
    .Q_N(_14218_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1597),
    .D(_00805_),
    .Q_N(_14217_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1598),
    .D(_00806_),
    .Q_N(_14216_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1599),
    .D(_00807_),
    .Q_N(_14215_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1600),
    .D(_00808_),
    .Q_N(_14214_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1601),
    .D(_00809_),
    .Q_N(_14213_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1602),
    .D(_00810_),
    .Q_N(_14212_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1603),
    .D(_00811_),
    .Q_N(_14211_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1604),
    .D(_00812_),
    .Q_N(_14210_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1605),
    .D(_00813_),
    .Q_N(_14209_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1606),
    .D(_00814_),
    .Q_N(_14208_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1607),
    .D(_00815_),
    .Q_N(_14207_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1608),
    .D(_00816_),
    .Q_N(_14206_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1609),
    .D(_00817_),
    .Q_N(_14205_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1610),
    .D(_00818_),
    .Q_N(_14204_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1611),
    .D(_00819_),
    .Q_N(_14203_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1612),
    .D(_00820_),
    .Q_N(_14202_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1613),
    .D(_00821_),
    .Q_N(_14201_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1614),
    .D(_00822_),
    .Q_N(_14200_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1615),
    .D(_00823_),
    .Q_N(_14199_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1616),
    .D(_00824_),
    .Q_N(_14198_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1617),
    .D(_00825_),
    .Q_N(_14197_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1618),
    .D(_00826_),
    .Q_N(_14196_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1619),
    .D(_00827_),
    .Q_N(_14195_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1620),
    .D(_00828_),
    .Q_N(_14194_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1621),
    .D(_00829_),
    .Q_N(_14193_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1622),
    .D(_00830_),
    .Q_N(_14192_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1623),
    .D(_00831_),
    .Q_N(_14191_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1624),
    .D(_00832_),
    .Q_N(_14190_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1625),
    .D(_00833_),
    .Q_N(_14189_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1626),
    .D(_00834_),
    .Q_N(_14188_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1627),
    .D(_00835_),
    .Q_N(_14187_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1628),
    .D(_00836_),
    .Q_N(_14186_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1629),
    .D(_00837_),
    .Q_N(_14185_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1630),
    .D(_00838_),
    .Q_N(_14184_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1631),
    .D(_00839_),
    .Q_N(_14183_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1632),
    .D(_00840_),
    .Q_N(_14182_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1633),
    .D(_00841_),
    .Q_N(_14181_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1634),
    .D(_00842_),
    .Q_N(_14180_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1635),
    .D(_00843_),
    .Q_N(_14179_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1636),
    .D(_00844_),
    .Q_N(_14178_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1637),
    .D(_00845_),
    .Q_N(_14177_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1638),
    .D(_00846_),
    .Q_N(_14176_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1639),
    .D(_00847_),
    .Q_N(_14175_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1640),
    .D(_00848_),
    .Q_N(_14174_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1641),
    .D(_00849_),
    .Q_N(_14173_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1642),
    .D(_00850_),
    .Q_N(_14172_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1643),
    .D(_00851_),
    .Q_N(_14171_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1644),
    .D(_00852_),
    .Q_N(_14170_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1645),
    .D(_00853_),
    .Q_N(_14169_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1646),
    .D(_00854_),
    .Q_N(_14168_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1647),
    .D(_00855_),
    .Q_N(_14167_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1648),
    .D(_00856_),
    .Q_N(_14166_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1649),
    .D(_00857_),
    .Q_N(_14165_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1650),
    .D(_00858_),
    .Q_N(_14164_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1651),
    .D(_00859_),
    .Q_N(_14163_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1652),
    .D(_00860_),
    .Q_N(_14162_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1653),
    .D(_00861_),
    .Q_N(_14161_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1654),
    .D(_00862_),
    .Q_N(_14160_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1655),
    .D(_00863_),
    .Q_N(_14159_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1656),
    .D(_00864_),
    .Q_N(_14158_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1657),
    .D(_00865_),
    .Q_N(_14157_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1658),
    .D(_00866_),
    .Q_N(_14156_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1659),
    .D(_00867_),
    .Q_N(_14155_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1660),
    .D(_00868_),
    .Q_N(_14154_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1661),
    .D(_00869_),
    .Q_N(_14153_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1662),
    .D(_00870_),
    .Q_N(_14152_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1663),
    .D(_00871_),
    .Q_N(_14151_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1664),
    .D(_00872_),
    .Q_N(_14150_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1665),
    .D(_00873_),
    .Q_N(_14149_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1666),
    .D(_00874_),
    .Q_N(_14148_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1667),
    .D(_00875_),
    .Q_N(_14147_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1668),
    .D(_00876_),
    .Q_N(_14146_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1669),
    .D(_00877_),
    .Q_N(_14145_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1670),
    .D(_00878_),
    .Q_N(_14144_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1671),
    .D(_00879_),
    .Q_N(_14143_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1672),
    .D(_00880_),
    .Q_N(_14142_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1673),
    .D(_00881_),
    .Q_N(_14141_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1674),
    .D(_00882_),
    .Q_N(_00268_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1675),
    .D(_00883_),
    .Q_N(_00269_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1676),
    .D(_00884_),
    .Q_N(_00270_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1677),
    .D(_00885_),
    .Q_N(_00271_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1678),
    .D(_00886_),
    .Q_N(_00272_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1679),
    .D(_00887_),
    .Q_N(_14140_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1680),
    .D(_00888_),
    .Q_N(_00259_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1681),
    .D(_00889_),
    .Q_N(_00260_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1682),
    .D(_00890_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1683),
    .D(_00891_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1684),
    .D(_00892_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1685),
    .D(_00893_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1686),
    .D(_00894_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1687),
    .D(_00895_),
    .Q_N(_00266_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1688),
    .D(_00896_),
    .Q_N(_00267_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1689),
    .D(_00897_),
    .Q_N(_14139_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1690),
    .D(_00898_),
    .Q_N(_14138_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1691),
    .D(_00899_),
    .Q_N(_14137_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1692),
    .D(_00900_),
    .Q_N(_14136_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1693),
    .D(_00901_),
    .Q_N(_14135_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1694),
    .D(_00902_),
    .Q_N(_14134_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1695),
    .D(_00903_),
    .Q_N(_14133_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1696),
    .D(_00904_),
    .Q_N(_14132_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1697),
    .D(_00905_),
    .Q_N(_14131_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1698),
    .D(_00906_),
    .Q_N(_14130_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1699),
    .D(_00907_),
    .Q_N(_14129_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1700),
    .D(_00908_),
    .Q_N(_14128_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1701),
    .D(_00909_),
    .Q_N(_14127_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1702),
    .D(_00910_),
    .Q_N(_14126_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1703),
    .D(_00911_),
    .Q_N(_14125_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1704),
    .D(_00912_),
    .Q_N(_14124_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1705),
    .D(_00913_),
    .Q_N(_14123_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1706),
    .D(_00914_),
    .Q_N(_14122_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1707),
    .D(_00915_),
    .Q_N(_14121_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1708),
    .D(_00916_),
    .Q_N(_14120_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1709),
    .D(_00917_),
    .Q_N(_14119_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1710),
    .D(_00918_),
    .Q_N(_14118_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1711),
    .D(_00919_),
    .Q_N(_14117_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1712),
    .D(_00920_),
    .Q_N(_14116_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1713),
    .D(_00921_),
    .Q_N(_14115_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1714),
    .D(_00922_),
    .Q_N(_14114_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1715),
    .D(_00923_),
    .Q_N(_14113_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1716),
    .D(_00924_),
    .Q_N(_14112_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1717),
    .D(_00925_),
    .Q_N(_14111_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1718),
    .D(_00926_),
    .Q_N(_14110_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1719),
    .D(_00927_),
    .Q_N(_14109_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1720),
    .D(_00928_),
    .Q_N(_14666_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1721),
    .D(_00053_),
    .Q_N(_14108_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1722),
    .D(_00929_),
    .Q_N(_14107_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1723),
    .D(_00930_),
    .Q_N(_14667_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1724),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14106_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1725),
    .D(_00931_),
    .Q_N(_14105_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1726),
    .D(_00932_),
    .Q_N(_14104_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1727),
    .D(_00933_),
    .Q_N(_14103_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1728),
    .D(_00934_),
    .Q_N(_14102_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1729),
    .D(_00935_),
    .Q_N(_14101_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1730),
    .D(_00936_),
    .Q_N(_14100_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1731),
    .D(_00937_),
    .Q_N(_14099_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1732),
    .D(_00938_),
    .Q_N(_14098_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1733),
    .D(_00939_),
    .Q_N(_14097_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1734),
    .D(_00940_),
    .Q_N(_14096_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1735),
    .D(_00941_),
    .Q_N(_14095_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1736),
    .D(_00942_),
    .Q_N(_14094_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1737),
    .D(_00943_),
    .Q_N(_14093_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1738),
    .D(_00944_),
    .Q_N(_14092_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1739),
    .D(_00945_),
    .Q_N(_14091_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1740),
    .D(_00946_),
    .Q_N(_00189_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1741),
    .D(_00947_),
    .Q_N(_14090_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1742),
    .D(_00948_),
    .Q_N(_14089_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1743),
    .D(_00949_),
    .Q_N(_14088_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1744),
    .D(_00950_),
    .Q_N(_00197_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1745),
    .D(_00951_),
    .Q_N(_14087_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1746),
    .D(_00952_),
    .Q_N(_14086_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1747),
    .D(_00953_),
    .Q_N(_14085_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1748),
    .D(_00954_),
    .Q_N(_14084_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1749),
    .D(_00955_),
    .Q_N(_14083_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1750),
    .D(_00956_),
    .Q_N(_14082_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1751),
    .D(_00957_),
    .Q_N(_14081_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1752),
    .D(_00958_),
    .Q_N(_14080_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1753),
    .D(_00959_),
    .Q_N(_14079_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1754),
    .D(_00960_),
    .Q_N(_14078_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1755),
    .D(_00961_),
    .Q_N(_14077_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1756),
    .D(_00962_),
    .Q_N(_14076_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1757),
    .D(_00963_),
    .Q_N(_14075_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1758),
    .D(_00964_),
    .Q_N(_14074_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1759),
    .D(_00965_),
    .Q_N(_14668_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1760),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14669_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1761),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00167_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1762),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00168_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1763),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00169_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1764),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00170_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1765),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00171_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1766),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14073_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1767),
    .D(_00966_),
    .Q_N(_00309_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1768),
    .D(_00967_),
    .Q_N(_00308_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1769),
    .D(_00968_),
    .Q_N(_00307_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1770),
    .D(_00969_),
    .Q_N(_00306_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1771),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14072_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1772),
    .D(_00970_),
    .Q_N(_00305_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1773),
    .D(_00971_),
    .Q_N(_00304_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1774),
    .D(_00972_),
    .Q_N(_14071_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1775),
    .D(_00973_),
    .Q_N(_00303_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1776),
    .D(_00974_),
    .Q_N(_00302_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1777),
    .D(_00975_),
    .Q_N(_00301_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1778),
    .D(_00976_),
    .Q_N(_14070_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1779),
    .D(_00977_),
    .Q_N(_00300_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1780),
    .D(_00978_),
    .Q_N(_14069_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1781),
    .D(_00979_),
    .Q_N(_14670_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1782),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1783),
    .D(_00980_),
    .Q_N(_00299_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1784),
    .D(_00981_),
    .Q_N(_14671_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1785),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00127_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1786),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00139_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1787),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00151_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1788),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1789),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00164_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1790),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00165_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1791),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00166_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1792),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14672_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1793),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14673_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1794),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14674_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1795),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14675_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1796),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00199_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1797),
    .D(_00982_),
    .Q_N(_00200_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1798),
    .D(_00983_),
    .Q_N(_00290_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1799),
    .D(_00984_),
    .Q_N(_00289_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1800),
    .D(_00985_),
    .Q_N(_00196_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1801),
    .D(_00986_),
    .Q_N(_00195_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1802),
    .D(_00987_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1803),
    .D(_00988_),
    .Q_N(_00297_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1804),
    .D(_00989_),
    .Q_N(_00191_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1805),
    .D(_00990_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1806),
    .D(_00991_),
    .Q_N(_00296_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1807),
    .D(_00992_),
    .Q_N(_00295_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1808),
    .D(_00993_),
    .Q_N(_00294_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1809),
    .D(_00994_),
    .Q_N(_00293_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1810),
    .D(_00995_),
    .Q_N(_00292_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1811),
    .D(_00996_),
    .Q_N(_00291_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1812),
    .D(_00997_),
    .Q_N(_14068_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1813),
    .D(_00998_),
    .Q_N(_00198_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1814),
    .D(_00999_),
    .Q_N(_14067_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1815),
    .D(_01000_),
    .Q_N(_14066_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1816),
    .D(_01001_),
    .Q_N(_14065_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1817),
    .D(_01002_),
    .Q_N(_14064_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1818),
    .D(_01003_),
    .Q_N(_14063_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1819),
    .D(_01004_),
    .Q_N(_14062_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1820),
    .D(_01005_),
    .Q_N(_14061_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1821),
    .D(_01006_),
    .Q_N(_14060_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1822),
    .D(_01007_),
    .Q_N(_14059_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1823),
    .D(_01008_),
    .Q_N(_14058_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1824),
    .D(_01009_),
    .Q_N(_14057_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1825),
    .D(_01010_),
    .Q_N(_14056_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1826),
    .D(_01011_),
    .Q_N(_14055_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1827),
    .D(_01012_),
    .Q_N(_14054_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1828),
    .D(_01013_),
    .Q_N(_14053_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1829),
    .D(_01014_),
    .Q_N(_14052_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1830),
    .D(_01015_),
    .Q_N(_14051_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1831),
    .D(_01016_),
    .Q_N(_14050_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1832),
    .D(_01017_),
    .Q_N(_14049_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1833),
    .D(_01018_),
    .Q_N(_14048_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1834),
    .D(_01019_),
    .Q_N(_14047_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1835),
    .D(_01020_),
    .Q_N(_14046_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1836),
    .D(_01021_),
    .Q_N(_14045_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1837),
    .D(_01022_),
    .Q_N(_14044_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1838),
    .D(_01023_),
    .Q_N(_14043_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1839),
    .D(_01024_),
    .Q_N(_14042_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1840),
    .D(_01025_),
    .Q_N(_14041_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1841),
    .D(_01026_),
    .Q_N(_14040_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1842),
    .D(_01027_),
    .Q_N(_14039_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1843),
    .D(_01028_),
    .Q_N(_14038_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1844),
    .D(_01029_),
    .Q_N(_14037_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1845),
    .D(_01030_),
    .Q_N(_14036_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1846),
    .D(_01031_),
    .Q_N(_00257_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1847),
    .D(_01032_),
    .Q_N(_00239_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1848),
    .D(_01033_),
    .Q_N(_00241_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1849),
    .D(_01034_),
    .Q_N(_14035_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1850),
    .D(_01035_),
    .Q_N(_14034_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1851),
    .D(_01036_),
    .Q_N(_14033_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1852),
    .D(_01037_),
    .Q_N(_14032_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1853),
    .D(_01038_),
    .Q_N(_00275_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1854),
    .D(_01039_),
    .Q_N(_14031_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1855),
    .D(_01040_),
    .Q_N(_00228_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1856),
    .D(_01041_),
    .Q_N(_00227_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1857),
    .D(_01042_),
    .Q_N(_00229_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1858),
    .D(_01043_),
    .Q_N(_00231_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1859),
    .D(_01044_),
    .Q_N(_00233_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1860),
    .D(_01045_),
    .Q_N(_00235_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1861),
    .D(_01046_),
    .Q_N(_00237_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1862),
    .D(_01047_),
    .Q_N(_14030_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1863),
    .D(_01048_),
    .Q_N(_14029_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1864),
    .D(_01049_),
    .Q_N(_14028_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1865),
    .D(_01050_),
    .Q_N(_14027_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1866),
    .D(_01051_),
    .Q_N(_14676_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1867),
    .D(_00054_),
    .Q_N(_00256_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1868),
    .D(_01052_),
    .Q_N(_00223_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1869),
    .D(_01053_),
    .Q_N(_14026_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1870),
    .D(_01054_),
    .Q_N(_14025_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1871),
    .D(_01055_),
    .Q_N(_14024_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1872),
    .D(_01056_),
    .Q_N(_14023_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1873),
    .D(_01057_),
    .Q_N(_14022_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1874),
    .D(_01058_),
    .Q_N(_14021_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1875),
    .D(_01059_),
    .Q_N(_00178_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1876),
    .D(_01060_),
    .Q_N(_00179_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1877),
    .D(_01061_),
    .Q_N(_00287_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1878),
    .D(_01062_),
    .Q_N(_00180_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1879),
    .D(_01063_),
    .Q_N(_00181_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1880),
    .D(_01064_),
    .Q_N(_00182_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1881),
    .D(_01065_),
    .Q_N(_00281_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1882),
    .D(_01066_),
    .Q_N(_14020_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1883),
    .D(_01067_),
    .Q_N(_14019_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1884),
    .D(_01068_),
    .Q_N(_14018_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1885),
    .D(_01069_),
    .Q_N(_14017_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1886),
    .D(_01070_),
    .Q_N(_00288_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1887),
    .D(_01071_),
    .Q_N(_14016_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1888),
    .D(_01072_),
    .Q_N(_00188_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1889),
    .D(_01073_),
    .Q_N(_14015_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1890),
    .D(_01074_),
    .Q_N(_00255_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1891),
    .D(_01075_),
    .Q_N(_14014_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1892),
    .D(_01076_),
    .Q_N(_14013_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1893),
    .D(_01077_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1894),
    .D(_01078_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1895),
    .D(_01079_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1896),
    .D(_01080_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1897),
    .D(_01081_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1898),
    .D(_01082_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1899),
    .D(_01083_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1900),
    .D(_01084_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1901),
    .D(_01085_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1902),
    .D(_01086_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1903),
    .D(_01087_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1904),
    .D(_01088_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1905),
    .D(_01089_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1906),
    .D(_01090_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1907),
    .D(_01091_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1908),
    .D(_01092_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1909),
    .D(_01093_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1910),
    .D(_01094_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1911),
    .D(_01095_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1912),
    .D(_01096_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1913),
    .D(_01097_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1914),
    .D(_01098_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1915),
    .D(_01099_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1916),
    .D(_01100_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1917),
    .D(_01101_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1918),
    .D(_01102_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1919),
    .D(_01103_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1920),
    .D(_01104_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1921),
    .D(_01105_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1922),
    .D(_01106_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1923),
    .D(_01107_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1924),
    .D(_01108_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1925),
    .D(_01109_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1926),
    .D(_01110_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1927),
    .D(_01111_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1928),
    .D(_01112_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1929),
    .D(_01113_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1930),
    .D(_01114_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1931),
    .D(_01115_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1932),
    .D(_01116_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1933),
    .D(_01117_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1934),
    .D(_01118_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1935),
    .D(_01119_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1936),
    .D(_01120_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1937),
    .D(_01121_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1938),
    .D(_01122_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1939),
    .D(_01123_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1940),
    .D(_01124_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1941),
    .D(_01125_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1942),
    .D(_01126_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1943),
    .D(_01127_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1944),
    .D(_01128_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1945),
    .D(_01129_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1946),
    .D(_01130_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1947),
    .D(_01131_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1948),
    .D(_01132_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1949),
    .D(_01133_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1950),
    .D(_01134_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1951),
    .D(_01135_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1952),
    .D(_01136_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1953),
    .D(_01137_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1954),
    .D(_01138_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1955),
    .D(_01139_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1956),
    .D(_01140_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1957),
    .D(_01141_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1958),
    .D(_01142_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1959),
    .D(_01143_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1960),
    .D(_01144_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1961),
    .D(_01145_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1962),
    .D(_01146_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1963),
    .D(_01147_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1964),
    .D(_01148_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1965),
    .D(_01149_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1966),
    .D(_01150_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1967),
    .D(_01151_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1968),
    .D(_01152_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1969),
    .D(_01153_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1970),
    .D(_01154_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1971),
    .D(_01155_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1972),
    .D(_01156_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1973),
    .D(_01157_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1974),
    .D(_01158_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1975),
    .D(_01159_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1976),
    .D(_01160_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1977),
    .D(_01161_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1978),
    .D(_01162_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1979),
    .D(_01163_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1980),
    .D(_01164_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1981),
    .D(_01165_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1982),
    .D(_01166_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1983),
    .D(_01167_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1984),
    .D(_01168_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1985),
    .D(_01169_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1986),
    .D(_01170_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1987),
    .D(_01171_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1988),
    .D(_01172_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1989),
    .D(_01173_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1990),
    .D(_01174_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1991),
    .D(_01175_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1992),
    .D(_01176_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1993),
    .D(_01177_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1994),
    .D(_01178_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1995),
    .D(_01179_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1996),
    .D(_01180_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1997),
    .D(_01181_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1998),
    .D(_01182_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1999),
    .D(_01183_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2000),
    .D(_01184_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2001),
    .D(_01185_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2002),
    .D(_01186_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2003),
    .D(_01187_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2004),
    .D(_01188_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2005),
    .D(_01189_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2006),
    .D(_01190_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2007),
    .D(_01191_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2008),
    .D(_01192_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2009),
    .D(_01193_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2010),
    .D(_01194_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2011),
    .D(_01195_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2012),
    .D(_01196_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2013),
    .D(_01197_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2014),
    .D(_01198_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2015),
    .D(_01199_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2016),
    .D(_01200_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2017),
    .D(_01201_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2018),
    .D(_01202_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2019),
    .D(_01203_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2020),
    .D(_01204_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2021),
    .D(_01205_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2022),
    .D(_01206_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2023),
    .D(_01207_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2024),
    .D(_01208_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2025),
    .D(_01209_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2026),
    .D(_01210_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2027),
    .D(_01211_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2028),
    .D(_01212_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2029),
    .D(_01213_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2030),
    .D(_01214_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2031),
    .D(_01215_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2032),
    .D(_01216_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2033),
    .D(_01217_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2034),
    .D(_01218_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2035),
    .D(_01219_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2036),
    .D(_01220_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2037),
    .D(_01221_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2038),
    .D(_01222_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2039),
    .D(_01223_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2040),
    .D(_01224_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2041),
    .D(_01225_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2042),
    .D(_01226_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2043),
    .D(_01227_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2044),
    .D(_01228_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2045),
    .D(_01229_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2046),
    .D(_01230_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2047),
    .D(_01231_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2048),
    .D(_01232_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2049),
    .D(_01233_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2050),
    .D(_01234_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2051),
    .D(_01235_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2052),
    .D(_01236_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2053),
    .D(_01237_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2054),
    .D(_01238_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2055),
    .D(_01239_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2056),
    .D(_01240_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2057),
    .D(_01241_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2058),
    .D(_01242_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2059),
    .D(_01243_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2060),
    .D(_01244_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2061),
    .D(_01245_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2062),
    .D(_01246_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2063),
    .D(_01247_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2064),
    .D(_01248_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2065),
    .D(_01249_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2066),
    .D(_01250_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2067),
    .D(_01251_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2068),
    .D(_01252_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2069),
    .D(_01253_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2070),
    .D(_01254_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2071),
    .D(_01255_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2072),
    .D(_01256_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2073),
    .D(_01257_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2074),
    .D(_01258_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2075),
    .D(_01259_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2076),
    .D(_01260_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2077),
    .D(_01261_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2078),
    .D(_01262_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2079),
    .D(_01263_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2080),
    .D(_01264_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2081),
    .D(_01265_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2082),
    .D(_01266_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2083),
    .D(_01267_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2084),
    .D(_01268_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2085),
    .D(_01269_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2086),
    .D(_01270_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2087),
    .D(_01271_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2088),
    .D(_01272_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2089),
    .D(_01273_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2090),
    .D(_01274_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2091),
    .D(_01275_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2092),
    .D(_01276_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2093),
    .D(_01277_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2094),
    .D(_01278_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2095),
    .D(_01279_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2096),
    .D(_01280_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2097),
    .D(_01281_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2098),
    .D(_01282_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2099),
    .D(_01283_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2100),
    .D(_01284_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2101),
    .D(_01285_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2102),
    .D(_01286_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2103),
    .D(_01287_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2104),
    .D(_01288_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2105),
    .D(_01289_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2106),
    .D(_01290_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2107),
    .D(_01291_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2108),
    .D(_01292_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2109),
    .D(_01293_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2110),
    .D(_01294_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2111),
    .D(_01295_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2112),
    .D(_01296_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2113),
    .D(_01297_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2114),
    .D(_01298_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2115),
    .D(_01299_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2116),
    .D(_01300_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2117),
    .D(_01301_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2118),
    .D(_01302_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2119),
    .D(_01303_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2120),
    .D(_01304_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2121),
    .D(_01305_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2122),
    .D(_01306_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2123),
    .D(_01307_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2124),
    .D(_01308_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2125),
    .D(_01309_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2126),
    .D(_01310_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2127),
    .D(_01311_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2128),
    .D(_01312_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2129),
    .D(_01313_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2130),
    .D(_01314_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2131),
    .D(_01315_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2132),
    .D(_01316_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2133),
    .D(_01317_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2134),
    .D(_01318_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2135),
    .D(_01319_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2136),
    .D(_01320_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2137),
    .D(_01321_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2138),
    .D(_01322_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2139),
    .D(_01323_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2140),
    .D(_01324_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2141),
    .D(_01325_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2142),
    .D(_01326_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2143),
    .D(_01327_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2144),
    .D(_01328_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2145),
    .D(_01329_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2146),
    .D(_01330_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2147),
    .D(_01331_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2148),
    .D(_01332_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2149),
    .D(_01333_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2150),
    .D(_01334_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2151),
    .D(_01335_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2152),
    .D(_01336_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2153),
    .D(_01337_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2154),
    .D(_01338_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2155),
    .D(_01339_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2156),
    .D(_01340_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2157),
    .D(_01341_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2158),
    .D(_01342_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2159),
    .D(_01343_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2160),
    .D(_01344_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2161),
    .D(_01345_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2162),
    .D(_01346_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2163),
    .D(_01347_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2164),
    .D(_01348_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2165),
    .D(_01349_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2166),
    .D(_01350_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2167),
    .D(_01351_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2168),
    .D(_01352_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2169),
    .D(_01353_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2170),
    .D(_01354_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2171),
    .D(_01355_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2172),
    .D(_01356_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2173),
    .D(_01357_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2174),
    .D(_01358_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2175),
    .D(_01359_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2176),
    .D(_01360_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2177),
    .D(_01361_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2178),
    .D(_01362_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2179),
    .D(_01363_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2180),
    .D(_01364_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2181),
    .D(_01365_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2182),
    .D(_01366_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2183),
    .D(_01367_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2184),
    .D(_01368_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2185),
    .D(_01369_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2186),
    .D(_01370_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2187),
    .D(_01371_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2188),
    .D(_01372_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2189),
    .D(_01373_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2190),
    .D(_01374_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2191),
    .D(_01375_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2192),
    .D(_01376_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2193),
    .D(_01377_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2194),
    .D(_01378_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2195),
    .D(_01379_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2196),
    .D(_01380_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2197),
    .D(_01381_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2198),
    .D(_01382_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2199),
    .D(_01383_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2200),
    .D(_01384_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2201),
    .D(_01385_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2202),
    .D(_01386_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2203),
    .D(_01387_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2204),
    .D(_01388_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2205),
    .D(_01389_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2206),
    .D(_01390_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2207),
    .D(_01391_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2208),
    .D(_01392_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2209),
    .D(_01393_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2210),
    .D(_01394_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2211),
    .D(_01395_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2212),
    .D(_01396_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2213),
    .D(_01397_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2214),
    .D(_01398_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2215),
    .D(_01399_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2216),
    .D(_01400_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2217),
    .D(_01401_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2218),
    .D(_01402_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2219),
    .D(_01403_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2220),
    .D(_01404_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2221),
    .D(_01405_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2222),
    .D(_01406_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2223),
    .D(_01407_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2224),
    .D(_01408_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2225),
    .D(_01409_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2226),
    .D(_01410_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2227),
    .D(_01411_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2228),
    .D(_01412_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2229),
    .D(_01413_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2230),
    .D(_01414_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2231),
    .D(_01415_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2232),
    .D(_01416_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2233),
    .D(_01417_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2234),
    .D(_01418_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2235),
    .D(_01419_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2236),
    .D(_01420_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2237),
    .D(_01421_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2238),
    .D(_01422_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2239),
    .D(_01423_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2240),
    .D(_01424_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2241),
    .D(_01425_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2242),
    .D(_01426_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2243),
    .D(_01427_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2244),
    .D(_01428_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2245),
    .D(_01429_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2246),
    .D(_01430_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2247),
    .D(_01431_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2248),
    .D(_01432_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2249),
    .D(_01433_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2250),
    .D(_01434_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2251),
    .D(_01435_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2252),
    .D(_01436_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2253),
    .D(_01437_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2254),
    .D(_01438_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2255),
    .D(_01439_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2256),
    .D(_01440_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2257),
    .D(_01441_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2258),
    .D(_01442_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2259),
    .D(_01443_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2260),
    .D(_01444_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2261),
    .D(_01445_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2262),
    .D(_01446_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2263),
    .D(_01447_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2264),
    .D(_01448_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2265),
    .D(_01449_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2266),
    .D(_01450_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2267),
    .D(_01451_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2268),
    .D(_01452_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2269),
    .D(_01453_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2270),
    .D(_01454_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2271),
    .D(_01455_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2272),
    .D(_01456_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2273),
    .D(_01457_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2274),
    .D(_01458_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2275),
    .D(_01459_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2276),
    .D(_01460_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2277),
    .D(_01461_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2278),
    .D(_01462_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2279),
    .D(_01463_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2280),
    .D(_01464_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2281),
    .D(_01465_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2282),
    .D(_01466_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2283),
    .D(_01467_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2284),
    .D(_01468_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2285),
    .D(_01469_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2286),
    .D(_01470_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2287),
    .D(_01471_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2288),
    .D(_01472_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2289),
    .D(_01473_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2290),
    .D(_01474_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2291),
    .D(_01475_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2292),
    .D(_01476_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2293),
    .D(_01477_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2294),
    .D(_01478_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2295),
    .D(_01479_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2296),
    .D(_01480_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2297),
    .D(_01481_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2298),
    .D(_01482_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2299),
    .D(_01483_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2300),
    .D(_01484_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2301),
    .D(_01485_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2302),
    .D(_01486_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2303),
    .D(_01487_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2304),
    .D(_01488_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2305),
    .D(_01489_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2306),
    .D(_01490_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2307),
    .D(_01491_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2308),
    .D(_01492_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2309),
    .D(_01493_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2310),
    .D(_01494_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2311),
    .D(_01495_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2312),
    .D(_01496_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2313),
    .D(_01497_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2314),
    .D(_01498_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2315),
    .D(_01499_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2316),
    .D(_01500_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2317),
    .D(_01501_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2318),
    .D(_01502_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2319),
    .D(_01503_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2320),
    .D(_01504_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2321),
    .D(_01505_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2322),
    .D(_01506_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2323),
    .D(_01507_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2324),
    .D(_01508_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2325),
    .D(_01509_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2326),
    .D(_01510_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2327),
    .D(_01511_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2328),
    .D(_01512_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2329),
    .D(_01513_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2330),
    .D(_01514_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2331),
    .D(_01515_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2332),
    .D(_01516_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2333),
    .D(_01517_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2334),
    .D(_01518_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2335),
    .D(_01519_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2336),
    .D(_01520_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2337),
    .D(_01521_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2338),
    .D(_01522_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2339),
    .D(_01523_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2340),
    .D(_01524_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2341),
    .D(_01525_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2342),
    .D(_01526_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2343),
    .D(_01527_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2344),
    .D(_01528_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2345),
    .D(_01529_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2346),
    .D(_01530_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2347),
    .D(_01531_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2348),
    .D(_01532_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2349),
    .D(_01533_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2350),
    .D(_01534_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2351),
    .D(_01535_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2352),
    .D(_01536_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2353),
    .D(_01537_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2354),
    .D(_01538_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2355),
    .D(_01539_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2356),
    .D(_01540_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2357),
    .D(_01541_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2358),
    .D(_01542_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2359),
    .D(_01543_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2360),
    .D(_01544_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2361),
    .D(_01545_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2362),
    .D(_01546_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2363),
    .D(_01547_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2364),
    .D(_01548_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2365),
    .D(_01549_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2366),
    .D(_01550_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2367),
    .D(_01551_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2368),
    .D(_01552_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2369),
    .D(_01553_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2370),
    .D(_01554_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2371),
    .D(_01555_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2372),
    .D(_01556_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2373),
    .D(_01557_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2374),
    .D(_01558_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2375),
    .D(_01559_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2376),
    .D(_01560_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2377),
    .D(_01561_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2378),
    .D(_01562_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2379),
    .D(_01563_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2380),
    .D(_01564_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2381),
    .D(_01565_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2382),
    .D(_01566_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2383),
    .D(_01567_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2384),
    .D(_01568_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2385),
    .D(_01569_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2386),
    .D(_01570_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2387),
    .D(_01571_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2388),
    .D(_01572_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2389),
    .D(_01573_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2390),
    .D(_01574_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2391),
    .D(_01575_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2392),
    .D(_01576_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2393),
    .D(_01577_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2394),
    .D(_01578_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2395),
    .D(_01579_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2396),
    .D(_01580_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2397),
    .D(_01581_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2398),
    .D(_01582_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2399),
    .D(_01583_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2400),
    .D(_01584_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2401),
    .D(_01585_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2402),
    .D(_01586_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2403),
    .D(_01587_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2404),
    .D(_01588_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2405),
    .D(_01589_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2406),
    .D(_01590_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2407),
    .D(_01591_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2408),
    .D(_01592_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2409),
    .D(_01593_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2410),
    .D(_01594_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2411),
    .D(_01595_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2412),
    .D(_01596_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2413),
    .D(_01597_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2414),
    .D(_01598_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2415),
    .D(_01599_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2416),
    .D(_01600_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2417),
    .D(_01601_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2418),
    .D(_01602_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2419),
    .D(_01603_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2420),
    .D(_01604_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2421),
    .D(_01605_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2422),
    .D(_01606_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2423),
    .D(_01607_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2424),
    .D(_01608_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2425),
    .D(_01609_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2426),
    .D(_01610_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2427),
    .D(_01611_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2428),
    .D(_01612_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2429),
    .D(_01613_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2430),
    .D(_01614_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2431),
    .D(_01615_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2432),
    .D(_01616_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2433),
    .D(_01617_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2434),
    .D(_01618_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2435),
    .D(_01619_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2436),
    .D(_01620_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2437),
    .D(_01621_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2438),
    .D(_01622_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2439),
    .D(_01623_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2440),
    .D(_01624_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2441),
    .D(_01625_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2442),
    .D(_01626_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2443),
    .D(_01627_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2444),
    .D(_01628_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2445),
    .D(_01629_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2446),
    .D(_01630_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2447),
    .D(_01631_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2448),
    .D(_01632_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2449),
    .D(_01633_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2450),
    .D(_01634_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2451),
    .D(_01635_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2452),
    .D(_01636_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2453),
    .D(_01637_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2454),
    .D(_01638_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2455),
    .D(_01639_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2456),
    .D(_01640_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2457),
    .D(_01641_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2458),
    .D(_01642_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2459),
    .D(_01643_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2460),
    .D(_01644_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2461),
    .D(_01645_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2462),
    .D(_01646_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2463),
    .D(_01647_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2464),
    .D(_01648_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2465),
    .D(_01649_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2466),
    .D(_01650_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2467),
    .D(_01651_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2468),
    .D(_01652_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2469),
    .D(_01653_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2470),
    .D(_01654_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2471),
    .D(_01655_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2472),
    .D(_01656_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2473),
    .D(_01657_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2474),
    .D(_01658_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2475),
    .D(_01659_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2476),
    .D(_01660_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2477),
    .D(_01661_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2478),
    .D(_01662_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2479),
    .D(_01663_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2480),
    .D(_01664_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2481),
    .D(_01665_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2482),
    .D(_01666_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2483),
    .D(_01667_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2484),
    .D(_01668_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2485),
    .D(_01669_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2486),
    .D(_01670_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2487),
    .D(_01671_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2488),
    .D(_01672_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2489),
    .D(_01673_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2490),
    .D(_01674_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2491),
    .D(_01675_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2492),
    .D(_01676_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2493),
    .D(_01677_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2494),
    .D(_01678_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2495),
    .D(_01679_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2496),
    .D(_01680_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2497),
    .D(_01681_),
    .Q_N(_13408_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2498),
    .D(_01682_),
    .Q_N(_13407_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2499),
    .D(_01683_),
    .Q_N(_13406_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2500),
    .D(_01684_),
    .Q_N(_13405_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2501),
    .D(_01685_),
    .Q_N(_13404_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2502),
    .D(_01686_),
    .Q_N(_13403_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2503),
    .D(_01687_),
    .Q_N(_13402_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2504),
    .D(_01688_),
    .Q_N(_13401_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2505),
    .D(_01689_),
    .Q_N(_13400_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2506),
    .D(_01690_),
    .Q_N(_13399_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2507),
    .D(_01691_),
    .Q_N(_13398_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2508),
    .D(_01692_),
    .Q_N(_13397_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2509),
    .D(_01693_),
    .Q_N(_13396_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2510),
    .D(_01694_),
    .Q_N(_13395_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2511),
    .D(_01695_),
    .Q_N(_13394_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2512),
    .D(_01696_),
    .Q_N(_13393_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2513),
    .D(_01697_),
    .Q_N(_13392_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2514),
    .D(_01698_),
    .Q_N(_13391_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2515),
    .D(_01699_),
    .Q_N(_13390_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2516),
    .D(_01700_),
    .Q_N(_13389_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2517),
    .D(_01701_),
    .Q_N(_13388_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2518),
    .D(_01702_),
    .Q_N(_13387_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2519),
    .D(_01703_),
    .Q_N(_13386_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2520),
    .D(_01704_),
    .Q_N(_13385_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2521),
    .D(_01705_),
    .Q_N(_13384_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2522),
    .D(_01706_),
    .Q_N(_13383_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2523),
    .D(_01707_),
    .Q_N(_13382_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2524),
    .D(_01708_),
    .Q_N(_13381_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2525),
    .D(_01709_),
    .Q_N(_13380_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2526),
    .D(_01710_),
    .Q_N(_13379_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2527),
    .D(_01711_),
    .Q_N(_13378_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2528),
    .D(_01712_),
    .Q_N(_13377_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2529),
    .D(_01713_),
    .Q_N(_13376_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2530),
    .D(_01714_),
    .Q_N(_13375_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2531),
    .D(_01715_),
    .Q_N(_13374_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2532),
    .D(_01716_),
    .Q_N(_13373_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2533),
    .D(_01717_),
    .Q_N(_13372_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2534),
    .D(_01718_),
    .Q_N(_13371_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2535),
    .D(_01719_),
    .Q_N(_13370_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2536),
    .D(_01720_),
    .Q_N(_13369_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2537),
    .D(_01721_),
    .Q_N(_13368_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2538),
    .D(_01722_),
    .Q_N(_13367_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2539),
    .D(_01723_),
    .Q_N(_13366_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2540),
    .D(_01724_),
    .Q_N(_13365_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2541),
    .D(_01725_),
    .Q_N(_13364_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2542),
    .D(_01726_),
    .Q_N(_13363_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2543),
    .D(_01727_),
    .Q_N(_13362_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2544),
    .D(_01728_),
    .Q_N(_13361_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2545),
    .D(_01729_),
    .Q_N(_13360_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2546),
    .D(_01730_),
    .Q_N(_13359_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2547),
    .D(_01731_),
    .Q_N(_13358_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2548),
    .D(_01732_),
    .Q_N(_13357_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2549),
    .D(_01733_),
    .Q_N(_13356_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2550),
    .D(_01734_),
    .Q_N(_13355_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2551),
    .D(_01735_),
    .Q_N(_13354_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2552),
    .D(_01736_),
    .Q_N(_13353_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2553),
    .D(_01737_),
    .Q_N(_13352_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2554),
    .D(_01738_),
    .Q_N(_13351_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2555),
    .D(_01739_),
    .Q_N(_13350_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2556),
    .D(_01740_),
    .Q_N(_13349_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2557),
    .D(_01741_),
    .Q_N(_13348_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2558),
    .D(_01742_),
    .Q_N(_13347_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2559),
    .D(_01743_),
    .Q_N(_13346_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2560),
    .D(_01744_),
    .Q_N(_13345_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2561),
    .D(_01745_),
    .Q_N(_13344_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2562),
    .D(_01746_),
    .Q_N(_13343_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2563),
    .D(_01747_),
    .Q_N(_13342_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2564),
    .D(_01748_),
    .Q_N(_13341_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2565),
    .D(_01749_),
    .Q_N(_13340_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2566),
    .D(_01750_),
    .Q_N(_13339_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2567),
    .D(_01751_),
    .Q_N(_13338_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2568),
    .D(_01752_),
    .Q_N(_13337_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2569),
    .D(_01753_),
    .Q_N(_13336_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2570),
    .D(_01754_),
    .Q_N(_13335_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2571),
    .D(_01755_),
    .Q_N(_13334_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2572),
    .D(_01756_),
    .Q_N(_13333_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2573),
    .D(_01757_),
    .Q_N(_13332_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2574),
    .D(_01758_),
    .Q_N(_13331_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2575),
    .D(_01759_),
    .Q_N(_13330_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2576),
    .D(_01760_),
    .Q_N(_13329_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2577),
    .D(_01761_),
    .Q_N(_13328_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2578),
    .D(_01762_),
    .Q_N(_13327_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2579),
    .D(_01763_),
    .Q_N(_13326_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2580),
    .D(_01764_),
    .Q_N(_13325_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2581),
    .D(_01765_),
    .Q_N(_13324_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2582),
    .D(_01766_),
    .Q_N(_13323_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2583),
    .D(_01767_),
    .Q_N(_13322_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2584),
    .D(_01768_),
    .Q_N(_13321_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2585),
    .D(_01769_),
    .Q_N(_13320_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2586),
    .D(_01770_),
    .Q_N(_13319_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2587),
    .D(_01771_),
    .Q_N(_13318_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2588),
    .D(_01772_),
    .Q_N(_13317_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2589),
    .D(_01773_),
    .Q_N(_13316_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2590),
    .D(_01774_),
    .Q_N(_13315_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2591),
    .D(_01775_),
    .Q_N(_13314_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2592),
    .D(_01776_),
    .Q_N(_13313_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2593),
    .D(_01777_),
    .Q_N(_13312_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2594),
    .D(_01778_),
    .Q_N(_13311_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2595),
    .D(_01779_),
    .Q_N(_13310_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2596),
    .D(_01780_),
    .Q_N(_13309_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2597),
    .D(_01781_),
    .Q_N(_13308_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2598),
    .D(_01782_),
    .Q_N(_13307_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2599),
    .D(_01783_),
    .Q_N(_13306_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2600),
    .D(_01784_),
    .Q_N(_13305_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2601),
    .D(_01785_),
    .Q_N(_13304_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2602),
    .D(_01786_),
    .Q_N(_13303_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2603),
    .D(_01787_),
    .Q_N(_13302_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2604),
    .D(_01788_),
    .Q_N(_13301_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2605),
    .D(_01789_),
    .Q_N(_13300_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2606),
    .D(_01790_),
    .Q_N(_13299_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2607),
    .D(_01791_),
    .Q_N(_13298_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2608),
    .D(_01792_),
    .Q_N(_13297_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2609),
    .D(_01793_),
    .Q_N(_13296_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2610),
    .D(_01794_),
    .Q_N(_13295_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2611),
    .D(_01795_),
    .Q_N(_13294_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2612),
    .D(_01796_),
    .Q_N(_13293_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2613),
    .D(_01797_),
    .Q_N(_13292_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2614),
    .D(_01798_),
    .Q_N(_13291_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2615),
    .D(_01799_),
    .Q_N(_13290_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2616),
    .D(_01800_),
    .Q_N(_13289_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2617),
    .D(_01801_),
    .Q_N(_13288_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2618),
    .D(_01802_),
    .Q_N(_13287_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2619),
    .D(_01803_),
    .Q_N(_13286_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2620),
    .D(_01804_),
    .Q_N(_13285_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2621),
    .D(_01805_),
    .Q_N(_13284_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2622),
    .D(_01806_),
    .Q_N(_13283_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2623),
    .D(_01807_),
    .Q_N(_13282_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2624),
    .D(_01808_),
    .Q_N(_13281_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2625),
    .D(_01809_),
    .Q_N(_13280_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2626),
    .D(_01810_),
    .Q_N(_13279_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2627),
    .D(_01811_),
    .Q_N(_13278_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2628),
    .D(_01812_),
    .Q_N(_13277_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2629),
    .D(_01813_),
    .Q_N(_13276_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2630),
    .D(_01814_),
    .Q_N(_13275_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2631),
    .D(_01815_),
    .Q_N(_13274_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2632),
    .D(_01816_),
    .Q_N(_13273_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2633),
    .D(_01817_),
    .Q_N(_13272_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2634),
    .D(_01818_),
    .Q_N(_13271_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2635),
    .D(_01819_),
    .Q_N(_13270_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2636),
    .D(_01820_),
    .Q_N(_13269_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2637),
    .D(_01821_),
    .Q_N(_13268_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2638),
    .D(_01822_),
    .Q_N(_13267_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2639),
    .D(_01823_),
    .Q_N(_13266_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2640),
    .D(_01824_),
    .Q_N(_13265_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2641),
    .D(_01825_),
    .Q_N(_13264_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2642),
    .D(_01826_),
    .Q_N(_13263_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2643),
    .D(_01827_),
    .Q_N(_13262_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2644),
    .D(_01828_),
    .Q_N(_13261_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2645),
    .D(_01829_),
    .Q_N(_13260_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2646),
    .D(_01830_),
    .Q_N(_13259_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2647),
    .D(_01831_),
    .Q_N(_13258_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2648),
    .D(_01832_),
    .Q_N(_13257_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2649),
    .D(_01833_),
    .Q_N(_13256_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2650),
    .D(_01834_),
    .Q_N(_13255_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2651),
    .D(_01835_),
    .Q_N(_13254_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2652),
    .D(_01836_),
    .Q_N(_13253_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2653),
    .D(_01837_),
    .Q_N(_13252_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2654),
    .D(_01838_),
    .Q_N(_13251_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2655),
    .D(_01839_),
    .Q_N(_13250_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2656),
    .D(_01840_),
    .Q_N(_13249_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2657),
    .D(_01841_),
    .Q_N(_13248_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2658),
    .D(_01842_),
    .Q_N(_13247_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2659),
    .D(_01843_),
    .Q_N(_13246_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2660),
    .D(_01844_),
    .Q_N(_13245_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2661),
    .D(_01845_),
    .Q_N(_13244_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2662),
    .D(_01846_),
    .Q_N(_13243_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2663),
    .D(_01847_),
    .Q_N(_13242_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2664),
    .D(_01848_),
    .Q_N(_13241_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2665),
    .D(_01849_),
    .Q_N(_13240_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2666),
    .D(_01850_),
    .Q_N(_13239_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2667),
    .D(_01851_),
    .Q_N(_13238_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2668),
    .D(_01852_),
    .Q_N(_13237_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2669),
    .D(_01853_),
    .Q_N(_13236_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2670),
    .D(_01854_),
    .Q_N(_13235_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2671),
    .D(_01855_),
    .Q_N(_13234_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2672),
    .D(_01856_),
    .Q_N(_13233_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2673),
    .D(_01857_),
    .Q_N(_13232_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2674),
    .D(_01858_),
    .Q_N(_13231_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2675),
    .D(_01859_),
    .Q_N(_13230_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2676),
    .D(_01860_),
    .Q_N(_13229_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2677),
    .D(_01861_),
    .Q_N(_13228_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2678),
    .D(_01862_),
    .Q_N(_13227_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2679),
    .D(_01863_),
    .Q_N(_13226_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2680),
    .D(_01864_),
    .Q_N(_13225_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2681),
    .D(_01865_),
    .Q_N(_13224_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2682),
    .D(_01866_),
    .Q_N(_13223_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2683),
    .D(_01867_),
    .Q_N(_13222_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2684),
    .D(_01868_),
    .Q_N(_13221_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2685),
    .D(_01869_),
    .Q_N(_13220_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2686),
    .D(_01870_),
    .Q_N(_13219_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2687),
    .D(_01871_),
    .Q_N(_13218_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2688),
    .D(_01872_),
    .Q_N(_13217_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2689),
    .D(_01873_),
    .Q_N(_13216_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2690),
    .D(_01874_),
    .Q_N(_13215_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2691),
    .D(_01875_),
    .Q_N(_13214_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2692),
    .D(_01876_),
    .Q_N(_13213_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2693),
    .D(_01877_),
    .Q_N(_13212_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2694),
    .D(_01878_),
    .Q_N(_13211_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2695),
    .D(_01879_),
    .Q_N(_13210_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2696),
    .D(_01880_),
    .Q_N(_13209_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2697),
    .D(_01881_),
    .Q_N(_13208_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2698),
    .D(_01882_),
    .Q_N(_13207_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2699),
    .D(_01883_),
    .Q_N(_13206_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2700),
    .D(_01884_),
    .Q_N(_13205_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2701),
    .D(_01885_),
    .Q_N(_13204_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2702),
    .D(_01886_),
    .Q_N(_13203_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2703),
    .D(_01887_),
    .Q_N(_13202_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2704),
    .D(_01888_),
    .Q_N(_13201_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2705),
    .D(_01889_),
    .Q_N(_13200_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2706),
    .D(_01890_),
    .Q_N(_13199_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2707),
    .D(_01891_),
    .Q_N(_13198_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2708),
    .D(_01892_),
    .Q_N(_13197_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2709),
    .D(_01893_),
    .Q_N(_13196_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2710),
    .D(_01894_),
    .Q_N(_13195_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2711),
    .D(_01895_),
    .Q_N(_13194_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2712),
    .D(_01896_),
    .Q_N(_13193_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2713),
    .D(_01897_),
    .Q_N(_13192_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2714),
    .D(_01898_),
    .Q_N(_13191_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2715),
    .D(_01899_),
    .Q_N(_13190_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2716),
    .D(_01900_),
    .Q_N(_13189_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2717),
    .D(_01901_),
    .Q_N(_13188_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2718),
    .D(_01902_),
    .Q_N(_13187_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2719),
    .D(_01903_),
    .Q_N(_13186_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2720),
    .D(_01904_),
    .Q_N(_13185_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2721),
    .D(_01905_),
    .Q_N(_13184_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2722),
    .D(_01906_),
    .Q_N(_13183_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2723),
    .D(_01907_),
    .Q_N(_13182_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2724),
    .D(_01908_),
    .Q_N(_13181_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2725),
    .D(_01909_),
    .Q_N(_13180_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2726),
    .D(_01910_),
    .Q_N(_13179_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2727),
    .D(_01911_),
    .Q_N(_13178_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2728),
    .D(_01912_),
    .Q_N(_13177_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2729),
    .D(_01913_),
    .Q_N(_13176_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2730),
    .D(_01914_),
    .Q_N(_13175_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2731),
    .D(_01915_),
    .Q_N(_13174_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2732),
    .D(_01916_),
    .Q_N(_13173_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2733),
    .D(_01917_),
    .Q_N(_13172_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2734),
    .D(_01918_),
    .Q_N(_13171_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2735),
    .D(_01919_),
    .Q_N(_13170_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2736),
    .D(_01920_),
    .Q_N(_13169_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2737),
    .D(_01921_),
    .Q_N(_13168_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2738),
    .D(_01922_),
    .Q_N(_13167_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2739),
    .D(_01923_),
    .Q_N(_13166_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2740),
    .D(_01924_),
    .Q_N(_13165_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2741),
    .D(_01925_),
    .Q_N(_13164_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2742),
    .D(_01926_),
    .Q_N(_13163_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2743),
    .D(_01927_),
    .Q_N(_13162_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2744),
    .D(_01928_),
    .Q_N(_13161_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2745),
    .D(_01929_),
    .Q_N(_13160_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2746),
    .D(_01930_),
    .Q_N(_13159_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2747),
    .D(_01931_),
    .Q_N(_13158_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2748),
    .D(_01932_),
    .Q_N(_13157_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2749),
    .D(_01933_),
    .Q_N(_13156_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2750),
    .D(_01934_),
    .Q_N(_13155_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2751),
    .D(_01935_),
    .Q_N(_13154_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2752),
    .D(_01936_),
    .Q_N(_13153_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2753),
    .D(_01937_),
    .Q_N(_13152_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2754),
    .D(_01938_),
    .Q_N(_13151_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2755),
    .D(_01939_),
    .Q_N(_13150_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2756),
    .D(_01940_),
    .Q_N(_13149_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2757),
    .D(_01941_),
    .Q_N(_13148_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2758),
    .D(_01942_),
    .Q_N(_13147_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2759),
    .D(_01943_),
    .Q_N(_13146_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2760),
    .D(_01944_),
    .Q_N(_13145_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2761),
    .D(_01945_),
    .Q_N(_13144_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2762),
    .D(_01946_),
    .Q_N(_13143_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2763),
    .D(_01947_),
    .Q_N(_13142_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2764),
    .D(_01948_),
    .Q_N(_13141_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2765),
    .D(_01949_),
    .Q_N(_13140_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2766),
    .D(_01950_),
    .Q_N(_13139_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2767),
    .D(_01951_),
    .Q_N(_13138_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2768),
    .D(_01952_),
    .Q_N(_13137_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2769),
    .D(_01953_),
    .Q_N(_13136_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2770),
    .D(_01954_),
    .Q_N(_13135_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2771),
    .D(_01955_),
    .Q_N(_13134_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2772),
    .D(_01956_),
    .Q_N(_13133_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2773),
    .D(_01957_),
    .Q_N(_13132_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2774),
    .D(_01958_),
    .Q_N(_13131_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2775),
    .D(_01959_),
    .Q_N(_13130_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2776),
    .D(_01960_),
    .Q_N(_13129_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2777),
    .D(_01961_),
    .Q_N(_13128_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2778),
    .D(_01962_),
    .Q_N(_13127_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2779),
    .D(_01963_),
    .Q_N(_13126_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2780),
    .D(_01964_),
    .Q_N(_13125_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2781),
    .D(_01965_),
    .Q_N(_13124_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2782),
    .D(_01966_),
    .Q_N(_13123_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2783),
    .D(_01967_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2784),
    .D(_01968_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2785),
    .D(_01969_),
    .Q_N(_00119_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2786),
    .D(_01970_),
    .Q_N(_13122_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2787),
    .D(_01971_),
    .Q_N(_00138_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2788),
    .D(_01972_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2789),
    .D(_01973_),
    .Q_N(_00162_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2790),
    .D(_01974_),
    .Q_N(_13121_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2791),
    .D(_01975_),
    .Q_N(_13120_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2792),
    .D(_01976_),
    .Q_N(_00187_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2793),
    .D(_01977_),
    .Q_N(_13119_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2794),
    .D(_01978_),
    .Q_N(_13118_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2795),
    .D(_01979_),
    .Q_N(_13117_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2796),
    .D(_01980_),
    .Q_N(_00186_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2797),
    .D(_01981_),
    .Q_N(_13116_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2798),
    .D(_01982_),
    .Q_N(_13115_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2799),
    .D(_01983_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2800),
    .D(_01984_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2801),
    .D(_01985_),
    .Q_N(_00116_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2802),
    .D(_01986_),
    .Q_N(_13114_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2803),
    .D(_01987_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2804),
    .D(_01988_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2805),
    .D(_01989_),
    .Q_N(_00158_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2806),
    .D(_01990_),
    .Q_N(_13113_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2807),
    .D(_01991_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2808),
    .D(_01992_),
    .Q_N(_00149_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2809),
    .D(_01993_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2810),
    .D(_01994_),
    .Q_N(_13112_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2811),
    .D(_01995_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2812),
    .D(_01996_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2813),
    .D(_01997_),
    .Q_N(_00118_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2814),
    .D(_01998_),
    .Q_N(_13111_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2815),
    .D(_01999_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2816),
    .D(_02000_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2817),
    .D(_02001_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2818),
    .D(_02002_),
    .Q_N(_13110_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2819),
    .D(_02003_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2820),
    .D(_02004_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2821),
    .D(_02005_),
    .Q_N(_00117_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2822),
    .D(_02006_),
    .Q_N(_13109_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2823),
    .D(_02007_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2824),
    .D(_02008_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2825),
    .D(_02009_),
    .Q_N(_00159_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2826),
    .D(_02010_),
    .Q_N(_13108_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2827),
    .D(_02011_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net2828),
    .D(_02012_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2829),
    .D(_02013_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2830),
    .D(_02014_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2831),
    .D(_02015_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2832),
    .D(_02016_),
    .Q_N(_00213_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2833),
    .D(_02017_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2834),
    .D(_02018_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2835),
    .D(_02019_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2836),
    .D(_02020_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2837),
    .D(_02021_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2838),
    .D(_02022_),
    .Q_N(_00216_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2839),
    .D(_02023_),
    .Q_N(_00218_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2840),
    .D(_02024_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2841),
    .D(_02025_),
    .Q_N(_00220_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2842),
    .D(_02026_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2843),
    .D(_02027_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2844),
    .D(_02028_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2845),
    .D(_02029_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2846),
    .D(_02030_),
    .Q_N(_00177_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2847),
    .D(_02031_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2848),
    .D(_02032_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2849),
    .D(_02033_),
    .Q_N(_00214_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2850),
    .D(_02034_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2851),
    .D(_02035_),
    .Q_N(_00215_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2852),
    .D(_02036_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2853),
    .D(_02037_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2854),
    .D(_02038_),
    .Q_N(_00217_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2855),
    .D(_02039_),
    .Q_N(_00219_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2856),
    .D(_02040_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2857),
    .D(_02041_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2858),
    .D(_02042_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2859),
    .D(_02043_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2860),
    .D(_02044_),
    .Q_N(_00176_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2861),
    .D(_02045_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2862),
    .D(_02046_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2863),
    .D(_02047_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2864),
    .D(_02048_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2865),
    .D(_02049_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2866),
    .D(_02050_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2867),
    .D(_02051_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2868),
    .D(_02052_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2869),
    .D(_02053_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2870),
    .D(_02054_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2871),
    .D(_02055_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2872),
    .D(_02056_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2873),
    .D(_02057_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2874),
    .D(_02058_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2875),
    .D(_02059_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2876),
    .D(_02060_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2877),
    .D(_02061_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2878),
    .D(_02062_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2879),
    .D(_02063_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2880),
    .D(_02064_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2881),
    .D(_02065_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2882),
    .D(_02066_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2883),
    .D(_02067_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2884),
    .D(_02068_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2885),
    .D(_02069_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2886),
    .D(_02070_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2887),
    .D(_02071_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2888),
    .D(_02072_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2889),
    .D(_02073_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2890),
    .D(_02074_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2891),
    .D(_02075_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2892),
    .D(_02076_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2893),
    .D(_02077_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2894),
    .D(_02078_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2895),
    .D(_02079_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2896),
    .D(_02080_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2897),
    .D(_02081_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2898),
    .D(_02082_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2899),
    .D(_02083_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2900),
    .D(_02084_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2901),
    .D(_02085_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2902),
    .D(_02086_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2903),
    .D(_02087_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2904),
    .D(_02088_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2905),
    .D(_02089_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2906),
    .D(_02090_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2907),
    .D(_02091_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2908),
    .D(_02092_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2909),
    .D(_02093_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2910),
    .D(_02094_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2911),
    .D(_02095_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2912),
    .D(_02096_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2913),
    .D(_02097_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2914),
    .D(_02098_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2915),
    .D(_02099_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2916),
    .D(_02100_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2917),
    .D(_02101_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2918),
    .D(_02102_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2919),
    .D(_02103_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2920),
    .D(_02104_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2921),
    .D(_02105_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2922),
    .D(_02106_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2923),
    .D(_02107_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2924),
    .D(_02108_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2925),
    .D(_02109_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2926),
    .D(_02110_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2927),
    .D(_02111_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2928),
    .D(_02112_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2929),
    .D(_02113_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2930),
    .D(_02114_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2931),
    .D(_02115_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2932),
    .D(_02116_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2933),
    .D(_02117_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2934),
    .D(_02118_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2935),
    .D(_02119_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2936),
    .D(_02120_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2937),
    .D(_02121_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2938),
    .D(_02122_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2939),
    .D(_02123_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2940),
    .D(_02124_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2941),
    .D(_02125_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2942),
    .D(_02126_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2943),
    .D(_02127_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2944),
    .D(_02128_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2945),
    .D(_02129_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2946),
    .D(_02130_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2947),
    .D(_02131_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2948),
    .D(_02132_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2949),
    .D(_02133_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2950),
    .D(_02134_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2951),
    .D(_02135_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2952),
    .D(_02136_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2953),
    .D(_02137_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2954),
    .D(_02138_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2955),
    .D(_02139_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2956),
    .D(_02140_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2957),
    .D(_02141_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2958),
    .D(_02142_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2959),
    .D(_02143_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2960),
    .D(_02144_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2961),
    .D(_02145_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2962),
    .D(_02146_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2963),
    .D(_02147_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2964),
    .D(_02148_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2965),
    .D(_02149_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2966),
    .D(_02150_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2967),
    .D(_02151_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2968),
    .D(_02152_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2969),
    .D(_02153_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2970),
    .D(_02154_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2971),
    .D(_02155_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2972),
    .D(_02156_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2973),
    .D(_02157_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2974),
    .D(_02158_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2975),
    .D(_02159_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2976),
    .D(_02160_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2977),
    .D(_02161_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2978),
    .D(_02162_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2979),
    .D(_02163_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2980),
    .D(_02164_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2981),
    .D(_02165_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2982),
    .D(_02166_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2983),
    .D(_02167_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2984),
    .D(_02168_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2985),
    .D(_02169_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2986),
    .D(_02170_),
    .Q_N(_12976_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2987),
    .D(_02171_),
    .Q_N(_12975_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2988),
    .D(_02172_),
    .Q_N(_12974_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2989),
    .D(_02173_),
    .Q_N(_12973_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2990),
    .D(_02174_),
    .Q_N(_12972_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2991),
    .D(_02175_),
    .Q_N(_12971_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2992),
    .D(_02176_),
    .Q_N(_12970_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2993),
    .D(_02177_),
    .Q_N(_12969_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2994),
    .D(_02178_),
    .Q_N(_12968_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2995),
    .D(_02179_),
    .Q_N(_12967_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2996),
    .D(_02180_),
    .Q_N(_12966_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2997),
    .D(_02181_),
    .Q_N(_12965_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2998),
    .D(_02182_),
    .Q_N(_12964_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2999),
    .D(_02183_),
    .Q_N(_12963_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3000),
    .D(_02184_),
    .Q_N(_12962_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3001),
    .D(_02185_),
    .Q_N(_12961_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3002),
    .D(_02186_),
    .Q_N(_12960_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3003),
    .D(_02187_),
    .Q_N(_12959_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3004),
    .D(_02188_),
    .Q_N(_12958_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3005),
    .D(_02189_),
    .Q_N(_12957_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3006),
    .D(_02190_),
    .Q_N(_12956_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3007),
    .D(_02191_),
    .Q_N(_12955_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3008),
    .D(_02192_),
    .Q_N(_12954_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3009),
    .D(_02193_),
    .Q_N(_12953_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3010),
    .D(_02194_),
    .Q_N(_12952_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3011),
    .D(_02195_),
    .Q_N(_12951_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3012),
    .D(_02196_),
    .Q_N(_12950_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3013),
    .D(_02197_),
    .Q_N(_12949_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3014),
    .D(_02198_),
    .Q_N(_12948_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3015),
    .D(_02199_),
    .Q_N(_12947_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3016),
    .D(_02200_),
    .Q_N(_12946_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3017),
    .D(_02201_),
    .Q_N(_12945_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3018),
    .D(_02202_),
    .Q_N(_12944_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3019),
    .D(_02203_),
    .Q_N(_12943_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3020),
    .D(_02204_),
    .Q_N(_12942_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3021),
    .D(_02205_),
    .Q_N(_12941_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3022),
    .D(_02206_),
    .Q_N(_12940_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3023),
    .D(_02207_),
    .Q_N(_12939_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3024),
    .D(_02208_),
    .Q_N(_12938_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3025),
    .D(_02209_),
    .Q_N(_12937_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3026),
    .D(_02210_),
    .Q_N(_12936_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3027),
    .D(_02211_),
    .Q_N(_12935_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3028),
    .D(_02212_),
    .Q_N(_12934_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3029),
    .D(_02213_),
    .Q_N(_12933_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3030),
    .D(_02214_),
    .Q_N(_12932_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3031),
    .D(_02215_),
    .Q_N(_12931_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3032),
    .D(_02216_),
    .Q_N(_12930_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3033),
    .D(_02217_),
    .Q_N(_12929_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3034),
    .D(_02218_),
    .Q_N(_12928_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3035),
    .D(_02219_),
    .Q_N(_12927_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3036),
    .D(_02220_),
    .Q_N(_12926_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3037),
    .D(_02221_),
    .Q_N(_12925_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3038),
    .D(_02222_),
    .Q_N(_12924_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3039),
    .D(_02223_),
    .Q_N(_12923_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3040),
    .D(_02224_),
    .Q_N(_12922_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net3041),
    .D(_02225_),
    .Q_N(_12921_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3042),
    .D(_02226_),
    .Q_N(_12920_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net3043),
    .D(_02227_),
    .Q_N(_12919_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net3044),
    .D(_02228_),
    .Q_N(_12918_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3045),
    .D(_02229_),
    .Q_N(_12917_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3046),
    .D(_02230_),
    .Q_N(_12916_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3047),
    .D(_02231_),
    .Q_N(_12915_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3048),
    .D(_02232_),
    .Q_N(_12914_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3049),
    .D(_02233_),
    .Q_N(_12913_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3050),
    .D(_02234_),
    .Q_N(_12912_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3051),
    .D(_02235_),
    .Q_N(_12911_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3052),
    .D(_02236_),
    .Q_N(_12910_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3053),
    .D(_02237_),
    .Q_N(_12909_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3054),
    .D(_02238_),
    .Q_N(_12908_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3055),
    .D(_02239_),
    .Q_N(_12907_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3056),
    .D(_02240_),
    .Q_N(_12906_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3057),
    .D(_02241_),
    .Q_N(_12905_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3058),
    .D(_02242_),
    .Q_N(_12904_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3059),
    .D(_02243_),
    .Q_N(_12903_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3060),
    .D(_02244_),
    .Q_N(_12902_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3061),
    .D(_02245_),
    .Q_N(_12901_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net3062),
    .D(_02246_),
    .Q_N(_12900_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3063),
    .D(_02247_),
    .Q_N(_12899_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3064),
    .D(_02248_),
    .Q_N(_12898_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3065),
    .D(_02249_),
    .Q_N(_12897_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3066),
    .D(_02250_),
    .Q_N(_12896_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3067),
    .D(_02251_),
    .Q_N(_12895_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3068),
    .D(_02252_),
    .Q_N(_12894_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3069),
    .D(_02253_),
    .Q_N(_12893_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net3070),
    .D(_02254_),
    .Q_N(_12892_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3071),
    .D(_02255_),
    .Q_N(_12891_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3072),
    .D(_02256_),
    .Q_N(_12890_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3073),
    .D(_02257_),
    .Q_N(_12889_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3074),
    .D(_02258_),
    .Q_N(_12888_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net3075),
    .D(_02259_),
    .Q_N(_12887_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3076),
    .D(_02260_),
    .Q_N(_12886_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3077),
    .D(_02261_),
    .Q_N(_12885_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3078),
    .D(_02262_),
    .Q_N(_12884_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3079),
    .D(_02263_),
    .Q_N(_12883_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3080),
    .D(_02264_),
    .Q_N(_12882_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3081),
    .D(_02265_),
    .Q_N(_12881_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3082),
    .D(_02266_),
    .Q_N(_12880_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3083),
    .D(_02267_),
    .Q_N(_12879_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3084),
    .D(_02268_),
    .Q_N(_12878_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3085),
    .D(_02269_),
    .Q_N(_00316_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net3086),
    .D(_02270_),
    .Q_N(_12877_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net3087),
    .D(_02271_),
    .Q_N(_00254_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3088),
    .D(_02272_),
    .Q_N(_12876_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3089),
    .D(_02273_),
    .Q_N(_12875_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3090),
    .D(_02274_),
    .Q_N(_12874_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3091),
    .D(_02275_),
    .Q_N(_12873_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3092),
    .D(_02276_),
    .Q_N(_12872_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3093),
    .D(_02277_),
    .Q_N(_12871_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3094),
    .D(_02278_),
    .Q_N(_12870_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3095),
    .D(_02279_),
    .Q_N(_12869_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3096),
    .D(_02280_),
    .Q_N(_12868_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3097),
    .D(_02281_),
    .Q_N(_12867_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3098),
    .D(_02282_),
    .Q_N(_12866_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3099),
    .D(_02283_),
    .Q_N(_12865_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3100),
    .D(_02284_),
    .Q_N(_12864_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3101),
    .D(_02285_),
    .Q_N(_12863_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3102),
    .D(_02286_),
    .Q_N(_12862_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3103),
    .D(_02287_),
    .Q_N(_12861_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3104),
    .D(_02288_),
    .Q_N(_12860_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3105),
    .D(_02289_),
    .Q_N(_12859_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3106),
    .D(_02290_),
    .Q_N(_12858_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3107),
    .D(_02291_),
    .Q_N(_12857_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3108),
    .D(_02292_),
    .Q_N(_12856_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3109),
    .D(_02293_),
    .Q_N(_12855_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net3110),
    .D(_02294_),
    .Q_N(_12854_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net3111),
    .D(_02295_),
    .Q_N(_12853_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net3112),
    .D(_02296_),
    .Q_N(_12852_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3113),
    .D(_02297_),
    .Q_N(_12851_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3114),
    .D(_02298_),
    .Q_N(_12850_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3115),
    .D(_02299_),
    .Q_N(_12849_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3116),
    .D(_02300_),
    .Q_N(_12848_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3117),
    .D(_02301_),
    .Q_N(_12847_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3118),
    .D(_02302_),
    .Q_N(_12846_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3119),
    .D(_02303_),
    .Q_N(_12845_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3120),
    .D(_02304_),
    .Q_N(_12844_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3121),
    .D(_02305_),
    .Q_N(_12843_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3122),
    .D(_02306_),
    .Q_N(_12842_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3123),
    .D(_02307_),
    .Q_N(_12841_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3124),
    .D(_02308_),
    .Q_N(_12840_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3125),
    .D(_02309_),
    .Q_N(_12839_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3126),
    .D(_02310_),
    .Q_N(_12838_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3127),
    .D(_02311_),
    .Q_N(_12837_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net3128),
    .D(_02312_),
    .Q_N(_12836_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net3129),
    .D(_02313_),
    .Q_N(_12835_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3130),
    .D(_02314_),
    .Q_N(_12834_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3131),
    .D(_02315_),
    .Q_N(_12833_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3132),
    .D(_02316_),
    .Q_N(_12832_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3133),
    .D(_02317_),
    .Q_N(_12831_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3134),
    .D(_02318_),
    .Q_N(_12830_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net3135),
    .D(_02319_),
    .Q_N(_12829_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3136),
    .D(_02320_),
    .Q_N(_12828_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3137),
    .D(_02321_),
    .Q_N(_12827_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3138),
    .D(_02322_),
    .Q_N(_12826_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3139),
    .D(_02323_),
    .Q_N(_12825_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3140),
    .D(_02324_),
    .Q_N(_12824_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3141),
    .D(_02325_),
    .Q_N(_12823_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3142),
    .D(_02326_),
    .Q_N(_12822_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3143),
    .D(_02327_),
    .Q_N(_12821_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net3144),
    .D(_02328_),
    .Q_N(_12820_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3145),
    .D(_02329_),
    .Q_N(_12819_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3146),
    .D(_02330_),
    .Q_N(_12818_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net3147),
    .D(_02331_),
    .Q_N(_12817_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3148),
    .D(_02332_),
    .Q_N(_12816_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3149),
    .D(_02333_),
    .Q_N(_12815_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3150),
    .D(_02334_),
    .Q_N(_12814_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3151),
    .D(_02335_),
    .Q_N(_12813_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3152),
    .D(_02336_),
    .Q_N(_12812_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3153),
    .D(_02337_),
    .Q_N(_12811_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net3154),
    .D(_02338_),
    .Q_N(_12810_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3155),
    .D(_02339_),
    .Q_N(_12809_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3156),
    .D(_02340_),
    .Q_N(_12808_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3157),
    .D(_02341_),
    .Q_N(_12807_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3158),
    .D(_02342_),
    .Q_N(_12806_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3159),
    .D(_02343_),
    .Q_N(_12805_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3160),
    .D(_02344_),
    .Q_N(_12804_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3161),
    .D(_02345_),
    .Q_N(_12803_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3162),
    .D(_02346_),
    .Q_N(_12802_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3163),
    .D(_02347_),
    .Q_N(_12801_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3164),
    .D(_02348_),
    .Q_N(_12800_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3165),
    .D(_02349_),
    .Q_N(_12799_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3166),
    .D(_02350_),
    .Q_N(_12798_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3167),
    .D(_02351_),
    .Q_N(_12797_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net3168),
    .D(_02352_),
    .Q_N(_12796_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net3169),
    .D(_02353_),
    .Q_N(_12795_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3170),
    .D(_02354_),
    .Q_N(_12794_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net3171),
    .D(_02355_),
    .Q_N(_12793_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3172),
    .D(_02356_),
    .Q_N(_12792_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net3173),
    .D(_02357_),
    .Q_N(_12791_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3174),
    .D(_02358_),
    .Q_N(_12790_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3175),
    .D(_02359_),
    .Q_N(_12789_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3176),
    .D(_02360_),
    .Q_N(_12788_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3177),
    .D(_02361_),
    .Q_N(_12787_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3178),
    .D(_02362_),
    .Q_N(_12786_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3179),
    .D(_02363_),
    .Q_N(_12785_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3180),
    .D(_02364_),
    .Q_N(_12784_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3181),
    .D(_02365_),
    .Q_N(_12783_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3182),
    .D(_02366_),
    .Q_N(_12782_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3183),
    .D(_02367_),
    .Q_N(_12781_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3184),
    .D(_02368_),
    .Q_N(_12780_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3185),
    .D(_02369_),
    .Q_N(_12779_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3186),
    .D(_02370_),
    .Q_N(_12778_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3187),
    .D(_02371_),
    .Q_N(_12777_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3188),
    .D(_02372_),
    .Q_N(_12776_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3189),
    .D(_02373_),
    .Q_N(_12775_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3190),
    .D(_02374_),
    .Q_N(_12774_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3191),
    .D(_02375_),
    .Q_N(_12773_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net3192),
    .D(_02376_),
    .Q_N(_12772_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3193),
    .D(_02377_),
    .Q_N(_12771_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3194),
    .D(_02378_),
    .Q_N(_12770_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3195),
    .D(_02379_),
    .Q_N(_12769_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net3196),
    .D(_02380_),
    .Q_N(_12768_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3197),
    .D(_02381_),
    .Q_N(_12767_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3198),
    .D(_02382_),
    .Q_N(_12766_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3199),
    .D(_02383_),
    .Q_N(_12765_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3200),
    .D(_02384_),
    .Q_N(_12764_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net3201),
    .D(_02385_),
    .Q_N(_12763_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3202),
    .D(_02386_),
    .Q_N(_12762_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3203),
    .D(_02387_),
    .Q_N(_12761_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3204),
    .D(_02388_),
    .Q_N(_12760_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net3205),
    .D(_02389_),
    .Q_N(_12759_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net3206),
    .D(_02390_),
    .Q_N(_12758_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net3207),
    .D(_02391_),
    .Q_N(_12757_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3208),
    .D(_02392_),
    .Q_N(_12756_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3209),
    .D(_02393_),
    .Q_N(_12755_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3210),
    .D(_02394_),
    .Q_N(_12754_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net3211),
    .D(_02395_),
    .Q_N(_12753_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3212),
    .D(_02396_),
    .Q_N(_12752_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3213),
    .D(_02397_),
    .Q_N(_12751_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net3214),
    .D(_02398_),
    .Q_N(_12750_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3215),
    .D(_02399_),
    .Q_N(_12749_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3216),
    .D(_02400_),
    .Q_N(_12748_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net3217),
    .D(_02401_),
    .Q_N(_12747_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net3218),
    .D(_02402_),
    .Q_N(_12746_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3219),
    .D(_02403_),
    .Q_N(_12745_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3220),
    .D(_02404_),
    .Q_N(_12744_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3221),
    .D(_02405_),
    .Q_N(_12743_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3222),
    .D(_02406_),
    .Q_N(_12742_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net3223),
    .D(_02407_),
    .Q_N(_12741_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net3224),
    .D(_02408_),
    .Q_N(_12740_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3225),
    .D(_02409_),
    .Q_N(_12739_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3226),
    .D(_02410_),
    .Q_N(_12738_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3227),
    .D(_02411_),
    .Q_N(_12737_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net3228),
    .D(_02412_),
    .Q_N(_12736_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3229),
    .D(_02413_),
    .Q_N(_12735_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3230),
    .D(_02414_),
    .Q_N(_12734_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3231),
    .D(_02415_),
    .Q_N(_12733_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3232),
    .D(_02416_),
    .Q_N(_12732_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net3233),
    .D(_02417_),
    .Q_N(_12731_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net3234),
    .D(_02418_),
    .Q_N(_12730_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net3235),
    .D(_02419_),
    .Q_N(_12729_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net3236),
    .D(_02420_),
    .Q_N(_12728_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3237),
    .D(_02421_),
    .Q_N(_12727_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3238),
    .D(_02422_),
    .Q_N(_12726_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net3239),
    .D(_02423_),
    .Q_N(_12725_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3240),
    .D(_02424_),
    .Q_N(_12724_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3241),
    .D(_02425_),
    .Q_N(_12723_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3242),
    .D(_02426_),
    .Q_N(_12722_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net3243),
    .D(_02427_),
    .Q_N(_12721_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3244),
    .D(_02428_),
    .Q_N(_12720_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3245),
    .D(_02429_),
    .Q_N(_12719_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3246),
    .D(_02430_),
    .Q_N(_12718_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3247),
    .D(_02431_),
    .Q_N(_12717_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3248),
    .D(_02432_),
    .Q_N(_12716_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3249),
    .D(_02433_),
    .Q_N(_12715_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3250),
    .D(_02434_),
    .Q_N(_12714_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3251),
    .D(_02435_),
    .Q_N(_12713_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3252),
    .D(_02436_),
    .Q_N(_12712_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3253),
    .D(_02437_),
    .Q_N(_12711_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3254),
    .D(_02438_),
    .Q_N(_12710_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3255),
    .D(_02439_),
    .Q_N(_12709_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3256),
    .D(_02440_),
    .Q_N(_12708_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3257),
    .D(_02441_),
    .Q_N(_12707_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3258),
    .D(_02442_),
    .Q_N(_12706_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3259),
    .D(_02443_),
    .Q_N(_12705_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3260),
    .D(_02444_),
    .Q_N(_12704_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3261),
    .D(_02445_),
    .Q_N(_12703_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3262),
    .D(_02446_),
    .Q_N(_12702_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3263),
    .D(_02447_),
    .Q_N(_12701_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3264),
    .D(_02448_),
    .Q_N(_12700_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3265),
    .D(_02449_),
    .Q_N(_12699_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3266),
    .D(_02450_),
    .Q_N(_12698_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3267),
    .D(_02451_),
    .Q_N(_12697_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3268),
    .D(_02452_),
    .Q_N(_12696_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3269),
    .D(_02453_),
    .Q_N(_12695_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3270),
    .D(_02454_),
    .Q_N(_12694_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3271),
    .D(_02455_),
    .Q_N(_12693_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3272),
    .D(_02456_),
    .Q_N(_12692_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3273),
    .D(_02457_),
    .Q_N(_12691_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3274),
    .D(_02458_),
    .Q_N(_12690_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3275),
    .D(_02459_),
    .Q_N(_12689_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3276),
    .D(_02460_),
    .Q_N(_12688_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3277),
    .D(_02461_),
    .Q_N(_12687_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3278),
    .D(_02462_),
    .Q_N(_12686_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3279),
    .D(_02463_),
    .Q_N(_12685_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3280),
    .D(_02464_),
    .Q_N(_14677_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3281),
    .D(_00036_),
    .Q_N(_00286_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3282),
    .D(_00037_),
    .Q_N(_14678_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3283),
    .D(_00038_),
    .Q_N(_14679_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3284),
    .D(_00039_),
    .Q_N(_14680_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3285),
    .D(_00040_),
    .Q_N(_14681_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3286),
    .D(_00041_),
    .Q_N(_14682_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3287),
    .D(_00042_),
    .Q_N(_12684_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3288),
    .D(_02465_),
    .Q_N(_12683_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3289),
    .D(_02466_),
    .Q_N(_12682_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3290),
    .D(_02467_),
    .Q_N(_12681_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3291),
    .D(_02468_),
    .Q_N(_14683_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3292),
    .D(_00043_),
    .Q_N(_12680_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3293),
    .D(_02469_),
    .Q_N(_12679_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3294),
    .D(_02470_),
    .Q_N(_12678_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3295),
    .D(_02471_),
    .Q_N(_12677_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3296),
    .D(_02472_),
    .Q_N(_12676_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3297),
    .D(_02473_),
    .Q_N(_12675_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3298),
    .D(_02474_),
    .Q_N(_12674_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3299),
    .D(_02475_),
    .Q_N(_12673_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3300),
    .D(_02476_),
    .Q_N(_12672_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3301),
    .D(_02477_),
    .Q_N(_12671_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3302),
    .D(_02478_),
    .Q_N(_14684_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3303),
    .D(_00044_),
    .Q_N(_12670_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3304),
    .D(_02479_),
    .Q_N(_12669_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3305),
    .D(_02480_),
    .Q_N(_14685_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3306),
    .D(_00045_),
    .Q_N(_14686_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3307),
    .D(_00046_),
    .Q_N(_14687_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3308),
    .D(_00047_),
    .Q_N(_14688_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3309),
    .D(_00048_),
    .Q_N(_14689_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3310),
    .D(_00049_),
    .Q_N(_14690_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3311),
    .D(_00050_),
    .Q_N(_14691_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3312),
    .D(_00051_),
    .Q_N(_12668_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3313),
    .D(_02481_),
    .Q_N(_12667_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3314),
    .D(_02482_),
    .Q_N(_12666_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3315),
    .D(_02483_),
    .Q_N(_12665_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net3316),
    .D(_02484_),
    .Q_N(_12664_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net3317),
    .D(_02485_),
    .Q_N(_12663_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3318),
    .D(_02486_),
    .Q_N(_12662_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3319),
    .D(_02487_),
    .Q_N(_14692_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3320),
    .D(_00055_),
    .Q_N(_00285_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3321),
    .D(_00056_),
    .Q_N(_14693_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3322),
    .D(_00057_),
    .Q_N(_14694_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3323),
    .D(_00058_),
    .Q_N(_14695_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3324),
    .D(_00059_),
    .Q_N(_14696_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3325),
    .D(_00060_),
    .Q_N(_14697_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3326),
    .D(_00061_),
    .Q_N(_14698_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3327),
    .D(_00062_),
    .Q_N(_14699_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3328),
    .D(_00063_),
    .Q_N(_14700_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3329),
    .D(_00064_),
    .Q_N(_14701_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3330),
    .D(_00065_),
    .Q_N(_14702_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3331),
    .D(_00066_),
    .Q_N(_14703_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3332),
    .D(_00067_),
    .Q_N(_14704_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3333),
    .D(_00068_),
    .Q_N(_14705_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3334),
    .D(_00069_),
    .Q_N(_14706_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3335),
    .D(_00070_),
    .Q_N(_14707_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3336),
    .D(_00071_),
    .Q_N(_14708_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3337),
    .D(_00072_),
    .Q_N(_14709_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3338),
    .D(_00073_),
    .Q_N(_14710_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3339),
    .D(_00074_),
    .Q_N(_14711_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3340),
    .D(_00075_),
    .Q_N(_14712_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3341),
    .D(_00076_),
    .Q_N(_14713_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3342),
    .D(_00077_),
    .Q_N(_14714_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3343),
    .D(_00078_),
    .Q_N(_12661_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3344),
    .D(_02488_),
    .Q_N(_12660_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3345),
    .D(_02489_),
    .Q_N(_12659_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3346),
    .D(_02490_),
    .Q_N(_12658_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3347),
    .D(_02491_),
    .Q_N(_12657_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3348),
    .D(_02492_),
    .Q_N(_12656_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3349),
    .D(_02493_),
    .Q_N(_12655_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3350),
    .D(_02494_),
    .Q_N(_12654_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3351),
    .D(_02495_),
    .Q_N(_12653_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3352),
    .D(_02496_),
    .Q_N(_12652_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3353),
    .D(_02497_),
    .Q_N(_12651_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3354),
    .D(_02498_),
    .Q_N(_12650_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3355),
    .D(_02499_),
    .Q_N(_12649_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3356),
    .D(_02500_),
    .Q_N(_12648_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3357),
    .D(_02501_),
    .Q_N(_12647_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3358),
    .D(_02502_),
    .Q_N(_12646_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3359),
    .D(_02503_),
    .Q_N(_12645_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3360),
    .D(_02504_),
    .Q_N(_12644_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3361),
    .D(_02505_),
    .Q_N(_12643_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3362),
    .D(_02506_),
    .Q_N(_12642_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3363),
    .D(_02507_),
    .Q_N(_12641_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3364),
    .D(_02508_),
    .Q_N(_12640_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3365),
    .D(_02509_),
    .Q_N(_12639_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3366),
    .D(_02510_),
    .Q_N(_12638_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3367),
    .D(_02511_),
    .Q_N(_12637_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3368),
    .D(_02512_),
    .Q_N(_00183_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3369),
    .D(_02513_),
    .Q_N(_12636_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3370),
    .D(_02514_),
    .Q_N(_00184_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3371),
    .D(_02515_),
    .Q_N(_12635_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3372),
    .D(_02516_),
    .Q_N(_00252_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3373),
    .D(_02517_),
    .Q_N(_12634_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3374),
    .D(_02518_),
    .Q_N(_12633_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3375),
    .D(_02519_),
    .Q_N(_12632_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3376),
    .D(_02520_),
    .Q_N(_12631_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3377),
    .D(_02521_),
    .Q_N(_12630_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net3378),
    .D(_02522_),
    .Q_N(_12629_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3379),
    .D(_02523_),
    .Q_N(_12628_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3380),
    .D(_02524_),
    .Q_N(_12627_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net3381),
    .D(_02525_),
    .Q_N(_12626_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3382),
    .D(_02526_),
    .Q_N(_12625_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3383),
    .D(_02527_),
    .Q_N(_12624_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3384),
    .D(_02528_),
    .Q_N(_12623_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3385),
    .D(_02529_),
    .Q_N(_12622_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3386),
    .D(_02530_),
    .Q_N(_12621_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3387),
    .D(_02531_),
    .Q_N(_12620_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3388),
    .D(_02532_),
    .Q_N(_12619_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3389),
    .D(_02533_),
    .Q_N(_12618_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3390),
    .D(_02534_),
    .Q_N(_12617_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3391),
    .D(_02535_),
    .Q_N(_12616_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3392),
    .D(_02536_),
    .Q_N(_12615_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3393),
    .D(_02537_),
    .Q_N(_12614_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3394),
    .D(_02538_),
    .Q_N(_12613_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3395),
    .D(_02539_),
    .Q_N(_12612_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3396),
    .D(_02540_),
    .Q_N(_14715_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3397),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14716_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3398),
    .D(_00021_),
    .Q_N(_00277_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3399),
    .D(_00008_),
    .Q_N(_14717_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3400),
    .D(_00022_),
    .Q_N(_14718_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3401),
    .D(_00023_),
    .Q_N(_14719_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3402),
    .D(_00009_),
    .Q_N(_14720_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3403),
    .D(_00024_),
    .Q_N(_14721_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3404),
    .D(_00010_),
    .Q_N(_14722_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3405),
    .D(_00025_),
    .Q_N(_14723_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3406),
    .D(_00026_),
    .Q_N(_14724_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3407),
    .D(_00001_),
    .Q_N(_14725_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3408),
    .D(_00027_),
    .Q_N(_14726_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3409),
    .D(_00002_),
    .Q_N(_14727_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3410),
    .D(_00028_),
    .Q_N(_14728_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3411),
    .D(_00003_),
    .Q_N(_14729_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3412),
    .D(_00004_),
    .Q_N(_14730_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3413),
    .D(_00005_),
    .Q_N(_14731_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3414),
    .D(_00006_),
    .Q_N(_00185_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3415),
    .D(_00007_),
    .Q_N(_12611_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3416),
    .D(_02541_),
    .Q_N(_12610_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3417),
    .D(_02542_),
    .Q_N(_12609_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3418),
    .D(_02543_),
    .Q_N(_12608_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3419),
    .D(_02544_),
    .Q_N(_12607_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3420),
    .D(_02545_),
    .Q_N(_12606_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3421),
    .D(_02546_),
    .Q_N(_14732_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net3422),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14733_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3423),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00253_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3424),
    .D(_02547_),
    .Q_N(_12605_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3425),
    .D(_02548_),
    .Q_N(_12604_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3426),
    .D(_02549_),
    .Q_N(_12603_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3427),
    .D(_02550_),
    .Q_N(_12602_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3428),
    .D(_02551_),
    .Q_N(_00314_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3429),
    .D(_02552_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3430),
    .D(_02553_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3431),
    .D(_02554_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3432),
    .D(_02555_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3433),
    .D(_02556_),
    .Q_N(_00133_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3434),
    .D(_02557_),
    .Q_N(_00145_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3435),
    .D(_02558_),
    .Q_N(_00157_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3436),
    .D(_02559_),
    .Q_N(_00313_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3437),
    .D(_02560_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3438),
    .D(_02561_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3439),
    .D(_02562_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3440),
    .D(_02563_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3441),
    .D(_02564_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3442),
    .D(_02565_),
    .Q_N(_00144_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3443),
    .D(_02566_),
    .Q_N(_00156_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3444),
    .D(_02567_),
    .Q_N(_12601_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3445),
    .D(_02568_),
    .Q_N(_12600_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3446),
    .D(_02569_),
    .Q_N(_12599_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3447),
    .D(_02570_),
    .Q_N(_12598_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3448),
    .D(_02571_),
    .Q_N(_12597_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3449),
    .D(_02572_),
    .Q_N(_12596_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3450),
    .D(_02573_),
    .Q_N(_12595_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3451),
    .D(_02574_),
    .Q_N(_12594_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3452),
    .D(_02575_),
    .Q_N(_12593_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3453),
    .D(_02576_),
    .Q_N(_12592_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3454),
    .D(_02577_),
    .Q_N(_12591_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3455),
    .D(_02578_),
    .Q_N(_12590_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3456),
    .D(_02579_),
    .Q_N(_12589_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3457),
    .D(_02580_),
    .Q_N(_12588_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3458),
    .D(_02581_),
    .Q_N(_12587_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3459),
    .D(_02582_),
    .Q_N(_12586_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3460),
    .D(_02583_),
    .Q_N(_12585_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3461),
    .D(_02584_),
    .Q_N(_12584_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3462),
    .D(_02585_),
    .Q_N(_12583_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3463),
    .D(_02586_),
    .Q_N(_12582_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3464),
    .D(_02587_),
    .Q_N(_12581_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3465),
    .D(_02588_),
    .Q_N(_12580_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3466),
    .D(_02589_),
    .Q_N(_12579_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3467),
    .D(_02590_),
    .Q_N(_12578_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3468),
    .D(_02591_),
    .Q_N(_12577_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3469),
    .D(_02592_),
    .Q_N(_12576_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3470),
    .D(_02593_),
    .Q_N(_00222_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3471),
    .D(_02594_),
    .Q_N(_12575_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3472),
    .D(_02595_),
    .Q_N(_00224_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3473),
    .D(_02596_),
    .Q_N(_12574_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3474),
    .D(_02597_),
    .Q_N(_12573_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3475),
    .D(_02598_),
    .Q_N(_12572_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3476),
    .D(_02599_),
    .Q_N(_12571_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3477),
    .D(_02600_),
    .Q_N(_12570_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3478),
    .D(_02601_),
    .Q_N(_12569_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3479),
    .D(_02602_),
    .Q_N(_12568_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3480),
    .D(_02603_),
    .Q_N(_12567_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3481),
    .D(_02604_),
    .Q_N(_12566_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3482),
    .D(_02605_),
    .Q_N(_12565_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3483),
    .D(_02606_),
    .Q_N(_12564_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3484),
    .D(_02607_),
    .Q_N(_12563_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3485),
    .D(_02608_),
    .Q_N(_12562_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3486),
    .D(_02609_),
    .Q_N(_12561_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3487),
    .D(_02610_),
    .Q_N(_00221_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3488),
    .D(_02611_),
    .Q_N(_12560_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3489),
    .D(_02612_),
    .Q_N(_12559_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3490),
    .D(_02613_),
    .Q_N(_00282_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3491),
    .D(_02614_),
    .Q_N(_00283_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3492),
    .D(_02615_),
    .Q_N(_14734_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3493),
    .D(_00029_),
    .Q_N(_14735_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3494),
    .D(_00030_),
    .Q_N(_00225_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3495),
    .D(_00031_),
    .Q_N(_14736_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3496),
    .D(_00032_),
    .Q_N(_14737_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3497),
    .D(_00033_),
    .Q_N(_00278_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3498),
    .D(_00034_),
    .Q_N(_14738_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3499),
    .D(_00035_),
    .Q_N(_00226_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3500),
    .D(_02616_),
    .Q_N(_12558_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3501),
    .D(_02617_),
    .Q_N(_12557_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3502),
    .D(_02618_),
    .Q_N(_12556_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3503),
    .D(_02619_),
    .Q_N(_12555_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3504),
    .D(_02620_),
    .Q_N(_12554_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3505),
    .D(_02621_),
    .Q_N(_12553_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3506),
    .D(_02622_),
    .Q_N(_12552_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3507),
    .D(_02623_),
    .Q_N(_12551_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3508),
    .D(_02624_),
    .Q_N(_00284_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3509),
    .D(_02625_),
    .Q_N(_12550_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3510),
    .D(_02626_),
    .Q_N(_12549_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3511),
    .D(_02627_),
    .Q_N(_12548_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3512),
    .D(_02628_),
    .Q_N(_12547_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3513),
    .D(_02629_),
    .Q_N(_12546_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3514),
    .D(_02630_),
    .Q_N(_12545_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3515),
    .D(_02631_),
    .Q_N(_14739_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3516),
    .D(_00079_),
    .Q_N(_00279_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3517),
    .D(_00080_),
    .Q_N(_14740_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3518),
    .D(_00081_),
    .Q_N(_14741_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3519),
    .D(_00082_),
    .Q_N(_14742_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3520),
    .D(_00083_),
    .Q_N(_14743_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3521),
    .D(_00084_),
    .Q_N(_14744_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3522),
    .D(_00085_),
    .Q_N(_14745_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3523),
    .D(_00086_),
    .Q_N(_14746_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3524),
    .D(_00087_),
    .Q_N(_14747_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3525),
    .D(_00088_),
    .Q_N(_14748_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3526),
    .D(_00089_),
    .Q_N(_14749_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3527),
    .D(_00090_),
    .Q_N(_12544_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3528),
    .D(_02632_),
    .Q_N(_12543_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3529),
    .D(_02633_),
    .Q_N(_12542_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3530),
    .D(_02634_),
    .Q_N(_12541_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3531),
    .D(_02635_),
    .Q_N(_12540_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3532),
    .D(_02636_),
    .Q_N(_12539_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3533),
    .D(_02637_),
    .Q_N(_12538_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3534),
    .D(_02638_),
    .Q_N(_12537_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3535),
    .D(_02639_),
    .Q_N(_12536_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3536),
    .D(_02640_),
    .Q_N(_12535_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3537),
    .D(_02641_),
    .Q_N(_12534_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3538),
    .D(_02642_),
    .Q_N(_12533_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3539),
    .D(_02643_),
    .Q_N(_12532_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3540),
    .D(_02644_),
    .Q_N(_12531_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3541),
    .D(_02645_),
    .Q_N(_12530_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3542),
    .D(_02646_),
    .Q_N(_12529_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3543),
    .D(_02647_),
    .Q_N(_12528_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3544),
    .D(_02648_),
    .Q_N(_12527_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3545),
    .D(_02649_),
    .Q_N(_12526_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3546),
    .D(_02650_),
    .Q_N(_12525_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3547),
    .D(_02651_),
    .Q_N(_12524_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3548),
    .D(_02652_),
    .Q_N(_12523_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3549),
    .D(_02653_),
    .Q_N(_12522_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3550),
    .D(_02654_),
    .Q_N(_12521_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3551),
    .D(_02655_),
    .Q_N(_12520_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3552),
    .D(_02656_),
    .Q_N(_12519_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3553),
    .D(_02657_),
    .Q_N(_12518_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3554),
    .D(_02658_),
    .Q_N(_12517_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3555),
    .D(_02659_),
    .Q_N(_12516_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3556),
    .D(_02660_),
    .Q_N(_12515_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3557),
    .D(_02661_),
    .Q_N(_12514_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3558),
    .D(_02662_),
    .Q_N(_12513_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3559),
    .D(_02663_),
    .Q_N(_12512_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3560),
    .D(_02664_),
    .Q_N(_12511_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3561),
    .D(_02665_),
    .Q_N(_12510_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3562),
    .D(_02666_),
    .Q_N(_14750_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3563),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12509_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3564),
    .D(_02667_),
    .Q_N(_12508_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3565),
    .D(_02668_),
    .Q_N(_12507_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3566),
    .D(_02669_),
    .Q_N(_12506_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3567),
    .D(_02670_),
    .Q_N(_12505_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3568),
    .D(_02671_),
    .Q_N(_12504_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3569),
    .D(_02672_),
    .Q_N(_12503_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3570),
    .D(_02673_),
    .Q_N(_12502_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3571),
    .D(_02674_),
    .Q_N(_12501_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3572),
    .D(_02675_),
    .Q_N(_12500_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3573),
    .D(_02676_),
    .Q_N(_12499_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3574),
    .D(_02677_),
    .Q_N(_00280_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3575),
    .D(_02678_),
    .Q_N(_12498_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3576),
    .D(_02679_),
    .Q_N(_12497_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3577),
    .D(_02680_),
    .Q_N(_12496_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3578),
    .D(_02681_),
    .Q_N(_12495_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3579),
    .D(_02682_),
    .Q_N(_12494_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3580),
    .D(_02683_),
    .Q_N(_14751_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3581),
    .D(_00000_),
    .Q_N(_12493_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_06504_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_04021_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_06889_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_03914_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03618_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_04104_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_11164_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_07668_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_04010_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_03396_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02794_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02768_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02748_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02738_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02687_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12464_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12444_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12434_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12384_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12351_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12331_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12321_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12248_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12227_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12220_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12173_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12145_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12125_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12115_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12063_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12033_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12013_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12003_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_11949_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_11915_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_11891_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_11879_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_11827_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_11766_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_11692_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_11672_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_09784_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_09773_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_09772_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_06812_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_06764_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_06119_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_04805_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04626_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_12281_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_11372_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_06130_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_06107_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_11289_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_11235_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_07644_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_06980_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_05002_),
    .X(net84));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_04967_));
 sg13g2_buf_2 fanout86 (.A(_04625_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_11257_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_11192_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_09677_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_09630_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_08624_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_06800_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_06596_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_06486_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_06485_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_06469_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_06468_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_06461_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_06460_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04836_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04624_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_03429_),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(_02950_));
 sg13g2_buf_2 fanout104 (.A(_02912_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_11256_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_11223_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09865_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_09656_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_09636_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_09086_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_08853_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_08852_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_08623_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_07884_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_07434_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_06990_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04087_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04067_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_04025_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03976_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_03064_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_09909_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_09884_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_09875_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_09864_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_09645_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_09631_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_09597_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_09571_));
 sg13g2_buf_2 fanout130 (.A(_09043_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_09026_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_08851_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_07331_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_07224_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_07183_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_07171_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_06546_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_06095_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04965_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04204_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_04082_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_04077_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_04072_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_04064_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_03975_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_03968_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_03967_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_03505_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_03464_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_02927_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_11514_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_09874_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_09813_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_09812_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_08719_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_07383_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_07360_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_07351_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_07334_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_07262_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_07192_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_07182_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_06858_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_05098_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_04964_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_04169_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_04063_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_03964_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03952_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03928_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03494_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03473_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03402_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02936_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02934_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02914_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02913_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_11497_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_11476_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_11426_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_10368_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_10116_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_09862_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_07323_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_07164_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_05602_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_04141_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04085_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_03961_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_03919_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_03529_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03498_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03489_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03400_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03029_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02938_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02920_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02917_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_11472_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_11450_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_11282_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_11273_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_11184_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_11150_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_10365_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_10269_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_10188_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_10184_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_10154_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_09698_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_09679_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_09663_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_09632_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_08784_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_07335_),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_06050_));
 sg13g2_buf_2 fanout217 (.A(_06008_),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_05939_));
 sg13g2_buf_2 fanout219 (.A(_05858_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_05835_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_04079_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03997_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_03982_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03937_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_03926_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_03915_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_03672_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_03453_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_03407_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_03403_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_03398_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_03138_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_03061_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11373_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_11272_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_11186_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11181_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11167_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_10903_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_10402_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_10230_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_09697_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_09680_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_09657_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_09646_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_09638_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_08880_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_08856_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_08830_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_08783_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_08760_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_08699_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_08620_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_06078_),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_06071_));
 sg13g2_buf_2 fanout256 (.A(_06064_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_06057_));
 sg13g2_buf_2 fanout258 (.A(_06043_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_06036_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_06029_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_06022_),
    .X(net261));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_05996_));
 sg13g2_buf_2 fanout263 (.A(_05988_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_05967_),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_05960_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_05953_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_05924_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_05913_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_05891_));
 sg13g2_buf_2 fanout270 (.A(_05883_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_05875_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_05850_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_05843_),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_05825_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_05786_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_05760_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_05745_));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_05736_));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_05715_));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_05694_));
 sg13g2_buf_1 fanout281 (.A(_04699_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_03656_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_03617_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_03025_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_02933_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_02925_),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_02896_));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_02894_));
 sg13g2_buf_2 fanout289 (.A(_11258_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_11254_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_11202_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_11193_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_10680_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_10526_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_10460_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_10065_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06363_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06356_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06340_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_06338_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_06337_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_06246_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_06245_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06085_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06015_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_05974_),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_05946_));
 sg13g2_buf_2 fanout308 (.A(_05931_),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_05905_));
 sg13g2_buf_2 fanout310 (.A(_05867_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_05822_));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_05819_));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_05814_));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_05808_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_05799_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_05796_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_05793_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_05789_));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_05772_));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_05766_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_05757_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05753_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_05748_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_05731_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_05722_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05710_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_05703_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_05700_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_05681_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_05676_));
 sg13g2_buf_2 fanout331 (.A(_12278_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_11180_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_11083_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_11055_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_11025_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_10525_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_09695_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_09235_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_08716_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_06421_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_06419_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_06418_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_06301_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_06294_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_06182_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_06181_),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_05803_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_05781_));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_05741_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_05688_));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(_05662_));
 sg13g2_buf_2 fanout352 (.A(_04718_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_12441_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_11886_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_11819_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_11759_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_11741_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_11727_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_11722_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_11708_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_11240_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_11173_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_10768_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_09554_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_09527_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_09427_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_09306_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_09285_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_09254_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_09206_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_09049_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_06400_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_06398_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_06397_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_06319_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_06317_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_06316_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_05880_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_05840_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_04940_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_04793_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_04755_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_04740_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_04638_),
    .X(net384));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(_02908_));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(_02907_));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_02902_));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(_02859_));
 sg13g2_buf_4 fanout389 (.X(net389),
    .A(_02858_));
 sg13g2_buf_2 fanout390 (.A(_02745_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_12440_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_12328_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_12122_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_12010_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_11885_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_11830_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_11750_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_11239_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_09882_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_09860_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_09395_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_09371_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_09350_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_09329_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_09048_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_08940_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_08305_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_08228_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_08196_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_08104_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_08101_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_06442_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_06440_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_06439_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_06379_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_06377_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_06376_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_06004_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_06003_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_05998_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_05921_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_05920_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_05915_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_05697_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_05667_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_04937_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_04928_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_04785_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_04762_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_04739_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_04735_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_04637_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_04593_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_04590_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_03606_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_03605_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_03604_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_03390_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_03363_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_03358_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_03355_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_03353_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_03351_),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(_02903_));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(_02899_));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_02893_));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(_02892_));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(_02889_));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(_02883_));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(_02880_));
 sg13g2_buf_2 fanout451 (.A(_02796_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_02744_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_02690_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_12439_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_12327_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_12121_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_12009_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_11884_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_11821_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_11248_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_11238_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_10197_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_09975_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_09881_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_09859_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_08425_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_08403_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_08380_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_08353_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_08276_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_08253_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_08230_),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_08157_));
 sg13g2_buf_2 fanout474 (.A(_08152_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_08121_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_08103_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_08100_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_08087_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_07669_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_06092_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_06091_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_06090_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_05776_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_05767_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_05762_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_05761_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_05726_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_05716_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_05712_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_05711_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_05653_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_04927_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_04595_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_04583_),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_04577_));
 sg13g2_buf_2 fanout496 (.A(_03667_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_03598_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_03389_),
    .X(net498));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(_03388_));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(_03385_));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(_03378_));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(_03377_));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(_03362_));
 sg13g2_buf_2 fanout504 (.A(_03359_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_03357_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_03352_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_03350_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_03348_),
    .X(net508));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(_03346_));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(_02900_));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_02890_));
 sg13g2_buf_2 fanout512 (.A(_02879_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_02743_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_12386_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_12326_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_12175_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_12065_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_12008_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_11953_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_11638_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_11241_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_11237_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_11233_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_10709_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_10645_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_10282_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_10009_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_10001_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_09880_),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_09869_));
 sg13g2_buf_2 fanout531 (.A(_09858_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_09457_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_09208_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_09175_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_09161_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_09142_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_09121_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_08947_));
 sg13g2_buf_2 fanout539 (.A(_08447_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_08438_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_08362_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_08327_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_08229_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_08155_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_08133_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_08120_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_08102_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_08099_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_05999_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_05916_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_05749_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_05695_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_04977_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_04973_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_04933_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_04838_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_04737_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_04685_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_03622_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_03607_),
    .X(net560));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_03597_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_03382_));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(_03374_));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_03368_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_03356_));
 sg13g2_buf_2 fanout566 (.A(_02878_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_02735_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_11874_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_11718_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_11675_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_11617_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_11614_),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_11613_));
 sg13g2_buf_2 fanout574 (.A(_10629_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_10543_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_10316_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_10286_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_10262_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_10091_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_10000_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_09879_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_09868_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_09737_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_09595_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_09212_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_09181_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_09178_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_09174_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_09170_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_09160_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_09154_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_09147_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_09141_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_08946_),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(_08309_));
 sg13g2_buf_2 fanout596 (.A(_08208_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_08154_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_08132_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_08127_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_07897_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_07683_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_07636_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_07610_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_07524_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_07448_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_07423_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_07406_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_07382_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_07359_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_07320_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_07287_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_07251_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_07186_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_06893_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_06570_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_05993_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_05979_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_05977_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_05910_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_05896_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_05894_),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(_05644_));
 sg13g2_buf_2 fanout623 (.A(_05631_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_04968_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_04958_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_04709_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_04701_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_04670_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_04648_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_04042_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_03613_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_03609_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_03602_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_03601_),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(_02877_));
 sg13g2_buf_2 fanout636 (.A(_02864_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_02857_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_12318_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_12217_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_12112_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_12000_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_11687_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_11612_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_11604_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_11550_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_11385_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_10733_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_10685_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_10684_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_10662_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_10634_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_10626_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_10624_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_10608_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_10547_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_10136_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_10135_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10130_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10126_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_10083_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_10049_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10028_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10020_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10012_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_09867_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_09729_),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(_09592_));
 sg13g2_buf_2 fanout668 (.A(_09430_),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_09273_));
 sg13g2_buf_8 fanout670 (.A(_09271_),
    .X(net670));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(_09268_));
 sg13g2_buf_8 fanout672 (.A(_09267_),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_09242_));
 sg13g2_buf_8 fanout674 (.A(_09241_),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_09238_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_09237_));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(_09225_));
 sg13g2_buf_8 fanout678 (.A(_09223_),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_09220_));
 sg13g2_buf_2 fanout680 (.A(_09196_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_09194_));
 sg13g2_buf_8 fanout682 (.A(_09192_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_09186_),
    .X(net683));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_09184_));
 sg13g2_buf_2 fanout685 (.A(_09169_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_09166_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_09146_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_09104_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_09100_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_09097_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_09039_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_08961_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_08945_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_08650_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_08450_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_08236_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_08210_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_08207_),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_08205_));
 sg13g2_buf_2 fanout700 (.A(_08200_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_08162_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_08126_),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(_08113_));
 sg13g2_buf_2 fanout704 (.A(_05981_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_05898_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_05669_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_04669_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_03612_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_03339_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_03305_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_02909_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_02884_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_02882_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_02868_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_02863_),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_02856_));
 sg13g2_buf_2 fanout717 (.A(_12431_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_12379_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_12376_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_12362_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_12245_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_11813_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_11809_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_11785_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_11611_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_11603_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_10687_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_10635_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_10607_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_10567_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_10560_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_10549_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_10546_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_10125_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_10120_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_10097_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_10070_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_10053_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_10044_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_10038_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_10035_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10027_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_10016_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_09866_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_09811_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_09728_),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(_09591_));
 sg13g2_buf_2 fanout748 (.A(_09444_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_09376_),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(_09315_));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(_09272_));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(_09266_));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_09224_));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(_09222_));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_09193_));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(_09191_));
 sg13g2_buf_2 fanout757 (.A(_09185_),
    .X(net757));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(_09183_));
 sg13g2_buf_2 fanout759 (.A(_09093_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_09041_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_09038_),
    .X(net761));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(_08960_));
 sg13g2_buf_2 fanout763 (.A(_08944_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_08821_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_08654_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_08385_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_08306_),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_08292_));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(_08290_));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_08282_));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(_08258_));
 sg13g2_buf_2 fanout772 (.A(_08204_),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(_08183_));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_08178_));
 sg13g2_buf_2 fanout775 (.A(_08161_),
    .X(net775));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_08112_));
 sg13g2_buf_2 fanout777 (.A(_08107_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_06770_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_06662_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_06623_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_06595_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_06273_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_06242_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_06241_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_06239_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_06237_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_06227_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_06224_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_06207_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_06203_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_06202_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_06199_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_06194_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_06189_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_06167_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_06161_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_06155_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_06142_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_05985_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_05984_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_05983_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_05982_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_05902_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_05901_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_05900_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_05899_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_05782_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_05773_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_05750_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_05732_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_05723_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_05696_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_05682_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_05664_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_05663_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_05636_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_05632_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_05592_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_05591_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_05567_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_05565_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_05363_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_04627_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_04580_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_04579_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_04578_),
    .X(net826));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(_03379_));
 sg13g2_buf_2 fanout828 (.A(_03369_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_03354_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_03347_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_03338_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_02911_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_02910_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_02888_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_02887_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_02886_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_02885_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_02881_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_02876_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_02874_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_02872_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_02870_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_02867_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_12292_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_11808_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_11783_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_11778_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_11755_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_11716_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_11627_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_11607_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_11602_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_11587_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_10606_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_10556_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_10548_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_10545_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_10122_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_10077_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_10058_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_10055_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_10037_),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(_10034_));
 sg13g2_buf_2 fanout864 (.A(_10022_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_10010_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_10003_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_09984_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_09978_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_09889_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_09827_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_09820_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_09810_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_09727_),
    .X(net873));
 sg13g2_buf_8 fanout874 (.A(_09314_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_09262_),
    .X(net875));
 sg13g2_buf_4 fanout876 (.X(net876),
    .A(_09182_));
 sg13g2_buf_2 fanout877 (.A(_09095_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_09085_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_09037_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_08964_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_08959_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_08943_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_08841_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_08722_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_08627_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_08611_),
    .X(net886));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(_08602_));
 sg13g2_buf_2 fanout888 (.A(_08462_),
    .X(net888));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(_08337_));
 sg13g2_buf_8 fanout890 (.A(_08336_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(_08291_));
 sg13g2_buf_8 fanout892 (.A(_08289_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_08279_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_08257_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_08203_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_08193_),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(_08189_));
 sg13g2_buf_8 fanout898 (.A(_08188_),
    .X(net898));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_08184_));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(_08177_));
 sg13g2_buf_8 fanout901 (.A(_08175_),
    .X(net901));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_08163_));
 sg13g2_buf_2 fanout903 (.A(_08160_),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_08111_));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_08109_));
 sg13g2_buf_2 fanout906 (.A(_08106_),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(_08074_));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(_08071_));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_08067_));
 sg13g2_buf_8 fanout910 (.A(_08066_),
    .X(net910));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(_08064_));
 sg13g2_buf_8 fanout912 (.A(_08063_),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(_08060_));
 sg13g2_buf_8 fanout914 (.A(_08057_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_07678_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_07675_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_06864_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_06860_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_06848_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_06845_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_06277_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_06276_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_06275_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_06228_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_06226_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_06204_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_06198_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_06116_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_06100_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_05790_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_05783_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_05775_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_05774_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_05742_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_05733_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_05725_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_05724_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_05704_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_05647_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_05638_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_05625_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_05564_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_04924_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_04676_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_04628_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_04570_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_04447_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_04412_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_04178_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_04096_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_03337_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_02875_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_02873_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_02871_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_02869_),
    .X(net955));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(_02866_));
 sg13g2_buf_2 fanout957 (.A(_12473_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_12469_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_12263_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_12185_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_12150_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_12090_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_11988_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_11984_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_11932_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_11923_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_11870_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_11866_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_11806_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_11803_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_11801_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_11793_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_11786_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_11780_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_11775_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_11767_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_11760_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_11751_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_11730_),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(_11729_));
 sg13g2_buf_2 fanout981 (.A(_11712_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_11695_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_11688_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_11678_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_11676_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_11665_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_11586_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_11580_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_11196_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_10555_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_10544_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_10537_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_10535_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_10200_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_10195_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_10025_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_10021_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_10014_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_10013_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_09996_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_09983_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_09977_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_09964_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_09883_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_09857_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_09846_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_09840_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_09826_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_09819_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_09733_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_09673_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_09655_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_09155_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_09149_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_09130_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_09084_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_09046_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_09036_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_09030_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_08963_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_08958_),
    .X(net1021));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(_08949_));
 sg13g2_buf_2 fanout1023 (.A(_08942_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_08763_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_08626_),
    .X(net1025));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(_08538_));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(_08531_));
 sg13g2_buf_4 fanout1028 (.X(net1028),
    .A(_08522_));
 sg13g2_buf_2 fanout1029 (.A(_08500_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_08446_),
    .X(net1030));
 sg13g2_buf_4 fanout1031 (.X(net1031),
    .A(_08288_));
 sg13g2_buf_2 fanout1032 (.A(_08176_),
    .X(net1032));
 sg13g2_buf_8 fanout1033 (.A(_08174_),
    .X(net1033));
 sg13g2_buf_1 fanout1034 (.A(_08173_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_08159_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_08110_),
    .X(net1036));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(_08108_));
 sg13g2_buf_2 fanout1038 (.A(_08092_),
    .X(net1038));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(_08082_));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(_08073_));
 sg13g2_buf_2 fanout1041 (.A(_08059_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_08054_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_08052_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_07846_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_07844_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_07842_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_07548_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_06952_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_06861_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_06846_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_06844_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_05612_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_12116_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_11908_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_11903_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_11845_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_11833_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_11810_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_11792_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_11774_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_11743_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_11728_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_11711_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_11694_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_11674_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_11648_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_11632_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_11630_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_11623_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_11370_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_10321_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_10302_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_10240_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_10231_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_10156_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_09966_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_09962_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_09833_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_09672_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_09661_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_09635_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_09604_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_09092_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_09019_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_08951_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_08921_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_08839_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_08762_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_08625_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_08592_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_08558_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_08089_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_08088_),
    .X(net1093));
 sg13g2_buf_4 fanout1094 (.X(net1094),
    .A(_08069_));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(_08058_));
 sg13g2_buf_4 fanout1096 (.X(net1096),
    .A(_08053_));
 sg13g2_tiehi _27057__1097 (.L_HI(net1097));
 sg13g2_tiehi _27058__1098 (.L_HI(net1098));
 sg13g2_tiehi _27059__1099 (.L_HI(net1099));
 sg13g2_tiehi _27060__1100 (.L_HI(net1100));
 sg13g2_tiehi _27061__1101 (.L_HI(net1101));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_rs2_inv$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.spi.r_count[0]$_SDFFE_PN0P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.spi.r_count[1]$_SDFFE_PN0P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.spi.r_count[2]$_SDFFE_PN0P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.spi.r_count[3]$_SDFFE_PN0P__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.spi.r_count[4]$_SDFFE_PN0P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.spi.r_count[5]$_SDFFE_PN0P__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.spi.r_count[6]$_SDFFE_PN0P__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.spi.r_count[7]$_SDFFE_PN0P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_SDFFE_PN0P__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_SDFFE_PN0P__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_SDFFE_PN0P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_SDFFE_PN0P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_SDFFE_PN0P__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_SDFFE_PN0P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_src[0]$_SDFFE_PN0P__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_src[1]$_SDFFE_PN0P__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_src[2]$_SDFFE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3580  (.L_HI(net3580));
 sg13g2_tiehi \r_reset$_DFF_P__3581  (.L_HI(net3581));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_311_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_272_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_263_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_40_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_84_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_78_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_79_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_250_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2 (.A(_00930_));
 sg13g2_antennanp ANTENNA_3 (.A(_00948_));
 sg13g2_antennanp ANTENNA_4 (.A(_01052_));
 sg13g2_antennanp ANTENNA_5 (.A(_01057_));
 sg13g2_antennanp ANTENNA_6 (.A(_01057_));
 sg13g2_antennanp ANTENNA_7 (.A(_01071_));
 sg13g2_antennanp ANTENNA_8 (.A(_02856_));
 sg13g2_antennanp ANTENNA_9 (.A(_02856_));
 sg13g2_antennanp ANTENNA_10 (.A(_02856_));
 sg13g2_antennanp ANTENNA_11 (.A(_02856_));
 sg13g2_antennanp ANTENNA_12 (.A(_02856_));
 sg13g2_antennanp ANTENNA_13 (.A(_02856_));
 sg13g2_antennanp ANTENNA_14 (.A(_02856_));
 sg13g2_antennanp ANTENNA_15 (.A(_02856_));
 sg13g2_antennanp ANTENNA_16 (.A(_02856_));
 sg13g2_antennanp ANTENNA_17 (.A(_02856_));
 sg13g2_antennanp ANTENNA_18 (.A(_02866_));
 sg13g2_antennanp ANTENNA_19 (.A(_02866_));
 sg13g2_antennanp ANTENNA_20 (.A(_02866_));
 sg13g2_antennanp ANTENNA_21 (.A(_02866_));
 sg13g2_antennanp ANTENNA_22 (.A(_02866_));
 sg13g2_antennanp ANTENNA_23 (.A(_02866_));
 sg13g2_antennanp ANTENNA_24 (.A(_02866_));
 sg13g2_antennanp ANTENNA_25 (.A(_02866_));
 sg13g2_antennanp ANTENNA_26 (.A(_02866_));
 sg13g2_antennanp ANTENNA_27 (.A(_02866_));
 sg13g2_antennanp ANTENNA_28 (.A(_02873_));
 sg13g2_antennanp ANTENNA_29 (.A(_02873_));
 sg13g2_antennanp ANTENNA_30 (.A(_02877_));
 sg13g2_antennanp ANTENNA_31 (.A(_02877_));
 sg13g2_antennanp ANTENNA_32 (.A(_02877_));
 sg13g2_antennanp ANTENNA_33 (.A(_02877_));
 sg13g2_antennanp ANTENNA_34 (.A(_02877_));
 sg13g2_antennanp ANTENNA_35 (.A(_02877_));
 sg13g2_antennanp ANTENNA_36 (.A(_02877_));
 sg13g2_antennanp ANTENNA_37 (.A(_02877_));
 sg13g2_antennanp ANTENNA_38 (.A(_02877_));
 sg13g2_antennanp ANTENNA_39 (.A(_03350_));
 sg13g2_antennanp ANTENNA_40 (.A(_03350_));
 sg13g2_antennanp ANTENNA_41 (.A(_03350_));
 sg13g2_antennanp ANTENNA_42 (.A(_03350_));
 sg13g2_antennanp ANTENNA_43 (.A(_03350_));
 sg13g2_antennanp ANTENNA_44 (.A(_03350_));
 sg13g2_antennanp ANTENNA_45 (.A(_03356_));
 sg13g2_antennanp ANTENNA_46 (.A(_03356_));
 sg13g2_antennanp ANTENNA_47 (.A(_03356_));
 sg13g2_antennanp ANTENNA_48 (.A(_03356_));
 sg13g2_antennanp ANTENNA_49 (.A(_03356_));
 sg13g2_antennanp ANTENNA_50 (.A(_03356_));
 sg13g2_antennanp ANTENNA_51 (.A(_03356_));
 sg13g2_antennanp ANTENNA_52 (.A(_03356_));
 sg13g2_antennanp ANTENNA_53 (.A(_03356_));
 sg13g2_antennanp ANTENNA_54 (.A(_03356_));
 sg13g2_antennanp ANTENNA_55 (.A(_03369_));
 sg13g2_antennanp ANTENNA_56 (.A(_03369_));
 sg13g2_antennanp ANTENNA_57 (.A(_03369_));
 sg13g2_antennanp ANTENNA_58 (.A(_03369_));
 sg13g2_antennanp ANTENNA_59 (.A(_03612_));
 sg13g2_antennanp ANTENNA_60 (.A(_03612_));
 sg13g2_antennanp ANTENNA_61 (.A(_03612_));
 sg13g2_antennanp ANTENNA_62 (.A(_03612_));
 sg13g2_antennanp ANTENNA_63 (.A(_03612_));
 sg13g2_antennanp ANTENNA_64 (.A(_03612_));
 sg13g2_antennanp ANTENNA_65 (.A(_03612_));
 sg13g2_antennanp ANTENNA_66 (.A(_04578_));
 sg13g2_antennanp ANTENNA_67 (.A(_04578_));
 sg13g2_antennanp ANTENNA_68 (.A(_04578_));
 sg13g2_antennanp ANTENNA_69 (.A(_04578_));
 sg13g2_antennanp ANTENNA_70 (.A(_04628_));
 sg13g2_antennanp ANTENNA_71 (.A(_04628_));
 sg13g2_antennanp ANTENNA_72 (.A(_04628_));
 sg13g2_antennanp ANTENNA_73 (.A(_04628_));
 sg13g2_antennanp ANTENNA_74 (.A(_04628_));
 sg13g2_antennanp ANTENNA_75 (.A(_04628_));
 sg13g2_antennanp ANTENNA_76 (.A(_04646_));
 sg13g2_antennanp ANTENNA_77 (.A(_04952_));
 sg13g2_antennanp ANTENNA_78 (.A(_04980_));
 sg13g2_antennanp ANTENNA_79 (.A(_05022_));
 sg13g2_antennanp ANTENNA_80 (.A(_05032_));
 sg13g2_antennanp ANTENNA_81 (.A(_05046_));
 sg13g2_antennanp ANTENNA_82 (.A(_05117_));
 sg13g2_antennanp ANTENNA_83 (.A(_05581_));
 sg13g2_antennanp ANTENNA_84 (.A(_05584_));
 sg13g2_antennanp ANTENNA_85 (.A(_05589_));
 sg13g2_antennanp ANTENNA_86 (.A(_05589_));
 sg13g2_antennanp ANTENNA_87 (.A(_05589_));
 sg13g2_antennanp ANTENNA_88 (.A(_05590_));
 sg13g2_antennanp ANTENNA_89 (.A(_05631_));
 sg13g2_antennanp ANTENNA_90 (.A(_05631_));
 sg13g2_antennanp ANTENNA_91 (.A(_05631_));
 sg13g2_antennanp ANTENNA_92 (.A(_05631_));
 sg13g2_antennanp ANTENNA_93 (.A(_05644_));
 sg13g2_antennanp ANTENNA_94 (.A(_05644_));
 sg13g2_antennanp ANTENNA_95 (.A(_05644_));
 sg13g2_antennanp ANTENNA_96 (.A(_05644_));
 sg13g2_antennanp ANTENNA_97 (.A(_05644_));
 sg13g2_antennanp ANTENNA_98 (.A(_05644_));
 sg13g2_antennanp ANTENNA_99 (.A(_05644_));
 sg13g2_antennanp ANTENNA_100 (.A(_05644_));
 sg13g2_antennanp ANTENNA_101 (.A(_05644_));
 sg13g2_antennanp ANTENNA_102 (.A(_06275_));
 sg13g2_antennanp ANTENNA_103 (.A(_06275_));
 sg13g2_antennanp ANTENNA_104 (.A(_06275_));
 sg13g2_antennanp ANTENNA_105 (.A(_07137_));
 sg13g2_antennanp ANTENNA_106 (.A(_07138_));
 sg13g2_antennanp ANTENNA_107 (.A(_07163_));
 sg13g2_antennanp ANTENNA_108 (.A(_07163_));
 sg13g2_antennanp ANTENNA_109 (.A(_07163_));
 sg13g2_antennanp ANTENNA_110 (.A(_07166_));
 sg13g2_antennanp ANTENNA_111 (.A(_07222_));
 sg13g2_antennanp ANTENNA_112 (.A(_07222_));
 sg13g2_antennanp ANTENNA_113 (.A(_07326_));
 sg13g2_antennanp ANTENNA_114 (.A(_07326_));
 sg13g2_antennanp ANTENNA_115 (.A(_07349_));
 sg13g2_antennanp ANTENNA_116 (.A(_07349_));
 sg13g2_antennanp ANTENNA_117 (.A(_07976_));
 sg13g2_antennanp ANTENNA_118 (.A(_07976_));
 sg13g2_antennanp ANTENNA_119 (.A(_08081_));
 sg13g2_antennanp ANTENNA_120 (.A(_08081_));
 sg13g2_antennanp ANTENNA_121 (.A(_08081_));
 sg13g2_antennanp ANTENNA_122 (.A(_08081_));
 sg13g2_antennanp ANTENNA_123 (.A(_08081_));
 sg13g2_antennanp ANTENNA_124 (.A(_08081_));
 sg13g2_antennanp ANTENNA_125 (.A(_08081_));
 sg13g2_antennanp ANTENNA_126 (.A(_08081_));
 sg13g2_antennanp ANTENNA_127 (.A(_08081_));
 sg13g2_antennanp ANTENNA_128 (.A(_08081_));
 sg13g2_antennanp ANTENNA_129 (.A(_08081_));
 sg13g2_antennanp ANTENNA_130 (.A(_08081_));
 sg13g2_antennanp ANTENNA_131 (.A(_08081_));
 sg13g2_antennanp ANTENNA_132 (.A(_08081_));
 sg13g2_antennanp ANTENNA_133 (.A(_08081_));
 sg13g2_antennanp ANTENNA_134 (.A(_08081_));
 sg13g2_antennanp ANTENNA_135 (.A(_08087_));
 sg13g2_antennanp ANTENNA_136 (.A(_08087_));
 sg13g2_antennanp ANTENNA_137 (.A(_08087_));
 sg13g2_antennanp ANTENNA_138 (.A(_08092_));
 sg13g2_antennanp ANTENNA_139 (.A(_08092_));
 sg13g2_antennanp ANTENNA_140 (.A(_08092_));
 sg13g2_antennanp ANTENNA_141 (.A(_08173_));
 sg13g2_antennanp ANTENNA_142 (.A(_08173_));
 sg13g2_antennanp ANTENNA_143 (.A(_08173_));
 sg13g2_antennanp ANTENNA_144 (.A(_08173_));
 sg13g2_antennanp ANTENNA_145 (.A(_08184_));
 sg13g2_antennanp ANTENNA_146 (.A(_08184_));
 sg13g2_antennanp ANTENNA_147 (.A(_08184_));
 sg13g2_antennanp ANTENNA_148 (.A(_08184_));
 sg13g2_antennanp ANTENNA_149 (.A(_08184_));
 sg13g2_antennanp ANTENNA_150 (.A(_08184_));
 sg13g2_antennanp ANTENNA_151 (.A(_08184_));
 sg13g2_antennanp ANTENNA_152 (.A(_08184_));
 sg13g2_antennanp ANTENNA_153 (.A(_08257_));
 sg13g2_antennanp ANTENNA_154 (.A(_08257_));
 sg13g2_antennanp ANTENNA_155 (.A(_08257_));
 sg13g2_antennanp ANTENNA_156 (.A(_08257_));
 sg13g2_antennanp ANTENNA_157 (.A(_08327_));
 sg13g2_antennanp ANTENNA_158 (.A(_08327_));
 sg13g2_antennanp ANTENNA_159 (.A(_08327_));
 sg13g2_antennanp ANTENNA_160 (.A(_08327_));
 sg13g2_antennanp ANTENNA_161 (.A(_08345_));
 sg13g2_antennanp ANTENNA_162 (.A(_08345_));
 sg13g2_antennanp ANTENNA_163 (.A(_08345_));
 sg13g2_antennanp ANTENNA_164 (.A(_08345_));
 sg13g2_antennanp ANTENNA_165 (.A(_08345_));
 sg13g2_antennanp ANTENNA_166 (.A(_08345_));
 sg13g2_antennanp ANTENNA_167 (.A(_08380_));
 sg13g2_antennanp ANTENNA_168 (.A(_08380_));
 sg13g2_antennanp ANTENNA_169 (.A(_08380_));
 sg13g2_antennanp ANTENNA_170 (.A(_08380_));
 sg13g2_antennanp ANTENNA_171 (.A(_08403_));
 sg13g2_antennanp ANTENNA_172 (.A(_08403_));
 sg13g2_antennanp ANTENNA_173 (.A(_08403_));
 sg13g2_antennanp ANTENNA_174 (.A(_08403_));
 sg13g2_antennanp ANTENNA_175 (.A(_08517_));
 sg13g2_antennanp ANTENNA_176 (.A(_08556_));
 sg13g2_antennanp ANTENNA_177 (.A(_08614_));
 sg13g2_antennanp ANTENNA_178 (.A(_08947_));
 sg13g2_antennanp ANTENNA_179 (.A(_08947_));
 sg13g2_antennanp ANTENNA_180 (.A(_08947_));
 sg13g2_antennanp ANTENNA_181 (.A(_08947_));
 sg13g2_antennanp ANTENNA_182 (.A(_08951_));
 sg13g2_antennanp ANTENNA_183 (.A(_08951_));
 sg13g2_antennanp ANTENNA_184 (.A(_08951_));
 sg13g2_antennanp ANTENNA_185 (.A(_08951_));
 sg13g2_antennanp ANTENNA_186 (.A(_08951_));
 sg13g2_antennanp ANTENNA_187 (.A(_08951_));
 sg13g2_antennanp ANTENNA_188 (.A(_08951_));
 sg13g2_antennanp ANTENNA_189 (.A(_08951_));
 sg13g2_antennanp ANTENNA_190 (.A(_08951_));
 sg13g2_antennanp ANTENNA_191 (.A(_08962_));
 sg13g2_antennanp ANTENNA_192 (.A(_08962_));
 sg13g2_antennanp ANTENNA_193 (.A(_08962_));
 sg13g2_antennanp ANTENNA_194 (.A(_08962_));
 sg13g2_antennanp ANTENNA_195 (.A(_08962_));
 sg13g2_antennanp ANTENNA_196 (.A(_08993_));
 sg13g2_antennanp ANTENNA_197 (.A(_09005_));
 sg13g2_antennanp ANTENNA_198 (.A(_09030_));
 sg13g2_antennanp ANTENNA_199 (.A(_09030_));
 sg13g2_antennanp ANTENNA_200 (.A(_09030_));
 sg13g2_antennanp ANTENNA_201 (.A(_09037_));
 sg13g2_antennanp ANTENNA_202 (.A(_09037_));
 sg13g2_antennanp ANTENNA_203 (.A(_09037_));
 sg13g2_antennanp ANTENNA_204 (.A(_09039_));
 sg13g2_antennanp ANTENNA_205 (.A(_09039_));
 sg13g2_antennanp ANTENNA_206 (.A(_09039_));
 sg13g2_antennanp ANTENNA_207 (.A(_09039_));
 sg13g2_antennanp ANTENNA_208 (.A(_09039_));
 sg13g2_antennanp ANTENNA_209 (.A(_09039_));
 sg13g2_antennanp ANTENNA_210 (.A(_09039_));
 sg13g2_antennanp ANTENNA_211 (.A(_09039_));
 sg13g2_antennanp ANTENNA_212 (.A(_09039_));
 sg13g2_antennanp ANTENNA_213 (.A(_09095_));
 sg13g2_antennanp ANTENNA_214 (.A(_09095_));
 sg13g2_antennanp ANTENNA_215 (.A(_09095_));
 sg13g2_antennanp ANTENNA_216 (.A(_09095_));
 sg13g2_antennanp ANTENNA_217 (.A(_09205_));
 sg13g2_antennanp ANTENNA_218 (.A(_09234_));
 sg13g2_antennanp ANTENNA_219 (.A(_09253_));
 sg13g2_antennanp ANTENNA_220 (.A(_09284_));
 sg13g2_antennanp ANTENNA_221 (.A(_09305_));
 sg13g2_antennanp ANTENNA_222 (.A(_09328_));
 sg13g2_antennanp ANTENNA_223 (.A(_09349_));
 sg13g2_antennanp ANTENNA_224 (.A(_09370_));
 sg13g2_antennanp ANTENNA_225 (.A(_09394_));
 sg13g2_antennanp ANTENNA_226 (.A(_09426_));
 sg13g2_antennanp ANTENNA_227 (.A(_09440_));
 sg13g2_antennanp ANTENNA_228 (.A(_09440_));
 sg13g2_antennanp ANTENNA_229 (.A(_09440_));
 sg13g2_antennanp ANTENNA_230 (.A(_09440_));
 sg13g2_antennanp ANTENNA_231 (.A(_09440_));
 sg13g2_antennanp ANTENNA_232 (.A(_09440_));
 sg13g2_antennanp ANTENNA_233 (.A(_09440_));
 sg13g2_antennanp ANTENNA_234 (.A(_09440_));
 sg13g2_antennanp ANTENNA_235 (.A(_09440_));
 sg13g2_antennanp ANTENNA_236 (.A(_09440_));
 sg13g2_antennanp ANTENNA_237 (.A(_09440_));
 sg13g2_antennanp ANTENNA_238 (.A(_09440_));
 sg13g2_antennanp ANTENNA_239 (.A(_09440_));
 sg13g2_antennanp ANTENNA_240 (.A(_09470_));
 sg13g2_antennanp ANTENNA_241 (.A(_09470_));
 sg13g2_antennanp ANTENNA_242 (.A(_09470_));
 sg13g2_antennanp ANTENNA_243 (.A(_09470_));
 sg13g2_antennanp ANTENNA_244 (.A(_09470_));
 sg13g2_antennanp ANTENNA_245 (.A(_09526_));
 sg13g2_antennanp ANTENNA_246 (.A(_09553_));
 sg13g2_antennanp ANTENNA_247 (.A(_09591_));
 sg13g2_antennanp ANTENNA_248 (.A(_09591_));
 sg13g2_antennanp ANTENNA_249 (.A(_09591_));
 sg13g2_antennanp ANTENNA_250 (.A(_09591_));
 sg13g2_antennanp ANTENNA_251 (.A(_09845_));
 sg13g2_antennanp ANTENNA_252 (.A(_09845_));
 sg13g2_antennanp ANTENNA_253 (.A(_09845_));
 sg13g2_antennanp ANTENNA_254 (.A(_09845_));
 sg13g2_antennanp ANTENNA_255 (.A(_09845_));
 sg13g2_antennanp ANTENNA_256 (.A(_09845_));
 sg13g2_antennanp ANTENNA_257 (.A(_09845_));
 sg13g2_antennanp ANTENNA_258 (.A(_09880_));
 sg13g2_antennanp ANTENNA_259 (.A(_09880_));
 sg13g2_antennanp ANTENNA_260 (.A(_09880_));
 sg13g2_antennanp ANTENNA_261 (.A(_09880_));
 sg13g2_antennanp ANTENNA_262 (.A(_09880_));
 sg13g2_antennanp ANTENNA_263 (.A(_09880_));
 sg13g2_antennanp ANTENNA_264 (.A(_09880_));
 sg13g2_antennanp ANTENNA_265 (.A(_09880_));
 sg13g2_antennanp ANTENNA_266 (.A(_09880_));
 sg13g2_antennanp ANTENNA_267 (.A(_09882_));
 sg13g2_antennanp ANTENNA_268 (.A(_09882_));
 sg13g2_antennanp ANTENNA_269 (.A(_09882_));
 sg13g2_antennanp ANTENNA_270 (.A(_09882_));
 sg13g2_antennanp ANTENNA_271 (.A(_09958_));
 sg13g2_antennanp ANTENNA_272 (.A(_09958_));
 sg13g2_antennanp ANTENNA_273 (.A(_09958_));
 sg13g2_antennanp ANTENNA_274 (.A(_09958_));
 sg13g2_antennanp ANTENNA_275 (.A(_09958_));
 sg13g2_antennanp ANTENNA_276 (.A(_09958_));
 sg13g2_antennanp ANTENNA_277 (.A(_09958_));
 sg13g2_antennanp ANTENNA_278 (.A(_09958_));
 sg13g2_antennanp ANTENNA_279 (.A(_09958_));
 sg13g2_antennanp ANTENNA_280 (.A(_09958_));
 sg13g2_antennanp ANTENNA_281 (.A(_09958_));
 sg13g2_antennanp ANTENNA_282 (.A(_09958_));
 sg13g2_antennanp ANTENNA_283 (.A(_09958_));
 sg13g2_antennanp ANTENNA_284 (.A(_09958_));
 sg13g2_antennanp ANTENNA_285 (.A(_09958_));
 sg13g2_antennanp ANTENNA_286 (.A(_09958_));
 sg13g2_antennanp ANTENNA_287 (.A(_09958_));
 sg13g2_antennanp ANTENNA_288 (.A(_09985_));
 sg13g2_antennanp ANTENNA_289 (.A(_09985_));
 sg13g2_antennanp ANTENNA_290 (.A(_09985_));
 sg13g2_antennanp ANTENNA_291 (.A(_09985_));
 sg13g2_antennanp ANTENNA_292 (.A(_09985_));
 sg13g2_antennanp ANTENNA_293 (.A(_09985_));
 sg13g2_antennanp ANTENNA_294 (.A(_09985_));
 sg13g2_antennanp ANTENNA_295 (.A(_09985_));
 sg13g2_antennanp ANTENNA_296 (.A(_09985_));
 sg13g2_antennanp ANTENNA_297 (.A(_09985_));
 sg13g2_antennanp ANTENNA_298 (.A(_09985_));
 sg13g2_antennanp ANTENNA_299 (.A(_09985_));
 sg13g2_antennanp ANTENNA_300 (.A(_09985_));
 sg13g2_antennanp ANTENNA_301 (.A(_09985_));
 sg13g2_antennanp ANTENNA_302 (.A(_09985_));
 sg13g2_antennanp ANTENNA_303 (.A(_09985_));
 sg13g2_antennanp ANTENNA_304 (.A(_09985_));
 sg13g2_antennanp ANTENNA_305 (.A(_09985_));
 sg13g2_antennanp ANTENNA_306 (.A(_09985_));
 sg13g2_antennanp ANTENNA_307 (.A(_09985_));
 sg13g2_antennanp ANTENNA_308 (.A(_09985_));
 sg13g2_antennanp ANTENNA_309 (.A(_09985_));
 sg13g2_antennanp ANTENNA_310 (.A(_09985_));
 sg13g2_antennanp ANTENNA_311 (.A(_09985_));
 sg13g2_antennanp ANTENNA_312 (.A(_09985_));
 sg13g2_antennanp ANTENNA_313 (.A(_09985_));
 sg13g2_antennanp ANTENNA_314 (.A(_09985_));
 sg13g2_antennanp ANTENNA_315 (.A(_10147_));
 sg13g2_antennanp ANTENNA_316 (.A(_10147_));
 sg13g2_antennanp ANTENNA_317 (.A(_10147_));
 sg13g2_antennanp ANTENNA_318 (.A(_10147_));
 sg13g2_antennanp ANTENNA_319 (.A(_10147_));
 sg13g2_antennanp ANTENNA_320 (.A(_10147_));
 sg13g2_antennanp ANTENNA_321 (.A(_10147_));
 sg13g2_antennanp ANTENNA_322 (.A(_10147_));
 sg13g2_antennanp ANTENNA_323 (.A(_10147_));
 sg13g2_antennanp ANTENNA_324 (.A(_10147_));
 sg13g2_antennanp ANTENNA_325 (.A(_10147_));
 sg13g2_antennanp ANTENNA_326 (.A(_10147_));
 sg13g2_antennanp ANTENNA_327 (.A(_10147_));
 sg13g2_antennanp ANTENNA_328 (.A(_10147_));
 sg13g2_antennanp ANTENNA_329 (.A(_10147_));
 sg13g2_antennanp ANTENNA_330 (.A(_10147_));
 sg13g2_antennanp ANTENNA_331 (.A(_10147_));
 sg13g2_antennanp ANTENNA_332 (.A(_10147_));
 sg13g2_antennanp ANTENNA_333 (.A(_10147_));
 sg13g2_antennanp ANTENNA_334 (.A(_10147_));
 sg13g2_antennanp ANTENNA_335 (.A(_10156_));
 sg13g2_antennanp ANTENNA_336 (.A(_10156_));
 sg13g2_antennanp ANTENNA_337 (.A(_10156_));
 sg13g2_antennanp ANTENNA_338 (.A(_10156_));
 sg13g2_antennanp ANTENNA_339 (.A(_10241_));
 sg13g2_antennanp ANTENNA_340 (.A(_10241_));
 sg13g2_antennanp ANTENNA_341 (.A(_10241_));
 sg13g2_antennanp ANTENNA_342 (.A(_10482_));
 sg13g2_antennanp ANTENNA_343 (.A(_10482_));
 sg13g2_antennanp ANTENNA_344 (.A(_10482_));
 sg13g2_antennanp ANTENNA_345 (.A(_10482_));
 sg13g2_antennanp ANTENNA_346 (.A(_10653_));
 sg13g2_antennanp ANTENNA_347 (.A(_10653_));
 sg13g2_antennanp ANTENNA_348 (.A(_10653_));
 sg13g2_antennanp ANTENNA_349 (.A(_10653_));
 sg13g2_antennanp ANTENNA_350 (.A(_10892_));
 sg13g2_antennanp ANTENNA_351 (.A(_10892_));
 sg13g2_antennanp ANTENNA_352 (.A(_10892_));
 sg13g2_antennanp ANTENNA_353 (.A(_10892_));
 sg13g2_antennanp ANTENNA_354 (.A(_10892_));
 sg13g2_antennanp ANTENNA_355 (.A(_10892_));
 sg13g2_antennanp ANTENNA_356 (.A(_10892_));
 sg13g2_antennanp ANTENNA_357 (.A(_10892_));
 sg13g2_antennanp ANTENNA_358 (.A(_10892_));
 sg13g2_antennanp ANTENNA_359 (.A(_11550_));
 sg13g2_antennanp ANTENNA_360 (.A(_11550_));
 sg13g2_antennanp ANTENNA_361 (.A(_11550_));
 sg13g2_antennanp ANTENNA_362 (.A(_11550_));
 sg13g2_antennanp ANTENNA_363 (.A(_11550_));
 sg13g2_antennanp ANTENNA_364 (.A(_11550_));
 sg13g2_antennanp ANTENNA_365 (.A(_11550_));
 sg13g2_antennanp ANTENNA_366 (.A(_11550_));
 sg13g2_antennanp ANTENNA_367 (.A(_11613_));
 sg13g2_antennanp ANTENNA_368 (.A(_11613_));
 sg13g2_antennanp ANTENNA_369 (.A(_11613_));
 sg13g2_antennanp ANTENNA_370 (.A(_11613_));
 sg13g2_antennanp ANTENNA_371 (.A(_11613_));
 sg13g2_antennanp ANTENNA_372 (.A(_11613_));
 sg13g2_antennanp ANTENNA_373 (.A(_11613_));
 sg13g2_antennanp ANTENNA_374 (.A(_11613_));
 sg13g2_antennanp ANTENNA_375 (.A(_11613_));
 sg13g2_antennanp ANTENNA_376 (.A(_11613_));
 sg13g2_antennanp ANTENNA_377 (.A(_11613_));
 sg13g2_antennanp ANTENNA_378 (.A(_11613_));
 sg13g2_antennanp ANTENNA_379 (.A(_11613_));
 sg13g2_antennanp ANTENNA_380 (.A(_11613_));
 sg13g2_antennanp ANTENNA_381 (.A(_11613_));
 sg13g2_antennanp ANTENNA_382 (.A(_11613_));
 sg13g2_antennanp ANTENNA_383 (.A(_11613_));
 sg13g2_antennanp ANTENNA_384 (.A(_11613_));
 sg13g2_antennanp ANTENNA_385 (.A(_11688_));
 sg13g2_antennanp ANTENNA_386 (.A(_11688_));
 sg13g2_antennanp ANTENNA_387 (.A(_11688_));
 sg13g2_antennanp ANTENNA_388 (.A(_11688_));
 sg13g2_antennanp ANTENNA_389 (.A(_11688_));
 sg13g2_antennanp ANTENNA_390 (.A(_11688_));
 sg13g2_antennanp ANTENNA_391 (.A(_11688_));
 sg13g2_antennanp ANTENNA_392 (.A(_11688_));
 sg13g2_antennanp ANTENNA_393 (.A(_11688_));
 sg13g2_antennanp ANTENNA_394 (.A(_11695_));
 sg13g2_antennanp ANTENNA_395 (.A(_11695_));
 sg13g2_antennanp ANTENNA_396 (.A(_11695_));
 sg13g2_antennanp ANTENNA_397 (.A(_11695_));
 sg13g2_antennanp ANTENNA_398 (.A(_11695_));
 sg13g2_antennanp ANTENNA_399 (.A(_11695_));
 sg13g2_antennanp ANTENNA_400 (.A(_11712_));
 sg13g2_antennanp ANTENNA_401 (.A(_11712_));
 sg13g2_antennanp ANTENNA_402 (.A(_11712_));
 sg13g2_antennanp ANTENNA_403 (.A(_11712_));
 sg13g2_antennanp ANTENNA_404 (.A(_11712_));
 sg13g2_antennanp ANTENNA_405 (.A(_11712_));
 sg13g2_antennanp ANTENNA_406 (.A(_11743_));
 sg13g2_antennanp ANTENNA_407 (.A(_11743_));
 sg13g2_antennanp ANTENNA_408 (.A(_11743_));
 sg13g2_antennanp ANTENNA_409 (.A(_11743_));
 sg13g2_antennanp ANTENNA_410 (.A(_11743_));
 sg13g2_antennanp ANTENNA_411 (.A(_11743_));
 sg13g2_antennanp ANTENNA_412 (.A(_11743_));
 sg13g2_antennanp ANTENNA_413 (.A(_11743_));
 sg13g2_antennanp ANTENNA_414 (.A(_11743_));
 sg13g2_antennanp ANTENNA_415 (.A(_11833_));
 sg13g2_antennanp ANTENNA_416 (.A(_11833_));
 sg13g2_antennanp ANTENNA_417 (.A(_11833_));
 sg13g2_antennanp ANTENNA_418 (.A(_11833_));
 sg13g2_antennanp ANTENNA_419 (.A(_11833_));
 sg13g2_antennanp ANTENNA_420 (.A(_11833_));
 sg13g2_antennanp ANTENNA_421 (.A(_11833_));
 sg13g2_antennanp ANTENNA_422 (.A(_11833_));
 sg13g2_antennanp ANTENNA_423 (.A(_11833_));
 sg13g2_antennanp ANTENNA_424 (.A(_11866_));
 sg13g2_antennanp ANTENNA_425 (.A(_11866_));
 sg13g2_antennanp ANTENNA_426 (.A(_11866_));
 sg13g2_antennanp ANTENNA_427 (.A(_11866_));
 sg13g2_antennanp ANTENNA_428 (.A(_11866_));
 sg13g2_antennanp ANTENNA_429 (.A(_11866_));
 sg13g2_antennanp ANTENNA_430 (.A(_11866_));
 sg13g2_antennanp ANTENNA_431 (.A(_11866_));
 sg13g2_antennanp ANTENNA_432 (.A(_11866_));
 sg13g2_antennanp ANTENNA_433 (.A(_11866_));
 sg13g2_antennanp ANTENNA_434 (.A(_11870_));
 sg13g2_antennanp ANTENNA_435 (.A(_11870_));
 sg13g2_antennanp ANTENNA_436 (.A(_11870_));
 sg13g2_antennanp ANTENNA_437 (.A(_11870_));
 sg13g2_antennanp ANTENNA_438 (.A(_11870_));
 sg13g2_antennanp ANTENNA_439 (.A(_11870_));
 sg13g2_antennanp ANTENNA_440 (.A(_11870_));
 sg13g2_antennanp ANTENNA_441 (.A(_11870_));
 sg13g2_antennanp ANTENNA_442 (.A(_11870_));
 sg13g2_antennanp ANTENNA_443 (.A(_12009_));
 sg13g2_antennanp ANTENNA_444 (.A(_12009_));
 sg13g2_antennanp ANTENNA_445 (.A(_12009_));
 sg13g2_antennanp ANTENNA_446 (.A(_12185_));
 sg13g2_antennanp ANTENNA_447 (.A(_12185_));
 sg13g2_antennanp ANTENNA_448 (.A(_12185_));
 sg13g2_antennanp ANTENNA_449 (.A(_12185_));
 sg13g2_antennanp ANTENNA_450 (.A(_12185_));
 sg13g2_antennanp ANTENNA_451 (.A(_12185_));
 sg13g2_antennanp ANTENNA_452 (.A(_12469_));
 sg13g2_antennanp ANTENNA_453 (.A(_12469_));
 sg13g2_antennanp ANTENNA_454 (.A(_12469_));
 sg13g2_antennanp ANTENNA_455 (.A(_12469_));
 sg13g2_antennanp ANTENNA_456 (.A(_12469_));
 sg13g2_antennanp ANTENNA_457 (.A(_12469_));
 sg13g2_antennanp ANTENNA_458 (.A(_12473_));
 sg13g2_antennanp ANTENNA_459 (.A(_12473_));
 sg13g2_antennanp ANTENNA_460 (.A(_12473_));
 sg13g2_antennanp ANTENNA_461 (.A(_12473_));
 sg13g2_antennanp ANTENNA_462 (.A(clk));
 sg13g2_antennanp ANTENNA_463 (.A(clk));
 sg13g2_antennanp ANTENNA_464 (.A(\cpu.addr[14] ));
 sg13g2_antennanp ANTENNA_465 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_466 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_467 (.A(net3));
 sg13g2_antennanp ANTENNA_468 (.A(net3));
 sg13g2_antennanp ANTENNA_469 (.A(net3));
 sg13g2_antennanp ANTENNA_470 (.A(net11));
 sg13g2_antennanp ANTENNA_471 (.A(net11));
 sg13g2_antennanp ANTENNA_472 (.A(net11));
 sg13g2_antennanp ANTENNA_473 (.A(net12));
 sg13g2_antennanp ANTENNA_474 (.A(net12));
 sg13g2_antennanp ANTENNA_475 (.A(net12));
 sg13g2_antennanp ANTENNA_476 (.A(net14));
 sg13g2_antennanp ANTENNA_477 (.A(net14));
 sg13g2_antennanp ANTENNA_478 (.A(net14));
 sg13g2_antennanp ANTENNA_479 (.A(net18));
 sg13g2_antennanp ANTENNA_480 (.A(net19));
 sg13g2_antennanp ANTENNA_481 (.A(net19));
 sg13g2_antennanp ANTENNA_482 (.A(net20));
 sg13g2_antennanp ANTENNA_483 (.A(net20));
 sg13g2_antennanp ANTENNA_484 (.A(net464));
 sg13g2_antennanp ANTENNA_485 (.A(net464));
 sg13g2_antennanp ANTENNA_486 (.A(net464));
 sg13g2_antennanp ANTENNA_487 (.A(net464));
 sg13g2_antennanp ANTENNA_488 (.A(net464));
 sg13g2_antennanp ANTENNA_489 (.A(net464));
 sg13g2_antennanp ANTENNA_490 (.A(net464));
 sg13g2_antennanp ANTENNA_491 (.A(net464));
 sg13g2_antennanp ANTENNA_492 (.A(net464));
 sg13g2_antennanp ANTENNA_493 (.A(net464));
 sg13g2_antennanp ANTENNA_494 (.A(net464));
 sg13g2_antennanp ANTENNA_495 (.A(net464));
 sg13g2_antennanp ANTENNA_496 (.A(net464));
 sg13g2_antennanp ANTENNA_497 (.A(net464));
 sg13g2_antennanp ANTENNA_498 (.A(net464));
 sg13g2_antennanp ANTENNA_499 (.A(net464));
 sg13g2_antennanp ANTENNA_500 (.A(net464));
 sg13g2_antennanp ANTENNA_501 (.A(net464));
 sg13g2_antennanp ANTENNA_502 (.A(net464));
 sg13g2_antennanp ANTENNA_503 (.A(net464));
 sg13g2_antennanp ANTENNA_504 (.A(net464));
 sg13g2_antennanp ANTENNA_505 (.A(net464));
 sg13g2_antennanp ANTENNA_506 (.A(net464));
 sg13g2_antennanp ANTENNA_507 (.A(net464));
 sg13g2_antennanp ANTENNA_508 (.A(net464));
 sg13g2_antennanp ANTENNA_509 (.A(net464));
 sg13g2_antennanp ANTENNA_510 (.A(net464));
 sg13g2_antennanp ANTENNA_511 (.A(net464));
 sg13g2_antennanp ANTENNA_512 (.A(net464));
 sg13g2_antennanp ANTENNA_513 (.A(net464));
 sg13g2_antennanp ANTENNA_514 (.A(net464));
 sg13g2_antennanp ANTENNA_515 (.A(net464));
 sg13g2_antennanp ANTENNA_516 (.A(net464));
 sg13g2_antennanp ANTENNA_517 (.A(net464));
 sg13g2_antennanp ANTENNA_518 (.A(net464));
 sg13g2_antennanp ANTENNA_519 (.A(net464));
 sg13g2_antennanp ANTENNA_520 (.A(net464));
 sg13g2_antennanp ANTENNA_521 (.A(net464));
 sg13g2_antennanp ANTENNA_522 (.A(net464));
 sg13g2_antennanp ANTENNA_523 (.A(net464));
 sg13g2_antennanp ANTENNA_524 (.A(net464));
 sg13g2_antennanp ANTENNA_525 (.A(net464));
 sg13g2_antennanp ANTENNA_526 (.A(net464));
 sg13g2_antennanp ANTENNA_527 (.A(net464));
 sg13g2_antennanp ANTENNA_528 (.A(net464));
 sg13g2_antennanp ANTENNA_529 (.A(net464));
 sg13g2_antennanp ANTENNA_530 (.A(net464));
 sg13g2_antennanp ANTENNA_531 (.A(net464));
 sg13g2_antennanp ANTENNA_532 (.A(net498));
 sg13g2_antennanp ANTENNA_533 (.A(net498));
 sg13g2_antennanp ANTENNA_534 (.A(net498));
 sg13g2_antennanp ANTENNA_535 (.A(net498));
 sg13g2_antennanp ANTENNA_536 (.A(net498));
 sg13g2_antennanp ANTENNA_537 (.A(net498));
 sg13g2_antennanp ANTENNA_538 (.A(net498));
 sg13g2_antennanp ANTENNA_539 (.A(net498));
 sg13g2_antennanp ANTENNA_540 (.A(net498));
 sg13g2_antennanp ANTENNA_541 (.A(net532));
 sg13g2_antennanp ANTENNA_542 (.A(net532));
 sg13g2_antennanp ANTENNA_543 (.A(net532));
 sg13g2_antennanp ANTENNA_544 (.A(net532));
 sg13g2_antennanp ANTENNA_545 (.A(net532));
 sg13g2_antennanp ANTENNA_546 (.A(net532));
 sg13g2_antennanp ANTENNA_547 (.A(net532));
 sg13g2_antennanp ANTENNA_548 (.A(net532));
 sg13g2_antennanp ANTENNA_549 (.A(net532));
 sg13g2_antennanp ANTENNA_550 (.A(net573));
 sg13g2_antennanp ANTENNA_551 (.A(net573));
 sg13g2_antennanp ANTENNA_552 (.A(net573));
 sg13g2_antennanp ANTENNA_553 (.A(net573));
 sg13g2_antennanp ANTENNA_554 (.A(net573));
 sg13g2_antennanp ANTENNA_555 (.A(net573));
 sg13g2_antennanp ANTENNA_556 (.A(net573));
 sg13g2_antennanp ANTENNA_557 (.A(net573));
 sg13g2_antennanp ANTENNA_558 (.A(net573));
 sg13g2_antennanp ANTENNA_559 (.A(net573));
 sg13g2_antennanp ANTENNA_560 (.A(net573));
 sg13g2_antennanp ANTENNA_561 (.A(net573));
 sg13g2_antennanp ANTENNA_562 (.A(net573));
 sg13g2_antennanp ANTENNA_563 (.A(net573));
 sg13g2_antennanp ANTENNA_564 (.A(net573));
 sg13g2_antennanp ANTENNA_565 (.A(net573));
 sg13g2_antennanp ANTENNA_566 (.A(net573));
 sg13g2_antennanp ANTENNA_567 (.A(net573));
 sg13g2_antennanp ANTENNA_568 (.A(net573));
 sg13g2_antennanp ANTENNA_569 (.A(net573));
 sg13g2_antennanp ANTENNA_570 (.A(net573));
 sg13g2_antennanp ANTENNA_571 (.A(net573));
 sg13g2_antennanp ANTENNA_572 (.A(net573));
 sg13g2_antennanp ANTENNA_573 (.A(net573));
 sg13g2_antennanp ANTENNA_574 (.A(net573));
 sg13g2_antennanp ANTENNA_575 (.A(net573));
 sg13g2_antennanp ANTENNA_576 (.A(net573));
 sg13g2_antennanp ANTENNA_577 (.A(net573));
 sg13g2_antennanp ANTENNA_578 (.A(net573));
 sg13g2_antennanp ANTENNA_579 (.A(net573));
 sg13g2_antennanp ANTENNA_580 (.A(net573));
 sg13g2_antennanp ANTENNA_581 (.A(net573));
 sg13g2_antennanp ANTENNA_582 (.A(net573));
 sg13g2_antennanp ANTENNA_583 (.A(net573));
 sg13g2_antennanp ANTENNA_584 (.A(net573));
 sg13g2_antennanp ANTENNA_585 (.A(net573));
 sg13g2_antennanp ANTENNA_586 (.A(net573));
 sg13g2_antennanp ANTENNA_587 (.A(net573));
 sg13g2_antennanp ANTENNA_588 (.A(net573));
 sg13g2_antennanp ANTENNA_589 (.A(net573));
 sg13g2_antennanp ANTENNA_590 (.A(net573));
 sg13g2_antennanp ANTENNA_591 (.A(net573));
 sg13g2_antennanp ANTENNA_592 (.A(net573));
 sg13g2_antennanp ANTENNA_593 (.A(net573));
 sg13g2_antennanp ANTENNA_594 (.A(net573));
 sg13g2_antennanp ANTENNA_595 (.A(net573));
 sg13g2_antennanp ANTENNA_596 (.A(net573));
 sg13g2_antennanp ANTENNA_597 (.A(net573));
 sg13g2_antennanp ANTENNA_598 (.A(net573));
 sg13g2_antennanp ANTENNA_599 (.A(net573));
 sg13g2_antennanp ANTENNA_600 (.A(net573));
 sg13g2_antennanp ANTENNA_601 (.A(net573));
 sg13g2_antennanp ANTENNA_602 (.A(net573));
 sg13g2_antennanp ANTENNA_603 (.A(net573));
 sg13g2_antennanp ANTENNA_604 (.A(net573));
 sg13g2_antennanp ANTENNA_605 (.A(net573));
 sg13g2_antennanp ANTENNA_606 (.A(net573));
 sg13g2_antennanp ANTENNA_607 (.A(net573));
 sg13g2_antennanp ANTENNA_608 (.A(net573));
 sg13g2_antennanp ANTENNA_609 (.A(net573));
 sg13g2_antennanp ANTENNA_610 (.A(net573));
 sg13g2_antennanp ANTENNA_611 (.A(net573));
 sg13g2_antennanp ANTENNA_612 (.A(net573));
 sg13g2_antennanp ANTENNA_613 (.A(net573));
 sg13g2_antennanp ANTENNA_614 (.A(net573));
 sg13g2_antennanp ANTENNA_615 (.A(net576));
 sg13g2_antennanp ANTENNA_616 (.A(net576));
 sg13g2_antennanp ANTENNA_617 (.A(net576));
 sg13g2_antennanp ANTENNA_618 (.A(net576));
 sg13g2_antennanp ANTENNA_619 (.A(net576));
 sg13g2_antennanp ANTENNA_620 (.A(net576));
 sg13g2_antennanp ANTENNA_621 (.A(net576));
 sg13g2_antennanp ANTENNA_622 (.A(net576));
 sg13g2_antennanp ANTENNA_623 (.A(net576));
 sg13g2_antennanp ANTENNA_624 (.A(net576));
 sg13g2_antennanp ANTENNA_625 (.A(net576));
 sg13g2_antennanp ANTENNA_626 (.A(net576));
 sg13g2_antennanp ANTENNA_627 (.A(net576));
 sg13g2_antennanp ANTENNA_628 (.A(net576));
 sg13g2_antennanp ANTENNA_629 (.A(net576));
 sg13g2_antennanp ANTENNA_630 (.A(net576));
 sg13g2_antennanp ANTENNA_631 (.A(net576));
 sg13g2_antennanp ANTENNA_632 (.A(net576));
 sg13g2_antennanp ANTENNA_633 (.A(net576));
 sg13g2_antennanp ANTENNA_634 (.A(net576));
 sg13g2_antennanp ANTENNA_635 (.A(net577));
 sg13g2_antennanp ANTENNA_636 (.A(net577));
 sg13g2_antennanp ANTENNA_637 (.A(net577));
 sg13g2_antennanp ANTENNA_638 (.A(net577));
 sg13g2_antennanp ANTENNA_639 (.A(net577));
 sg13g2_antennanp ANTENNA_640 (.A(net577));
 sg13g2_antennanp ANTENNA_641 (.A(net577));
 sg13g2_antennanp ANTENNA_642 (.A(net577));
 sg13g2_antennanp ANTENNA_643 (.A(net577));
 sg13g2_antennanp ANTENNA_644 (.A(net577));
 sg13g2_antennanp ANTENNA_645 (.A(net577));
 sg13g2_antennanp ANTENNA_646 (.A(net577));
 sg13g2_antennanp ANTENNA_647 (.A(net577));
 sg13g2_antennanp ANTENNA_648 (.A(net577));
 sg13g2_antennanp ANTENNA_649 (.A(net577));
 sg13g2_antennanp ANTENNA_650 (.A(net577));
 sg13g2_antennanp ANTENNA_651 (.A(net578));
 sg13g2_antennanp ANTENNA_652 (.A(net578));
 sg13g2_antennanp ANTENNA_653 (.A(net578));
 sg13g2_antennanp ANTENNA_654 (.A(net578));
 sg13g2_antennanp ANTENNA_655 (.A(net578));
 sg13g2_antennanp ANTENNA_656 (.A(net578));
 sg13g2_antennanp ANTENNA_657 (.A(net578));
 sg13g2_antennanp ANTENNA_658 (.A(net578));
 sg13g2_antennanp ANTENNA_659 (.A(net578));
 sg13g2_antennanp ANTENNA_660 (.A(net578));
 sg13g2_antennanp ANTENNA_661 (.A(net578));
 sg13g2_antennanp ANTENNA_662 (.A(net578));
 sg13g2_antennanp ANTENNA_663 (.A(net578));
 sg13g2_antennanp ANTENNA_664 (.A(net578));
 sg13g2_antennanp ANTENNA_665 (.A(net578));
 sg13g2_antennanp ANTENNA_666 (.A(net578));
 sg13g2_antennanp ANTENNA_667 (.A(net578));
 sg13g2_antennanp ANTENNA_668 (.A(net578));
 sg13g2_antennanp ANTENNA_669 (.A(net578));
 sg13g2_antennanp ANTENNA_670 (.A(net578));
 sg13g2_antennanp ANTENNA_671 (.A(net714));
 sg13g2_antennanp ANTENNA_672 (.A(net714));
 sg13g2_antennanp ANTENNA_673 (.A(net714));
 sg13g2_antennanp ANTENNA_674 (.A(net714));
 sg13g2_antennanp ANTENNA_675 (.A(net714));
 sg13g2_antennanp ANTENNA_676 (.A(net714));
 sg13g2_antennanp ANTENNA_677 (.A(net714));
 sg13g2_antennanp ANTENNA_678 (.A(net714));
 sg13g2_antennanp ANTENNA_679 (.A(net714));
 sg13g2_antennanp ANTENNA_680 (.A(net716));
 sg13g2_antennanp ANTENNA_681 (.A(net716));
 sg13g2_antennanp ANTENNA_682 (.A(net716));
 sg13g2_antennanp ANTENNA_683 (.A(net716));
 sg13g2_antennanp ANTENNA_684 (.A(net716));
 sg13g2_antennanp ANTENNA_685 (.A(net716));
 sg13g2_antennanp ANTENNA_686 (.A(net716));
 sg13g2_antennanp ANTENNA_687 (.A(net716));
 sg13g2_antennanp ANTENNA_688 (.A(net716));
 sg13g2_antennanp ANTENNA_689 (.A(net716));
 sg13g2_antennanp ANTENNA_690 (.A(net716));
 sg13g2_antennanp ANTENNA_691 (.A(net716));
 sg13g2_antennanp ANTENNA_692 (.A(net716));
 sg13g2_antennanp ANTENNA_693 (.A(net716));
 sg13g2_antennanp ANTENNA_694 (.A(net716));
 sg13g2_antennanp ANTENNA_695 (.A(net716));
 sg13g2_antennanp ANTENNA_696 (.A(net716));
 sg13g2_antennanp ANTENNA_697 (.A(net716));
 sg13g2_antennanp ANTENNA_698 (.A(net716));
 sg13g2_antennanp ANTENNA_699 (.A(net716));
 sg13g2_antennanp ANTENNA_700 (.A(net716));
 sg13g2_antennanp ANTENNA_701 (.A(net716));
 sg13g2_antennanp ANTENNA_702 (.A(net716));
 sg13g2_antennanp ANTENNA_703 (.A(net747));
 sg13g2_antennanp ANTENNA_704 (.A(net747));
 sg13g2_antennanp ANTENNA_705 (.A(net747));
 sg13g2_antennanp ANTENNA_706 (.A(net747));
 sg13g2_antennanp ANTENNA_707 (.A(net747));
 sg13g2_antennanp ANTENNA_708 (.A(net747));
 sg13g2_antennanp ANTENNA_709 (.A(net747));
 sg13g2_antennanp ANTENNA_710 (.A(net747));
 sg13g2_antennanp ANTENNA_711 (.A(net749));
 sg13g2_antennanp ANTENNA_712 (.A(net749));
 sg13g2_antennanp ANTENNA_713 (.A(net749));
 sg13g2_antennanp ANTENNA_714 (.A(net749));
 sg13g2_antennanp ANTENNA_715 (.A(net749));
 sg13g2_antennanp ANTENNA_716 (.A(net749));
 sg13g2_antennanp ANTENNA_717 (.A(net749));
 sg13g2_antennanp ANTENNA_718 (.A(net749));
 sg13g2_antennanp ANTENNA_719 (.A(net749));
 sg13g2_antennanp ANTENNA_720 (.A(net827));
 sg13g2_antennanp ANTENNA_721 (.A(net827));
 sg13g2_antennanp ANTENNA_722 (.A(net827));
 sg13g2_antennanp ANTENNA_723 (.A(net827));
 sg13g2_antennanp ANTENNA_724 (.A(net827));
 sg13g2_antennanp ANTENNA_725 (.A(net827));
 sg13g2_antennanp ANTENNA_726 (.A(net827));
 sg13g2_antennanp ANTENNA_727 (.A(net827));
 sg13g2_antennanp ANTENNA_728 (.A(net827));
 sg13g2_antennanp ANTENNA_729 (.A(net831));
 sg13g2_antennanp ANTENNA_730 (.A(net831));
 sg13g2_antennanp ANTENNA_731 (.A(net831));
 sg13g2_antennanp ANTENNA_732 (.A(net831));
 sg13g2_antennanp ANTENNA_733 (.A(net831));
 sg13g2_antennanp ANTENNA_734 (.A(net831));
 sg13g2_antennanp ANTENNA_735 (.A(net831));
 sg13g2_antennanp ANTENNA_736 (.A(net831));
 sg13g2_antennanp ANTENNA_737 (.A(net831));
 sg13g2_antennanp ANTENNA_738 (.A(net834));
 sg13g2_antennanp ANTENNA_739 (.A(net834));
 sg13g2_antennanp ANTENNA_740 (.A(net834));
 sg13g2_antennanp ANTENNA_741 (.A(net834));
 sg13g2_antennanp ANTENNA_742 (.A(net834));
 sg13g2_antennanp ANTENNA_743 (.A(net834));
 sg13g2_antennanp ANTENNA_744 (.A(net834));
 sg13g2_antennanp ANTENNA_745 (.A(net834));
 sg13g2_antennanp ANTENNA_746 (.A(net834));
 sg13g2_antennanp ANTENNA_747 (.A(net836));
 sg13g2_antennanp ANTENNA_748 (.A(net836));
 sg13g2_antennanp ANTENNA_749 (.A(net836));
 sg13g2_antennanp ANTENNA_750 (.A(net836));
 sg13g2_antennanp ANTENNA_751 (.A(net836));
 sg13g2_antennanp ANTENNA_752 (.A(net836));
 sg13g2_antennanp ANTENNA_753 (.A(net836));
 sg13g2_antennanp ANTENNA_754 (.A(net836));
 sg13g2_antennanp ANTENNA_755 (.A(net836));
 sg13g2_antennanp ANTENNA_756 (.A(net837));
 sg13g2_antennanp ANTENNA_757 (.A(net837));
 sg13g2_antennanp ANTENNA_758 (.A(net837));
 sg13g2_antennanp ANTENNA_759 (.A(net837));
 sg13g2_antennanp ANTENNA_760 (.A(net837));
 sg13g2_antennanp ANTENNA_761 (.A(net837));
 sg13g2_antennanp ANTENNA_762 (.A(net837));
 sg13g2_antennanp ANTENNA_763 (.A(net837));
 sg13g2_antennanp ANTENNA_764 (.A(net837));
 sg13g2_antennanp ANTENNA_765 (.A(net841));
 sg13g2_antennanp ANTENNA_766 (.A(net841));
 sg13g2_antennanp ANTENNA_767 (.A(net841));
 sg13g2_antennanp ANTENNA_768 (.A(net841));
 sg13g2_antennanp ANTENNA_769 (.A(net841));
 sg13g2_antennanp ANTENNA_770 (.A(net841));
 sg13g2_antennanp ANTENNA_771 (.A(net841));
 sg13g2_antennanp ANTENNA_772 (.A(net841));
 sg13g2_antennanp ANTENNA_773 (.A(net841));
 sg13g2_antennanp ANTENNA_774 (.A(net871));
 sg13g2_antennanp ANTENNA_775 (.A(net871));
 sg13g2_antennanp ANTENNA_776 (.A(net871));
 sg13g2_antennanp ANTENNA_777 (.A(net871));
 sg13g2_antennanp ANTENNA_778 (.A(net871));
 sg13g2_antennanp ANTENNA_779 (.A(net871));
 sg13g2_antennanp ANTENNA_780 (.A(net871));
 sg13g2_antennanp ANTENNA_781 (.A(net871));
 sg13g2_antennanp ANTENNA_782 (.A(net879));
 sg13g2_antennanp ANTENNA_783 (.A(net879));
 sg13g2_antennanp ANTENNA_784 (.A(net879));
 sg13g2_antennanp ANTENNA_785 (.A(net879));
 sg13g2_antennanp ANTENNA_786 (.A(net879));
 sg13g2_antennanp ANTENNA_787 (.A(net879));
 sg13g2_antennanp ANTENNA_788 (.A(net879));
 sg13g2_antennanp ANTENNA_789 (.A(net879));
 sg13g2_antennanp ANTENNA_790 (.A(net879));
 sg13g2_antennanp ANTENNA_791 (.A(net879));
 sg13g2_antennanp ANTENNA_792 (.A(net879));
 sg13g2_antennanp ANTENNA_793 (.A(net879));
 sg13g2_antennanp ANTENNA_794 (.A(net896));
 sg13g2_antennanp ANTENNA_795 (.A(net896));
 sg13g2_antennanp ANTENNA_796 (.A(net896));
 sg13g2_antennanp ANTENNA_797 (.A(net896));
 sg13g2_antennanp ANTENNA_798 (.A(net896));
 sg13g2_antennanp ANTENNA_799 (.A(net896));
 sg13g2_antennanp ANTENNA_800 (.A(net896));
 sg13g2_antennanp ANTENNA_801 (.A(net896));
 sg13g2_antennanp ANTENNA_802 (.A(net896));
 sg13g2_antennanp ANTENNA_803 (.A(net896));
 sg13g2_antennanp ANTENNA_804 (.A(net896));
 sg13g2_antennanp ANTENNA_805 (.A(net896));
 sg13g2_antennanp ANTENNA_806 (.A(net896));
 sg13g2_antennanp ANTENNA_807 (.A(net896));
 sg13g2_antennanp ANTENNA_808 (.A(net896));
 sg13g2_antennanp ANTENNA_809 (.A(net896));
 sg13g2_antennanp ANTENNA_810 (.A(net896));
 sg13g2_antennanp ANTENNA_811 (.A(net896));
 sg13g2_antennanp ANTENNA_812 (.A(net896));
 sg13g2_antennanp ANTENNA_813 (.A(net896));
 sg13g2_antennanp ANTENNA_814 (.A(net896));
 sg13g2_antennanp ANTENNA_815 (.A(net905));
 sg13g2_antennanp ANTENNA_816 (.A(net905));
 sg13g2_antennanp ANTENNA_817 (.A(net905));
 sg13g2_antennanp ANTENNA_818 (.A(net905));
 sg13g2_antennanp ANTENNA_819 (.A(net905));
 sg13g2_antennanp ANTENNA_820 (.A(net905));
 sg13g2_antennanp ANTENNA_821 (.A(net905));
 sg13g2_antennanp ANTENNA_822 (.A(net905));
 sg13g2_antennanp ANTENNA_823 (.A(net905));
 sg13g2_antennanp ANTENNA_824 (.A(net953));
 sg13g2_antennanp ANTENNA_825 (.A(net953));
 sg13g2_antennanp ANTENNA_826 (.A(net953));
 sg13g2_antennanp ANTENNA_827 (.A(net953));
 sg13g2_antennanp ANTENNA_828 (.A(net953));
 sg13g2_antennanp ANTENNA_829 (.A(net953));
 sg13g2_antennanp ANTENNA_830 (.A(net953));
 sg13g2_antennanp ANTENNA_831 (.A(net953));
 sg13g2_antennanp ANTENNA_832 (.A(net953));
 sg13g2_antennanp ANTENNA_833 (.A(net953));
 sg13g2_antennanp ANTENNA_834 (.A(net953));
 sg13g2_antennanp ANTENNA_835 (.A(net953));
 sg13g2_antennanp ANTENNA_836 (.A(net953));
 sg13g2_antennanp ANTENNA_837 (.A(net953));
 sg13g2_antennanp ANTENNA_838 (.A(net967));
 sg13g2_antennanp ANTENNA_839 (.A(net967));
 sg13g2_antennanp ANTENNA_840 (.A(net967));
 sg13g2_antennanp ANTENNA_841 (.A(net967));
 sg13g2_antennanp ANTENNA_842 (.A(net967));
 sg13g2_antennanp ANTENNA_843 (.A(net967));
 sg13g2_antennanp ANTENNA_844 (.A(net967));
 sg13g2_antennanp ANTENNA_845 (.A(net967));
 sg13g2_antennanp ANTENNA_846 (.A(net967));
 sg13g2_antennanp ANTENNA_847 (.A(net967));
 sg13g2_antennanp ANTENNA_848 (.A(net967));
 sg13g2_antennanp ANTENNA_849 (.A(net967));
 sg13g2_antennanp ANTENNA_850 (.A(net967));
 sg13g2_antennanp ANTENNA_851 (.A(net967));
 sg13g2_antennanp ANTENNA_852 (.A(net967));
 sg13g2_antennanp ANTENNA_853 (.A(net967));
 sg13g2_antennanp ANTENNA_854 (.A(net968));
 sg13g2_antennanp ANTENNA_855 (.A(net968));
 sg13g2_antennanp ANTENNA_856 (.A(net968));
 sg13g2_antennanp ANTENNA_857 (.A(net968));
 sg13g2_antennanp ANTENNA_858 (.A(net968));
 sg13g2_antennanp ANTENNA_859 (.A(net968));
 sg13g2_antennanp ANTENNA_860 (.A(net968));
 sg13g2_antennanp ANTENNA_861 (.A(net968));
 sg13g2_antennanp ANTENNA_862 (.A(net968));
 sg13g2_antennanp ANTENNA_863 (.A(net968));
 sg13g2_antennanp ANTENNA_864 (.A(net968));
 sg13g2_antennanp ANTENNA_865 (.A(net968));
 sg13g2_antennanp ANTENNA_866 (.A(net968));
 sg13g2_antennanp ANTENNA_867 (.A(net968));
 sg13g2_antennanp ANTENNA_868 (.A(net968));
 sg13g2_antennanp ANTENNA_869 (.A(net968));
 sg13g2_antennanp ANTENNA_870 (.A(net968));
 sg13g2_antennanp ANTENNA_871 (.A(net968));
 sg13g2_antennanp ANTENNA_872 (.A(net968));
 sg13g2_antennanp ANTENNA_873 (.A(net968));
 sg13g2_antennanp ANTENNA_874 (.A(net968));
 sg13g2_antennanp ANTENNA_875 (.A(net981));
 sg13g2_antennanp ANTENNA_876 (.A(net981));
 sg13g2_antennanp ANTENNA_877 (.A(net981));
 sg13g2_antennanp ANTENNA_878 (.A(net981));
 sg13g2_antennanp ANTENNA_879 (.A(net981));
 sg13g2_antennanp ANTENNA_880 (.A(net981));
 sg13g2_antennanp ANTENNA_881 (.A(net981));
 sg13g2_antennanp ANTENNA_882 (.A(net981));
 sg13g2_antennanp ANTENNA_883 (.A(net981));
 sg13g2_antennanp ANTENNA_884 (.A(net981));
 sg13g2_antennanp ANTENNA_885 (.A(net981));
 sg13g2_antennanp ANTENNA_886 (.A(net981));
 sg13g2_antennanp ANTENNA_887 (.A(net981));
 sg13g2_antennanp ANTENNA_888 (.A(net981));
 sg13g2_antennanp ANTENNA_889 (.A(net981));
 sg13g2_antennanp ANTENNA_890 (.A(net981));
 sg13g2_antennanp ANTENNA_891 (.A(net981));
 sg13g2_antennanp ANTENNA_892 (.A(net994));
 sg13g2_antennanp ANTENNA_893 (.A(net994));
 sg13g2_antennanp ANTENNA_894 (.A(net994));
 sg13g2_antennanp ANTENNA_895 (.A(net994));
 sg13g2_antennanp ANTENNA_896 (.A(net994));
 sg13g2_antennanp ANTENNA_897 (.A(net994));
 sg13g2_antennanp ANTENNA_898 (.A(net994));
 sg13g2_antennanp ANTENNA_899 (.A(net994));
 sg13g2_antennanp ANTENNA_900 (.A(net994));
 sg13g2_antennanp ANTENNA_901 (.A(net994));
 sg13g2_antennanp ANTENNA_902 (.A(net994));
 sg13g2_antennanp ANTENNA_903 (.A(net994));
 sg13g2_antennanp ANTENNA_904 (.A(net994));
 sg13g2_antennanp ANTENNA_905 (.A(net994));
 sg13g2_antennanp ANTENNA_906 (.A(net994));
 sg13g2_antennanp ANTENNA_907 (.A(net994));
 sg13g2_antennanp ANTENNA_908 (.A(net994));
 sg13g2_antennanp ANTENNA_909 (.A(net994));
 sg13g2_antennanp ANTENNA_910 (.A(net994));
 sg13g2_antennanp ANTENNA_911 (.A(net994));
 sg13g2_antennanp ANTENNA_912 (.A(net994));
 sg13g2_antennanp ANTENNA_913 (.A(net994));
 sg13g2_antennanp ANTENNA_914 (.A(net994));
 sg13g2_antennanp ANTENNA_915 (.A(net1019));
 sg13g2_antennanp ANTENNA_916 (.A(net1019));
 sg13g2_antennanp ANTENNA_917 (.A(net1019));
 sg13g2_antennanp ANTENNA_918 (.A(net1019));
 sg13g2_antennanp ANTENNA_919 (.A(net1019));
 sg13g2_antennanp ANTENNA_920 (.A(net1019));
 sg13g2_antennanp ANTENNA_921 (.A(net1019));
 sg13g2_antennanp ANTENNA_922 (.A(net1019));
 sg13g2_antennanp ANTENNA_923 (.A(net1019));
 sg13g2_antennanp ANTENNA_924 (.A(net1019));
 sg13g2_antennanp ANTENNA_925 (.A(net1019));
 sg13g2_antennanp ANTENNA_926 (.A(net1019));
 sg13g2_antennanp ANTENNA_927 (.A(net1019));
 sg13g2_antennanp ANTENNA_928 (.A(net1019));
 sg13g2_antennanp ANTENNA_929 (.A(net1019));
 sg13g2_antennanp ANTENNA_930 (.A(net1019));
 sg13g2_antennanp ANTENNA_931 (.A(net1019));
 sg13g2_antennanp ANTENNA_932 (.A(net1019));
 sg13g2_antennanp ANTENNA_933 (.A(net1019));
 sg13g2_antennanp ANTENNA_934 (.A(net1019));
 sg13g2_antennanp ANTENNA_935 (.A(net1022));
 sg13g2_antennanp ANTENNA_936 (.A(net1022));
 sg13g2_antennanp ANTENNA_937 (.A(net1022));
 sg13g2_antennanp ANTENNA_938 (.A(net1022));
 sg13g2_antennanp ANTENNA_939 (.A(net1022));
 sg13g2_antennanp ANTENNA_940 (.A(net1022));
 sg13g2_antennanp ANTENNA_941 (.A(net1022));
 sg13g2_antennanp ANTENNA_942 (.A(net1022));
 sg13g2_antennanp ANTENNA_943 (.A(net1022));
 sg13g2_antennanp ANTENNA_944 (.A(net1022));
 sg13g2_antennanp ANTENNA_945 (.A(net1022));
 sg13g2_antennanp ANTENNA_946 (.A(net1022));
 sg13g2_antennanp ANTENNA_947 (.A(net1022));
 sg13g2_antennanp ANTENNA_948 (.A(net1022));
 sg13g2_antennanp ANTENNA_949 (.A(net1022));
 sg13g2_antennanp ANTENNA_950 (.A(net1022));
 sg13g2_antennanp ANTENNA_951 (.A(net1022));
 sg13g2_antennanp ANTENNA_952 (.A(net1022));
 sg13g2_antennanp ANTENNA_953 (.A(net1022));
 sg13g2_antennanp ANTENNA_954 (.A(net1022));
 sg13g2_antennanp ANTENNA_955 (.A(net1085));
 sg13g2_antennanp ANTENNA_956 (.A(net1085));
 sg13g2_antennanp ANTENNA_957 (.A(net1085));
 sg13g2_antennanp ANTENNA_958 (.A(net1085));
 sg13g2_antennanp ANTENNA_959 (.A(net1085));
 sg13g2_antennanp ANTENNA_960 (.A(net1085));
 sg13g2_antennanp ANTENNA_961 (.A(net1085));
 sg13g2_antennanp ANTENNA_962 (.A(net1085));
 sg13g2_antennanp ANTENNA_963 (.A(net1096));
 sg13g2_antennanp ANTENNA_964 (.A(net1096));
 sg13g2_antennanp ANTENNA_965 (.A(net1096));
 sg13g2_antennanp ANTENNA_966 (.A(net1096));
 sg13g2_antennanp ANTENNA_967 (.A(net1096));
 sg13g2_antennanp ANTENNA_968 (.A(net1096));
 sg13g2_antennanp ANTENNA_969 (.A(net1096));
 sg13g2_antennanp ANTENNA_970 (.A(net1096));
 sg13g2_antennanp ANTENNA_971 (.A(_00930_));
 sg13g2_antennanp ANTENNA_972 (.A(_00930_));
 sg13g2_antennanp ANTENNA_973 (.A(_01052_));
 sg13g2_antennanp ANTENNA_974 (.A(_01052_));
 sg13g2_antennanp ANTENNA_975 (.A(_01057_));
 sg13g2_antennanp ANTENNA_976 (.A(_01057_));
 sg13g2_antennanp ANTENNA_977 (.A(_01071_));
 sg13g2_antennanp ANTENNA_978 (.A(_02855_));
 sg13g2_antennanp ANTENNA_979 (.A(_02855_));
 sg13g2_antennanp ANTENNA_980 (.A(_02855_));
 sg13g2_antennanp ANTENNA_981 (.A(_02855_));
 sg13g2_antennanp ANTENNA_982 (.A(_02855_));
 sg13g2_antennanp ANTENNA_983 (.A(_02855_));
 sg13g2_antennanp ANTENNA_984 (.A(_02855_));
 sg13g2_antennanp ANTENNA_985 (.A(_02855_));
 sg13g2_antennanp ANTENNA_986 (.A(_02856_));
 sg13g2_antennanp ANTENNA_987 (.A(_02856_));
 sg13g2_antennanp ANTENNA_988 (.A(_02856_));
 sg13g2_antennanp ANTENNA_989 (.A(_02856_));
 sg13g2_antennanp ANTENNA_990 (.A(_02856_));
 sg13g2_antennanp ANTENNA_991 (.A(_02856_));
 sg13g2_antennanp ANTENNA_992 (.A(_02856_));
 sg13g2_antennanp ANTENNA_993 (.A(_02856_));
 sg13g2_antennanp ANTENNA_994 (.A(_02856_));
 sg13g2_antennanp ANTENNA_995 (.A(_02856_));
 sg13g2_antennanp ANTENNA_996 (.A(_02866_));
 sg13g2_antennanp ANTENNA_997 (.A(_02866_));
 sg13g2_antennanp ANTENNA_998 (.A(_02866_));
 sg13g2_antennanp ANTENNA_999 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1000 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1001 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1002 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1003 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1004 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1005 (.A(_02873_));
 sg13g2_antennanp ANTENNA_1006 (.A(_02873_));
 sg13g2_antennanp ANTENNA_1007 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1008 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1009 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1010 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1011 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1012 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1013 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1014 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1015 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1016 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1017 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1018 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1019 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1020 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1021 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1022 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1023 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1024 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1025 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1026 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1027 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1028 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1029 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1030 (.A(_03369_));
 sg13g2_antennanp ANTENNA_1031 (.A(_03369_));
 sg13g2_antennanp ANTENNA_1032 (.A(_03369_));
 sg13g2_antennanp ANTENNA_1033 (.A(_03369_));
 sg13g2_antennanp ANTENNA_1034 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1035 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1036 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1037 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1038 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1039 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1040 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1041 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1042 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1043 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1044 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1045 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1046 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1047 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1048 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1049 (.A(_04646_));
 sg13g2_antennanp ANTENNA_1050 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1051 (.A(_05022_));
 sg13g2_antennanp ANTENNA_1052 (.A(_05046_));
 sg13g2_antennanp ANTENNA_1053 (.A(_05581_));
 sg13g2_antennanp ANTENNA_1054 (.A(_05584_));
 sg13g2_antennanp ANTENNA_1055 (.A(_05593_));
 sg13g2_antennanp ANTENNA_1056 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1057 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1058 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1059 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1060 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1061 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1062 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1063 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1064 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1065 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1066 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1067 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1068 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1069 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1070 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1071 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1072 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1073 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1074 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1075 (.A(_07137_));
 sg13g2_antennanp ANTENNA_1076 (.A(_07138_));
 sg13g2_antennanp ANTENNA_1077 (.A(_07166_));
 sg13g2_antennanp ANTENNA_1078 (.A(_07166_));
 sg13g2_antennanp ANTENNA_1079 (.A(_07222_));
 sg13g2_antennanp ANTENNA_1080 (.A(_07326_));
 sg13g2_antennanp ANTENNA_1081 (.A(_07326_));
 sg13g2_antennanp ANTENNA_1082 (.A(_07976_));
 sg13g2_antennanp ANTENNA_1083 (.A(_07976_));
 sg13g2_antennanp ANTENNA_1084 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1085 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1086 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1087 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1088 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1089 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1090 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1091 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1092 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1093 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1094 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1095 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1096 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1097 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1098 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1099 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1100 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1101 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1102 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1103 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1104 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1105 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1106 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1107 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1108 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1109 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1110 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1111 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1112 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1113 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1114 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1115 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1116 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1117 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1118 (.A(_08345_));
 sg13g2_antennanp ANTENNA_1119 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1120 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1121 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1122 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1123 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1124 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1125 (.A(_08517_));
 sg13g2_antennanp ANTENNA_1126 (.A(_08556_));
 sg13g2_antennanp ANTENNA_1127 (.A(_08614_));
 sg13g2_antennanp ANTENNA_1128 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1129 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1130 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1131 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1132 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1133 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1134 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1135 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1136 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1137 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1138 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1139 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1140 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1141 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1142 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1143 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1144 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1145 (.A(_08993_));
 sg13g2_antennanp ANTENNA_1146 (.A(_09005_));
 sg13g2_antennanp ANTENNA_1147 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1148 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1149 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1150 (.A(_09037_));
 sg13g2_antennanp ANTENNA_1151 (.A(_09037_));
 sg13g2_antennanp ANTENNA_1152 (.A(_09037_));
 sg13g2_antennanp ANTENNA_1153 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1154 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1155 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1156 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1157 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1158 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1159 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1160 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1161 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1162 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1163 (.A(_09234_));
 sg13g2_antennanp ANTENNA_1164 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1165 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1166 (.A(_09305_));
 sg13g2_antennanp ANTENNA_1167 (.A(_09328_));
 sg13g2_antennanp ANTENNA_1168 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1169 (.A(_09370_));
 sg13g2_antennanp ANTENNA_1170 (.A(_09394_));
 sg13g2_antennanp ANTENNA_1171 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1172 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1173 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1174 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1175 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1176 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1177 (.A(_09526_));
 sg13g2_antennanp ANTENNA_1178 (.A(_09553_));
 sg13g2_antennanp ANTENNA_1179 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1180 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1181 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1182 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1183 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1184 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1185 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1186 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1187 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1188 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1189 (.A(_09839_));
 sg13g2_antennanp ANTENNA_1190 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1191 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1192 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1193 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1194 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1195 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1196 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1197 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1198 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1199 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1200 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1201 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1202 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1203 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1204 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1205 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1206 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1207 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1208 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1209 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1210 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1211 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1212 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1213 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1214 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1215 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1216 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1217 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1218 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1219 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1220 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1221 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1222 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1223 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1224 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1225 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1226 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1227 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1228 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1229 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1230 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1231 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1232 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1233 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1234 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1235 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1236 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1237 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1238 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1239 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1240 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1241 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1242 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1243 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1244 (.A(_09985_));
 sg13g2_antennanp ANTENNA_1245 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1246 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1247 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1248 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1249 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1250 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1251 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1252 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1253 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1254 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1255 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1256 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1257 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1258 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1259 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1260 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1261 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1262 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1263 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1264 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1265 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1266 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1267 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1268 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1269 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1270 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1271 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1272 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1273 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1274 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1275 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1276 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1277 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1278 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1279 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1280 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1281 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1282 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1283 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1284 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1285 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1286 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1287 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1288 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1289 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1290 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1291 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1292 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1293 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1294 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1295 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1296 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1297 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1298 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1299 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1300 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1301 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1302 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1303 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1304 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1305 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1306 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1307 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1308 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1309 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1310 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1311 (.A(_11712_));
 sg13g2_antennanp ANTENNA_1312 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1313 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1314 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1315 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1316 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1317 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1318 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1319 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1320 (.A(_11743_));
 sg13g2_antennanp ANTENNA_1321 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1322 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1323 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1324 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1325 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1326 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1327 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1328 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1329 (.A(_11833_));
 sg13g2_antennanp ANTENNA_1330 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1331 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1332 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1333 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1334 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1335 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1336 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1337 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1338 (.A(_11866_));
 sg13g2_antennanp ANTENNA_1339 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1340 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1341 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1342 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1343 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1344 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1345 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1346 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1347 (.A(_11870_));
 sg13g2_antennanp ANTENNA_1348 (.A(_12009_));
 sg13g2_antennanp ANTENNA_1349 (.A(_12009_));
 sg13g2_antennanp ANTENNA_1350 (.A(_12009_));
 sg13g2_antennanp ANTENNA_1351 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1352 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1353 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1354 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1355 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1356 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1357 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1358 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1359 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1360 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1361 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1362 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1363 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1364 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1365 (.A(_12469_));
 sg13g2_antennanp ANTENNA_1366 (.A(_12473_));
 sg13g2_antennanp ANTENNA_1367 (.A(_12473_));
 sg13g2_antennanp ANTENNA_1368 (.A(_12473_));
 sg13g2_antennanp ANTENNA_1369 (.A(_12473_));
 sg13g2_antennanp ANTENNA_1370 (.A(clk));
 sg13g2_antennanp ANTENNA_1371 (.A(clk));
 sg13g2_antennanp ANTENNA_1372 (.A(\cpu.addr[14] ));
 sg13g2_antennanp ANTENNA_1373 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1374 (.A(net3));
 sg13g2_antennanp ANTENNA_1375 (.A(net3));
 sg13g2_antennanp ANTENNA_1376 (.A(net3));
 sg13g2_antennanp ANTENNA_1377 (.A(net11));
 sg13g2_antennanp ANTENNA_1378 (.A(net11));
 sg13g2_antennanp ANTENNA_1379 (.A(net11));
 sg13g2_antennanp ANTENNA_1380 (.A(net12));
 sg13g2_antennanp ANTENNA_1381 (.A(net12));
 sg13g2_antennanp ANTENNA_1382 (.A(net12));
 sg13g2_antennanp ANTENNA_1383 (.A(net14));
 sg13g2_antennanp ANTENNA_1384 (.A(net14));
 sg13g2_antennanp ANTENNA_1385 (.A(net14));
 sg13g2_antennanp ANTENNA_1386 (.A(net18));
 sg13g2_antennanp ANTENNA_1387 (.A(net19));
 sg13g2_antennanp ANTENNA_1388 (.A(net19));
 sg13g2_antennanp ANTENNA_1389 (.A(net20));
 sg13g2_antennanp ANTENNA_1390 (.A(net20));
 sg13g2_antennanp ANTENNA_1391 (.A(net464));
 sg13g2_antennanp ANTENNA_1392 (.A(net464));
 sg13g2_antennanp ANTENNA_1393 (.A(net464));
 sg13g2_antennanp ANTENNA_1394 (.A(net464));
 sg13g2_antennanp ANTENNA_1395 (.A(net464));
 sg13g2_antennanp ANTENNA_1396 (.A(net464));
 sg13g2_antennanp ANTENNA_1397 (.A(net464));
 sg13g2_antennanp ANTENNA_1398 (.A(net464));
 sg13g2_antennanp ANTENNA_1399 (.A(net464));
 sg13g2_antennanp ANTENNA_1400 (.A(net464));
 sg13g2_antennanp ANTENNA_1401 (.A(net464));
 sg13g2_antennanp ANTENNA_1402 (.A(net464));
 sg13g2_antennanp ANTENNA_1403 (.A(net464));
 sg13g2_antennanp ANTENNA_1404 (.A(net464));
 sg13g2_antennanp ANTENNA_1405 (.A(net464));
 sg13g2_antennanp ANTENNA_1406 (.A(net464));
 sg13g2_antennanp ANTENNA_1407 (.A(net464));
 sg13g2_antennanp ANTENNA_1408 (.A(net464));
 sg13g2_antennanp ANTENNA_1409 (.A(net464));
 sg13g2_antennanp ANTENNA_1410 (.A(net464));
 sg13g2_antennanp ANTENNA_1411 (.A(net498));
 sg13g2_antennanp ANTENNA_1412 (.A(net498));
 sg13g2_antennanp ANTENNA_1413 (.A(net498));
 sg13g2_antennanp ANTENNA_1414 (.A(net498));
 sg13g2_antennanp ANTENNA_1415 (.A(net498));
 sg13g2_antennanp ANTENNA_1416 (.A(net498));
 sg13g2_antennanp ANTENNA_1417 (.A(net498));
 sg13g2_antennanp ANTENNA_1418 (.A(net498));
 sg13g2_antennanp ANTENNA_1419 (.A(net498));
 sg13g2_antennanp ANTENNA_1420 (.A(net573));
 sg13g2_antennanp ANTENNA_1421 (.A(net573));
 sg13g2_antennanp ANTENNA_1422 (.A(net573));
 sg13g2_antennanp ANTENNA_1423 (.A(net573));
 sg13g2_antennanp ANTENNA_1424 (.A(net573));
 sg13g2_antennanp ANTENNA_1425 (.A(net573));
 sg13g2_antennanp ANTENNA_1426 (.A(net573));
 sg13g2_antennanp ANTENNA_1427 (.A(net573));
 sg13g2_antennanp ANTENNA_1428 (.A(net573));
 sg13g2_antennanp ANTENNA_1429 (.A(net573));
 sg13g2_antennanp ANTENNA_1430 (.A(net573));
 sg13g2_antennanp ANTENNA_1431 (.A(net573));
 sg13g2_antennanp ANTENNA_1432 (.A(net573));
 sg13g2_antennanp ANTENNA_1433 (.A(net573));
 sg13g2_antennanp ANTENNA_1434 (.A(net573));
 sg13g2_antennanp ANTENNA_1435 (.A(net573));
 sg13g2_antennanp ANTENNA_1436 (.A(net573));
 sg13g2_antennanp ANTENNA_1437 (.A(net573));
 sg13g2_antennanp ANTENNA_1438 (.A(net573));
 sg13g2_antennanp ANTENNA_1439 (.A(net573));
 sg13g2_antennanp ANTENNA_1440 (.A(net576));
 sg13g2_antennanp ANTENNA_1441 (.A(net576));
 sg13g2_antennanp ANTENNA_1442 (.A(net576));
 sg13g2_antennanp ANTENNA_1443 (.A(net576));
 sg13g2_antennanp ANTENNA_1444 (.A(net576));
 sg13g2_antennanp ANTENNA_1445 (.A(net576));
 sg13g2_antennanp ANTENNA_1446 (.A(net576));
 sg13g2_antennanp ANTENNA_1447 (.A(net576));
 sg13g2_antennanp ANTENNA_1448 (.A(net576));
 sg13g2_antennanp ANTENNA_1449 (.A(net576));
 sg13g2_antennanp ANTENNA_1450 (.A(net576));
 sg13g2_antennanp ANTENNA_1451 (.A(net576));
 sg13g2_antennanp ANTENNA_1452 (.A(net576));
 sg13g2_antennanp ANTENNA_1453 (.A(net576));
 sg13g2_antennanp ANTENNA_1454 (.A(net576));
 sg13g2_antennanp ANTENNA_1455 (.A(net576));
 sg13g2_antennanp ANTENNA_1456 (.A(net576));
 sg13g2_antennanp ANTENNA_1457 (.A(net576));
 sg13g2_antennanp ANTENNA_1458 (.A(net576));
 sg13g2_antennanp ANTENNA_1459 (.A(net576));
 sg13g2_antennanp ANTENNA_1460 (.A(net578));
 sg13g2_antennanp ANTENNA_1461 (.A(net578));
 sg13g2_antennanp ANTENNA_1462 (.A(net578));
 sg13g2_antennanp ANTENNA_1463 (.A(net578));
 sg13g2_antennanp ANTENNA_1464 (.A(net578));
 sg13g2_antennanp ANTENNA_1465 (.A(net578));
 sg13g2_antennanp ANTENNA_1466 (.A(net578));
 sg13g2_antennanp ANTENNA_1467 (.A(net578));
 sg13g2_antennanp ANTENNA_1468 (.A(net578));
 sg13g2_antennanp ANTENNA_1469 (.A(net578));
 sg13g2_antennanp ANTENNA_1470 (.A(net578));
 sg13g2_antennanp ANTENNA_1471 (.A(net578));
 sg13g2_antennanp ANTENNA_1472 (.A(net578));
 sg13g2_antennanp ANTENNA_1473 (.A(net578));
 sg13g2_antennanp ANTENNA_1474 (.A(net578));
 sg13g2_antennanp ANTENNA_1475 (.A(net578));
 sg13g2_antennanp ANTENNA_1476 (.A(net578));
 sg13g2_antennanp ANTENNA_1477 (.A(net578));
 sg13g2_antennanp ANTENNA_1478 (.A(net578));
 sg13g2_antennanp ANTENNA_1479 (.A(net578));
 sg13g2_antennanp ANTENNA_1480 (.A(net714));
 sg13g2_antennanp ANTENNA_1481 (.A(net714));
 sg13g2_antennanp ANTENNA_1482 (.A(net714));
 sg13g2_antennanp ANTENNA_1483 (.A(net714));
 sg13g2_antennanp ANTENNA_1484 (.A(net714));
 sg13g2_antennanp ANTENNA_1485 (.A(net714));
 sg13g2_antennanp ANTENNA_1486 (.A(net714));
 sg13g2_antennanp ANTENNA_1487 (.A(net714));
 sg13g2_antennanp ANTENNA_1488 (.A(net714));
 sg13g2_antennanp ANTENNA_1489 (.A(net747));
 sg13g2_antennanp ANTENNA_1490 (.A(net747));
 sg13g2_antennanp ANTENNA_1491 (.A(net747));
 sg13g2_antennanp ANTENNA_1492 (.A(net747));
 sg13g2_antennanp ANTENNA_1493 (.A(net747));
 sg13g2_antennanp ANTENNA_1494 (.A(net747));
 sg13g2_antennanp ANTENNA_1495 (.A(net747));
 sg13g2_antennanp ANTENNA_1496 (.A(net747));
 sg13g2_antennanp ANTENNA_1497 (.A(net760));
 sg13g2_antennanp ANTENNA_1498 (.A(net760));
 sg13g2_antennanp ANTENNA_1499 (.A(net760));
 sg13g2_antennanp ANTENNA_1500 (.A(net760));
 sg13g2_antennanp ANTENNA_1501 (.A(net760));
 sg13g2_antennanp ANTENNA_1502 (.A(net760));
 sg13g2_antennanp ANTENNA_1503 (.A(net760));
 sg13g2_antennanp ANTENNA_1504 (.A(net760));
 sg13g2_antennanp ANTENNA_1505 (.A(net760));
 sg13g2_antennanp ANTENNA_1506 (.A(net760));
 sg13g2_antennanp ANTENNA_1507 (.A(net760));
 sg13g2_antennanp ANTENNA_1508 (.A(net760));
 sg13g2_antennanp ANTENNA_1509 (.A(net760));
 sg13g2_antennanp ANTENNA_1510 (.A(net760));
 sg13g2_antennanp ANTENNA_1511 (.A(net760));
 sg13g2_antennanp ANTENNA_1512 (.A(net760));
 sg13g2_antennanp ANTENNA_1513 (.A(net760));
 sg13g2_antennanp ANTENNA_1514 (.A(net827));
 sg13g2_antennanp ANTENNA_1515 (.A(net827));
 sg13g2_antennanp ANTENNA_1516 (.A(net827));
 sg13g2_antennanp ANTENNA_1517 (.A(net827));
 sg13g2_antennanp ANTENNA_1518 (.A(net827));
 sg13g2_antennanp ANTENNA_1519 (.A(net827));
 sg13g2_antennanp ANTENNA_1520 (.A(net827));
 sg13g2_antennanp ANTENNA_1521 (.A(net827));
 sg13g2_antennanp ANTENNA_1522 (.A(net827));
 sg13g2_antennanp ANTENNA_1523 (.A(net831));
 sg13g2_antennanp ANTENNA_1524 (.A(net831));
 sg13g2_antennanp ANTENNA_1525 (.A(net831));
 sg13g2_antennanp ANTENNA_1526 (.A(net831));
 sg13g2_antennanp ANTENNA_1527 (.A(net831));
 sg13g2_antennanp ANTENNA_1528 (.A(net831));
 sg13g2_antennanp ANTENNA_1529 (.A(net831));
 sg13g2_antennanp ANTENNA_1530 (.A(net831));
 sg13g2_antennanp ANTENNA_1531 (.A(net831));
 sg13g2_antennanp ANTENNA_1532 (.A(net834));
 sg13g2_antennanp ANTENNA_1533 (.A(net834));
 sg13g2_antennanp ANTENNA_1534 (.A(net834));
 sg13g2_antennanp ANTENNA_1535 (.A(net834));
 sg13g2_antennanp ANTENNA_1536 (.A(net834));
 sg13g2_antennanp ANTENNA_1537 (.A(net834));
 sg13g2_antennanp ANTENNA_1538 (.A(net834));
 sg13g2_antennanp ANTENNA_1539 (.A(net834));
 sg13g2_antennanp ANTENNA_1540 (.A(net834));
 sg13g2_antennanp ANTENNA_1541 (.A(net836));
 sg13g2_antennanp ANTENNA_1542 (.A(net836));
 sg13g2_antennanp ANTENNA_1543 (.A(net836));
 sg13g2_antennanp ANTENNA_1544 (.A(net836));
 sg13g2_antennanp ANTENNA_1545 (.A(net836));
 sg13g2_antennanp ANTENNA_1546 (.A(net836));
 sg13g2_antennanp ANTENNA_1547 (.A(net836));
 sg13g2_antennanp ANTENNA_1548 (.A(net836));
 sg13g2_antennanp ANTENNA_1549 (.A(net836));
 sg13g2_antennanp ANTENNA_1550 (.A(net837));
 sg13g2_antennanp ANTENNA_1551 (.A(net837));
 sg13g2_antennanp ANTENNA_1552 (.A(net837));
 sg13g2_antennanp ANTENNA_1553 (.A(net837));
 sg13g2_antennanp ANTENNA_1554 (.A(net837));
 sg13g2_antennanp ANTENNA_1555 (.A(net837));
 sg13g2_antennanp ANTENNA_1556 (.A(net837));
 sg13g2_antennanp ANTENNA_1557 (.A(net837));
 sg13g2_antennanp ANTENNA_1558 (.A(net837));
 sg13g2_antennanp ANTENNA_1559 (.A(net871));
 sg13g2_antennanp ANTENNA_1560 (.A(net871));
 sg13g2_antennanp ANTENNA_1561 (.A(net871));
 sg13g2_antennanp ANTENNA_1562 (.A(net871));
 sg13g2_antennanp ANTENNA_1563 (.A(net871));
 sg13g2_antennanp ANTENNA_1564 (.A(net871));
 sg13g2_antennanp ANTENNA_1565 (.A(net871));
 sg13g2_antennanp ANTENNA_1566 (.A(net871));
 sg13g2_antennanp ANTENNA_1567 (.A(net871));
 sg13g2_antennanp ANTENNA_1568 (.A(net953));
 sg13g2_antennanp ANTENNA_1569 (.A(net953));
 sg13g2_antennanp ANTENNA_1570 (.A(net953));
 sg13g2_antennanp ANTENNA_1571 (.A(net953));
 sg13g2_antennanp ANTENNA_1572 (.A(net953));
 sg13g2_antennanp ANTENNA_1573 (.A(net953));
 sg13g2_antennanp ANTENNA_1574 (.A(net953));
 sg13g2_antennanp ANTENNA_1575 (.A(net953));
 sg13g2_antennanp ANTENNA_1576 (.A(net953));
 sg13g2_antennanp ANTENNA_1577 (.A(net953));
 sg13g2_antennanp ANTENNA_1578 (.A(net953));
 sg13g2_antennanp ANTENNA_1579 (.A(net953));
 sg13g2_antennanp ANTENNA_1580 (.A(net953));
 sg13g2_antennanp ANTENNA_1581 (.A(net953));
 sg13g2_antennanp ANTENNA_1582 (.A(net967));
 sg13g2_antennanp ANTENNA_1583 (.A(net967));
 sg13g2_antennanp ANTENNA_1584 (.A(net967));
 sg13g2_antennanp ANTENNA_1585 (.A(net967));
 sg13g2_antennanp ANTENNA_1586 (.A(net967));
 sg13g2_antennanp ANTENNA_1587 (.A(net967));
 sg13g2_antennanp ANTENNA_1588 (.A(net967));
 sg13g2_antennanp ANTENNA_1589 (.A(net967));
 sg13g2_antennanp ANTENNA_1590 (.A(net967));
 sg13g2_antennanp ANTENNA_1591 (.A(net967));
 sg13g2_antennanp ANTENNA_1592 (.A(net967));
 sg13g2_antennanp ANTENNA_1593 (.A(net967));
 sg13g2_antennanp ANTENNA_1594 (.A(net967));
 sg13g2_antennanp ANTENNA_1595 (.A(net967));
 sg13g2_antennanp ANTENNA_1596 (.A(net967));
 sg13g2_antennanp ANTENNA_1597 (.A(net967));
 sg13g2_antennanp ANTENNA_1598 (.A(net968));
 sg13g2_antennanp ANTENNA_1599 (.A(net968));
 sg13g2_antennanp ANTENNA_1600 (.A(net968));
 sg13g2_antennanp ANTENNA_1601 (.A(net968));
 sg13g2_antennanp ANTENNA_1602 (.A(net968));
 sg13g2_antennanp ANTENNA_1603 (.A(net968));
 sg13g2_antennanp ANTENNA_1604 (.A(net968));
 sg13g2_antennanp ANTENNA_1605 (.A(net968));
 sg13g2_antennanp ANTENNA_1606 (.A(net968));
 sg13g2_antennanp ANTENNA_1607 (.A(net981));
 sg13g2_antennanp ANTENNA_1608 (.A(net981));
 sg13g2_antennanp ANTENNA_1609 (.A(net981));
 sg13g2_antennanp ANTENNA_1610 (.A(net981));
 sg13g2_antennanp ANTENNA_1611 (.A(net981));
 sg13g2_antennanp ANTENNA_1612 (.A(net981));
 sg13g2_antennanp ANTENNA_1613 (.A(net981));
 sg13g2_antennanp ANTENNA_1614 (.A(net981));
 sg13g2_antennanp ANTENNA_1615 (.A(net981));
 sg13g2_antennanp ANTENNA_1616 (.A(net994));
 sg13g2_antennanp ANTENNA_1617 (.A(net994));
 sg13g2_antennanp ANTENNA_1618 (.A(net994));
 sg13g2_antennanp ANTENNA_1619 (.A(net994));
 sg13g2_antennanp ANTENNA_1620 (.A(net994));
 sg13g2_antennanp ANTENNA_1621 (.A(net994));
 sg13g2_antennanp ANTENNA_1622 (.A(net994));
 sg13g2_antennanp ANTENNA_1623 (.A(net994));
 sg13g2_antennanp ANTENNA_1624 (.A(net994));
 sg13g2_antennanp ANTENNA_1625 (.A(net1022));
 sg13g2_antennanp ANTENNA_1626 (.A(net1022));
 sg13g2_antennanp ANTENNA_1627 (.A(net1022));
 sg13g2_antennanp ANTENNA_1628 (.A(net1022));
 sg13g2_antennanp ANTENNA_1629 (.A(net1022));
 sg13g2_antennanp ANTENNA_1630 (.A(net1022));
 sg13g2_antennanp ANTENNA_1631 (.A(net1022));
 sg13g2_antennanp ANTENNA_1632 (.A(net1022));
 sg13g2_antennanp ANTENNA_1633 (.A(net1022));
 sg13g2_antennanp ANTENNA_1634 (.A(net1022));
 sg13g2_antennanp ANTENNA_1635 (.A(net1022));
 sg13g2_antennanp ANTENNA_1636 (.A(net1022));
 sg13g2_antennanp ANTENNA_1637 (.A(net1022));
 sg13g2_antennanp ANTENNA_1638 (.A(net1022));
 sg13g2_antennanp ANTENNA_1639 (.A(net1022));
 sg13g2_antennanp ANTENNA_1640 (.A(net1022));
 sg13g2_antennanp ANTENNA_1641 (.A(net1057));
 sg13g2_antennanp ANTENNA_1642 (.A(net1057));
 sg13g2_antennanp ANTENNA_1643 (.A(net1057));
 sg13g2_antennanp ANTENNA_1644 (.A(net1057));
 sg13g2_antennanp ANTENNA_1645 (.A(net1057));
 sg13g2_antennanp ANTENNA_1646 (.A(net1057));
 sg13g2_antennanp ANTENNA_1647 (.A(net1057));
 sg13g2_antennanp ANTENNA_1648 (.A(net1057));
 sg13g2_antennanp ANTENNA_1649 (.A(net1057));
 sg13g2_antennanp ANTENNA_1650 (.A(net1057));
 sg13g2_antennanp ANTENNA_1651 (.A(net1057));
 sg13g2_antennanp ANTENNA_1652 (.A(net1057));
 sg13g2_antennanp ANTENNA_1653 (.A(net1057));
 sg13g2_antennanp ANTENNA_1654 (.A(net1057));
 sg13g2_antennanp ANTENNA_1655 (.A(net1057));
 sg13g2_antennanp ANTENNA_1656 (.A(net1057));
 sg13g2_antennanp ANTENNA_1657 (.A(net1057));
 sg13g2_antennanp ANTENNA_1658 (.A(net1057));
 sg13g2_antennanp ANTENNA_1659 (.A(net1057));
 sg13g2_antennanp ANTENNA_1660 (.A(net1057));
 sg13g2_antennanp ANTENNA_1661 (.A(net1057));
 sg13g2_antennanp ANTENNA_1662 (.A(net1057));
 sg13g2_antennanp ANTENNA_1663 (.A(net1057));
 sg13g2_antennanp ANTENNA_1664 (.A(net1057));
 sg13g2_antennanp ANTENNA_1665 (.A(net1057));
 sg13g2_antennanp ANTENNA_1666 (.A(net1057));
 sg13g2_antennanp ANTENNA_1667 (.A(net1057));
 sg13g2_antennanp ANTENNA_1668 (.A(net1057));
 sg13g2_antennanp ANTENNA_1669 (.A(net1057));
 sg13g2_antennanp ANTENNA_1670 (.A(net1057));
 sg13g2_antennanp ANTENNA_1671 (.A(net1057));
 sg13g2_antennanp ANTENNA_1672 (.A(net1057));
 sg13g2_antennanp ANTENNA_1673 (.A(net1057));
 sg13g2_antennanp ANTENNA_1674 (.A(net1057));
 sg13g2_antennanp ANTENNA_1675 (.A(net1057));
 sg13g2_antennanp ANTENNA_1676 (.A(net1057));
 sg13g2_antennanp ANTENNA_1677 (.A(net1057));
 sg13g2_antennanp ANTENNA_1678 (.A(net1057));
 sg13g2_antennanp ANTENNA_1679 (.A(net1057));
 sg13g2_antennanp ANTENNA_1680 (.A(net1057));
 sg13g2_antennanp ANTENNA_1681 (.A(net1057));
 sg13g2_antennanp ANTENNA_1682 (.A(net1057));
 sg13g2_antennanp ANTENNA_1683 (.A(net1057));
 sg13g2_antennanp ANTENNA_1684 (.A(net1057));
 sg13g2_antennanp ANTENNA_1685 (.A(net1075));
 sg13g2_antennanp ANTENNA_1686 (.A(net1075));
 sg13g2_antennanp ANTENNA_1687 (.A(net1075));
 sg13g2_antennanp ANTENNA_1688 (.A(net1075));
 sg13g2_antennanp ANTENNA_1689 (.A(net1075));
 sg13g2_antennanp ANTENNA_1690 (.A(net1075));
 sg13g2_antennanp ANTENNA_1691 (.A(net1075));
 sg13g2_antennanp ANTENNA_1692 (.A(net1075));
 sg13g2_antennanp ANTENNA_1693 (.A(net1075));
 sg13g2_antennanp ANTENNA_1694 (.A(net1085));
 sg13g2_antennanp ANTENNA_1695 (.A(net1085));
 sg13g2_antennanp ANTENNA_1696 (.A(net1085));
 sg13g2_antennanp ANTENNA_1697 (.A(net1085));
 sg13g2_antennanp ANTENNA_1698 (.A(net1085));
 sg13g2_antennanp ANTENNA_1699 (.A(net1085));
 sg13g2_antennanp ANTENNA_1700 (.A(net1085));
 sg13g2_antennanp ANTENNA_1701 (.A(net1085));
 sg13g2_antennanp ANTENNA_1702 (.A(net1085));
 sg13g2_antennanp ANTENNA_1703 (.A(net1085));
 sg13g2_antennanp ANTENNA_1704 (.A(net1085));
 sg13g2_antennanp ANTENNA_1705 (.A(net1085));
 sg13g2_antennanp ANTENNA_1706 (.A(net1085));
 sg13g2_antennanp ANTENNA_1707 (.A(net1096));
 sg13g2_antennanp ANTENNA_1708 (.A(net1096));
 sg13g2_antennanp ANTENNA_1709 (.A(net1096));
 sg13g2_antennanp ANTENNA_1710 (.A(net1096));
 sg13g2_antennanp ANTENNA_1711 (.A(net1096));
 sg13g2_antennanp ANTENNA_1712 (.A(net1096));
 sg13g2_antennanp ANTENNA_1713 (.A(net1096));
 sg13g2_antennanp ANTENNA_1714 (.A(net1096));
 sg13g2_antennanp ANTENNA_1715 (.A(net1096));
 sg13g2_antennanp ANTENNA_1716 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1717 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1718 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1719 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1720 (.A(_01057_));
 sg13g2_antennanp ANTENNA_1721 (.A(_01057_));
 sg13g2_antennanp ANTENNA_1722 (.A(_01071_));
 sg13g2_antennanp ANTENNA_1723 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1724 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1725 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1726 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1727 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1728 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1729 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1730 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1731 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1732 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1733 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1734 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1735 (.A(_02855_));
 sg13g2_antennanp ANTENNA_1736 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1737 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1738 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1739 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1740 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1741 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1742 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1743 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1744 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1745 (.A(_02856_));
 sg13g2_antennanp ANTENNA_1746 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1747 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1748 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1749 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1750 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1751 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1752 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1753 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1754 (.A(_02866_));
 sg13g2_antennanp ANTENNA_1755 (.A(_02873_));
 sg13g2_antennanp ANTENNA_1756 (.A(_02873_));
 sg13g2_antennanp ANTENNA_1757 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1758 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1759 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1760 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1761 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1762 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1763 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1764 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1765 (.A(_02877_));
 sg13g2_antennanp ANTENNA_1766 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1767 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1768 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1769 (.A(_03350_));
 sg13g2_antennanp ANTENNA_1770 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1771 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1772 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1773 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1774 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1775 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1776 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1777 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1778 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1779 (.A(_03356_));
 sg13g2_antennanp ANTENNA_1780 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1781 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1782 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1783 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1784 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1785 (.A(_03612_));
 sg13g2_antennanp ANTENNA_1786 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1787 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1788 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1789 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1790 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1791 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1792 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1793 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1794 (.A(_04628_));
 sg13g2_antennanp ANTENNA_1795 (.A(_04646_));
 sg13g2_antennanp ANTENNA_1796 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1797 (.A(_05022_));
 sg13g2_antennanp ANTENNA_1798 (.A(_05046_));
 sg13g2_antennanp ANTENNA_1799 (.A(_05581_));
 sg13g2_antennanp ANTENNA_1800 (.A(_05584_));
 sg13g2_antennanp ANTENNA_1801 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1802 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1803 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1804 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1805 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1806 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1807 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1808 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1809 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1810 (.A(_05644_));
 sg13g2_antennanp ANTENNA_1811 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1812 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1813 (.A(_06275_));
 sg13g2_antennanp ANTENNA_1814 (.A(_07137_));
 sg13g2_antennanp ANTENNA_1815 (.A(_07138_));
 sg13g2_antennanp ANTENNA_1816 (.A(_07166_));
 sg13g2_antennanp ANTENNA_1817 (.A(_07166_));
 sg13g2_antennanp ANTENNA_1818 (.A(_07222_));
 sg13g2_antennanp ANTENNA_1819 (.A(_07326_));
 sg13g2_antennanp ANTENNA_1820 (.A(_07326_));
 sg13g2_antennanp ANTENNA_1821 (.A(_07976_));
 sg13g2_antennanp ANTENNA_1822 (.A(_07976_));
 sg13g2_antennanp ANTENNA_1823 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1824 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1825 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1826 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1827 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1828 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1829 (.A(_08081_));
 sg13g2_antennanp ANTENNA_1830 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1831 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1832 (.A(_08087_));
 sg13g2_antennanp ANTENNA_1833 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1834 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1835 (.A(_08092_));
 sg13g2_antennanp ANTENNA_1836 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1837 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1838 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1839 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1840 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1841 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1842 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1843 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1844 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1845 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1846 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1847 (.A(_08257_));
 sg13g2_antennanp ANTENNA_1848 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1849 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1850 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1851 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1852 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1853 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1854 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1855 (.A(_08403_));
 sg13g2_antennanp ANTENNA_1856 (.A(_08517_));
 sg13g2_antennanp ANTENNA_1857 (.A(_08556_));
 sg13g2_antennanp ANTENNA_1858 (.A(_08614_));
 sg13g2_antennanp ANTENNA_1859 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1860 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1861 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1862 (.A(_08620_));
 sg13g2_antennanp ANTENNA_1863 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1864 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1865 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1866 (.A(_08947_));
 sg13g2_antennanp ANTENNA_1867 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1868 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1869 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1870 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1871 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1872 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1873 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1874 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1875 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1876 (.A(_08951_));
 sg13g2_antennanp ANTENNA_1877 (.A(_08993_));
 sg13g2_antennanp ANTENNA_1878 (.A(_09005_));
 sg13g2_antennanp ANTENNA_1879 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1880 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1881 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1882 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1883 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1884 (.A(_09030_));
 sg13g2_antennanp ANTENNA_1885 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1886 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1887 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1888 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1889 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1890 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1891 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1892 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1893 (.A(_09039_));
 sg13g2_antennanp ANTENNA_1894 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1895 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1896 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1897 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1898 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1899 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1900 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1901 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1902 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1903 (.A(_09234_));
 sg13g2_antennanp ANTENNA_1904 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1905 (.A(_09284_));
 sg13g2_antennanp ANTENNA_1906 (.A(_09305_));
 sg13g2_antennanp ANTENNA_1907 (.A(_09328_));
 sg13g2_antennanp ANTENNA_1908 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1909 (.A(_09370_));
 sg13g2_antennanp ANTENNA_1910 (.A(_09394_));
 sg13g2_antennanp ANTENNA_1911 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1912 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1913 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1914 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1915 (.A(_09470_));
 sg13g2_antennanp ANTENNA_1916 (.A(_09526_));
 sg13g2_antennanp ANTENNA_1917 (.A(_09553_));
 sg13g2_antennanp ANTENNA_1918 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1919 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1920 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1921 (.A(_09591_));
 sg13g2_antennanp ANTENNA_1922 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1923 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1924 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1925 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1926 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1927 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1928 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1929 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1930 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1931 (.A(_09869_));
 sg13g2_antennanp ANTENNA_1932 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1933 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1934 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1935 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1936 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1937 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1938 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1939 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1940 (.A(_09880_));
 sg13g2_antennanp ANTENNA_1941 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1942 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1943 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1944 (.A(_09882_));
 sg13g2_antennanp ANTENNA_1945 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1946 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1947 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1948 (.A(_10156_));
 sg13g2_antennanp ANTENNA_1949 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1950 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1951 (.A(_10241_));
 sg13g2_antennanp ANTENNA_1952 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1953 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1954 (.A(_10482_));
 sg13g2_antennanp ANTENNA_1955 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1956 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1957 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1958 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1959 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1960 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1961 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1962 (.A(_10576_));
 sg13g2_antennanp ANTENNA_1963 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1964 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1965 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1966 (.A(_10653_));
 sg13g2_antennanp ANTENNA_1967 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1968 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1969 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1970 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1971 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1972 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1973 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1974 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1975 (.A(_10892_));
 sg13g2_antennanp ANTENNA_1976 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1977 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1978 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1979 (.A(_11550_));
 sg13g2_antennanp ANTENNA_1980 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1981 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1982 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1983 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1984 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1985 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1986 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1987 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1988 (.A(_11613_));
 sg13g2_antennanp ANTENNA_1989 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1990 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1991 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1992 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1993 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1994 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1995 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1996 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1997 (.A(_11688_));
 sg13g2_antennanp ANTENNA_1998 (.A(_11695_));
 sg13g2_antennanp ANTENNA_1999 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2000 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2001 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2002 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2003 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2004 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2005 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2006 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2007 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2008 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2009 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2010 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2011 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2012 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2013 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2014 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2015 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2016 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2017 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2018 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2019 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2020 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2021 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2022 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2023 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2024 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2025 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2026 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2027 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2028 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2029 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2030 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2031 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2032 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2033 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2034 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2035 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2036 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2037 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2038 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2039 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2040 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2041 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2042 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2043 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2044 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2045 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2046 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2047 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2048 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2049 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2050 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2051 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2052 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2053 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2054 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2055 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2056 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2057 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2058 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2059 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2060 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2061 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2062 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2063 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2064 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2065 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2066 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2067 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2068 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2069 (.A(\cpu.addr[14] ));
 sg13g2_antennanp ANTENNA_2070 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2071 (.A(net3));
 sg13g2_antennanp ANTENNA_2072 (.A(net3));
 sg13g2_antennanp ANTENNA_2073 (.A(net3));
 sg13g2_antennanp ANTENNA_2074 (.A(net11));
 sg13g2_antennanp ANTENNA_2075 (.A(net11));
 sg13g2_antennanp ANTENNA_2076 (.A(net11));
 sg13g2_antennanp ANTENNA_2077 (.A(net12));
 sg13g2_antennanp ANTENNA_2078 (.A(net12));
 sg13g2_antennanp ANTENNA_2079 (.A(net12));
 sg13g2_antennanp ANTENNA_2080 (.A(net14));
 sg13g2_antennanp ANTENNA_2081 (.A(net14));
 sg13g2_antennanp ANTENNA_2082 (.A(net14));
 sg13g2_antennanp ANTENNA_2083 (.A(net18));
 sg13g2_antennanp ANTENNA_2084 (.A(net18));
 sg13g2_antennanp ANTENNA_2085 (.A(net19));
 sg13g2_antennanp ANTENNA_2086 (.A(net19));
 sg13g2_antennanp ANTENNA_2087 (.A(net19));
 sg13g2_antennanp ANTENNA_2088 (.A(net20));
 sg13g2_antennanp ANTENNA_2089 (.A(net20));
 sg13g2_antennanp ANTENNA_2090 (.A(net20));
 sg13g2_antennanp ANTENNA_2091 (.A(net464));
 sg13g2_antennanp ANTENNA_2092 (.A(net464));
 sg13g2_antennanp ANTENNA_2093 (.A(net464));
 sg13g2_antennanp ANTENNA_2094 (.A(net464));
 sg13g2_antennanp ANTENNA_2095 (.A(net464));
 sg13g2_antennanp ANTENNA_2096 (.A(net464));
 sg13g2_antennanp ANTENNA_2097 (.A(net464));
 sg13g2_antennanp ANTENNA_2098 (.A(net464));
 sg13g2_antennanp ANTENNA_2099 (.A(net464));
 sg13g2_antennanp ANTENNA_2100 (.A(net464));
 sg13g2_antennanp ANTENNA_2101 (.A(net464));
 sg13g2_antennanp ANTENNA_2102 (.A(net464));
 sg13g2_antennanp ANTENNA_2103 (.A(net464));
 sg13g2_antennanp ANTENNA_2104 (.A(net464));
 sg13g2_antennanp ANTENNA_2105 (.A(net464));
 sg13g2_antennanp ANTENNA_2106 (.A(net464));
 sg13g2_antennanp ANTENNA_2107 (.A(net464));
 sg13g2_antennanp ANTENNA_2108 (.A(net464));
 sg13g2_antennanp ANTENNA_2109 (.A(net464));
 sg13g2_antennanp ANTENNA_2110 (.A(net464));
 sg13g2_antennanp ANTENNA_2111 (.A(net498));
 sg13g2_antennanp ANTENNA_2112 (.A(net498));
 sg13g2_antennanp ANTENNA_2113 (.A(net498));
 sg13g2_antennanp ANTENNA_2114 (.A(net498));
 sg13g2_antennanp ANTENNA_2115 (.A(net498));
 sg13g2_antennanp ANTENNA_2116 (.A(net498));
 sg13g2_antennanp ANTENNA_2117 (.A(net498));
 sg13g2_antennanp ANTENNA_2118 (.A(net498));
 sg13g2_antennanp ANTENNA_2119 (.A(net498));
 sg13g2_antennanp ANTENNA_2120 (.A(net573));
 sg13g2_antennanp ANTENNA_2121 (.A(net573));
 sg13g2_antennanp ANTENNA_2122 (.A(net573));
 sg13g2_antennanp ANTENNA_2123 (.A(net573));
 sg13g2_antennanp ANTENNA_2124 (.A(net573));
 sg13g2_antennanp ANTENNA_2125 (.A(net573));
 sg13g2_antennanp ANTENNA_2126 (.A(net573));
 sg13g2_antennanp ANTENNA_2127 (.A(net573));
 sg13g2_antennanp ANTENNA_2128 (.A(net573));
 sg13g2_antennanp ANTENNA_2129 (.A(net573));
 sg13g2_antennanp ANTENNA_2130 (.A(net573));
 sg13g2_antennanp ANTENNA_2131 (.A(net573));
 sg13g2_antennanp ANTENNA_2132 (.A(net573));
 sg13g2_antennanp ANTENNA_2133 (.A(net573));
 sg13g2_antennanp ANTENNA_2134 (.A(net573));
 sg13g2_antennanp ANTENNA_2135 (.A(net573));
 sg13g2_antennanp ANTENNA_2136 (.A(net573));
 sg13g2_antennanp ANTENNA_2137 (.A(net573));
 sg13g2_antennanp ANTENNA_2138 (.A(net573));
 sg13g2_antennanp ANTENNA_2139 (.A(net573));
 sg13g2_antennanp ANTENNA_2140 (.A(net576));
 sg13g2_antennanp ANTENNA_2141 (.A(net576));
 sg13g2_antennanp ANTENNA_2142 (.A(net576));
 sg13g2_antennanp ANTENNA_2143 (.A(net576));
 sg13g2_antennanp ANTENNA_2144 (.A(net576));
 sg13g2_antennanp ANTENNA_2145 (.A(net576));
 sg13g2_antennanp ANTENNA_2146 (.A(net576));
 sg13g2_antennanp ANTENNA_2147 (.A(net576));
 sg13g2_antennanp ANTENNA_2148 (.A(net576));
 sg13g2_antennanp ANTENNA_2149 (.A(net576));
 sg13g2_antennanp ANTENNA_2150 (.A(net576));
 sg13g2_antennanp ANTENNA_2151 (.A(net576));
 sg13g2_antennanp ANTENNA_2152 (.A(net576));
 sg13g2_antennanp ANTENNA_2153 (.A(net576));
 sg13g2_antennanp ANTENNA_2154 (.A(net576));
 sg13g2_antennanp ANTENNA_2155 (.A(net576));
 sg13g2_antennanp ANTENNA_2156 (.A(net576));
 sg13g2_antennanp ANTENNA_2157 (.A(net576));
 sg13g2_antennanp ANTENNA_2158 (.A(net576));
 sg13g2_antennanp ANTENNA_2159 (.A(net576));
 sg13g2_antennanp ANTENNA_2160 (.A(net714));
 sg13g2_antennanp ANTENNA_2161 (.A(net714));
 sg13g2_antennanp ANTENNA_2162 (.A(net714));
 sg13g2_antennanp ANTENNA_2163 (.A(net714));
 sg13g2_antennanp ANTENNA_2164 (.A(net714));
 sg13g2_antennanp ANTENNA_2165 (.A(net714));
 sg13g2_antennanp ANTENNA_2166 (.A(net714));
 sg13g2_antennanp ANTENNA_2167 (.A(net714));
 sg13g2_antennanp ANTENNA_2168 (.A(net714));
 sg13g2_antennanp ANTENNA_2169 (.A(net716));
 sg13g2_antennanp ANTENNA_2170 (.A(net716));
 sg13g2_antennanp ANTENNA_2171 (.A(net716));
 sg13g2_antennanp ANTENNA_2172 (.A(net716));
 sg13g2_antennanp ANTENNA_2173 (.A(net716));
 sg13g2_antennanp ANTENNA_2174 (.A(net716));
 sg13g2_antennanp ANTENNA_2175 (.A(net716));
 sg13g2_antennanp ANTENNA_2176 (.A(net716));
 sg13g2_antennanp ANTENNA_2177 (.A(net716));
 sg13g2_antennanp ANTENNA_2178 (.A(net747));
 sg13g2_antennanp ANTENNA_2179 (.A(net747));
 sg13g2_antennanp ANTENNA_2180 (.A(net747));
 sg13g2_antennanp ANTENNA_2181 (.A(net747));
 sg13g2_antennanp ANTENNA_2182 (.A(net747));
 sg13g2_antennanp ANTENNA_2183 (.A(net747));
 sg13g2_antennanp ANTENNA_2184 (.A(net747));
 sg13g2_antennanp ANTENNA_2185 (.A(net747));
 sg13g2_antennanp ANTENNA_2186 (.A(net760));
 sg13g2_antennanp ANTENNA_2187 (.A(net760));
 sg13g2_antennanp ANTENNA_2188 (.A(net760));
 sg13g2_antennanp ANTENNA_2189 (.A(net760));
 sg13g2_antennanp ANTENNA_2190 (.A(net760));
 sg13g2_antennanp ANTENNA_2191 (.A(net760));
 sg13g2_antennanp ANTENNA_2192 (.A(net760));
 sg13g2_antennanp ANTENNA_2193 (.A(net760));
 sg13g2_antennanp ANTENNA_2194 (.A(net834));
 sg13g2_antennanp ANTENNA_2195 (.A(net834));
 sg13g2_antennanp ANTENNA_2196 (.A(net834));
 sg13g2_antennanp ANTENNA_2197 (.A(net834));
 sg13g2_antennanp ANTENNA_2198 (.A(net834));
 sg13g2_antennanp ANTENNA_2199 (.A(net834));
 sg13g2_antennanp ANTENNA_2200 (.A(net834));
 sg13g2_antennanp ANTENNA_2201 (.A(net834));
 sg13g2_antennanp ANTENNA_2202 (.A(net834));
 sg13g2_antennanp ANTENNA_2203 (.A(net836));
 sg13g2_antennanp ANTENNA_2204 (.A(net836));
 sg13g2_antennanp ANTENNA_2205 (.A(net836));
 sg13g2_antennanp ANTENNA_2206 (.A(net836));
 sg13g2_antennanp ANTENNA_2207 (.A(net836));
 sg13g2_antennanp ANTENNA_2208 (.A(net836));
 sg13g2_antennanp ANTENNA_2209 (.A(net836));
 sg13g2_antennanp ANTENNA_2210 (.A(net836));
 sg13g2_antennanp ANTENNA_2211 (.A(net836));
 sg13g2_antennanp ANTENNA_2212 (.A(net837));
 sg13g2_antennanp ANTENNA_2213 (.A(net837));
 sg13g2_antennanp ANTENNA_2214 (.A(net837));
 sg13g2_antennanp ANTENNA_2215 (.A(net837));
 sg13g2_antennanp ANTENNA_2216 (.A(net837));
 sg13g2_antennanp ANTENNA_2217 (.A(net837));
 sg13g2_antennanp ANTENNA_2218 (.A(net837));
 sg13g2_antennanp ANTENNA_2219 (.A(net837));
 sg13g2_antennanp ANTENNA_2220 (.A(net837));
 sg13g2_antennanp ANTENNA_2221 (.A(net871));
 sg13g2_antennanp ANTENNA_2222 (.A(net871));
 sg13g2_antennanp ANTENNA_2223 (.A(net871));
 sg13g2_antennanp ANTENNA_2224 (.A(net871));
 sg13g2_antennanp ANTENNA_2225 (.A(net871));
 sg13g2_antennanp ANTENNA_2226 (.A(net871));
 sg13g2_antennanp ANTENNA_2227 (.A(net871));
 sg13g2_antennanp ANTENNA_2228 (.A(net871));
 sg13g2_antennanp ANTENNA_2229 (.A(net871));
 sg13g2_antennanp ANTENNA_2230 (.A(net953));
 sg13g2_antennanp ANTENNA_2231 (.A(net953));
 sg13g2_antennanp ANTENNA_2232 (.A(net953));
 sg13g2_antennanp ANTENNA_2233 (.A(net953));
 sg13g2_antennanp ANTENNA_2234 (.A(net953));
 sg13g2_antennanp ANTENNA_2235 (.A(net953));
 sg13g2_antennanp ANTENNA_2236 (.A(net953));
 sg13g2_antennanp ANTENNA_2237 (.A(net953));
 sg13g2_antennanp ANTENNA_2238 (.A(net953));
 sg13g2_antennanp ANTENNA_2239 (.A(net958));
 sg13g2_antennanp ANTENNA_2240 (.A(net958));
 sg13g2_antennanp ANTENNA_2241 (.A(net958));
 sg13g2_antennanp ANTENNA_2242 (.A(net958));
 sg13g2_antennanp ANTENNA_2243 (.A(net958));
 sg13g2_antennanp ANTENNA_2244 (.A(net958));
 sg13g2_antennanp ANTENNA_2245 (.A(net958));
 sg13g2_antennanp ANTENNA_2246 (.A(net958));
 sg13g2_antennanp ANTENNA_2247 (.A(net967));
 sg13g2_antennanp ANTENNA_2248 (.A(net967));
 sg13g2_antennanp ANTENNA_2249 (.A(net967));
 sg13g2_antennanp ANTENNA_2250 (.A(net967));
 sg13g2_antennanp ANTENNA_2251 (.A(net967));
 sg13g2_antennanp ANTENNA_2252 (.A(net967));
 sg13g2_antennanp ANTENNA_2253 (.A(net967));
 sg13g2_antennanp ANTENNA_2254 (.A(net967));
 sg13g2_antennanp ANTENNA_2255 (.A(net967));
 sg13g2_antennanp ANTENNA_2256 (.A(net968));
 sg13g2_antennanp ANTENNA_2257 (.A(net968));
 sg13g2_antennanp ANTENNA_2258 (.A(net968));
 sg13g2_antennanp ANTENNA_2259 (.A(net968));
 sg13g2_antennanp ANTENNA_2260 (.A(net968));
 sg13g2_antennanp ANTENNA_2261 (.A(net968));
 sg13g2_antennanp ANTENNA_2262 (.A(net968));
 sg13g2_antennanp ANTENNA_2263 (.A(net968));
 sg13g2_antennanp ANTENNA_2264 (.A(net968));
 sg13g2_antennanp ANTENNA_2265 (.A(net981));
 sg13g2_antennanp ANTENNA_2266 (.A(net981));
 sg13g2_antennanp ANTENNA_2267 (.A(net981));
 sg13g2_antennanp ANTENNA_2268 (.A(net981));
 sg13g2_antennanp ANTENNA_2269 (.A(net981));
 sg13g2_antennanp ANTENNA_2270 (.A(net981));
 sg13g2_antennanp ANTENNA_2271 (.A(net981));
 sg13g2_antennanp ANTENNA_2272 (.A(net981));
 sg13g2_antennanp ANTENNA_2273 (.A(net981));
 sg13g2_antennanp ANTENNA_2274 (.A(net994));
 sg13g2_antennanp ANTENNA_2275 (.A(net994));
 sg13g2_antennanp ANTENNA_2276 (.A(net994));
 sg13g2_antennanp ANTENNA_2277 (.A(net994));
 sg13g2_antennanp ANTENNA_2278 (.A(net994));
 sg13g2_antennanp ANTENNA_2279 (.A(net994));
 sg13g2_antennanp ANTENNA_2280 (.A(net994));
 sg13g2_antennanp ANTENNA_2281 (.A(net994));
 sg13g2_antennanp ANTENNA_2282 (.A(net994));
 sg13g2_antennanp ANTENNA_2283 (.A(net1022));
 sg13g2_antennanp ANTENNA_2284 (.A(net1022));
 sg13g2_antennanp ANTENNA_2285 (.A(net1022));
 sg13g2_antennanp ANTENNA_2286 (.A(net1022));
 sg13g2_antennanp ANTENNA_2287 (.A(net1022));
 sg13g2_antennanp ANTENNA_2288 (.A(net1022));
 sg13g2_antennanp ANTENNA_2289 (.A(net1022));
 sg13g2_antennanp ANTENNA_2290 (.A(net1022));
 sg13g2_antennanp ANTENNA_2291 (.A(net1022));
 sg13g2_antennanp ANTENNA_2292 (.A(net1022));
 sg13g2_antennanp ANTENNA_2293 (.A(net1022));
 sg13g2_antennanp ANTENNA_2294 (.A(net1022));
 sg13g2_antennanp ANTENNA_2295 (.A(net1022));
 sg13g2_antennanp ANTENNA_2296 (.A(net1022));
 sg13g2_antennanp ANTENNA_2297 (.A(net1022));
 sg13g2_antennanp ANTENNA_2298 (.A(net1022));
 sg13g2_antennanp ANTENNA_2299 (.A(net1022));
 sg13g2_antennanp ANTENNA_2300 (.A(net1022));
 sg13g2_antennanp ANTENNA_2301 (.A(net1022));
 sg13g2_antennanp ANTENNA_2302 (.A(net1022));
 sg13g2_antennanp ANTENNA_2303 (.A(net1057));
 sg13g2_antennanp ANTENNA_2304 (.A(net1057));
 sg13g2_antennanp ANTENNA_2305 (.A(net1057));
 sg13g2_antennanp ANTENNA_2306 (.A(net1057));
 sg13g2_antennanp ANTENNA_2307 (.A(net1057));
 sg13g2_antennanp ANTENNA_2308 (.A(net1057));
 sg13g2_antennanp ANTENNA_2309 (.A(net1057));
 sg13g2_antennanp ANTENNA_2310 (.A(net1057));
 sg13g2_antennanp ANTENNA_2311 (.A(net1057));
 sg13g2_antennanp ANTENNA_2312 (.A(net1057));
 sg13g2_antennanp ANTENNA_2313 (.A(net1057));
 sg13g2_antennanp ANTENNA_2314 (.A(net1057));
 sg13g2_antennanp ANTENNA_2315 (.A(net1057));
 sg13g2_antennanp ANTENNA_2316 (.A(net1057));
 sg13g2_antennanp ANTENNA_2317 (.A(net1057));
 sg13g2_antennanp ANTENNA_2318 (.A(net1057));
 sg13g2_antennanp ANTENNA_2319 (.A(net1057));
 sg13g2_antennanp ANTENNA_2320 (.A(net1057));
 sg13g2_antennanp ANTENNA_2321 (.A(net1057));
 sg13g2_antennanp ANTENNA_2322 (.A(net1057));
 sg13g2_antennanp ANTENNA_2323 (.A(net1075));
 sg13g2_antennanp ANTENNA_2324 (.A(net1075));
 sg13g2_antennanp ANTENNA_2325 (.A(net1075));
 sg13g2_antennanp ANTENNA_2326 (.A(net1075));
 sg13g2_antennanp ANTENNA_2327 (.A(net1075));
 sg13g2_antennanp ANTENNA_2328 (.A(net1075));
 sg13g2_antennanp ANTENNA_2329 (.A(net1075));
 sg13g2_antennanp ANTENNA_2330 (.A(net1075));
 sg13g2_antennanp ANTENNA_2331 (.A(net1075));
 sg13g2_antennanp ANTENNA_2332 (.A(net1085));
 sg13g2_antennanp ANTENNA_2333 (.A(net1085));
 sg13g2_antennanp ANTENNA_2334 (.A(net1085));
 sg13g2_antennanp ANTENNA_2335 (.A(net1085));
 sg13g2_antennanp ANTENNA_2336 (.A(net1085));
 sg13g2_antennanp ANTENNA_2337 (.A(net1085));
 sg13g2_antennanp ANTENNA_2338 (.A(net1085));
 sg13g2_antennanp ANTENNA_2339 (.A(net1085));
 sg13g2_antennanp ANTENNA_2340 (.A(net1085));
 sg13g2_antennanp ANTENNA_2341 (.A(net1085));
 sg13g2_antennanp ANTENNA_2342 (.A(net1085));
 sg13g2_antennanp ANTENNA_2343 (.A(net1085));
 sg13g2_antennanp ANTENNA_2344 (.A(net1085));
 sg13g2_antennanp ANTENNA_2345 (.A(net1085));
 sg13g2_antennanp ANTENNA_2346 (.A(net1085));
 sg13g2_antennanp ANTENNA_2347 (.A(net1085));
 sg13g2_antennanp ANTENNA_2348 (.A(net1085));
 sg13g2_antennanp ANTENNA_2349 (.A(net1085));
 sg13g2_antennanp ANTENNA_2350 (.A(net1085));
 sg13g2_antennanp ANTENNA_2351 (.A(net1085));
 sg13g2_antennanp ANTENNA_2352 (.A(net1085));
 sg13g2_antennanp ANTENNA_2353 (.A(net1085));
 sg13g2_antennanp ANTENNA_2354 (.A(net1085));
 sg13g2_antennanp ANTENNA_2355 (.A(net1085));
 sg13g2_antennanp ANTENNA_2356 (.A(net1085));
 sg13g2_antennanp ANTENNA_2357 (.A(net1085));
 sg13g2_antennanp ANTENNA_2358 (.A(net1085));
 sg13g2_antennanp ANTENNA_2359 (.A(net1085));
 sg13g2_antennanp ANTENNA_2360 (.A(net1085));
 sg13g2_antennanp ANTENNA_2361 (.A(net1085));
 sg13g2_antennanp ANTENNA_2362 (.A(net1085));
 sg13g2_antennanp ANTENNA_2363 (.A(net1085));
 sg13g2_antennanp ANTENNA_2364 (.A(net1085));
 sg13g2_antennanp ANTENNA_2365 (.A(net1085));
 sg13g2_antennanp ANTENNA_2366 (.A(net1085));
 sg13g2_antennanp ANTENNA_2367 (.A(net1085));
 sg13g2_antennanp ANTENNA_2368 (.A(net1085));
 sg13g2_antennanp ANTENNA_2369 (.A(net1085));
 sg13g2_antennanp ANTENNA_2370 (.A(net1085));
 sg13g2_antennanp ANTENNA_2371 (.A(net1085));
 sg13g2_antennanp ANTENNA_2372 (.A(net1085));
 sg13g2_antennanp ANTENNA_2373 (.A(net1085));
 sg13g2_antennanp ANTENNA_2374 (.A(net1085));
 sg13g2_antennanp ANTENNA_2375 (.A(net1085));
 sg13g2_antennanp ANTENNA_2376 (.A(net1085));
 sg13g2_antennanp ANTENNA_2377 (.A(net1085));
 sg13g2_antennanp ANTENNA_2378 (.A(net1085));
 sg13g2_antennanp ANTENNA_2379 (.A(net1085));
 sg13g2_antennanp ANTENNA_2380 (.A(net1096));
 sg13g2_antennanp ANTENNA_2381 (.A(net1096));
 sg13g2_antennanp ANTENNA_2382 (.A(net1096));
 sg13g2_antennanp ANTENNA_2383 (.A(net1096));
 sg13g2_antennanp ANTENNA_2384 (.A(net1096));
 sg13g2_antennanp ANTENNA_2385 (.A(net1096));
 sg13g2_antennanp ANTENNA_2386 (.A(net1096));
 sg13g2_antennanp ANTENNA_2387 (.A(net1096));
 sg13g2_antennanp ANTENNA_2388 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2389 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2390 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2391 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2392 (.A(_01057_));
 sg13g2_antennanp ANTENNA_2393 (.A(_01057_));
 sg13g2_antennanp ANTENNA_2394 (.A(_01071_));
 sg13g2_antennanp ANTENNA_2395 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2396 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2397 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2398 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2399 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2400 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2401 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2402 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2403 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2404 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2405 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2406 (.A(_02855_));
 sg13g2_antennanp ANTENNA_2407 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2408 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2409 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2410 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2411 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2412 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2413 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2414 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2415 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2416 (.A(_02856_));
 sg13g2_antennanp ANTENNA_2417 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2418 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2419 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2420 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2421 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2422 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2423 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2424 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2425 (.A(_02866_));
 sg13g2_antennanp ANTENNA_2426 (.A(_02873_));
 sg13g2_antennanp ANTENNA_2427 (.A(_02873_));
 sg13g2_antennanp ANTENNA_2428 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2429 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2430 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2431 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2432 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2433 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2434 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2435 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2436 (.A(_02877_));
 sg13g2_antennanp ANTENNA_2437 (.A(_03350_));
 sg13g2_antennanp ANTENNA_2438 (.A(_03350_));
 sg13g2_antennanp ANTENNA_2439 (.A(_03350_));
 sg13g2_antennanp ANTENNA_2440 (.A(_03350_));
 sg13g2_antennanp ANTENNA_2441 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2442 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2443 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2444 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2445 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2446 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2447 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2448 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2449 (.A(_03356_));
 sg13g2_antennanp ANTENNA_2450 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2451 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2452 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2453 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2454 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2455 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2456 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2457 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2458 (.A(_03612_));
 sg13g2_antennanp ANTENNA_2459 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2460 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2461 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2462 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2463 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2464 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2465 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2466 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2467 (.A(_04628_));
 sg13g2_antennanp ANTENNA_2468 (.A(_04646_));
 sg13g2_antennanp ANTENNA_2469 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2470 (.A(_05022_));
 sg13g2_antennanp ANTENNA_2471 (.A(_05046_));
 sg13g2_antennanp ANTENNA_2472 (.A(_05581_));
 sg13g2_antennanp ANTENNA_2473 (.A(_05584_));
 sg13g2_antennanp ANTENNA_2474 (.A(_05589_));
 sg13g2_antennanp ANTENNA_2475 (.A(_05589_));
 sg13g2_antennanp ANTENNA_2476 (.A(_05589_));
 sg13g2_antennanp ANTENNA_2477 (.A(_05631_));
 sg13g2_antennanp ANTENNA_2478 (.A(_05631_));
 sg13g2_antennanp ANTENNA_2479 (.A(_05631_));
 sg13g2_antennanp ANTENNA_2480 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2481 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2482 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2483 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2484 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2485 (.A(_05644_));
 sg13g2_antennanp ANTENNA_2486 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2487 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2488 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2489 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2490 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2491 (.A(_06275_));
 sg13g2_antennanp ANTENNA_2492 (.A(_07137_));
 sg13g2_antennanp ANTENNA_2493 (.A(_07138_));
 sg13g2_antennanp ANTENNA_2494 (.A(_07163_));
 sg13g2_antennanp ANTENNA_2495 (.A(_07163_));
 sg13g2_antennanp ANTENNA_2496 (.A(_07166_));
 sg13g2_antennanp ANTENNA_2497 (.A(_07166_));
 sg13g2_antennanp ANTENNA_2498 (.A(_07222_));
 sg13g2_antennanp ANTENNA_2499 (.A(_07326_));
 sg13g2_antennanp ANTENNA_2500 (.A(_07326_));
 sg13g2_antennanp ANTENNA_2501 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2502 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2503 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2504 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2505 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2506 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2507 (.A(_08081_));
 sg13g2_antennanp ANTENNA_2508 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2509 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2510 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2511 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2512 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2513 (.A(_08087_));
 sg13g2_antennanp ANTENNA_2514 (.A(_08092_));
 sg13g2_antennanp ANTENNA_2515 (.A(_08092_));
 sg13g2_antennanp ANTENNA_2516 (.A(_08092_));
 sg13g2_antennanp ANTENNA_2517 (.A(_08092_));
 sg13g2_antennanp ANTENNA_2518 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2519 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2520 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2521 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2522 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2523 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2524 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2525 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2526 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2527 (.A(_08184_));
 sg13g2_antennanp ANTENNA_2528 (.A(_08257_));
 sg13g2_antennanp ANTENNA_2529 (.A(_08257_));
 sg13g2_antennanp ANTENNA_2530 (.A(_08257_));
 sg13g2_antennanp ANTENNA_2531 (.A(_08257_));
 sg13g2_antennanp ANTENNA_2532 (.A(_08345_));
 sg13g2_antennanp ANTENNA_2533 (.A(_08345_));
 sg13g2_antennanp ANTENNA_2534 (.A(_08345_));
 sg13g2_antennanp ANTENNA_2535 (.A(_08345_));
 sg13g2_antennanp ANTENNA_2536 (.A(_08345_));
 sg13g2_antennanp ANTENNA_2537 (.A(_08403_));
 sg13g2_antennanp ANTENNA_2538 (.A(_08403_));
 sg13g2_antennanp ANTENNA_2539 (.A(_08403_));
 sg13g2_antennanp ANTENNA_2540 (.A(_08403_));
 sg13g2_antennanp ANTENNA_2541 (.A(_08517_));
 sg13g2_antennanp ANTENNA_2542 (.A(_08556_));
 sg13g2_antennanp ANTENNA_2543 (.A(_08614_));
 sg13g2_antennanp ANTENNA_2544 (.A(_08620_));
 sg13g2_antennanp ANTENNA_2545 (.A(_08620_));
 sg13g2_antennanp ANTENNA_2546 (.A(_08620_));
 sg13g2_antennanp ANTENNA_2547 (.A(_08620_));
 sg13g2_antennanp ANTENNA_2548 (.A(_08947_));
 sg13g2_antennanp ANTENNA_2549 (.A(_08947_));
 sg13g2_antennanp ANTENNA_2550 (.A(_08947_));
 sg13g2_antennanp ANTENNA_2551 (.A(_08947_));
 sg13g2_antennanp ANTENNA_2552 (.A(_08951_));
 sg13g2_antennanp ANTENNA_2553 (.A(_08951_));
 sg13g2_antennanp ANTENNA_2554 (.A(_08951_));
 sg13g2_antennanp ANTENNA_2555 (.A(_08951_));
 sg13g2_antennanp ANTENNA_2556 (.A(_08993_));
 sg13g2_antennanp ANTENNA_2557 (.A(_09005_));
 sg13g2_antennanp ANTENNA_2558 (.A(_09030_));
 sg13g2_antennanp ANTENNA_2559 (.A(_09030_));
 sg13g2_antennanp ANTENNA_2560 (.A(_09030_));
 sg13g2_antennanp ANTENNA_2561 (.A(_09037_));
 sg13g2_antennanp ANTENNA_2562 (.A(_09037_));
 sg13g2_antennanp ANTENNA_2563 (.A(_09037_));
 sg13g2_antennanp ANTENNA_2564 (.A(_09037_));
 sg13g2_antennanp ANTENNA_2565 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2566 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2567 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2568 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2569 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2570 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2571 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2572 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2573 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2574 (.A(_09039_));
 sg13g2_antennanp ANTENNA_2575 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2576 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2577 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2578 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2579 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2580 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2581 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2582 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2583 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2584 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2585 (.A(_09234_));
 sg13g2_antennanp ANTENNA_2586 (.A(_09253_));
 sg13g2_antennanp ANTENNA_2587 (.A(_09284_));
 sg13g2_antennanp ANTENNA_2588 (.A(_09305_));
 sg13g2_antennanp ANTENNA_2589 (.A(_09328_));
 sg13g2_antennanp ANTENNA_2590 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2591 (.A(_09370_));
 sg13g2_antennanp ANTENNA_2592 (.A(_09394_));
 sg13g2_antennanp ANTENNA_2593 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2594 (.A(_09470_));
 sg13g2_antennanp ANTENNA_2595 (.A(_09470_));
 sg13g2_antennanp ANTENNA_2596 (.A(_09470_));
 sg13g2_antennanp ANTENNA_2597 (.A(_09470_));
 sg13g2_antennanp ANTENNA_2598 (.A(_09470_));
 sg13g2_antennanp ANTENNA_2599 (.A(_09526_));
 sg13g2_antennanp ANTENNA_2600 (.A(_09553_));
 sg13g2_antennanp ANTENNA_2601 (.A(_09591_));
 sg13g2_antennanp ANTENNA_2602 (.A(_09591_));
 sg13g2_antennanp ANTENNA_2603 (.A(_09591_));
 sg13g2_antennanp ANTENNA_2604 (.A(_09591_));
 sg13g2_antennanp ANTENNA_2605 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2606 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2607 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2608 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2609 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2610 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2611 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2612 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2613 (.A(_09880_));
 sg13g2_antennanp ANTENNA_2614 (.A(_09882_));
 sg13g2_antennanp ANTENNA_2615 (.A(_09882_));
 sg13g2_antennanp ANTENNA_2616 (.A(_09882_));
 sg13g2_antennanp ANTENNA_2617 (.A(_09882_));
 sg13g2_antennanp ANTENNA_2618 (.A(_10156_));
 sg13g2_antennanp ANTENNA_2619 (.A(_10156_));
 sg13g2_antennanp ANTENNA_2620 (.A(_10156_));
 sg13g2_antennanp ANTENNA_2621 (.A(_10156_));
 sg13g2_antennanp ANTENNA_2622 (.A(_10241_));
 sg13g2_antennanp ANTENNA_2623 (.A(_10241_));
 sg13g2_antennanp ANTENNA_2624 (.A(_10241_));
 sg13g2_antennanp ANTENNA_2625 (.A(_10653_));
 sg13g2_antennanp ANTENNA_2626 (.A(_10653_));
 sg13g2_antennanp ANTENNA_2627 (.A(_10653_));
 sg13g2_antennanp ANTENNA_2628 (.A(_10653_));
 sg13g2_antennanp ANTENNA_2629 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2630 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2631 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2632 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2633 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2634 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2635 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2636 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2637 (.A(_10892_));
 sg13g2_antennanp ANTENNA_2638 (.A(_11550_));
 sg13g2_antennanp ANTENNA_2639 (.A(_11550_));
 sg13g2_antennanp ANTENNA_2640 (.A(_11550_));
 sg13g2_antennanp ANTENNA_2641 (.A(_11550_));
 sg13g2_antennanp ANTENNA_2642 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2643 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2644 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2645 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2646 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2647 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2648 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2649 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2650 (.A(_11613_));
 sg13g2_antennanp ANTENNA_2651 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2652 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2653 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2654 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2655 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2656 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2657 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2658 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2659 (.A(_11688_));
 sg13g2_antennanp ANTENNA_2660 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2661 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2662 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2663 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2664 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2665 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2666 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2667 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2668 (.A(_11695_));
 sg13g2_antennanp ANTENNA_2669 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2670 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2671 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2672 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2673 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2674 (.A(_11712_));
 sg13g2_antennanp ANTENNA_2675 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2676 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2677 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2678 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2679 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2680 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2681 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2682 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2683 (.A(_11743_));
 sg13g2_antennanp ANTENNA_2684 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2685 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2686 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2687 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2688 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2689 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2690 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2691 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2692 (.A(_11833_));
 sg13g2_antennanp ANTENNA_2693 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2694 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2695 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2696 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2697 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2698 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2699 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2700 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2701 (.A(_11866_));
 sg13g2_antennanp ANTENNA_2702 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2703 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2704 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2705 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2706 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2707 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2708 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2709 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2710 (.A(_11870_));
 sg13g2_antennanp ANTENNA_2711 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2712 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2713 (.A(_12009_));
 sg13g2_antennanp ANTENNA_2714 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2715 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2716 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2717 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2718 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2719 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2720 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2721 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2722 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2723 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2724 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2725 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2726 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2727 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2728 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2729 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2730 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2731 (.A(_12469_));
 sg13g2_antennanp ANTENNA_2732 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2733 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2734 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2735 (.A(_12473_));
 sg13g2_antennanp ANTENNA_2736 (.A(\cpu.addr[14] ));
 sg13g2_antennanp ANTENNA_2737 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2738 (.A(net3));
 sg13g2_antennanp ANTENNA_2739 (.A(net3));
 sg13g2_antennanp ANTENNA_2740 (.A(net3));
 sg13g2_antennanp ANTENNA_2741 (.A(net11));
 sg13g2_antennanp ANTENNA_2742 (.A(net11));
 sg13g2_antennanp ANTENNA_2743 (.A(net11));
 sg13g2_antennanp ANTENNA_2744 (.A(net12));
 sg13g2_antennanp ANTENNA_2745 (.A(net12));
 sg13g2_antennanp ANTENNA_2746 (.A(net12));
 sg13g2_antennanp ANTENNA_2747 (.A(net14));
 sg13g2_antennanp ANTENNA_2748 (.A(net14));
 sg13g2_antennanp ANTENNA_2749 (.A(net14));
 sg13g2_antennanp ANTENNA_2750 (.A(net19));
 sg13g2_antennanp ANTENNA_2751 (.A(net19));
 sg13g2_antennanp ANTENNA_2752 (.A(net19));
 sg13g2_antennanp ANTENNA_2753 (.A(net20));
 sg13g2_antennanp ANTENNA_2754 (.A(net20));
 sg13g2_antennanp ANTENNA_2755 (.A(net20));
 sg13g2_antennanp ANTENNA_2756 (.A(net464));
 sg13g2_antennanp ANTENNA_2757 (.A(net464));
 sg13g2_antennanp ANTENNA_2758 (.A(net464));
 sg13g2_antennanp ANTENNA_2759 (.A(net464));
 sg13g2_antennanp ANTENNA_2760 (.A(net464));
 sg13g2_antennanp ANTENNA_2761 (.A(net464));
 sg13g2_antennanp ANTENNA_2762 (.A(net464));
 sg13g2_antennanp ANTENNA_2763 (.A(net464));
 sg13g2_antennanp ANTENNA_2764 (.A(net464));
 sg13g2_antennanp ANTENNA_2765 (.A(net464));
 sg13g2_antennanp ANTENNA_2766 (.A(net464));
 sg13g2_antennanp ANTENNA_2767 (.A(net464));
 sg13g2_antennanp ANTENNA_2768 (.A(net464));
 sg13g2_antennanp ANTENNA_2769 (.A(net464));
 sg13g2_antennanp ANTENNA_2770 (.A(net464));
 sg13g2_antennanp ANTENNA_2771 (.A(net464));
 sg13g2_antennanp ANTENNA_2772 (.A(net464));
 sg13g2_antennanp ANTENNA_2773 (.A(net464));
 sg13g2_antennanp ANTENNA_2774 (.A(net464));
 sg13g2_antennanp ANTENNA_2775 (.A(net464));
 sg13g2_antennanp ANTENNA_2776 (.A(net498));
 sg13g2_antennanp ANTENNA_2777 (.A(net498));
 sg13g2_antennanp ANTENNA_2778 (.A(net498));
 sg13g2_antennanp ANTENNA_2779 (.A(net498));
 sg13g2_antennanp ANTENNA_2780 (.A(net498));
 sg13g2_antennanp ANTENNA_2781 (.A(net498));
 sg13g2_antennanp ANTENNA_2782 (.A(net498));
 sg13g2_antennanp ANTENNA_2783 (.A(net498));
 sg13g2_antennanp ANTENNA_2784 (.A(net498));
 sg13g2_antennanp ANTENNA_2785 (.A(net573));
 sg13g2_antennanp ANTENNA_2786 (.A(net573));
 sg13g2_antennanp ANTENNA_2787 (.A(net573));
 sg13g2_antennanp ANTENNA_2788 (.A(net573));
 sg13g2_antennanp ANTENNA_2789 (.A(net573));
 sg13g2_antennanp ANTENNA_2790 (.A(net573));
 sg13g2_antennanp ANTENNA_2791 (.A(net573));
 sg13g2_antennanp ANTENNA_2792 (.A(net573));
 sg13g2_antennanp ANTENNA_2793 (.A(net573));
 sg13g2_antennanp ANTENNA_2794 (.A(net576));
 sg13g2_antennanp ANTENNA_2795 (.A(net576));
 sg13g2_antennanp ANTENNA_2796 (.A(net576));
 sg13g2_antennanp ANTENNA_2797 (.A(net576));
 sg13g2_antennanp ANTENNA_2798 (.A(net576));
 sg13g2_antennanp ANTENNA_2799 (.A(net576));
 sg13g2_antennanp ANTENNA_2800 (.A(net576));
 sg13g2_antennanp ANTENNA_2801 (.A(net576));
 sg13g2_antennanp ANTENNA_2802 (.A(net576));
 sg13g2_antennanp ANTENNA_2803 (.A(net576));
 sg13g2_antennanp ANTENNA_2804 (.A(net576));
 sg13g2_antennanp ANTENNA_2805 (.A(net576));
 sg13g2_antennanp ANTENNA_2806 (.A(net576));
 sg13g2_antennanp ANTENNA_2807 (.A(net576));
 sg13g2_antennanp ANTENNA_2808 (.A(net576));
 sg13g2_antennanp ANTENNA_2809 (.A(net576));
 sg13g2_antennanp ANTENNA_2810 (.A(net576));
 sg13g2_antennanp ANTENNA_2811 (.A(net576));
 sg13g2_antennanp ANTENNA_2812 (.A(net576));
 sg13g2_antennanp ANTENNA_2813 (.A(net576));
 sg13g2_antennanp ANTENNA_2814 (.A(net714));
 sg13g2_antennanp ANTENNA_2815 (.A(net714));
 sg13g2_antennanp ANTENNA_2816 (.A(net714));
 sg13g2_antennanp ANTENNA_2817 (.A(net714));
 sg13g2_antennanp ANTENNA_2818 (.A(net714));
 sg13g2_antennanp ANTENNA_2819 (.A(net714));
 sg13g2_antennanp ANTENNA_2820 (.A(net714));
 sg13g2_antennanp ANTENNA_2821 (.A(net714));
 sg13g2_antennanp ANTENNA_2822 (.A(net714));
 sg13g2_antennanp ANTENNA_2823 (.A(net747));
 sg13g2_antennanp ANTENNA_2824 (.A(net747));
 sg13g2_antennanp ANTENNA_2825 (.A(net747));
 sg13g2_antennanp ANTENNA_2826 (.A(net747));
 sg13g2_antennanp ANTENNA_2827 (.A(net747));
 sg13g2_antennanp ANTENNA_2828 (.A(net747));
 sg13g2_antennanp ANTENNA_2829 (.A(net747));
 sg13g2_antennanp ANTENNA_2830 (.A(net747));
 sg13g2_antennanp ANTENNA_2831 (.A(net831));
 sg13g2_antennanp ANTENNA_2832 (.A(net831));
 sg13g2_antennanp ANTENNA_2833 (.A(net831));
 sg13g2_antennanp ANTENNA_2834 (.A(net831));
 sg13g2_antennanp ANTENNA_2835 (.A(net831));
 sg13g2_antennanp ANTENNA_2836 (.A(net831));
 sg13g2_antennanp ANTENNA_2837 (.A(net831));
 sg13g2_antennanp ANTENNA_2838 (.A(net831));
 sg13g2_antennanp ANTENNA_2839 (.A(net831));
 sg13g2_antennanp ANTENNA_2840 (.A(net834));
 sg13g2_antennanp ANTENNA_2841 (.A(net834));
 sg13g2_antennanp ANTENNA_2842 (.A(net834));
 sg13g2_antennanp ANTENNA_2843 (.A(net834));
 sg13g2_antennanp ANTENNA_2844 (.A(net834));
 sg13g2_antennanp ANTENNA_2845 (.A(net834));
 sg13g2_antennanp ANTENNA_2846 (.A(net834));
 sg13g2_antennanp ANTENNA_2847 (.A(net834));
 sg13g2_antennanp ANTENNA_2848 (.A(net834));
 sg13g2_antennanp ANTENNA_2849 (.A(net836));
 sg13g2_antennanp ANTENNA_2850 (.A(net836));
 sg13g2_antennanp ANTENNA_2851 (.A(net836));
 sg13g2_antennanp ANTENNA_2852 (.A(net836));
 sg13g2_antennanp ANTENNA_2853 (.A(net836));
 sg13g2_antennanp ANTENNA_2854 (.A(net836));
 sg13g2_antennanp ANTENNA_2855 (.A(net836));
 sg13g2_antennanp ANTENNA_2856 (.A(net836));
 sg13g2_antennanp ANTENNA_2857 (.A(net836));
 sg13g2_antennanp ANTENNA_2858 (.A(net837));
 sg13g2_antennanp ANTENNA_2859 (.A(net837));
 sg13g2_antennanp ANTENNA_2860 (.A(net837));
 sg13g2_antennanp ANTENNA_2861 (.A(net837));
 sg13g2_antennanp ANTENNA_2862 (.A(net837));
 sg13g2_antennanp ANTENNA_2863 (.A(net837));
 sg13g2_antennanp ANTENNA_2864 (.A(net837));
 sg13g2_antennanp ANTENNA_2865 (.A(net837));
 sg13g2_antennanp ANTENNA_2866 (.A(net837));
 sg13g2_antennanp ANTENNA_2867 (.A(net871));
 sg13g2_antennanp ANTENNA_2868 (.A(net871));
 sg13g2_antennanp ANTENNA_2869 (.A(net871));
 sg13g2_antennanp ANTENNA_2870 (.A(net871));
 sg13g2_antennanp ANTENNA_2871 (.A(net871));
 sg13g2_antennanp ANTENNA_2872 (.A(net871));
 sg13g2_antennanp ANTENNA_2873 (.A(net871));
 sg13g2_antennanp ANTENNA_2874 (.A(net871));
 sg13g2_antennanp ANTENNA_2875 (.A(net871));
 sg13g2_antennanp ANTENNA_2876 (.A(net905));
 sg13g2_antennanp ANTENNA_2877 (.A(net905));
 sg13g2_antennanp ANTENNA_2878 (.A(net905));
 sg13g2_antennanp ANTENNA_2879 (.A(net905));
 sg13g2_antennanp ANTENNA_2880 (.A(net905));
 sg13g2_antennanp ANTENNA_2881 (.A(net905));
 sg13g2_antennanp ANTENNA_2882 (.A(net905));
 sg13g2_antennanp ANTENNA_2883 (.A(net905));
 sg13g2_antennanp ANTENNA_2884 (.A(net905));
 sg13g2_antennanp ANTENNA_2885 (.A(net953));
 sg13g2_antennanp ANTENNA_2886 (.A(net953));
 sg13g2_antennanp ANTENNA_2887 (.A(net953));
 sg13g2_antennanp ANTENNA_2888 (.A(net953));
 sg13g2_antennanp ANTENNA_2889 (.A(net953));
 sg13g2_antennanp ANTENNA_2890 (.A(net953));
 sg13g2_antennanp ANTENNA_2891 (.A(net953));
 sg13g2_antennanp ANTENNA_2892 (.A(net953));
 sg13g2_antennanp ANTENNA_2893 (.A(net953));
 sg13g2_antennanp ANTENNA_2894 (.A(net958));
 sg13g2_antennanp ANTENNA_2895 (.A(net958));
 sg13g2_antennanp ANTENNA_2896 (.A(net958));
 sg13g2_antennanp ANTENNA_2897 (.A(net958));
 sg13g2_antennanp ANTENNA_2898 (.A(net958));
 sg13g2_antennanp ANTENNA_2899 (.A(net958));
 sg13g2_antennanp ANTENNA_2900 (.A(net958));
 sg13g2_antennanp ANTENNA_2901 (.A(net958));
 sg13g2_antennanp ANTENNA_2902 (.A(net967));
 sg13g2_antennanp ANTENNA_2903 (.A(net967));
 sg13g2_antennanp ANTENNA_2904 (.A(net967));
 sg13g2_antennanp ANTENNA_2905 (.A(net967));
 sg13g2_antennanp ANTENNA_2906 (.A(net967));
 sg13g2_antennanp ANTENNA_2907 (.A(net967));
 sg13g2_antennanp ANTENNA_2908 (.A(net967));
 sg13g2_antennanp ANTENNA_2909 (.A(net967));
 sg13g2_antennanp ANTENNA_2910 (.A(net967));
 sg13g2_antennanp ANTENNA_2911 (.A(net981));
 sg13g2_antennanp ANTENNA_2912 (.A(net981));
 sg13g2_antennanp ANTENNA_2913 (.A(net981));
 sg13g2_antennanp ANTENNA_2914 (.A(net981));
 sg13g2_antennanp ANTENNA_2915 (.A(net981));
 sg13g2_antennanp ANTENNA_2916 (.A(net981));
 sg13g2_antennanp ANTENNA_2917 (.A(net981));
 sg13g2_antennanp ANTENNA_2918 (.A(net981));
 sg13g2_antennanp ANTENNA_2919 (.A(net981));
 sg13g2_antennanp ANTENNA_2920 (.A(net994));
 sg13g2_antennanp ANTENNA_2921 (.A(net994));
 sg13g2_antennanp ANTENNA_2922 (.A(net994));
 sg13g2_antennanp ANTENNA_2923 (.A(net994));
 sg13g2_antennanp ANTENNA_2924 (.A(net994));
 sg13g2_antennanp ANTENNA_2925 (.A(net994));
 sg13g2_antennanp ANTENNA_2926 (.A(net994));
 sg13g2_antennanp ANTENNA_2927 (.A(net994));
 sg13g2_antennanp ANTENNA_2928 (.A(net994));
 sg13g2_antennanp ANTENNA_2929 (.A(net1022));
 sg13g2_antennanp ANTENNA_2930 (.A(net1022));
 sg13g2_antennanp ANTENNA_2931 (.A(net1022));
 sg13g2_antennanp ANTENNA_2932 (.A(net1022));
 sg13g2_antennanp ANTENNA_2933 (.A(net1022));
 sg13g2_antennanp ANTENNA_2934 (.A(net1022));
 sg13g2_antennanp ANTENNA_2935 (.A(net1022));
 sg13g2_antennanp ANTENNA_2936 (.A(net1022));
 sg13g2_antennanp ANTENNA_2937 (.A(net1022));
 sg13g2_antennanp ANTENNA_2938 (.A(net1022));
 sg13g2_antennanp ANTENNA_2939 (.A(net1022));
 sg13g2_antennanp ANTENNA_2940 (.A(net1022));
 sg13g2_antennanp ANTENNA_2941 (.A(net1022));
 sg13g2_antennanp ANTENNA_2942 (.A(net1022));
 sg13g2_antennanp ANTENNA_2943 (.A(net1022));
 sg13g2_antennanp ANTENNA_2944 (.A(net1022));
 sg13g2_antennanp ANTENNA_2945 (.A(net1022));
 sg13g2_antennanp ANTENNA_2946 (.A(net1022));
 sg13g2_antennanp ANTENNA_2947 (.A(net1022));
 sg13g2_antennanp ANTENNA_2948 (.A(net1022));
 sg13g2_antennanp ANTENNA_2949 (.A(net1075));
 sg13g2_antennanp ANTENNA_2950 (.A(net1075));
 sg13g2_antennanp ANTENNA_2951 (.A(net1075));
 sg13g2_antennanp ANTENNA_2952 (.A(net1075));
 sg13g2_antennanp ANTENNA_2953 (.A(net1075));
 sg13g2_antennanp ANTENNA_2954 (.A(net1075));
 sg13g2_antennanp ANTENNA_2955 (.A(net1075));
 sg13g2_antennanp ANTENNA_2956 (.A(net1075));
 sg13g2_antennanp ANTENNA_2957 (.A(net1075));
 sg13g2_antennanp ANTENNA_2958 (.A(net1085));
 sg13g2_antennanp ANTENNA_2959 (.A(net1085));
 sg13g2_antennanp ANTENNA_2960 (.A(net1085));
 sg13g2_antennanp ANTENNA_2961 (.A(net1085));
 sg13g2_antennanp ANTENNA_2962 (.A(net1085));
 sg13g2_antennanp ANTENNA_2963 (.A(net1085));
 sg13g2_antennanp ANTENNA_2964 (.A(net1085));
 sg13g2_antennanp ANTENNA_2965 (.A(net1085));
 sg13g2_antennanp ANTENNA_2966 (.A(net1085));
 sg13g2_antennanp ANTENNA_2967 (.A(net1085));
 sg13g2_antennanp ANTENNA_2968 (.A(net1085));
 sg13g2_antennanp ANTENNA_2969 (.A(net1085));
 sg13g2_antennanp ANTENNA_2970 (.A(net1085));
 sg13g2_antennanp ANTENNA_2971 (.A(net1085));
 sg13g2_antennanp ANTENNA_2972 (.A(net1085));
 sg13g2_antennanp ANTENNA_2973 (.A(net1085));
 sg13g2_antennanp ANTENNA_2974 (.A(net1085));
 sg13g2_antennanp ANTENNA_2975 (.A(net1085));
 sg13g2_antennanp ANTENNA_2976 (.A(net1085));
 sg13g2_antennanp ANTENNA_2977 (.A(net1085));
 sg13g2_antennanp ANTENNA_2978 (.A(net1085));
 sg13g2_antennanp ANTENNA_2979 (.A(net1085));
 sg13g2_antennanp ANTENNA_2980 (.A(net1085));
 sg13g2_antennanp ANTENNA_2981 (.A(net1085));
 sg13g2_antennanp ANTENNA_2982 (.A(net1085));
 sg13g2_antennanp ANTENNA_2983 (.A(net1085));
 sg13g2_antennanp ANTENNA_2984 (.A(net1085));
 sg13g2_antennanp ANTENNA_2985 (.A(net1085));
 sg13g2_antennanp ANTENNA_2986 (.A(net1085));
 sg13g2_antennanp ANTENNA_2987 (.A(net1096));
 sg13g2_antennanp ANTENNA_2988 (.A(net1096));
 sg13g2_antennanp ANTENNA_2989 (.A(net1096));
 sg13g2_antennanp ANTENNA_2990 (.A(net1096));
 sg13g2_antennanp ANTENNA_2991 (.A(net1096));
 sg13g2_antennanp ANTENNA_2992 (.A(net1096));
 sg13g2_antennanp ANTENNA_2993 (.A(net1096));
 sg13g2_antennanp ANTENNA_2994 (.A(net1096));
 sg13g2_antennanp ANTENNA_2995 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2996 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2997 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2998 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2999 (.A(_01057_));
 sg13g2_antennanp ANTENNA_3000 (.A(_01057_));
 sg13g2_antennanp ANTENNA_3001 (.A(_01071_));
 sg13g2_antennanp ANTENNA_3002 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3003 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3004 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3005 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3006 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3007 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3008 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3009 (.A(_02855_));
 sg13g2_antennanp ANTENNA_3010 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3011 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3012 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3013 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3014 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3015 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3016 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3017 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3018 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3019 (.A(_02856_));
 sg13g2_antennanp ANTENNA_3020 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3021 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3022 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3023 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3024 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3025 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3026 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3027 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3028 (.A(_02866_));
 sg13g2_antennanp ANTENNA_3029 (.A(_02873_));
 sg13g2_antennanp ANTENNA_3030 (.A(_02873_));
 sg13g2_antennanp ANTENNA_3031 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3032 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3033 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3034 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3035 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3036 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3037 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3038 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3039 (.A(_02877_));
 sg13g2_antennanp ANTENNA_3040 (.A(_03350_));
 sg13g2_antennanp ANTENNA_3041 (.A(_03350_));
 sg13g2_antennanp ANTENNA_3042 (.A(_03350_));
 sg13g2_antennanp ANTENNA_3043 (.A(_03350_));
 sg13g2_antennanp ANTENNA_3044 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3045 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3046 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3047 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3048 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3049 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3050 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3051 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3052 (.A(_03356_));
 sg13g2_antennanp ANTENNA_3053 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3054 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3055 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3056 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3057 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3058 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3059 (.A(_03612_));
 sg13g2_antennanp ANTENNA_3060 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3061 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3062 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3063 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3064 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3065 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3066 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3067 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3068 (.A(_04628_));
 sg13g2_antennanp ANTENNA_3069 (.A(_04646_));
 sg13g2_antennanp ANTENNA_3070 (.A(_04980_));
 sg13g2_antennanp ANTENNA_3071 (.A(_05022_));
 sg13g2_antennanp ANTENNA_3072 (.A(_05046_));
 sg13g2_antennanp ANTENNA_3073 (.A(_05581_));
 sg13g2_antennanp ANTENNA_3074 (.A(_05584_));
 sg13g2_antennanp ANTENNA_3075 (.A(_05589_));
 sg13g2_antennanp ANTENNA_3076 (.A(_05589_));
 sg13g2_antennanp ANTENNA_3077 (.A(_05589_));
 sg13g2_antennanp ANTENNA_3078 (.A(_05631_));
 sg13g2_antennanp ANTENNA_3079 (.A(_05631_));
 sg13g2_antennanp ANTENNA_3080 (.A(_05631_));
 sg13g2_antennanp ANTENNA_3081 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3082 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3083 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3084 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3085 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3086 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3087 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3088 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3089 (.A(_05644_));
 sg13g2_antennanp ANTENNA_3090 (.A(_07138_));
 sg13g2_antennanp ANTENNA_3091 (.A(_07163_));
 sg13g2_antennanp ANTENNA_3092 (.A(_07163_));
 sg13g2_antennanp ANTENNA_3093 (.A(_07166_));
 sg13g2_antennanp ANTENNA_3094 (.A(_07222_));
 sg13g2_antennanp ANTENNA_3095 (.A(_07326_));
 sg13g2_antennanp ANTENNA_3096 (.A(_07326_));
 sg13g2_antennanp ANTENNA_3097 (.A(_08092_));
 sg13g2_antennanp ANTENNA_3098 (.A(_08092_));
 sg13g2_antennanp ANTENNA_3099 (.A(_08092_));
 sg13g2_antennanp ANTENNA_3100 (.A(_08092_));
 sg13g2_antennanp ANTENNA_3101 (.A(_08403_));
 sg13g2_antennanp ANTENNA_3102 (.A(_08403_));
 sg13g2_antennanp ANTENNA_3103 (.A(_08403_));
 sg13g2_antennanp ANTENNA_3104 (.A(_08403_));
 sg13g2_antennanp ANTENNA_3105 (.A(_08517_));
 sg13g2_antennanp ANTENNA_3106 (.A(_08556_));
 sg13g2_antennanp ANTENNA_3107 (.A(_08556_));
 sg13g2_antennanp ANTENNA_3108 (.A(_08614_));
 sg13g2_antennanp ANTENNA_3109 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3110 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3111 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3112 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3113 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3114 (.A(_08947_));
 sg13g2_antennanp ANTENNA_3115 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3116 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3117 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3118 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3119 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3120 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3121 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3122 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3123 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3124 (.A(_08951_));
 sg13g2_antennanp ANTENNA_3125 (.A(_08993_));
 sg13g2_antennanp ANTENNA_3126 (.A(_08993_));
 sg13g2_antennanp ANTENNA_3127 (.A(_09005_));
 sg13g2_antennanp ANTENNA_3128 (.A(_09005_));
 sg13g2_antennanp ANTENNA_3129 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3130 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3131 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3132 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3133 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3134 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3135 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3136 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3137 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3138 (.A(_09037_));
 sg13g2_antennanp ANTENNA_3139 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3140 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3141 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3142 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3143 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3144 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3145 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3146 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3147 (.A(_09039_));
 sg13g2_antennanp ANTENNA_3148 (.A(_09095_));
 sg13g2_antennanp ANTENNA_3149 (.A(_09095_));
 sg13g2_antennanp ANTENNA_3150 (.A(_09095_));
 sg13g2_antennanp ANTENNA_3151 (.A(_09095_));
 sg13g2_antennanp ANTENNA_3152 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3153 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3154 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3155 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3156 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3157 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3158 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3159 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3160 (.A(_09151_));
 sg13g2_antennanp ANTENNA_3161 (.A(_09205_));
 sg13g2_antennanp ANTENNA_3162 (.A(_09234_));
 sg13g2_antennanp ANTENNA_3163 (.A(_09253_));
 sg13g2_antennanp ANTENNA_3164 (.A(_09305_));
 sg13g2_antennanp ANTENNA_3165 (.A(_09328_));
 sg13g2_antennanp ANTENNA_3166 (.A(_09349_));
 sg13g2_antennanp ANTENNA_3167 (.A(_09370_));
 sg13g2_antennanp ANTENNA_3168 (.A(_09394_));
 sg13g2_antennanp ANTENNA_3169 (.A(_09426_));
 sg13g2_antennanp ANTENNA_3170 (.A(_09526_));
 sg13g2_antennanp ANTENNA_3171 (.A(_09553_));
 sg13g2_antennanp ANTENNA_3172 (.A(_09591_));
 sg13g2_antennanp ANTENNA_3173 (.A(_09591_));
 sg13g2_antennanp ANTENNA_3174 (.A(_09591_));
 sg13g2_antennanp ANTENNA_3175 (.A(_09591_));
 sg13g2_antennanp ANTENNA_3176 (.A(_09869_));
 sg13g2_antennanp ANTENNA_3177 (.A(_09869_));
 sg13g2_antennanp ANTENNA_3178 (.A(_09869_));
 sg13g2_antennanp ANTENNA_3179 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3180 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3181 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3182 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3183 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3184 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3185 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3186 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3187 (.A(_09880_));
 sg13g2_antennanp ANTENNA_3188 (.A(_09882_));
 sg13g2_antennanp ANTENNA_3189 (.A(_09882_));
 sg13g2_antennanp ANTENNA_3190 (.A(_09882_));
 sg13g2_antennanp ANTENNA_3191 (.A(_09882_));
 sg13g2_antennanp ANTENNA_3192 (.A(_10156_));
 sg13g2_antennanp ANTENNA_3193 (.A(_10156_));
 sg13g2_antennanp ANTENNA_3194 (.A(_10156_));
 sg13g2_antennanp ANTENNA_3195 (.A(_10156_));
 sg13g2_antennanp ANTENNA_3196 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3197 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3198 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3199 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3200 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3201 (.A(_10241_));
 sg13g2_antennanp ANTENNA_3202 (.A(_10653_));
 sg13g2_antennanp ANTENNA_3203 (.A(_10653_));
 sg13g2_antennanp ANTENNA_3204 (.A(_10653_));
 sg13g2_antennanp ANTENNA_3205 (.A(_10653_));
 sg13g2_antennanp ANTENNA_3206 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3207 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3208 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3209 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3210 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3211 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3212 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3213 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3214 (.A(_10892_));
 sg13g2_antennanp ANTENNA_3215 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3216 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3217 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3218 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3219 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3220 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3221 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3222 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3223 (.A(_11613_));
 sg13g2_antennanp ANTENNA_3224 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3225 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3226 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3227 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3228 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3229 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3230 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3231 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3232 (.A(_11688_));
 sg13g2_antennanp ANTENNA_3233 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3234 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3235 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3236 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3237 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3238 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3239 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3240 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3241 (.A(_11695_));
 sg13g2_antennanp ANTENNA_3242 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3243 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3244 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3245 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3246 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3247 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3248 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3249 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3250 (.A(_11712_));
 sg13g2_antennanp ANTENNA_3251 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3252 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3253 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3254 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3255 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3256 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3257 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3258 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3259 (.A(_11743_));
 sg13g2_antennanp ANTENNA_3260 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3261 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3262 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3263 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3264 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3265 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3266 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3267 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3268 (.A(_11833_));
 sg13g2_antennanp ANTENNA_3269 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3270 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3271 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3272 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3273 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3274 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3275 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3276 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3277 (.A(_11866_));
 sg13g2_antennanp ANTENNA_3278 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3279 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3280 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3281 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3282 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3283 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3284 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3285 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3286 (.A(_11870_));
 sg13g2_antennanp ANTENNA_3287 (.A(_12009_));
 sg13g2_antennanp ANTENNA_3288 (.A(_12009_));
 sg13g2_antennanp ANTENNA_3289 (.A(_12009_));
 sg13g2_antennanp ANTENNA_3290 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3291 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3292 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3293 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3294 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3295 (.A(_12185_));
 sg13g2_antennanp ANTENNA_3296 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3297 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3298 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3299 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3300 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3301 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3302 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3303 (.A(_12469_));
 sg13g2_antennanp ANTENNA_3304 (.A(_12473_));
 sg13g2_antennanp ANTENNA_3305 (.A(_12473_));
 sg13g2_antennanp ANTENNA_3306 (.A(_12473_));
 sg13g2_antennanp ANTENNA_3307 (.A(_12473_));
 sg13g2_antennanp ANTENNA_3308 (.A(\cpu.addr[14] ));
 sg13g2_antennanp ANTENNA_3309 (.A(net3));
 sg13g2_antennanp ANTENNA_3310 (.A(net3));
 sg13g2_antennanp ANTENNA_3311 (.A(net3));
 sg13g2_antennanp ANTENNA_3312 (.A(net11));
 sg13g2_antennanp ANTENNA_3313 (.A(net11));
 sg13g2_antennanp ANTENNA_3314 (.A(net11));
 sg13g2_antennanp ANTENNA_3315 (.A(net12));
 sg13g2_antennanp ANTENNA_3316 (.A(net12));
 sg13g2_antennanp ANTENNA_3317 (.A(net12));
 sg13g2_antennanp ANTENNA_3318 (.A(net14));
 sg13g2_antennanp ANTENNA_3319 (.A(net14));
 sg13g2_antennanp ANTENNA_3320 (.A(net14));
 sg13g2_antennanp ANTENNA_3321 (.A(net19));
 sg13g2_antennanp ANTENNA_3322 (.A(net19));
 sg13g2_antennanp ANTENNA_3323 (.A(net19));
 sg13g2_antennanp ANTENNA_3324 (.A(net20));
 sg13g2_antennanp ANTENNA_3325 (.A(net20));
 sg13g2_antennanp ANTENNA_3326 (.A(net20));
 sg13g2_antennanp ANTENNA_3327 (.A(net464));
 sg13g2_antennanp ANTENNA_3328 (.A(net464));
 sg13g2_antennanp ANTENNA_3329 (.A(net464));
 sg13g2_antennanp ANTENNA_3330 (.A(net464));
 sg13g2_antennanp ANTENNA_3331 (.A(net464));
 sg13g2_antennanp ANTENNA_3332 (.A(net464));
 sg13g2_antennanp ANTENNA_3333 (.A(net464));
 sg13g2_antennanp ANTENNA_3334 (.A(net464));
 sg13g2_antennanp ANTENNA_3335 (.A(net464));
 sg13g2_antennanp ANTENNA_3336 (.A(net464));
 sg13g2_antennanp ANTENNA_3337 (.A(net464));
 sg13g2_antennanp ANTENNA_3338 (.A(net464));
 sg13g2_antennanp ANTENNA_3339 (.A(net464));
 sg13g2_antennanp ANTENNA_3340 (.A(net464));
 sg13g2_antennanp ANTENNA_3341 (.A(net464));
 sg13g2_antennanp ANTENNA_3342 (.A(net464));
 sg13g2_antennanp ANTENNA_3343 (.A(net464));
 sg13g2_antennanp ANTENNA_3344 (.A(net464));
 sg13g2_antennanp ANTENNA_3345 (.A(net464));
 sg13g2_antennanp ANTENNA_3346 (.A(net464));
 sg13g2_antennanp ANTENNA_3347 (.A(net498));
 sg13g2_antennanp ANTENNA_3348 (.A(net498));
 sg13g2_antennanp ANTENNA_3349 (.A(net498));
 sg13g2_antennanp ANTENNA_3350 (.A(net498));
 sg13g2_antennanp ANTENNA_3351 (.A(net498));
 sg13g2_antennanp ANTENNA_3352 (.A(net498));
 sg13g2_antennanp ANTENNA_3353 (.A(net498));
 sg13g2_antennanp ANTENNA_3354 (.A(net498));
 sg13g2_antennanp ANTENNA_3355 (.A(net498));
 sg13g2_antennanp ANTENNA_3356 (.A(net573));
 sg13g2_antennanp ANTENNA_3357 (.A(net573));
 sg13g2_antennanp ANTENNA_3358 (.A(net573));
 sg13g2_antennanp ANTENNA_3359 (.A(net573));
 sg13g2_antennanp ANTENNA_3360 (.A(net573));
 sg13g2_antennanp ANTENNA_3361 (.A(net573));
 sg13g2_antennanp ANTENNA_3362 (.A(net573));
 sg13g2_antennanp ANTENNA_3363 (.A(net573));
 sg13g2_antennanp ANTENNA_3364 (.A(net573));
 sg13g2_antennanp ANTENNA_3365 (.A(net576));
 sg13g2_antennanp ANTENNA_3366 (.A(net576));
 sg13g2_antennanp ANTENNA_3367 (.A(net576));
 sg13g2_antennanp ANTENNA_3368 (.A(net576));
 sg13g2_antennanp ANTENNA_3369 (.A(net576));
 sg13g2_antennanp ANTENNA_3370 (.A(net576));
 sg13g2_antennanp ANTENNA_3371 (.A(net576));
 sg13g2_antennanp ANTENNA_3372 (.A(net576));
 sg13g2_antennanp ANTENNA_3373 (.A(net576));
 sg13g2_antennanp ANTENNA_3374 (.A(net576));
 sg13g2_antennanp ANTENNA_3375 (.A(net576));
 sg13g2_antennanp ANTENNA_3376 (.A(net576));
 sg13g2_antennanp ANTENNA_3377 (.A(net576));
 sg13g2_antennanp ANTENNA_3378 (.A(net576));
 sg13g2_antennanp ANTENNA_3379 (.A(net576));
 sg13g2_antennanp ANTENNA_3380 (.A(net576));
 sg13g2_antennanp ANTENNA_3381 (.A(net576));
 sg13g2_antennanp ANTENNA_3382 (.A(net576));
 sg13g2_antennanp ANTENNA_3383 (.A(net576));
 sg13g2_antennanp ANTENNA_3384 (.A(net576));
 sg13g2_antennanp ANTENNA_3385 (.A(net714));
 sg13g2_antennanp ANTENNA_3386 (.A(net714));
 sg13g2_antennanp ANTENNA_3387 (.A(net714));
 sg13g2_antennanp ANTENNA_3388 (.A(net714));
 sg13g2_antennanp ANTENNA_3389 (.A(net714));
 sg13g2_antennanp ANTENNA_3390 (.A(net714));
 sg13g2_antennanp ANTENNA_3391 (.A(net714));
 sg13g2_antennanp ANTENNA_3392 (.A(net714));
 sg13g2_antennanp ANTENNA_3393 (.A(net714));
 sg13g2_antennanp ANTENNA_3394 (.A(net747));
 sg13g2_antennanp ANTENNA_3395 (.A(net747));
 sg13g2_antennanp ANTENNA_3396 (.A(net747));
 sg13g2_antennanp ANTENNA_3397 (.A(net747));
 sg13g2_antennanp ANTENNA_3398 (.A(net747));
 sg13g2_antennanp ANTENNA_3399 (.A(net747));
 sg13g2_antennanp ANTENNA_3400 (.A(net747));
 sg13g2_antennanp ANTENNA_3401 (.A(net747));
 sg13g2_antennanp ANTENNA_3402 (.A(net831));
 sg13g2_antennanp ANTENNA_3403 (.A(net831));
 sg13g2_antennanp ANTENNA_3404 (.A(net831));
 sg13g2_antennanp ANTENNA_3405 (.A(net831));
 sg13g2_antennanp ANTENNA_3406 (.A(net831));
 sg13g2_antennanp ANTENNA_3407 (.A(net831));
 sg13g2_antennanp ANTENNA_3408 (.A(net831));
 sg13g2_antennanp ANTENNA_3409 (.A(net831));
 sg13g2_antennanp ANTENNA_3410 (.A(net831));
 sg13g2_antennanp ANTENNA_3411 (.A(net834));
 sg13g2_antennanp ANTENNA_3412 (.A(net834));
 sg13g2_antennanp ANTENNA_3413 (.A(net834));
 sg13g2_antennanp ANTENNA_3414 (.A(net834));
 sg13g2_antennanp ANTENNA_3415 (.A(net834));
 sg13g2_antennanp ANTENNA_3416 (.A(net834));
 sg13g2_antennanp ANTENNA_3417 (.A(net834));
 sg13g2_antennanp ANTENNA_3418 (.A(net834));
 sg13g2_antennanp ANTENNA_3419 (.A(net834));
 sg13g2_antennanp ANTENNA_3420 (.A(net836));
 sg13g2_antennanp ANTENNA_3421 (.A(net836));
 sg13g2_antennanp ANTENNA_3422 (.A(net836));
 sg13g2_antennanp ANTENNA_3423 (.A(net836));
 sg13g2_antennanp ANTENNA_3424 (.A(net836));
 sg13g2_antennanp ANTENNA_3425 (.A(net836));
 sg13g2_antennanp ANTENNA_3426 (.A(net836));
 sg13g2_antennanp ANTENNA_3427 (.A(net836));
 sg13g2_antennanp ANTENNA_3428 (.A(net836));
 sg13g2_antennanp ANTENNA_3429 (.A(net837));
 sg13g2_antennanp ANTENNA_3430 (.A(net837));
 sg13g2_antennanp ANTENNA_3431 (.A(net837));
 sg13g2_antennanp ANTENNA_3432 (.A(net837));
 sg13g2_antennanp ANTENNA_3433 (.A(net837));
 sg13g2_antennanp ANTENNA_3434 (.A(net837));
 sg13g2_antennanp ANTENNA_3435 (.A(net837));
 sg13g2_antennanp ANTENNA_3436 (.A(net837));
 sg13g2_antennanp ANTENNA_3437 (.A(net837));
 sg13g2_antennanp ANTENNA_3438 (.A(net953));
 sg13g2_antennanp ANTENNA_3439 (.A(net953));
 sg13g2_antennanp ANTENNA_3440 (.A(net953));
 sg13g2_antennanp ANTENNA_3441 (.A(net953));
 sg13g2_antennanp ANTENNA_3442 (.A(net953));
 sg13g2_antennanp ANTENNA_3443 (.A(net953));
 sg13g2_antennanp ANTENNA_3444 (.A(net953));
 sg13g2_antennanp ANTENNA_3445 (.A(net953));
 sg13g2_antennanp ANTENNA_3446 (.A(net953));
 sg13g2_antennanp ANTENNA_3447 (.A(net953));
 sg13g2_antennanp ANTENNA_3448 (.A(net953));
 sg13g2_antennanp ANTENNA_3449 (.A(net953));
 sg13g2_antennanp ANTENNA_3450 (.A(net953));
 sg13g2_antennanp ANTENNA_3451 (.A(net953));
 sg13g2_antennanp ANTENNA_3452 (.A(net958));
 sg13g2_antennanp ANTENNA_3453 (.A(net958));
 sg13g2_antennanp ANTENNA_3454 (.A(net958));
 sg13g2_antennanp ANTENNA_3455 (.A(net958));
 sg13g2_antennanp ANTENNA_3456 (.A(net958));
 sg13g2_antennanp ANTENNA_3457 (.A(net958));
 sg13g2_antennanp ANTENNA_3458 (.A(net958));
 sg13g2_antennanp ANTENNA_3459 (.A(net958));
 sg13g2_antennanp ANTENNA_3460 (.A(net958));
 sg13g2_antennanp ANTENNA_3461 (.A(net958));
 sg13g2_antennanp ANTENNA_3462 (.A(net967));
 sg13g2_antennanp ANTENNA_3463 (.A(net967));
 sg13g2_antennanp ANTENNA_3464 (.A(net967));
 sg13g2_antennanp ANTENNA_3465 (.A(net967));
 sg13g2_antennanp ANTENNA_3466 (.A(net967));
 sg13g2_antennanp ANTENNA_3467 (.A(net967));
 sg13g2_antennanp ANTENNA_3468 (.A(net967));
 sg13g2_antennanp ANTENNA_3469 (.A(net967));
 sg13g2_antennanp ANTENNA_3470 (.A(net967));
 sg13g2_antennanp ANTENNA_3471 (.A(net981));
 sg13g2_antennanp ANTENNA_3472 (.A(net981));
 sg13g2_antennanp ANTENNA_3473 (.A(net981));
 sg13g2_antennanp ANTENNA_3474 (.A(net981));
 sg13g2_antennanp ANTENNA_3475 (.A(net981));
 sg13g2_antennanp ANTENNA_3476 (.A(net981));
 sg13g2_antennanp ANTENNA_3477 (.A(net981));
 sg13g2_antennanp ANTENNA_3478 (.A(net981));
 sg13g2_antennanp ANTENNA_3479 (.A(net981));
 sg13g2_antennanp ANTENNA_3480 (.A(net994));
 sg13g2_antennanp ANTENNA_3481 (.A(net994));
 sg13g2_antennanp ANTENNA_3482 (.A(net994));
 sg13g2_antennanp ANTENNA_3483 (.A(net994));
 sg13g2_antennanp ANTENNA_3484 (.A(net994));
 sg13g2_antennanp ANTENNA_3485 (.A(net994));
 sg13g2_antennanp ANTENNA_3486 (.A(net994));
 sg13g2_antennanp ANTENNA_3487 (.A(net994));
 sg13g2_antennanp ANTENNA_3488 (.A(net994));
 sg13g2_antennanp ANTENNA_3489 (.A(net1022));
 sg13g2_antennanp ANTENNA_3490 (.A(net1022));
 sg13g2_antennanp ANTENNA_3491 (.A(net1022));
 sg13g2_antennanp ANTENNA_3492 (.A(net1022));
 sg13g2_antennanp ANTENNA_3493 (.A(net1022));
 sg13g2_antennanp ANTENNA_3494 (.A(net1022));
 sg13g2_antennanp ANTENNA_3495 (.A(net1022));
 sg13g2_antennanp ANTENNA_3496 (.A(net1022));
 sg13g2_antennanp ANTENNA_3497 (.A(net1022));
 sg13g2_antennanp ANTENNA_3498 (.A(net1022));
 sg13g2_antennanp ANTENNA_3499 (.A(net1022));
 sg13g2_antennanp ANTENNA_3500 (.A(net1022));
 sg13g2_antennanp ANTENNA_3501 (.A(net1022));
 sg13g2_antennanp ANTENNA_3502 (.A(net1022));
 sg13g2_antennanp ANTENNA_3503 (.A(net1022));
 sg13g2_antennanp ANTENNA_3504 (.A(net1022));
 sg13g2_antennanp ANTENNA_3505 (.A(net1022));
 sg13g2_antennanp ANTENNA_3506 (.A(net1022));
 sg13g2_antennanp ANTENNA_3507 (.A(net1022));
 sg13g2_antennanp ANTENNA_3508 (.A(net1022));
 sg13g2_antennanp ANTENNA_3509 (.A(net1075));
 sg13g2_antennanp ANTENNA_3510 (.A(net1075));
 sg13g2_antennanp ANTENNA_3511 (.A(net1075));
 sg13g2_antennanp ANTENNA_3512 (.A(net1075));
 sg13g2_antennanp ANTENNA_3513 (.A(net1075));
 sg13g2_antennanp ANTENNA_3514 (.A(net1075));
 sg13g2_antennanp ANTENNA_3515 (.A(net1075));
 sg13g2_antennanp ANTENNA_3516 (.A(net1075));
 sg13g2_antennanp ANTENNA_3517 (.A(net1075));
 sg13g2_antennanp ANTENNA_3518 (.A(net1085));
 sg13g2_antennanp ANTENNA_3519 (.A(net1085));
 sg13g2_antennanp ANTENNA_3520 (.A(net1085));
 sg13g2_antennanp ANTENNA_3521 (.A(net1085));
 sg13g2_antennanp ANTENNA_3522 (.A(net1085));
 sg13g2_antennanp ANTENNA_3523 (.A(net1085));
 sg13g2_antennanp ANTENNA_3524 (.A(net1085));
 sg13g2_antennanp ANTENNA_3525 (.A(net1085));
 sg13g2_antennanp ANTENNA_3526 (.A(net1085));
 sg13g2_antennanp ANTENNA_3527 (.A(net1085));
 sg13g2_antennanp ANTENNA_3528 (.A(net1085));
 sg13g2_antennanp ANTENNA_3529 (.A(net1085));
 sg13g2_antennanp ANTENNA_3530 (.A(net1085));
 sg13g2_antennanp ANTENNA_3531 (.A(net1085));
 sg13g2_antennanp ANTENNA_3532 (.A(net1085));
 sg13g2_antennanp ANTENNA_3533 (.A(net1085));
 sg13g2_antennanp ANTENNA_3534 (.A(net1085));
 sg13g2_antennanp ANTENNA_3535 (.A(net1085));
 sg13g2_antennanp ANTENNA_3536 (.A(net1085));
 sg13g2_antennanp ANTENNA_3537 (.A(net1085));
 sg13g2_antennanp ANTENNA_3538 (.A(net1085));
 sg13g2_antennanp ANTENNA_3539 (.A(net1085));
 sg13g2_antennanp ANTENNA_3540 (.A(net1085));
 sg13g2_antennanp ANTENNA_3541 (.A(net1085));
 sg13g2_antennanp ANTENNA_3542 (.A(net1085));
 sg13g2_antennanp ANTENNA_3543 (.A(net1085));
 sg13g2_antennanp ANTENNA_3544 (.A(net1085));
 sg13g2_antennanp ANTENNA_3545 (.A(net1085));
 sg13g2_antennanp ANTENNA_3546 (.A(net1085));
 sg13g2_antennanp ANTENNA_3547 (.A(net1096));
 sg13g2_antennanp ANTENNA_3548 (.A(net1096));
 sg13g2_antennanp ANTENNA_3549 (.A(net1096));
 sg13g2_antennanp ANTENNA_3550 (.A(net1096));
 sg13g2_antennanp ANTENNA_3551 (.A(net1096));
 sg13g2_antennanp ANTENNA_3552 (.A(net1096));
 sg13g2_antennanp ANTENNA_3553 (.A(net1096));
 sg13g2_antennanp ANTENNA_3554 (.A(net1096));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_fill_2 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_160 ();
 sg13g2_fill_2 FILLER_0_167 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_4 FILLER_0_289 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_fill_2 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_4 FILLER_0_381 ();
 sg13g2_fill_1 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_fill_1 FILLER_0_426 ();
 sg13g2_fill_2 FILLER_0_453 ();
 sg13g2_fill_1 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_460 ();
 sg13g2_fill_1 FILLER_0_467 ();
 sg13g2_decap_8 FILLER_0_472 ();
 sg13g2_decap_8 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_486 ();
 sg13g2_decap_8 FILLER_0_493 ();
 sg13g2_fill_2 FILLER_0_500 ();
 sg13g2_decap_8 FILLER_0_506 ();
 sg13g2_fill_2 FILLER_0_513 ();
 sg13g2_fill_1 FILLER_0_515 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_552 ();
 sg13g2_decap_4 FILLER_0_559 ();
 sg13g2_fill_2 FILLER_0_563 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_4 FILLER_0_576 ();
 sg13g2_fill_2 FILLER_0_580 ();
 sg13g2_fill_2 FILLER_0_586 ();
 sg13g2_decap_4 FILLER_0_601 ();
 sg13g2_fill_2 FILLER_0_605 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_fill_1 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_739 ();
 sg13g2_fill_1 FILLER_0_746 ();
 sg13g2_fill_1 FILLER_0_757 ();
 sg13g2_decap_4 FILLER_0_784 ();
 sg13g2_fill_2 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_fill_2 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_832 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_fill_1 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_4 FILLER_0_866 ();
 sg13g2_fill_2 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_fill_1 FILLER_0_883 ();
 sg13g2_decap_4 FILLER_0_888 ();
 sg13g2_fill_1 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_fill_1 FILLER_0_950 ();
 sg13g2_fill_2 FILLER_0_955 ();
 sg13g2_fill_1 FILLER_0_973 ();
 sg13g2_fill_1 FILLER_0_1006 ();
 sg13g2_fill_1 FILLER_0_1019 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_4 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1199 ();
 sg13g2_decap_8 FILLER_0_1206 ();
 sg13g2_decap_4 FILLER_0_1213 ();
 sg13g2_decap_8 FILLER_0_1221 ();
 sg13g2_decap_8 FILLER_0_1228 ();
 sg13g2_fill_1 FILLER_0_1235 ();
 sg13g2_fill_2 FILLER_0_1240 ();
 sg13g2_fill_1 FILLER_0_1242 ();
 sg13g2_fill_2 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1257 ();
 sg13g2_decap_8 FILLER_0_1264 ();
 sg13g2_fill_1 FILLER_0_1271 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_4 FILLER_0_1283 ();
 sg13g2_fill_1 FILLER_0_1287 ();
 sg13g2_decap_4 FILLER_0_1298 ();
 sg13g2_decap_8 FILLER_0_1310 ();
 sg13g2_decap_8 FILLER_0_1343 ();
 sg13g2_decap_8 FILLER_0_1350 ();
 sg13g2_decap_8 FILLER_0_1357 ();
 sg13g2_fill_2 FILLER_0_1364 ();
 sg13g2_fill_1 FILLER_0_1366 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_4 FILLER_0_1449 ();
 sg13g2_fill_1 FILLER_0_1453 ();
 sg13g2_decap_8 FILLER_0_1480 ();
 sg13g2_decap_8 FILLER_0_1487 ();
 sg13g2_decap_8 FILLER_0_1494 ();
 sg13g2_decap_4 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1515 ();
 sg13g2_decap_4 FILLER_0_1522 ();
 sg13g2_fill_2 FILLER_0_1536 ();
 sg13g2_decap_8 FILLER_0_1548 ();
 sg13g2_decap_8 FILLER_0_1555 ();
 sg13g2_decap_8 FILLER_0_1562 ();
 sg13g2_decap_8 FILLER_0_1569 ();
 sg13g2_decap_8 FILLER_0_1576 ();
 sg13g2_decap_8 FILLER_0_1583 ();
 sg13g2_decap_8 FILLER_0_1590 ();
 sg13g2_decap_8 FILLER_0_1597 ();
 sg13g2_decap_8 FILLER_0_1604 ();
 sg13g2_decap_4 FILLER_0_1611 ();
 sg13g2_decap_8 FILLER_0_1641 ();
 sg13g2_decap_8 FILLER_0_1648 ();
 sg13g2_decap_8 FILLER_0_1655 ();
 sg13g2_decap_8 FILLER_0_1662 ();
 sg13g2_decap_8 FILLER_0_1669 ();
 sg13g2_decap_4 FILLER_0_1676 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_fill_2 FILLER_0_1727 ();
 sg13g2_fill_1 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1760 ();
 sg13g2_decap_4 FILLER_0_1767 ();
 sg13g2_fill_2 FILLER_0_1771 ();
 sg13g2_decap_8 FILLER_0_1803 ();
 sg13g2_decap_8 FILLER_0_1810 ();
 sg13g2_decap_8 FILLER_0_1817 ();
 sg13g2_fill_1 FILLER_0_1824 ();
 sg13g2_decap_8 FILLER_0_1851 ();
 sg13g2_decap_8 FILLER_0_1858 ();
 sg13g2_decap_8 FILLER_0_1865 ();
 sg13g2_decap_8 FILLER_0_1898 ();
 sg13g2_decap_8 FILLER_0_1905 ();
 sg13g2_decap_8 FILLER_0_1912 ();
 sg13g2_decap_8 FILLER_0_1953 ();
 sg13g2_fill_2 FILLER_0_1960 ();
 sg13g2_fill_1 FILLER_0_1962 ();
 sg13g2_decap_8 FILLER_0_1989 ();
 sg13g2_decap_8 FILLER_0_1996 ();
 sg13g2_decap_8 FILLER_0_2003 ();
 sg13g2_decap_8 FILLER_0_2010 ();
 sg13g2_fill_2 FILLER_0_2017 ();
 sg13g2_fill_1 FILLER_0_2045 ();
 sg13g2_decap_8 FILLER_0_2067 ();
 sg13g2_decap_8 FILLER_0_2074 ();
 sg13g2_fill_2 FILLER_0_2081 ();
 sg13g2_fill_1 FILLER_0_2083 ();
 sg13g2_decap_8 FILLER_0_2107 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_fill_2 FILLER_0_2121 ();
 sg13g2_decap_8 FILLER_0_2127 ();
 sg13g2_decap_8 FILLER_0_2134 ();
 sg13g2_decap_8 FILLER_0_2141 ();
 sg13g2_decap_4 FILLER_0_2148 ();
 sg13g2_fill_1 FILLER_0_2152 ();
 sg13g2_decap_8 FILLER_0_2183 ();
 sg13g2_fill_2 FILLER_0_2190 ();
 sg13g2_fill_1 FILLER_0_2192 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_4 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2273 ();
 sg13g2_decap_8 FILLER_0_2280 ();
 sg13g2_decap_8 FILLER_0_2287 ();
 sg13g2_decap_8 FILLER_0_2294 ();
 sg13g2_decap_8 FILLER_0_2301 ();
 sg13g2_decap_8 FILLER_0_2308 ();
 sg13g2_decap_8 FILLER_0_2315 ();
 sg13g2_decap_8 FILLER_0_2322 ();
 sg13g2_decap_8 FILLER_0_2329 ();
 sg13g2_decap_8 FILLER_0_2336 ();
 sg13g2_decap_8 FILLER_0_2343 ();
 sg13g2_decap_8 FILLER_0_2350 ();
 sg13g2_decap_8 FILLER_0_2357 ();
 sg13g2_decap_8 FILLER_0_2364 ();
 sg13g2_decap_8 FILLER_0_2371 ();
 sg13g2_decap_8 FILLER_0_2378 ();
 sg13g2_decap_8 FILLER_0_2385 ();
 sg13g2_decap_8 FILLER_0_2392 ();
 sg13g2_decap_8 FILLER_0_2399 ();
 sg13g2_decap_8 FILLER_0_2406 ();
 sg13g2_decap_8 FILLER_0_2413 ();
 sg13g2_decap_8 FILLER_0_2420 ();
 sg13g2_decap_8 FILLER_0_2427 ();
 sg13g2_decap_8 FILLER_0_2434 ();
 sg13g2_decap_8 FILLER_0_2441 ();
 sg13g2_decap_8 FILLER_0_2448 ();
 sg13g2_decap_8 FILLER_0_2455 ();
 sg13g2_decap_8 FILLER_0_2462 ();
 sg13g2_decap_8 FILLER_0_2469 ();
 sg13g2_decap_8 FILLER_0_2476 ();
 sg13g2_decap_8 FILLER_0_2483 ();
 sg13g2_decap_8 FILLER_0_2490 ();
 sg13g2_decap_8 FILLER_0_2497 ();
 sg13g2_decap_8 FILLER_0_2504 ();
 sg13g2_decap_8 FILLER_0_2511 ();
 sg13g2_decap_8 FILLER_0_2518 ();
 sg13g2_decap_8 FILLER_0_2525 ();
 sg13g2_decap_8 FILLER_0_2532 ();
 sg13g2_decap_8 FILLER_0_2539 ();
 sg13g2_decap_8 FILLER_0_2546 ();
 sg13g2_decap_8 FILLER_0_2553 ();
 sg13g2_decap_8 FILLER_0_2560 ();
 sg13g2_decap_8 FILLER_0_2567 ();
 sg13g2_decap_8 FILLER_0_2574 ();
 sg13g2_decap_8 FILLER_0_2581 ();
 sg13g2_decap_8 FILLER_0_2588 ();
 sg13g2_decap_8 FILLER_0_2595 ();
 sg13g2_decap_8 FILLER_0_2602 ();
 sg13g2_decap_8 FILLER_0_2609 ();
 sg13g2_decap_8 FILLER_0_2616 ();
 sg13g2_decap_8 FILLER_0_2623 ();
 sg13g2_decap_8 FILLER_0_2630 ();
 sg13g2_decap_8 FILLER_0_2637 ();
 sg13g2_decap_8 FILLER_0_2644 ();
 sg13g2_decap_8 FILLER_0_2651 ();
 sg13g2_decap_8 FILLER_0_2658 ();
 sg13g2_decap_4 FILLER_0_2665 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_64 ();
 sg13g2_decap_8 FILLER_1_71 ();
 sg13g2_decap_8 FILLER_1_78 ();
 sg13g2_decap_8 FILLER_1_85 ();
 sg13g2_fill_2 FILLER_1_92 ();
 sg13g2_fill_1 FILLER_1_94 ();
 sg13g2_fill_2 FILLER_1_135 ();
 sg13g2_decap_8 FILLER_1_163 ();
 sg13g2_decap_4 FILLER_1_170 ();
 sg13g2_fill_2 FILLER_1_178 ();
 sg13g2_fill_1 FILLER_1_180 ();
 sg13g2_fill_2 FILLER_1_229 ();
 sg13g2_fill_2 FILLER_1_257 ();
 sg13g2_fill_1 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_286 ();
 sg13g2_decap_4 FILLER_1_318 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_2 FILLER_1_332 ();
 sg13g2_fill_1 FILLER_1_334 ();
 sg13g2_fill_2 FILLER_1_339 ();
 sg13g2_fill_2 FILLER_1_367 ();
 sg13g2_fill_1 FILLER_1_369 ();
 sg13g2_decap_4 FILLER_1_374 ();
 sg13g2_fill_2 FILLER_1_378 ();
 sg13g2_fill_2 FILLER_1_454 ();
 sg13g2_decap_8 FILLER_1_487 ();
 sg13g2_decap_8 FILLER_1_550 ();
 sg13g2_fill_1 FILLER_1_557 ();
 sg13g2_fill_2 FILLER_1_584 ();
 sg13g2_fill_1 FILLER_1_586 ();
 sg13g2_fill_2 FILLER_1_687 ();
 sg13g2_fill_2 FILLER_1_710 ();
 sg13g2_fill_1 FILLER_1_712 ();
 sg13g2_decap_8 FILLER_1_717 ();
 sg13g2_decap_4 FILLER_1_754 ();
 sg13g2_fill_1 FILLER_1_758 ();
 sg13g2_decap_8 FILLER_1_792 ();
 sg13g2_decap_4 FILLER_1_813 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_fill_1 FILLER_1_866 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_fill_1 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_922 ();
 sg13g2_decap_4 FILLER_1_929 ();
 sg13g2_fill_1 FILLER_1_933 ();
 sg13g2_fill_1 FILLER_1_970 ();
 sg13g2_fill_1 FILLER_1_977 ();
 sg13g2_fill_2 FILLER_1_1014 ();
 sg13g2_fill_1 FILLER_1_1039 ();
 sg13g2_decap_4 FILLER_1_1057 ();
 sg13g2_fill_2 FILLER_1_1065 ();
 sg13g2_fill_1 FILLER_1_1067 ();
 sg13g2_decap_4 FILLER_1_1082 ();
 sg13g2_fill_1 FILLER_1_1086 ();
 sg13g2_decap_8 FILLER_1_1097 ();
 sg13g2_decap_8 FILLER_1_1104 ();
 sg13g2_fill_2 FILLER_1_1111 ();
 sg13g2_fill_1 FILLER_1_1139 ();
 sg13g2_fill_1 FILLER_1_1166 ();
 sg13g2_fill_2 FILLER_1_1177 ();
 sg13g2_fill_1 FILLER_1_1205 ();
 sg13g2_fill_2 FILLER_1_1210 ();
 sg13g2_fill_1 FILLER_1_1222 ();
 sg13g2_fill_2 FILLER_1_1227 ();
 sg13g2_decap_4 FILLER_1_1321 ();
 sg13g2_decap_8 FILLER_1_1339 ();
 sg13g2_decap_8 FILLER_1_1346 ();
 sg13g2_decap_4 FILLER_1_1353 ();
 sg13g2_fill_1 FILLER_1_1357 ();
 sg13g2_decap_8 FILLER_1_1368 ();
 sg13g2_decap_4 FILLER_1_1441 ();
 sg13g2_fill_1 FILLER_1_1445 ();
 sg13g2_decap_4 FILLER_1_1450 ();
 sg13g2_fill_1 FILLER_1_1454 ();
 sg13g2_fill_2 FILLER_1_1465 ();
 sg13g2_fill_1 FILLER_1_1467 ();
 sg13g2_decap_8 FILLER_1_1472 ();
 sg13g2_decap_8 FILLER_1_1479 ();
 sg13g2_fill_2 FILLER_1_1486 ();
 sg13g2_fill_1 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1571 ();
 sg13g2_decap_8 FILLER_1_1578 ();
 sg13g2_decap_8 FILLER_1_1585 ();
 sg13g2_decap_8 FILLER_1_1592 ();
 sg13g2_fill_1 FILLER_1_1599 ();
 sg13g2_decap_4 FILLER_1_1640 ();
 sg13g2_fill_1 FILLER_1_1674 ();
 sg13g2_decap_8 FILLER_1_1701 ();
 sg13g2_decap_4 FILLER_1_1718 ();
 sg13g2_fill_2 FILLER_1_1722 ();
 sg13g2_decap_4 FILLER_1_1750 ();
 sg13g2_fill_1 FILLER_1_1754 ();
 sg13g2_fill_2 FILLER_1_1765 ();
 sg13g2_decap_8 FILLER_1_1803 ();
 sg13g2_fill_2 FILLER_1_1810 ();
 sg13g2_fill_1 FILLER_1_1816 ();
 sg13g2_fill_1 FILLER_1_1847 ();
 sg13g2_fill_2 FILLER_1_1874 ();
 sg13g2_fill_2 FILLER_1_1880 ();
 sg13g2_fill_2 FILLER_1_1903 ();
 sg13g2_fill_1 FILLER_1_1905 ();
 sg13g2_fill_1 FILLER_1_1932 ();
 sg13g2_decap_8 FILLER_1_1995 ();
 sg13g2_decap_4 FILLER_1_2002 ();
 sg13g2_fill_2 FILLER_1_2006 ();
 sg13g2_fill_2 FILLER_1_2018 ();
 sg13g2_fill_1 FILLER_1_2020 ();
 sg13g2_decap_8 FILLER_1_2047 ();
 sg13g2_decap_4 FILLER_1_2054 ();
 sg13g2_fill_2 FILLER_1_2058 ();
 sg13g2_decap_4 FILLER_1_2142 ();
 sg13g2_fill_1 FILLER_1_2146 ();
 sg13g2_fill_2 FILLER_1_2203 ();
 sg13g2_decap_4 FILLER_1_2231 ();
 sg13g2_fill_1 FILLER_1_2235 ();
 sg13g2_decap_4 FILLER_1_2257 ();
 sg13g2_fill_1 FILLER_1_2261 ();
 sg13g2_decap_8 FILLER_1_2288 ();
 sg13g2_decap_8 FILLER_1_2295 ();
 sg13g2_decap_8 FILLER_1_2302 ();
 sg13g2_decap_8 FILLER_1_2309 ();
 sg13g2_decap_8 FILLER_1_2316 ();
 sg13g2_decap_8 FILLER_1_2323 ();
 sg13g2_decap_8 FILLER_1_2330 ();
 sg13g2_decap_8 FILLER_1_2337 ();
 sg13g2_decap_8 FILLER_1_2344 ();
 sg13g2_decap_8 FILLER_1_2351 ();
 sg13g2_decap_8 FILLER_1_2358 ();
 sg13g2_decap_8 FILLER_1_2365 ();
 sg13g2_decap_8 FILLER_1_2372 ();
 sg13g2_decap_8 FILLER_1_2379 ();
 sg13g2_decap_8 FILLER_1_2386 ();
 sg13g2_decap_8 FILLER_1_2393 ();
 sg13g2_decap_8 FILLER_1_2400 ();
 sg13g2_decap_8 FILLER_1_2407 ();
 sg13g2_decap_8 FILLER_1_2414 ();
 sg13g2_decap_8 FILLER_1_2421 ();
 sg13g2_decap_8 FILLER_1_2428 ();
 sg13g2_decap_8 FILLER_1_2435 ();
 sg13g2_decap_8 FILLER_1_2442 ();
 sg13g2_decap_8 FILLER_1_2449 ();
 sg13g2_decap_8 FILLER_1_2456 ();
 sg13g2_decap_8 FILLER_1_2463 ();
 sg13g2_decap_8 FILLER_1_2470 ();
 sg13g2_decap_8 FILLER_1_2477 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_decap_8 FILLER_1_2491 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_decap_8 FILLER_1_2505 ();
 sg13g2_decap_8 FILLER_1_2512 ();
 sg13g2_decap_8 FILLER_1_2519 ();
 sg13g2_decap_8 FILLER_1_2526 ();
 sg13g2_decap_8 FILLER_1_2533 ();
 sg13g2_decap_8 FILLER_1_2540 ();
 sg13g2_decap_8 FILLER_1_2547 ();
 sg13g2_decap_8 FILLER_1_2554 ();
 sg13g2_decap_8 FILLER_1_2561 ();
 sg13g2_decap_8 FILLER_1_2568 ();
 sg13g2_decap_8 FILLER_1_2575 ();
 sg13g2_decap_8 FILLER_1_2582 ();
 sg13g2_decap_8 FILLER_1_2589 ();
 sg13g2_decap_8 FILLER_1_2596 ();
 sg13g2_decap_8 FILLER_1_2603 ();
 sg13g2_decap_8 FILLER_1_2610 ();
 sg13g2_decap_8 FILLER_1_2617 ();
 sg13g2_decap_8 FILLER_1_2624 ();
 sg13g2_decap_8 FILLER_1_2631 ();
 sg13g2_decap_8 FILLER_1_2638 ();
 sg13g2_decap_8 FILLER_1_2645 ();
 sg13g2_decap_8 FILLER_1_2652 ();
 sg13g2_decap_8 FILLER_1_2659 ();
 sg13g2_decap_4 FILLER_1_2666 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_decap_4 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_83 ();
 sg13g2_fill_2 FILLER_2_132 ();
 sg13g2_fill_1 FILLER_2_134 ();
 sg13g2_decap_4 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_170 ();
 sg13g2_fill_1 FILLER_2_211 ();
 sg13g2_fill_2 FILLER_2_216 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_decap_4 FILLER_2_254 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_fill_1 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_352 ();
 sg13g2_fill_2 FILLER_2_396 ();
 sg13g2_fill_1 FILLER_2_398 ();
 sg13g2_fill_1 FILLER_2_413 ();
 sg13g2_fill_2 FILLER_2_424 ();
 sg13g2_fill_1 FILLER_2_426 ();
 sg13g2_fill_1 FILLER_2_432 ();
 sg13g2_fill_1 FILLER_2_437 ();
 sg13g2_fill_2 FILLER_2_474 ();
 sg13g2_fill_2 FILLER_2_520 ();
 sg13g2_fill_1 FILLER_2_522 ();
 sg13g2_fill_1 FILLER_2_528 ();
 sg13g2_fill_1 FILLER_2_534 ();
 sg13g2_fill_1 FILLER_2_539 ();
 sg13g2_fill_2 FILLER_2_550 ();
 sg13g2_fill_2 FILLER_2_583 ();
 sg13g2_fill_1 FILLER_2_585 ();
 sg13g2_fill_2 FILLER_2_621 ();
 sg13g2_fill_1 FILLER_2_635 ();
 sg13g2_fill_2 FILLER_2_642 ();
 sg13g2_fill_1 FILLER_2_648 ();
 sg13g2_fill_1 FILLER_2_653 ();
 sg13g2_fill_2 FILLER_2_668 ();
 sg13g2_decap_4 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_4 FILLER_2_725 ();
 sg13g2_fill_1 FILLER_2_729 ();
 sg13g2_fill_1 FILLER_2_756 ();
 sg13g2_fill_2 FILLER_2_767 ();
 sg13g2_fill_2 FILLER_2_773 ();
 sg13g2_fill_1 FILLER_2_775 ();
 sg13g2_fill_1 FILLER_2_821 ();
 sg13g2_fill_1 FILLER_2_848 ();
 sg13g2_fill_2 FILLER_2_853 ();
 sg13g2_fill_2 FILLER_2_891 ();
 sg13g2_fill_2 FILLER_2_945 ();
 sg13g2_fill_1 FILLER_2_951 ();
 sg13g2_fill_1 FILLER_2_1017 ();
 sg13g2_fill_2 FILLER_2_1050 ();
 sg13g2_fill_2 FILLER_2_1078 ();
 sg13g2_fill_2 FILLER_2_1097 ();
 sg13g2_fill_1 FILLER_2_1099 ();
 sg13g2_fill_1 FILLER_2_1156 ();
 sg13g2_fill_2 FILLER_2_1167 ();
 sg13g2_fill_1 FILLER_2_1169 ();
 sg13g2_fill_1 FILLER_2_1193 ();
 sg13g2_fill_1 FILLER_2_1324 ();
 sg13g2_decap_4 FILLER_2_1351 ();
 sg13g2_fill_1 FILLER_2_1385 ();
 sg13g2_fill_1 FILLER_2_1396 ();
 sg13g2_fill_2 FILLER_2_1466 ();
 sg13g2_fill_1 FILLER_2_1482 ();
 sg13g2_fill_1 FILLER_2_1493 ();
 sg13g2_fill_1 FILLER_2_1498 ();
 sg13g2_fill_1 FILLER_2_1525 ();
 sg13g2_decap_8 FILLER_2_1566 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_decap_8 FILLER_2_1580 ();
 sg13g2_decap_8 FILLER_2_1587 ();
 sg13g2_fill_2 FILLER_2_1594 ();
 sg13g2_fill_1 FILLER_2_1596 ();
 sg13g2_decap_8 FILLER_2_1633 ();
 sg13g2_fill_1 FILLER_2_1680 ();
 sg13g2_fill_2 FILLER_2_1707 ();
 sg13g2_fill_1 FILLER_2_1709 ();
 sg13g2_fill_2 FILLER_2_1713 ();
 sg13g2_fill_1 FILLER_2_1715 ();
 sg13g2_fill_1 FILLER_2_1786 ();
 sg13g2_fill_1 FILLER_2_1797 ();
 sg13g2_decap_4 FILLER_2_1860 ();
 sg13g2_fill_1 FILLER_2_1864 ();
 sg13g2_fill_2 FILLER_2_1925 ();
 sg13g2_fill_2 FILLER_2_1997 ();
 sg13g2_fill_2 FILLER_2_2029 ();
 sg13g2_fill_2 FILLER_2_2035 ();
 sg13g2_fill_2 FILLER_2_2073 ();
 sg13g2_fill_1 FILLER_2_2129 ();
 sg13g2_fill_1 FILLER_2_2207 ();
 sg13g2_decap_4 FILLER_2_2233 ();
 sg13g2_fill_2 FILLER_2_2237 ();
 sg13g2_fill_2 FILLER_2_2249 ();
 sg13g2_fill_1 FILLER_2_2251 ();
 sg13g2_fill_1 FILLER_2_2262 ();
 sg13g2_fill_2 FILLER_2_2267 ();
 sg13g2_decap_8 FILLER_2_2273 ();
 sg13g2_decap_8 FILLER_2_2280 ();
 sg13g2_decap_8 FILLER_2_2287 ();
 sg13g2_decap_8 FILLER_2_2294 ();
 sg13g2_decap_8 FILLER_2_2301 ();
 sg13g2_decap_8 FILLER_2_2308 ();
 sg13g2_decap_8 FILLER_2_2315 ();
 sg13g2_decap_8 FILLER_2_2322 ();
 sg13g2_decap_8 FILLER_2_2329 ();
 sg13g2_decap_8 FILLER_2_2336 ();
 sg13g2_decap_8 FILLER_2_2343 ();
 sg13g2_decap_8 FILLER_2_2350 ();
 sg13g2_decap_8 FILLER_2_2357 ();
 sg13g2_decap_8 FILLER_2_2364 ();
 sg13g2_decap_8 FILLER_2_2371 ();
 sg13g2_decap_8 FILLER_2_2378 ();
 sg13g2_decap_8 FILLER_2_2385 ();
 sg13g2_decap_8 FILLER_2_2392 ();
 sg13g2_decap_8 FILLER_2_2399 ();
 sg13g2_decap_8 FILLER_2_2406 ();
 sg13g2_decap_8 FILLER_2_2413 ();
 sg13g2_decap_8 FILLER_2_2420 ();
 sg13g2_decap_8 FILLER_2_2427 ();
 sg13g2_decap_8 FILLER_2_2434 ();
 sg13g2_decap_8 FILLER_2_2441 ();
 sg13g2_decap_8 FILLER_2_2448 ();
 sg13g2_decap_8 FILLER_2_2455 ();
 sg13g2_decap_8 FILLER_2_2462 ();
 sg13g2_decap_8 FILLER_2_2469 ();
 sg13g2_decap_8 FILLER_2_2476 ();
 sg13g2_decap_8 FILLER_2_2483 ();
 sg13g2_decap_8 FILLER_2_2490 ();
 sg13g2_decap_8 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2504 ();
 sg13g2_decap_8 FILLER_2_2511 ();
 sg13g2_decap_8 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_61 ();
 sg13g2_fill_1 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_76 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_108 ();
 sg13g2_fill_1 FILLER_3_123 ();
 sg13g2_fill_2 FILLER_3_132 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_166 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_201 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_fill_2 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_246 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_fill_2 FILLER_3_292 ();
 sg13g2_fill_1 FILLER_3_304 ();
 sg13g2_fill_1 FILLER_3_310 ();
 sg13g2_fill_1 FILLER_3_316 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_4 FILLER_3_379 ();
 sg13g2_fill_1 FILLER_3_383 ();
 sg13g2_fill_2 FILLER_3_447 ();
 sg13g2_decap_8 FILLER_3_454 ();
 sg13g2_fill_2 FILLER_3_461 ();
 sg13g2_fill_1 FILLER_3_463 ();
 sg13g2_fill_2 FILLER_3_469 ();
 sg13g2_decap_4 FILLER_3_476 ();
 sg13g2_fill_2 FILLER_3_484 ();
 sg13g2_fill_2 FILLER_3_512 ();
 sg13g2_fill_1 FILLER_3_514 ();
 sg13g2_fill_2 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_527 ();
 sg13g2_fill_2 FILLER_3_554 ();
 sg13g2_fill_1 FILLER_3_556 ();
 sg13g2_decap_4 FILLER_3_566 ();
 sg13g2_fill_2 FILLER_3_594 ();
 sg13g2_fill_1 FILLER_3_596 ();
 sg13g2_fill_2 FILLER_3_610 ();
 sg13g2_fill_1 FILLER_3_622 ();
 sg13g2_fill_2 FILLER_3_637 ();
 sg13g2_fill_2 FILLER_3_644 ();
 sg13g2_fill_1 FILLER_3_670 ();
 sg13g2_decap_4 FILLER_3_676 ();
 sg13g2_fill_1 FILLER_3_688 ();
 sg13g2_fill_1 FILLER_3_708 ();
 sg13g2_fill_1 FILLER_3_714 ();
 sg13g2_fill_2 FILLER_3_784 ();
 sg13g2_fill_1 FILLER_3_786 ();
 sg13g2_decap_4 FILLER_3_823 ();
 sg13g2_fill_1 FILLER_3_827 ();
 sg13g2_decap_8 FILLER_3_832 ();
 sg13g2_decap_8 FILLER_3_932 ();
 sg13g2_fill_1 FILLER_3_939 ();
 sg13g2_fill_1 FILLER_3_970 ();
 sg13g2_fill_1 FILLER_3_1035 ();
 sg13g2_fill_2 FILLER_3_1040 ();
 sg13g2_decap_8 FILLER_3_1068 ();
 sg13g2_decap_8 FILLER_3_1075 ();
 sg13g2_fill_1 FILLER_3_1082 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_fill_1 FILLER_3_1134 ();
 sg13g2_decap_8 FILLER_3_1153 ();
 sg13g2_fill_2 FILLER_3_1160 ();
 sg13g2_fill_2 FILLER_3_1212 ();
 sg13g2_fill_1 FILLER_3_1246 ();
 sg13g2_fill_2 FILLER_3_1290 ();
 sg13g2_decap_4 FILLER_3_1328 ();
 sg13g2_decap_8 FILLER_3_1336 ();
 sg13g2_decap_8 FILLER_3_1343 ();
 sg13g2_fill_2 FILLER_3_1350 ();
 sg13g2_fill_1 FILLER_3_1352 ();
 sg13g2_decap_8 FILLER_3_1357 ();
 sg13g2_fill_1 FILLER_3_1364 ();
 sg13g2_fill_2 FILLER_3_1375 ();
 sg13g2_fill_2 FILLER_3_1381 ();
 sg13g2_fill_1 FILLER_3_1387 ();
 sg13g2_fill_1 FILLER_3_1392 ();
 sg13g2_fill_2 FILLER_3_1403 ();
 sg13g2_fill_2 FILLER_3_1409 ();
 sg13g2_fill_2 FILLER_3_1447 ();
 sg13g2_decap_4 FILLER_3_1485 ();
 sg13g2_fill_1 FILLER_3_1493 ();
 sg13g2_fill_2 FILLER_3_1504 ();
 sg13g2_fill_1 FILLER_3_1516 ();
 sg13g2_fill_2 FILLER_3_1521 ();
 sg13g2_fill_1 FILLER_3_1527 ();
 sg13g2_fill_1 FILLER_3_1545 ();
 sg13g2_decap_8 FILLER_3_1572 ();
 sg13g2_fill_2 FILLER_3_1579 ();
 sg13g2_decap_4 FILLER_3_1611 ();
 sg13g2_fill_2 FILLER_3_1619 ();
 sg13g2_fill_2 FILLER_3_1642 ();
 sg13g2_decap_8 FILLER_3_1648 ();
 sg13g2_decap_4 FILLER_3_1665 ();
 sg13g2_decap_4 FILLER_3_1714 ();
 sg13g2_fill_1 FILLER_3_1718 ();
 sg13g2_fill_2 FILLER_3_1750 ();
 sg13g2_fill_2 FILLER_3_1778 ();
 sg13g2_fill_1 FILLER_3_1780 ();
 sg13g2_fill_1 FILLER_3_1825 ();
 sg13g2_fill_2 FILLER_3_1836 ();
 sg13g2_fill_2 FILLER_3_1859 ();
 sg13g2_fill_1 FILLER_3_1913 ();
 sg13g2_decap_8 FILLER_3_1949 ();
 sg13g2_decap_8 FILLER_3_1956 ();
 sg13g2_decap_4 FILLER_3_1963 ();
 sg13g2_fill_2 FILLER_3_1967 ();
 sg13g2_fill_1 FILLER_3_2010 ();
 sg13g2_decap_4 FILLER_3_2015 ();
 sg13g2_fill_2 FILLER_3_2029 ();
 sg13g2_fill_1 FILLER_3_2031 ();
 sg13g2_fill_2 FILLER_3_2042 ();
 sg13g2_decap_4 FILLER_3_2080 ();
 sg13g2_fill_1 FILLER_3_2084 ();
 sg13g2_decap_4 FILLER_3_2106 ();
 sg13g2_fill_1 FILLER_3_2140 ();
 sg13g2_decap_4 FILLER_3_2151 ();
 sg13g2_fill_1 FILLER_3_2155 ();
 sg13g2_decap_4 FILLER_3_2179 ();
 sg13g2_fill_1 FILLER_3_2183 ();
 sg13g2_decap_8 FILLER_3_2231 ();
 sg13g2_fill_2 FILLER_3_2238 ();
 sg13g2_fill_1 FILLER_3_2240 ();
 sg13g2_decap_8 FILLER_3_2277 ();
 sg13g2_decap_8 FILLER_3_2284 ();
 sg13g2_decap_8 FILLER_3_2291 ();
 sg13g2_decap_8 FILLER_3_2298 ();
 sg13g2_decap_8 FILLER_3_2305 ();
 sg13g2_decap_8 FILLER_3_2312 ();
 sg13g2_decap_8 FILLER_3_2319 ();
 sg13g2_decap_8 FILLER_3_2326 ();
 sg13g2_decap_8 FILLER_3_2333 ();
 sg13g2_decap_8 FILLER_3_2340 ();
 sg13g2_decap_8 FILLER_3_2347 ();
 sg13g2_decap_8 FILLER_3_2354 ();
 sg13g2_decap_8 FILLER_3_2361 ();
 sg13g2_decap_8 FILLER_3_2368 ();
 sg13g2_decap_8 FILLER_3_2375 ();
 sg13g2_decap_8 FILLER_3_2382 ();
 sg13g2_decap_8 FILLER_3_2389 ();
 sg13g2_decap_8 FILLER_3_2396 ();
 sg13g2_decap_8 FILLER_3_2403 ();
 sg13g2_decap_8 FILLER_3_2410 ();
 sg13g2_decap_8 FILLER_3_2417 ();
 sg13g2_decap_8 FILLER_3_2424 ();
 sg13g2_decap_8 FILLER_3_2431 ();
 sg13g2_decap_8 FILLER_3_2438 ();
 sg13g2_decap_8 FILLER_3_2445 ();
 sg13g2_decap_8 FILLER_3_2452 ();
 sg13g2_decap_8 FILLER_3_2459 ();
 sg13g2_decap_8 FILLER_3_2466 ();
 sg13g2_decap_8 FILLER_3_2473 ();
 sg13g2_decap_8 FILLER_3_2480 ();
 sg13g2_decap_8 FILLER_3_2487 ();
 sg13g2_decap_8 FILLER_3_2494 ();
 sg13g2_decap_8 FILLER_3_2501 ();
 sg13g2_decap_8 FILLER_3_2508 ();
 sg13g2_decap_8 FILLER_3_2515 ();
 sg13g2_decap_8 FILLER_3_2522 ();
 sg13g2_decap_8 FILLER_3_2529 ();
 sg13g2_decap_8 FILLER_3_2536 ();
 sg13g2_decap_8 FILLER_3_2543 ();
 sg13g2_decap_8 FILLER_3_2550 ();
 sg13g2_decap_8 FILLER_3_2557 ();
 sg13g2_decap_8 FILLER_3_2564 ();
 sg13g2_decap_8 FILLER_3_2571 ();
 sg13g2_decap_8 FILLER_3_2578 ();
 sg13g2_decap_8 FILLER_3_2585 ();
 sg13g2_decap_8 FILLER_3_2592 ();
 sg13g2_decap_8 FILLER_3_2599 ();
 sg13g2_decap_8 FILLER_3_2606 ();
 sg13g2_decap_8 FILLER_3_2613 ();
 sg13g2_decap_8 FILLER_3_2620 ();
 sg13g2_decap_8 FILLER_3_2627 ();
 sg13g2_decap_8 FILLER_3_2634 ();
 sg13g2_decap_8 FILLER_3_2641 ();
 sg13g2_decap_8 FILLER_3_2648 ();
 sg13g2_decap_8 FILLER_3_2655 ();
 sg13g2_decap_8 FILLER_3_2662 ();
 sg13g2_fill_1 FILLER_3_2669 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_46 ();
 sg13g2_fill_1 FILLER_4_78 ();
 sg13g2_fill_1 FILLER_4_88 ();
 sg13g2_fill_1 FILLER_4_102 ();
 sg13g2_decap_4 FILLER_4_108 ();
 sg13g2_fill_2 FILLER_4_112 ();
 sg13g2_decap_4 FILLER_4_128 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_fill_2 FILLER_4_142 ();
 sg13g2_decap_4 FILLER_4_170 ();
 sg13g2_fill_1 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_298 ();
 sg13g2_fill_1 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_315 ();
 sg13g2_fill_1 FILLER_4_336 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_365 ();
 sg13g2_fill_2 FILLER_4_377 ();
 sg13g2_fill_1 FILLER_4_379 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_fill_2 FILLER_4_412 ();
 sg13g2_fill_1 FILLER_4_414 ();
 sg13g2_decap_4 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_fill_1 FILLER_4_430 ();
 sg13g2_decap_4 FILLER_4_436 ();
 sg13g2_fill_2 FILLER_4_440 ();
 sg13g2_fill_2 FILLER_4_447 ();
 sg13g2_decap_4 FILLER_4_463 ();
 sg13g2_fill_1 FILLER_4_477 ();
 sg13g2_decap_8 FILLER_4_484 ();
 sg13g2_fill_2 FILLER_4_491 ();
 sg13g2_fill_1 FILLER_4_493 ();
 sg13g2_decap_8 FILLER_4_498 ();
 sg13g2_fill_1 FILLER_4_505 ();
 sg13g2_fill_2 FILLER_4_541 ();
 sg13g2_decap_8 FILLER_4_552 ();
 sg13g2_decap_4 FILLER_4_559 ();
 sg13g2_fill_2 FILLER_4_563 ();
 sg13g2_fill_1 FILLER_4_587 ();
 sg13g2_fill_1 FILLER_4_597 ();
 sg13g2_fill_1 FILLER_4_643 ();
 sg13g2_decap_4 FILLER_4_668 ();
 sg13g2_fill_1 FILLER_4_672 ();
 sg13g2_fill_1 FILLER_4_679 ();
 sg13g2_fill_1 FILLER_4_685 ();
 sg13g2_decap_4 FILLER_4_723 ();
 sg13g2_fill_1 FILLER_4_727 ();
 sg13g2_fill_2 FILLER_4_755 ();
 sg13g2_fill_1 FILLER_4_757 ();
 sg13g2_fill_2 FILLER_4_768 ();
 sg13g2_fill_1 FILLER_4_770 ();
 sg13g2_fill_1 FILLER_4_777 ();
 sg13g2_fill_1 FILLER_4_784 ();
 sg13g2_fill_2 FILLER_4_795 ();
 sg13g2_fill_1 FILLER_4_797 ();
 sg13g2_fill_2 FILLER_4_828 ();
 sg13g2_fill_2 FILLER_4_878 ();
 sg13g2_fill_1 FILLER_4_890 ();
 sg13g2_fill_1 FILLER_4_901 ();
 sg13g2_decap_8 FILLER_4_906 ();
 sg13g2_fill_1 FILLER_4_913 ();
 sg13g2_fill_1 FILLER_4_920 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_decap_4 FILLER_4_941 ();
 sg13g2_fill_1 FILLER_4_1052 ();
 sg13g2_decap_8 FILLER_4_1080 ();
 sg13g2_fill_2 FILLER_4_1087 ();
 sg13g2_decap_4 FILLER_4_1093 ();
 sg13g2_fill_1 FILLER_4_1109 ();
 sg13g2_fill_2 FILLER_4_1119 ();
 sg13g2_fill_1 FILLER_4_1121 ();
 sg13g2_fill_1 FILLER_4_1132 ();
 sg13g2_fill_2 FILLER_4_1205 ();
 sg13g2_fill_1 FILLER_4_1207 ();
 sg13g2_fill_2 FILLER_4_1218 ();
 sg13g2_fill_2 FILLER_4_1238 ();
 sg13g2_fill_2 FILLER_4_1304 ();
 sg13g2_fill_1 FILLER_4_1306 ();
 sg13g2_decap_8 FILLER_4_1311 ();
 sg13g2_fill_1 FILLER_4_1318 ();
 sg13g2_fill_1 FILLER_4_1329 ();
 sg13g2_decap_4 FILLER_4_1340 ();
 sg13g2_decap_8 FILLER_4_1370 ();
 sg13g2_decap_4 FILLER_4_1377 ();
 sg13g2_fill_2 FILLER_4_1381 ();
 sg13g2_fill_1 FILLER_4_1393 ();
 sg13g2_decap_8 FILLER_4_1398 ();
 sg13g2_fill_2 FILLER_4_1405 ();
 sg13g2_fill_1 FILLER_4_1480 ();
 sg13g2_fill_1 FILLER_4_1507 ();
 sg13g2_decap_8 FILLER_4_1534 ();
 sg13g2_decap_8 FILLER_4_1571 ();
 sg13g2_decap_8 FILLER_4_1578 ();
 sg13g2_decap_4 FILLER_4_1585 ();
 sg13g2_fill_1 FILLER_4_1589 ();
 sg13g2_fill_2 FILLER_4_1594 ();
 sg13g2_fill_2 FILLER_4_1606 ();
 sg13g2_fill_1 FILLER_4_1618 ();
 sg13g2_fill_1 FILLER_4_1632 ();
 sg13g2_decap_8 FILLER_4_1667 ();
 sg13g2_decap_4 FILLER_4_1674 ();
 sg13g2_fill_1 FILLER_4_1682 ();
 sg13g2_fill_1 FILLER_4_1693 ();
 sg13g2_decap_8 FILLER_4_1724 ();
 sg13g2_fill_2 FILLER_4_1731 ();
 sg13g2_fill_1 FILLER_4_1777 ();
 sg13g2_decap_8 FILLER_4_1782 ();
 sg13g2_fill_2 FILLER_4_1789 ();
 sg13g2_decap_4 FILLER_4_1841 ();
 sg13g2_fill_1 FILLER_4_1845 ();
 sg13g2_decap_4 FILLER_4_1856 ();
 sg13g2_fill_2 FILLER_4_1889 ();
 sg13g2_fill_1 FILLER_4_1899 ();
 sg13g2_fill_1 FILLER_4_1919 ();
 sg13g2_decap_8 FILLER_4_1946 ();
 sg13g2_fill_1 FILLER_4_1953 ();
 sg13g2_decap_4 FILLER_4_2077 ();
 sg13g2_fill_1 FILLER_4_2081 ();
 sg13g2_decap_4 FILLER_4_2092 ();
 sg13g2_fill_2 FILLER_4_2096 ();
 sg13g2_decap_4 FILLER_4_2112 ();
 sg13g2_fill_1 FILLER_4_2116 ();
 sg13g2_decap_8 FILLER_4_2122 ();
 sg13g2_decap_8 FILLER_4_2129 ();
 sg13g2_fill_2 FILLER_4_2136 ();
 sg13g2_fill_1 FILLER_4_2138 ();
 sg13g2_decap_4 FILLER_4_2143 ();
 sg13g2_decap_4 FILLER_4_2167 ();
 sg13g2_fill_2 FILLER_4_2171 ();
 sg13g2_decap_4 FILLER_4_2209 ();
 sg13g2_fill_2 FILLER_4_2213 ();
 sg13g2_fill_2 FILLER_4_2255 ();
 sg13g2_decap_8 FILLER_4_2287 ();
 sg13g2_decap_8 FILLER_4_2294 ();
 sg13g2_decap_8 FILLER_4_2301 ();
 sg13g2_decap_8 FILLER_4_2308 ();
 sg13g2_decap_8 FILLER_4_2315 ();
 sg13g2_decap_8 FILLER_4_2322 ();
 sg13g2_decap_8 FILLER_4_2329 ();
 sg13g2_decap_8 FILLER_4_2336 ();
 sg13g2_decap_8 FILLER_4_2343 ();
 sg13g2_decap_8 FILLER_4_2350 ();
 sg13g2_decap_8 FILLER_4_2357 ();
 sg13g2_decap_8 FILLER_4_2364 ();
 sg13g2_decap_8 FILLER_4_2371 ();
 sg13g2_decap_8 FILLER_4_2378 ();
 sg13g2_decap_8 FILLER_4_2385 ();
 sg13g2_decap_8 FILLER_4_2392 ();
 sg13g2_decap_8 FILLER_4_2399 ();
 sg13g2_decap_8 FILLER_4_2406 ();
 sg13g2_decap_8 FILLER_4_2413 ();
 sg13g2_decap_8 FILLER_4_2420 ();
 sg13g2_decap_8 FILLER_4_2427 ();
 sg13g2_decap_8 FILLER_4_2434 ();
 sg13g2_decap_8 FILLER_4_2441 ();
 sg13g2_decap_8 FILLER_4_2448 ();
 sg13g2_decap_8 FILLER_4_2455 ();
 sg13g2_decap_8 FILLER_4_2462 ();
 sg13g2_decap_8 FILLER_4_2469 ();
 sg13g2_decap_8 FILLER_4_2476 ();
 sg13g2_decap_8 FILLER_4_2483 ();
 sg13g2_decap_8 FILLER_4_2490 ();
 sg13g2_decap_8 FILLER_4_2497 ();
 sg13g2_decap_8 FILLER_4_2504 ();
 sg13g2_decap_8 FILLER_4_2511 ();
 sg13g2_decap_8 FILLER_4_2518 ();
 sg13g2_decap_8 FILLER_4_2525 ();
 sg13g2_decap_8 FILLER_4_2532 ();
 sg13g2_decap_8 FILLER_4_2539 ();
 sg13g2_decap_8 FILLER_4_2546 ();
 sg13g2_decap_8 FILLER_4_2553 ();
 sg13g2_decap_8 FILLER_4_2560 ();
 sg13g2_decap_8 FILLER_4_2567 ();
 sg13g2_decap_8 FILLER_4_2574 ();
 sg13g2_decap_8 FILLER_4_2581 ();
 sg13g2_decap_8 FILLER_4_2588 ();
 sg13g2_decap_8 FILLER_4_2595 ();
 sg13g2_decap_8 FILLER_4_2602 ();
 sg13g2_decap_8 FILLER_4_2609 ();
 sg13g2_decap_8 FILLER_4_2616 ();
 sg13g2_decap_8 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_4 FILLER_4_2665 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_60 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_4 FILLER_5_99 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_114 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_146 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_fill_2 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_decap_4 FILLER_5_290 ();
 sg13g2_fill_2 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_332 ();
 sg13g2_fill_1 FILLER_5_334 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_fill_1 FILLER_5_355 ();
 sg13g2_fill_1 FILLER_5_361 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_decap_4 FILLER_5_375 ();
 sg13g2_fill_1 FILLER_5_387 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_5_440 ();
 sg13g2_fill_1 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_467 ();
 sg13g2_fill_1 FILLER_5_472 ();
 sg13g2_fill_1 FILLER_5_477 ();
 sg13g2_fill_2 FILLER_5_488 ();
 sg13g2_fill_1 FILLER_5_490 ();
 sg13g2_fill_2 FILLER_5_501 ();
 sg13g2_fill_1 FILLER_5_503 ();
 sg13g2_fill_2 FILLER_5_530 ();
 sg13g2_fill_1 FILLER_5_542 ();
 sg13g2_fill_2 FILLER_5_553 ();
 sg13g2_fill_2 FILLER_5_587 ();
 sg13g2_fill_1 FILLER_5_593 ();
 sg13g2_decap_4 FILLER_5_598 ();
 sg13g2_fill_2 FILLER_5_602 ();
 sg13g2_fill_1 FILLER_5_612 ();
 sg13g2_decap_4 FILLER_5_617 ();
 sg13g2_fill_2 FILLER_5_621 ();
 sg13g2_fill_2 FILLER_5_627 ();
 sg13g2_fill_1 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_678 ();
 sg13g2_decap_4 FILLER_5_685 ();
 sg13g2_fill_1 FILLER_5_689 ();
 sg13g2_fill_1 FILLER_5_703 ();
 sg13g2_fill_2 FILLER_5_730 ();
 sg13g2_fill_1 FILLER_5_736 ();
 sg13g2_fill_2 FILLER_5_763 ();
 sg13g2_fill_2 FILLER_5_797 ();
 sg13g2_fill_2 FILLER_5_803 ();
 sg13g2_fill_1 FILLER_5_805 ();
 sg13g2_fill_2 FILLER_5_810 ();
 sg13g2_fill_1 FILLER_5_812 ();
 sg13g2_decap_4 FILLER_5_823 ();
 sg13g2_fill_2 FILLER_5_827 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_4 FILLER_5_851 ();
 sg13g2_fill_1 FILLER_5_865 ();
 sg13g2_decap_4 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_882 ();
 sg13g2_decap_4 FILLER_5_889 ();
 sg13g2_fill_2 FILLER_5_903 ();
 sg13g2_fill_1 FILLER_5_905 ();
 sg13g2_fill_2 FILLER_5_917 ();
 sg13g2_decap_4 FILLER_5_935 ();
 sg13g2_fill_1 FILLER_5_939 ();
 sg13g2_fill_1 FILLER_5_1013 ();
 sg13g2_fill_2 FILLER_5_1022 ();
 sg13g2_decap_4 FILLER_5_1074 ();
 sg13g2_fill_1 FILLER_5_1078 ();
 sg13g2_fill_1 FILLER_5_1105 ();
 sg13g2_decap_4 FILLER_5_1136 ();
 sg13g2_decap_8 FILLER_5_1144 ();
 sg13g2_fill_2 FILLER_5_1151 ();
 sg13g2_decap_8 FILLER_5_1156 ();
 sg13g2_decap_8 FILLER_5_1163 ();
 sg13g2_decap_4 FILLER_5_1170 ();
 sg13g2_decap_4 FILLER_5_1179 ();
 sg13g2_fill_1 FILLER_5_1183 ();
 sg13g2_decap_8 FILLER_5_1192 ();
 sg13g2_decap_8 FILLER_5_1199 ();
 sg13g2_decap_8 FILLER_5_1206 ();
 sg13g2_fill_1 FILLER_5_1227 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_decap_8 FILLER_5_1312 ();
 sg13g2_decap_4 FILLER_5_1319 ();
 sg13g2_fill_1 FILLER_5_1333 ();
 sg13g2_decap_8 FILLER_5_1342 ();
 sg13g2_fill_1 FILLER_5_1349 ();
 sg13g2_fill_2 FILLER_5_1354 ();
 sg13g2_fill_1 FILLER_5_1356 ();
 sg13g2_fill_1 FILLER_5_1367 ();
 sg13g2_decap_4 FILLER_5_1372 ();
 sg13g2_fill_1 FILLER_5_1376 ();
 sg13g2_fill_2 FILLER_5_1413 ();
 sg13g2_fill_2 FILLER_5_1486 ();
 sg13g2_fill_1 FILLER_5_1488 ();
 sg13g2_fill_2 FILLER_5_1515 ();
 sg13g2_fill_1 FILLER_5_1517 ();
 sg13g2_fill_2 FILLER_5_1522 ();
 sg13g2_fill_1 FILLER_5_1524 ();
 sg13g2_fill_1 FILLER_5_1535 ();
 sg13g2_fill_1 FILLER_5_1555 ();
 sg13g2_fill_2 FILLER_5_1598 ();
 sg13g2_fill_1 FILLER_5_1600 ();
 sg13g2_decap_8 FILLER_5_1692 ();
 sg13g2_fill_1 FILLER_5_1699 ();
 sg13g2_decap_4 FILLER_5_1736 ();
 sg13g2_decap_8 FILLER_5_1776 ();
 sg13g2_fill_1 FILLER_5_1783 ();
 sg13g2_fill_1 FILLER_5_1819 ();
 sg13g2_fill_1 FILLER_5_1830 ();
 sg13g2_fill_2 FILLER_5_1835 ();
 sg13g2_fill_2 FILLER_5_1867 ();
 sg13g2_fill_1 FILLER_5_1885 ();
 sg13g2_decap_8 FILLER_5_1949 ();
 sg13g2_decap_8 FILLER_5_1956 ();
 sg13g2_decap_8 FILLER_5_1973 ();
 sg13g2_decap_8 FILLER_5_1980 ();
 sg13g2_decap_8 FILLER_5_1987 ();
 sg13g2_decap_8 FILLER_5_1994 ();
 sg13g2_decap_4 FILLER_5_2001 ();
 sg13g2_fill_1 FILLER_5_2005 ();
 sg13g2_decap_8 FILLER_5_2041 ();
 sg13g2_decap_8 FILLER_5_2048 ();
 sg13g2_fill_1 FILLER_5_2055 ();
 sg13g2_decap_8 FILLER_5_2064 ();
 sg13g2_fill_2 FILLER_5_2071 ();
 sg13g2_fill_2 FILLER_5_2094 ();
 sg13g2_fill_1 FILLER_5_2096 ();
 sg13g2_decap_4 FILLER_5_2128 ();
 sg13g2_fill_2 FILLER_5_2136 ();
 sg13g2_fill_1 FILLER_5_2138 ();
 sg13g2_fill_1 FILLER_5_2236 ();
 sg13g2_decap_8 FILLER_5_2254 ();
 sg13g2_decap_8 FILLER_5_2261 ();
 sg13g2_decap_8 FILLER_5_2268 ();
 sg13g2_decap_8 FILLER_5_2275 ();
 sg13g2_decap_8 FILLER_5_2282 ();
 sg13g2_decap_8 FILLER_5_2289 ();
 sg13g2_decap_8 FILLER_5_2296 ();
 sg13g2_decap_8 FILLER_5_2303 ();
 sg13g2_decap_8 FILLER_5_2310 ();
 sg13g2_decap_8 FILLER_5_2317 ();
 sg13g2_decap_8 FILLER_5_2324 ();
 sg13g2_decap_8 FILLER_5_2331 ();
 sg13g2_decap_8 FILLER_5_2338 ();
 sg13g2_decap_8 FILLER_5_2345 ();
 sg13g2_decap_8 FILLER_5_2352 ();
 sg13g2_decap_8 FILLER_5_2359 ();
 sg13g2_decap_8 FILLER_5_2366 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_decap_8 FILLER_5_2387 ();
 sg13g2_decap_8 FILLER_5_2394 ();
 sg13g2_decap_8 FILLER_5_2401 ();
 sg13g2_decap_8 FILLER_5_2408 ();
 sg13g2_decap_8 FILLER_5_2415 ();
 sg13g2_decap_8 FILLER_5_2422 ();
 sg13g2_decap_8 FILLER_5_2429 ();
 sg13g2_decap_8 FILLER_5_2436 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_decap_8 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2478 ();
 sg13g2_decap_8 FILLER_5_2485 ();
 sg13g2_decap_8 FILLER_5_2492 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_decap_8 FILLER_5_2513 ();
 sg13g2_decap_8 FILLER_5_2520 ();
 sg13g2_decap_8 FILLER_5_2527 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2569 ();
 sg13g2_decap_8 FILLER_5_2576 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_8 FILLER_5_2590 ();
 sg13g2_decap_8 FILLER_5_2597 ();
 sg13g2_decap_8 FILLER_5_2604 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_fill_2 FILLER_5_2667 ();
 sg13g2_fill_1 FILLER_5_2669 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_18 ();
 sg13g2_fill_1 FILLER_6_23 ();
 sg13g2_fill_2 FILLER_6_50 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_66 ();
 sg13g2_fill_1 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_decap_4 FILLER_6_156 ();
 sg13g2_fill_1 FILLER_6_203 ();
 sg13g2_fill_1 FILLER_6_213 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_4 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_265 ();
 sg13g2_decap_4 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_4 FILLER_6_298 ();
 sg13g2_decap_4 FILLER_6_332 ();
 sg13g2_decap_4 FILLER_6_341 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_fill_1 FILLER_6_395 ();
 sg13g2_fill_1 FILLER_6_411 ();
 sg13g2_fill_2 FILLER_6_473 ();
 sg13g2_fill_2 FILLER_6_486 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_fill_2 FILLER_6_504 ();
 sg13g2_fill_2 FILLER_6_510 ();
 sg13g2_fill_1 FILLER_6_534 ();
 sg13g2_fill_1 FILLER_6_541 ();
 sg13g2_decap_4 FILLER_6_552 ();
 sg13g2_fill_1 FILLER_6_571 ();
 sg13g2_fill_1 FILLER_6_603 ();
 sg13g2_fill_1 FILLER_6_617 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_fill_1 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_639 ();
 sg13g2_fill_1 FILLER_6_660 ();
 sg13g2_decap_8 FILLER_6_678 ();
 sg13g2_decap_8 FILLER_6_685 ();
 sg13g2_decap_4 FILLER_6_692 ();
 sg13g2_fill_1 FILLER_6_696 ();
 sg13g2_decap_4 FILLER_6_706 ();
 sg13g2_fill_1 FILLER_6_710 ();
 sg13g2_decap_8 FILLER_6_720 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_decap_8 FILLER_6_745 ();
 sg13g2_decap_8 FILLER_6_752 ();
 sg13g2_decap_8 FILLER_6_759 ();
 sg13g2_decap_4 FILLER_6_766 ();
 sg13g2_fill_2 FILLER_6_770 ();
 sg13g2_fill_2 FILLER_6_780 ();
 sg13g2_fill_1 FILLER_6_782 ();
 sg13g2_decap_4 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_813 ();
 sg13g2_fill_2 FILLER_6_820 ();
 sg13g2_decap_4 FILLER_6_848 ();
 sg13g2_fill_2 FILLER_6_856 ();
 sg13g2_decap_4 FILLER_6_889 ();
 sg13g2_fill_1 FILLER_6_893 ();
 sg13g2_fill_1 FILLER_6_920 ();
 sg13g2_fill_1 FILLER_6_931 ();
 sg13g2_fill_1 FILLER_6_958 ();
 sg13g2_fill_1 FILLER_6_999 ();
 sg13g2_fill_1 FILLER_6_1109 ();
 sg13g2_fill_2 FILLER_6_1132 ();
 sg13g2_fill_1 FILLER_6_1160 ();
 sg13g2_decap_4 FILLER_6_1223 ();
 sg13g2_fill_2 FILLER_6_1237 ();
 sg13g2_fill_1 FILLER_6_1239 ();
 sg13g2_fill_2 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_fill_2 FILLER_6_1318 ();
 sg13g2_fill_1 FILLER_6_1320 ();
 sg13g2_fill_1 FILLER_6_1325 ();
 sg13g2_fill_1 FILLER_6_1352 ();
 sg13g2_fill_1 FILLER_6_1357 ();
 sg13g2_fill_2 FILLER_6_1434 ();
 sg13g2_fill_2 FILLER_6_1468 ();
 sg13g2_fill_1 FILLER_6_1470 ();
 sg13g2_decap_4 FILLER_6_1481 ();
 sg13g2_fill_2 FILLER_6_1485 ();
 sg13g2_decap_4 FILLER_6_1491 ();
 sg13g2_fill_2 FILLER_6_1495 ();
 sg13g2_decap_4 FILLER_6_1501 ();
 sg13g2_fill_1 FILLER_6_1505 ();
 sg13g2_decap_8 FILLER_6_1546 ();
 sg13g2_decap_8 FILLER_6_1553 ();
 sg13g2_fill_2 FILLER_6_1560 ();
 sg13g2_fill_1 FILLER_6_1562 ();
 sg13g2_decap_8 FILLER_6_1567 ();
 sg13g2_decap_8 FILLER_6_1574 ();
 sg13g2_decap_4 FILLER_6_1581 ();
 sg13g2_decap_4 FILLER_6_1589 ();
 sg13g2_fill_2 FILLER_6_1593 ();
 sg13g2_fill_2 FILLER_6_1605 ();
 sg13g2_fill_2 FILLER_6_1620 ();
 sg13g2_fill_2 FILLER_6_1643 ();
 sg13g2_fill_1 FILLER_6_1645 ();
 sg13g2_fill_2 FILLER_6_1650 ();
 sg13g2_fill_1 FILLER_6_1652 ();
 sg13g2_decap_8 FILLER_6_1657 ();
 sg13g2_fill_2 FILLER_6_1674 ();
 sg13g2_fill_2 FILLER_6_1702 ();
 sg13g2_fill_1 FILLER_6_1763 ();
 sg13g2_fill_2 FILLER_6_1811 ();
 sg13g2_fill_2 FILLER_6_1878 ();
 sg13g2_fill_1 FILLER_6_1883 ();
 sg13g2_decap_4 FILLER_6_1928 ();
 sg13g2_fill_2 FILLER_6_1932 ();
 sg13g2_fill_1 FILLER_6_1942 ();
 sg13g2_decap_4 FILLER_6_1947 ();
 sg13g2_decap_8 FILLER_6_1961 ();
 sg13g2_fill_1 FILLER_6_1968 ();
 sg13g2_decap_4 FILLER_6_1979 ();
 sg13g2_decap_8 FILLER_6_1993 ();
 sg13g2_decap_4 FILLER_6_2000 ();
 sg13g2_fill_1 FILLER_6_2004 ();
 sg13g2_decap_4 FILLER_6_2031 ();
 sg13g2_decap_4 FILLER_6_2045 ();
 sg13g2_decap_8 FILLER_6_2053 ();
 sg13g2_decap_4 FILLER_6_2060 ();
 sg13g2_fill_1 FILLER_6_2085 ();
 sg13g2_fill_2 FILLER_6_2099 ();
 sg13g2_fill_2 FILLER_6_2106 ();
 sg13g2_decap_8 FILLER_6_2165 ();
 sg13g2_fill_1 FILLER_6_2172 ();
 sg13g2_decap_4 FILLER_6_2177 ();
 sg13g2_fill_1 FILLER_6_2181 ();
 sg13g2_decap_4 FILLER_6_2196 ();
 sg13g2_fill_2 FILLER_6_2204 ();
 sg13g2_fill_1 FILLER_6_2206 ();
 sg13g2_decap_8 FILLER_6_2243 ();
 sg13g2_fill_2 FILLER_6_2291 ();
 sg13g2_fill_1 FILLER_6_2293 ();
 sg13g2_decap_8 FILLER_6_2298 ();
 sg13g2_decap_8 FILLER_6_2305 ();
 sg13g2_decap_8 FILLER_6_2312 ();
 sg13g2_decap_8 FILLER_6_2319 ();
 sg13g2_decap_8 FILLER_6_2326 ();
 sg13g2_decap_8 FILLER_6_2333 ();
 sg13g2_decap_8 FILLER_6_2340 ();
 sg13g2_decap_8 FILLER_6_2347 ();
 sg13g2_decap_8 FILLER_6_2354 ();
 sg13g2_decap_8 FILLER_6_2361 ();
 sg13g2_decap_8 FILLER_6_2368 ();
 sg13g2_decap_8 FILLER_6_2375 ();
 sg13g2_decap_8 FILLER_6_2382 ();
 sg13g2_decap_8 FILLER_6_2389 ();
 sg13g2_decap_8 FILLER_6_2396 ();
 sg13g2_decap_8 FILLER_6_2403 ();
 sg13g2_decap_8 FILLER_6_2410 ();
 sg13g2_decap_8 FILLER_6_2417 ();
 sg13g2_decap_8 FILLER_6_2424 ();
 sg13g2_decap_8 FILLER_6_2431 ();
 sg13g2_decap_8 FILLER_6_2438 ();
 sg13g2_decap_8 FILLER_6_2445 ();
 sg13g2_decap_8 FILLER_6_2452 ();
 sg13g2_decap_8 FILLER_6_2459 ();
 sg13g2_decap_8 FILLER_6_2466 ();
 sg13g2_decap_8 FILLER_6_2473 ();
 sg13g2_decap_8 FILLER_6_2480 ();
 sg13g2_decap_8 FILLER_6_2487 ();
 sg13g2_decap_8 FILLER_6_2494 ();
 sg13g2_decap_8 FILLER_6_2501 ();
 sg13g2_decap_8 FILLER_6_2508 ();
 sg13g2_decap_8 FILLER_6_2515 ();
 sg13g2_decap_8 FILLER_6_2522 ();
 sg13g2_decap_8 FILLER_6_2529 ();
 sg13g2_decap_8 FILLER_6_2536 ();
 sg13g2_decap_8 FILLER_6_2543 ();
 sg13g2_decap_8 FILLER_6_2550 ();
 sg13g2_decap_8 FILLER_6_2557 ();
 sg13g2_decap_8 FILLER_6_2564 ();
 sg13g2_decap_8 FILLER_6_2571 ();
 sg13g2_decap_8 FILLER_6_2578 ();
 sg13g2_decap_8 FILLER_6_2585 ();
 sg13g2_decap_8 FILLER_6_2592 ();
 sg13g2_decap_8 FILLER_6_2599 ();
 sg13g2_decap_8 FILLER_6_2606 ();
 sg13g2_decap_8 FILLER_6_2613 ();
 sg13g2_decap_8 FILLER_6_2620 ();
 sg13g2_decap_8 FILLER_6_2627 ();
 sg13g2_decap_8 FILLER_6_2634 ();
 sg13g2_decap_8 FILLER_6_2641 ();
 sg13g2_decap_8 FILLER_6_2648 ();
 sg13g2_decap_8 FILLER_6_2655 ();
 sg13g2_decap_8 FILLER_6_2662 ();
 sg13g2_fill_1 FILLER_6_2669 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_fill_1 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_59 ();
 sg13g2_fill_2 FILLER_7_80 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_1 FILLER_7_198 ();
 sg13g2_decap_4 FILLER_7_240 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_4 FILLER_7_278 ();
 sg13g2_fill_2 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_7_413 ();
 sg13g2_fill_1 FILLER_7_415 ();
 sg13g2_fill_2 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_430 ();
 sg13g2_fill_1 FILLER_7_432 ();
 sg13g2_fill_1 FILLER_7_468 ();
 sg13g2_decap_8 FILLER_7_505 ();
 sg13g2_decap_8 FILLER_7_512 ();
 sg13g2_decap_4 FILLER_7_523 ();
 sg13g2_decap_8 FILLER_7_557 ();
 sg13g2_fill_2 FILLER_7_564 ();
 sg13g2_fill_1 FILLER_7_566 ();
 sg13g2_fill_1 FILLER_7_581 ();
 sg13g2_fill_2 FILLER_7_598 ();
 sg13g2_decap_8 FILLER_7_606 ();
 sg13g2_fill_2 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_682 ();
 sg13g2_decap_8 FILLER_7_689 ();
 sg13g2_fill_2 FILLER_7_696 ();
 sg13g2_fill_1 FILLER_7_698 ();
 sg13g2_decap_8 FILLER_7_725 ();
 sg13g2_decap_8 FILLER_7_732 ();
 sg13g2_fill_2 FILLER_7_739 ();
 sg13g2_decap_8 FILLER_7_745 ();
 sg13g2_decap_4 FILLER_7_752 ();
 sg13g2_fill_1 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_fill_2 FILLER_7_768 ();
 sg13g2_decap_4 FILLER_7_780 ();
 sg13g2_fill_2 FILLER_7_784 ();
 sg13g2_fill_2 FILLER_7_800 ();
 sg13g2_fill_1 FILLER_7_807 ();
 sg13g2_fill_1 FILLER_7_850 ();
 sg13g2_decap_8 FILLER_7_887 ();
 sg13g2_decap_4 FILLER_7_920 ();
 sg13g2_fill_1 FILLER_7_924 ();
 sg13g2_fill_2 FILLER_7_1004 ();
 sg13g2_fill_1 FILLER_7_1035 ();
 sg13g2_decap_4 FILLER_7_1072 ();
 sg13g2_fill_2 FILLER_7_1076 ();
 sg13g2_fill_1 FILLER_7_1116 ();
 sg13g2_fill_1 FILLER_7_1136 ();
 sg13g2_fill_2 FILLER_7_1167 ();
 sg13g2_decap_4 FILLER_7_1174 ();
 sg13g2_fill_1 FILLER_7_1178 ();
 sg13g2_fill_1 FILLER_7_1189 ();
 sg13g2_decap_8 FILLER_7_1212 ();
 sg13g2_fill_1 FILLER_7_1219 ();
 sg13g2_fill_2 FILLER_7_1246 ();
 sg13g2_fill_1 FILLER_7_1248 ();
 sg13g2_decap_8 FILLER_7_1324 ();
 sg13g2_fill_1 FILLER_7_1331 ();
 sg13g2_decap_8 FILLER_7_1362 ();
 sg13g2_fill_1 FILLER_7_1369 ();
 sg13g2_decap_4 FILLER_7_1406 ();
 sg13g2_fill_1 FILLER_7_1410 ();
 sg13g2_fill_1 FILLER_7_1418 ();
 sg13g2_fill_1 FILLER_7_1432 ();
 sg13g2_fill_1 FILLER_7_1453 ();
 sg13g2_decap_8 FILLER_7_1462 ();
 sg13g2_fill_2 FILLER_7_1469 ();
 sg13g2_decap_4 FILLER_7_1507 ();
 sg13g2_fill_2 FILLER_7_1511 ();
 sg13g2_decap_8 FILLER_7_1523 ();
 sg13g2_decap_8 FILLER_7_1530 ();
 sg13g2_decap_8 FILLER_7_1537 ();
 sg13g2_decap_8 FILLER_7_1544 ();
 sg13g2_decap_8 FILLER_7_1551 ();
 sg13g2_decap_8 FILLER_7_1558 ();
 sg13g2_decap_8 FILLER_7_1565 ();
 sg13g2_fill_1 FILLER_7_1572 ();
 sg13g2_decap_8 FILLER_7_1661 ();
 sg13g2_decap_4 FILLER_7_1668 ();
 sg13g2_fill_2 FILLER_7_1682 ();
 sg13g2_fill_1 FILLER_7_1684 ();
 sg13g2_decap_4 FILLER_7_1689 ();
 sg13g2_fill_1 FILLER_7_1693 ();
 sg13g2_fill_2 FILLER_7_1720 ();
 sg13g2_decap_8 FILLER_7_1726 ();
 sg13g2_fill_2 FILLER_7_1748 ();
 sg13g2_fill_1 FILLER_7_1750 ();
 sg13g2_fill_1 FILLER_7_1788 ();
 sg13g2_fill_1 FILLER_7_1815 ();
 sg13g2_fill_1 FILLER_7_1827 ();
 sg13g2_decap_4 FILLER_7_1847 ();
 sg13g2_fill_1 FILLER_7_1851 ();
 sg13g2_fill_2 FILLER_7_1962 ();
 sg13g2_decap_4 FILLER_7_1974 ();
 sg13g2_decap_8 FILLER_7_2004 ();
 sg13g2_fill_2 FILLER_7_2011 ();
 sg13g2_decap_8 FILLER_7_2017 ();
 sg13g2_fill_2 FILLER_7_2024 ();
 sg13g2_fill_1 FILLER_7_2026 ();
 sg13g2_decap_4 FILLER_7_2068 ();
 sg13g2_fill_2 FILLER_7_2072 ();
 sg13g2_decap_8 FILLER_7_2126 ();
 sg13g2_decap_8 FILLER_7_2137 ();
 sg13g2_fill_2 FILLER_7_2144 ();
 sg13g2_fill_1 FILLER_7_2146 ();
 sg13g2_fill_2 FILLER_7_2151 ();
 sg13g2_decap_8 FILLER_7_2186 ();
 sg13g2_decap_4 FILLER_7_2193 ();
 sg13g2_fill_2 FILLER_7_2197 ();
 sg13g2_decap_8 FILLER_7_2220 ();
 sg13g2_decap_4 FILLER_7_2248 ();
 sg13g2_fill_2 FILLER_7_2252 ();
 sg13g2_decap_8 FILLER_7_2294 ();
 sg13g2_decap_8 FILLER_7_2301 ();
 sg13g2_decap_8 FILLER_7_2308 ();
 sg13g2_decap_8 FILLER_7_2315 ();
 sg13g2_decap_8 FILLER_7_2322 ();
 sg13g2_decap_8 FILLER_7_2329 ();
 sg13g2_decap_8 FILLER_7_2336 ();
 sg13g2_decap_8 FILLER_7_2343 ();
 sg13g2_decap_8 FILLER_7_2350 ();
 sg13g2_decap_8 FILLER_7_2357 ();
 sg13g2_decap_8 FILLER_7_2364 ();
 sg13g2_decap_8 FILLER_7_2371 ();
 sg13g2_decap_8 FILLER_7_2378 ();
 sg13g2_decap_8 FILLER_7_2385 ();
 sg13g2_decap_8 FILLER_7_2392 ();
 sg13g2_decap_8 FILLER_7_2399 ();
 sg13g2_decap_8 FILLER_7_2406 ();
 sg13g2_decap_8 FILLER_7_2413 ();
 sg13g2_decap_8 FILLER_7_2420 ();
 sg13g2_decap_8 FILLER_7_2427 ();
 sg13g2_decap_8 FILLER_7_2434 ();
 sg13g2_decap_8 FILLER_7_2441 ();
 sg13g2_decap_8 FILLER_7_2448 ();
 sg13g2_decap_8 FILLER_7_2455 ();
 sg13g2_decap_8 FILLER_7_2462 ();
 sg13g2_decap_8 FILLER_7_2469 ();
 sg13g2_decap_8 FILLER_7_2476 ();
 sg13g2_decap_8 FILLER_7_2483 ();
 sg13g2_decap_8 FILLER_7_2490 ();
 sg13g2_decap_8 FILLER_7_2497 ();
 sg13g2_decap_8 FILLER_7_2504 ();
 sg13g2_decap_8 FILLER_7_2511 ();
 sg13g2_decap_8 FILLER_7_2518 ();
 sg13g2_decap_8 FILLER_7_2525 ();
 sg13g2_decap_8 FILLER_7_2532 ();
 sg13g2_decap_8 FILLER_7_2539 ();
 sg13g2_decap_8 FILLER_7_2546 ();
 sg13g2_decap_8 FILLER_7_2553 ();
 sg13g2_decap_8 FILLER_7_2560 ();
 sg13g2_decap_8 FILLER_7_2567 ();
 sg13g2_decap_8 FILLER_7_2574 ();
 sg13g2_decap_8 FILLER_7_2581 ();
 sg13g2_decap_8 FILLER_7_2588 ();
 sg13g2_decap_8 FILLER_7_2595 ();
 sg13g2_decap_8 FILLER_7_2602 ();
 sg13g2_decap_8 FILLER_7_2609 ();
 sg13g2_decap_8 FILLER_7_2616 ();
 sg13g2_decap_8 FILLER_7_2623 ();
 sg13g2_decap_8 FILLER_7_2630 ();
 sg13g2_decap_8 FILLER_7_2637 ();
 sg13g2_decap_8 FILLER_7_2644 ();
 sg13g2_decap_8 FILLER_7_2651 ();
 sg13g2_decap_8 FILLER_7_2658 ();
 sg13g2_decap_4 FILLER_7_2665 ();
 sg13g2_fill_1 FILLER_7_2669 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_9 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_decap_4 FILLER_8_40 ();
 sg13g2_fill_2 FILLER_8_44 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_2 FILLER_8_156 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_4 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_2 FILLER_8_343 ();
 sg13g2_decap_4 FILLER_8_381 ();
 sg13g2_fill_1 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_1 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_402 ();
 sg13g2_fill_2 FILLER_8_410 ();
 sg13g2_fill_1 FILLER_8_421 ();
 sg13g2_decap_8 FILLER_8_433 ();
 sg13g2_fill_1 FILLER_8_440 ();
 sg13g2_fill_1 FILLER_8_493 ();
 sg13g2_decap_4 FILLER_8_504 ();
 sg13g2_fill_1 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_513 ();
 sg13g2_fill_2 FILLER_8_520 ();
 sg13g2_decap_4 FILLER_8_532 ();
 sg13g2_decap_4 FILLER_8_545 ();
 sg13g2_fill_1 FILLER_8_549 ();
 sg13g2_decap_4 FILLER_8_560 ();
 sg13g2_fill_1 FILLER_8_564 ();
 sg13g2_decap_4 FILLER_8_617 ();
 sg13g2_fill_1 FILLER_8_621 ();
 sg13g2_fill_1 FILLER_8_626 ();
 sg13g2_fill_1 FILLER_8_647 ();
 sg13g2_decap_4 FILLER_8_730 ();
 sg13g2_fill_1 FILLER_8_734 ();
 sg13g2_fill_1 FILLER_8_796 ();
 sg13g2_fill_2 FILLER_8_883 ();
 sg13g2_fill_1 FILLER_8_885 ();
 sg13g2_fill_2 FILLER_8_896 ();
 sg13g2_decap_4 FILLER_8_906 ();
 sg13g2_fill_2 FILLER_8_910 ();
 sg13g2_fill_1 FILLER_8_960 ();
 sg13g2_fill_2 FILLER_8_991 ();
 sg13g2_fill_1 FILLER_8_996 ();
 sg13g2_fill_1 FILLER_8_1023 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_4 FILLER_8_1068 ();
 sg13g2_decap_8 FILLER_8_1168 ();
 sg13g2_decap_8 FILLER_8_1175 ();
 sg13g2_decap_4 FILLER_8_1182 ();
 sg13g2_fill_2 FILLER_8_1186 ();
 sg13g2_fill_2 FILLER_8_1196 ();
 sg13g2_fill_1 FILLER_8_1198 ();
 sg13g2_fill_1 FILLER_8_1204 ();
 sg13g2_fill_1 FILLER_8_1210 ();
 sg13g2_fill_1 FILLER_8_1218 ();
 sg13g2_fill_2 FILLER_8_1229 ();
 sg13g2_decap_4 FILLER_8_1235 ();
 sg13g2_fill_1 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1244 ();
 sg13g2_fill_2 FILLER_8_1275 ();
 sg13g2_fill_2 FILLER_8_1299 ();
 sg13g2_fill_1 FILLER_8_1301 ();
 sg13g2_decap_8 FILLER_8_1336 ();
 sg13g2_decap_8 FILLER_8_1343 ();
 sg13g2_decap_4 FILLER_8_1368 ();
 sg13g2_fill_2 FILLER_8_1372 ();
 sg13g2_fill_2 FILLER_8_1378 ();
 sg13g2_fill_2 FILLER_8_1385 ();
 sg13g2_decap_8 FILLER_8_1395 ();
 sg13g2_fill_1 FILLER_8_1402 ();
 sg13g2_fill_1 FILLER_8_1414 ();
 sg13g2_fill_2 FILLER_8_1422 ();
 sg13g2_decap_8 FILLER_8_1447 ();
 sg13g2_fill_2 FILLER_8_1454 ();
 sg13g2_fill_2 FILLER_8_1466 ();
 sg13g2_fill_1 FILLER_8_1478 ();
 sg13g2_fill_2 FILLER_8_1505 ();
 sg13g2_fill_2 FILLER_8_1517 ();
 sg13g2_fill_2 FILLER_8_1545 ();
 sg13g2_decap_8 FILLER_8_1583 ();
 sg13g2_decap_8 FILLER_8_1590 ();
 sg13g2_fill_2 FILLER_8_1597 ();
 sg13g2_fill_1 FILLER_8_1610 ();
 sg13g2_fill_2 FILLER_8_1637 ();
 sg13g2_fill_1 FILLER_8_1639 ();
 sg13g2_decap_8 FILLER_8_1644 ();
 sg13g2_fill_2 FILLER_8_1651 ();
 sg13g2_fill_1 FILLER_8_1653 ();
 sg13g2_decap_8 FILLER_8_1694 ();
 sg13g2_fill_1 FILLER_8_1701 ();
 sg13g2_fill_2 FILLER_8_1747 ();
 sg13g2_decap_8 FILLER_8_1834 ();
 sg13g2_decap_8 FILLER_8_1841 ();
 sg13g2_fill_1 FILLER_8_1879 ();
 sg13g2_fill_2 FILLER_8_1947 ();
 sg13g2_fill_1 FILLER_8_1975 ();
 sg13g2_decap_4 FILLER_8_2016 ();
 sg13g2_fill_1 FILLER_8_2020 ();
 sg13g2_fill_1 FILLER_8_2096 ();
 sg13g2_fill_2 FILLER_8_2111 ();
 sg13g2_decap_4 FILLER_8_2211 ();
 sg13g2_decap_4 FILLER_8_2251 ();
 sg13g2_fill_2 FILLER_8_2255 ();
 sg13g2_fill_2 FILLER_8_2267 ();
 sg13g2_decap_8 FILLER_8_2295 ();
 sg13g2_decap_8 FILLER_8_2302 ();
 sg13g2_decap_8 FILLER_8_2309 ();
 sg13g2_decap_8 FILLER_8_2316 ();
 sg13g2_fill_2 FILLER_8_2323 ();
 sg13g2_fill_1 FILLER_8_2325 ();
 sg13g2_decap_4 FILLER_8_2332 ();
 sg13g2_decap_8 FILLER_8_2365 ();
 sg13g2_fill_2 FILLER_8_2372 ();
 sg13g2_fill_1 FILLER_8_2374 ();
 sg13g2_fill_1 FILLER_8_2432 ();
 sg13g2_decap_8 FILLER_8_2459 ();
 sg13g2_decap_8 FILLER_8_2466 ();
 sg13g2_decap_8 FILLER_8_2473 ();
 sg13g2_decap_8 FILLER_8_2480 ();
 sg13g2_decap_8 FILLER_8_2487 ();
 sg13g2_decap_8 FILLER_8_2494 ();
 sg13g2_decap_8 FILLER_8_2501 ();
 sg13g2_decap_8 FILLER_8_2508 ();
 sg13g2_decap_8 FILLER_8_2515 ();
 sg13g2_decap_8 FILLER_8_2522 ();
 sg13g2_decap_8 FILLER_8_2529 ();
 sg13g2_decap_8 FILLER_8_2536 ();
 sg13g2_decap_8 FILLER_8_2543 ();
 sg13g2_decap_8 FILLER_8_2550 ();
 sg13g2_decap_8 FILLER_8_2557 ();
 sg13g2_decap_8 FILLER_8_2564 ();
 sg13g2_decap_8 FILLER_8_2571 ();
 sg13g2_decap_8 FILLER_8_2578 ();
 sg13g2_decap_8 FILLER_8_2585 ();
 sg13g2_decap_8 FILLER_8_2592 ();
 sg13g2_decap_8 FILLER_8_2599 ();
 sg13g2_decap_8 FILLER_8_2606 ();
 sg13g2_decap_8 FILLER_8_2613 ();
 sg13g2_decap_8 FILLER_8_2620 ();
 sg13g2_decap_8 FILLER_8_2627 ();
 sg13g2_decap_8 FILLER_8_2634 ();
 sg13g2_decap_8 FILLER_8_2641 ();
 sg13g2_decap_8 FILLER_8_2648 ();
 sg13g2_decap_8 FILLER_8_2655 ();
 sg13g2_decap_8 FILLER_8_2662 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_2 FILLER_9_73 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_1 FILLER_9_111 ();
 sg13g2_decap_4 FILLER_9_117 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_decap_8 FILLER_9_160 ();
 sg13g2_fill_2 FILLER_9_181 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_fill_2 FILLER_9_217 ();
 sg13g2_decap_4 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_4 FILLER_9_238 ();
 sg13g2_fill_1 FILLER_9_242 ();
 sg13g2_fill_2 FILLER_9_257 ();
 sg13g2_fill_1 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_303 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_353 ();
 sg13g2_decap_4 FILLER_9_380 ();
 sg13g2_fill_2 FILLER_9_384 ();
 sg13g2_fill_1 FILLER_9_453 ();
 sg13g2_fill_2 FILLER_9_459 ();
 sg13g2_fill_1 FILLER_9_465 ();
 sg13g2_fill_1 FILLER_9_502 ();
 sg13g2_decap_4 FILLER_9_559 ();
 sg13g2_fill_1 FILLER_9_563 ();
 sg13g2_fill_2 FILLER_9_581 ();
 sg13g2_fill_2 FILLER_9_602 ();
 sg13g2_fill_1 FILLER_9_604 ();
 sg13g2_fill_1 FILLER_9_621 ();
 sg13g2_fill_1 FILLER_9_626 ();
 sg13g2_fill_1 FILLER_9_662 ();
 sg13g2_fill_2 FILLER_9_697 ();
 sg13g2_fill_1 FILLER_9_699 ();
 sg13g2_fill_2 FILLER_9_705 ();
 sg13g2_fill_2 FILLER_9_711 ();
 sg13g2_decap_4 FILLER_9_739 ();
 sg13g2_fill_2 FILLER_9_743 ();
 sg13g2_fill_2 FILLER_9_778 ();
 sg13g2_fill_2 FILLER_9_806 ();
 sg13g2_decap_8 FILLER_9_857 ();
 sg13g2_fill_2 FILLER_9_864 ();
 sg13g2_decap_8 FILLER_9_871 ();
 sg13g2_decap_8 FILLER_9_878 ();
 sg13g2_decap_8 FILLER_9_885 ();
 sg13g2_decap_8 FILLER_9_892 ();
 sg13g2_decap_4 FILLER_9_899 ();
 sg13g2_fill_2 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_922 ();
 sg13g2_fill_2 FILLER_9_965 ();
 sg13g2_fill_1 FILLER_9_1003 ();
 sg13g2_fill_1 FILLER_9_1008 ();
 sg13g2_fill_1 FILLER_9_1025 ();
 sg13g2_fill_1 FILLER_9_1039 ();
 sg13g2_fill_2 FILLER_9_1046 ();
 sg13g2_fill_2 FILLER_9_1099 ();
 sg13g2_fill_2 FILLER_9_1122 ();
 sg13g2_decap_4 FILLER_9_1164 ();
 sg13g2_fill_1 FILLER_9_1168 ();
 sg13g2_fill_2 FILLER_9_1216 ();
 sg13g2_fill_1 FILLER_9_1236 ();
 sg13g2_decap_8 FILLER_9_1251 ();
 sg13g2_fill_2 FILLER_9_1258 ();
 sg13g2_decap_8 FILLER_9_1272 ();
 sg13g2_decap_8 FILLER_9_1279 ();
 sg13g2_fill_2 FILLER_9_1286 ();
 sg13g2_fill_2 FILLER_9_1310 ();
 sg13g2_fill_1 FILLER_9_1312 ();
 sg13g2_fill_2 FILLER_9_1317 ();
 sg13g2_fill_1 FILLER_9_1319 ();
 sg13g2_fill_2 FILLER_9_1327 ();
 sg13g2_fill_1 FILLER_9_1329 ();
 sg13g2_decap_8 FILLER_9_1343 ();
 sg13g2_decap_4 FILLER_9_1350 ();
 sg13g2_fill_2 FILLER_9_1354 ();
 sg13g2_decap_8 FILLER_9_1388 ();
 sg13g2_decap_8 FILLER_9_1395 ();
 sg13g2_fill_1 FILLER_9_1402 ();
 sg13g2_fill_1 FILLER_9_1406 ();
 sg13g2_fill_1 FILLER_9_1417 ();
 sg13g2_decap_4 FILLER_9_1440 ();
 sg13g2_fill_1 FILLER_9_1444 ();
 sg13g2_fill_2 FILLER_9_1450 ();
 sg13g2_decap_8 FILLER_9_1476 ();
 sg13g2_decap_4 FILLER_9_1483 ();
 sg13g2_fill_1 FILLER_9_1487 ();
 sg13g2_decap_8 FILLER_9_1492 ();
 sg13g2_fill_1 FILLER_9_1499 ();
 sg13g2_fill_1 FILLER_9_1514 ();
 sg13g2_fill_2 FILLER_9_1541 ();
 sg13g2_fill_1 FILLER_9_1547 ();
 sg13g2_fill_2 FILLER_9_1574 ();
 sg13g2_fill_2 FILLER_9_1602 ();
 sg13g2_fill_1 FILLER_9_1617 ();
 sg13g2_fill_1 FILLER_9_1622 ();
 sg13g2_fill_2 FILLER_9_1633 ();
 sg13g2_fill_1 FILLER_9_1635 ();
 sg13g2_fill_1 FILLER_9_1655 ();
 sg13g2_fill_2 FILLER_9_1686 ();
 sg13g2_fill_1 FILLER_9_1688 ();
 sg13g2_fill_2 FILLER_9_1720 ();
 sg13g2_fill_2 FILLER_9_1791 ();
 sg13g2_fill_1 FILLER_9_1925 ();
 sg13g2_fill_2 FILLER_9_1993 ();
 sg13g2_fill_2 FILLER_9_1999 ();
 sg13g2_fill_2 FILLER_9_2027 ();
 sg13g2_fill_1 FILLER_9_2029 ();
 sg13g2_fill_1 FILLER_9_2056 ();
 sg13g2_fill_1 FILLER_9_2061 ();
 sg13g2_fill_1 FILLER_9_2072 ();
 sg13g2_decap_4 FILLER_9_2091 ();
 sg13g2_decap_4 FILLER_9_2131 ();
 sg13g2_fill_2 FILLER_9_2135 ();
 sg13g2_decap_4 FILLER_9_2141 ();
 sg13g2_fill_1 FILLER_9_2145 ();
 sg13g2_fill_2 FILLER_9_2168 ();
 sg13g2_decap_8 FILLER_9_2200 ();
 sg13g2_decap_8 FILLER_9_2207 ();
 sg13g2_fill_1 FILLER_9_2214 ();
 sg13g2_decap_8 FILLER_9_2291 ();
 sg13g2_decap_8 FILLER_9_2298 ();
 sg13g2_decap_8 FILLER_9_2305 ();
 sg13g2_decap_8 FILLER_9_2312 ();
 sg13g2_fill_2 FILLER_9_2323 ();
 sg13g2_fill_1 FILLER_9_2325 ();
 sg13g2_fill_1 FILLER_9_2336 ();
 sg13g2_decap_4 FILLER_9_2392 ();
 sg13g2_fill_1 FILLER_9_2396 ();
 sg13g2_fill_2 FILLER_9_2454 ();
 sg13g2_decap_8 FILLER_9_2482 ();
 sg13g2_decap_8 FILLER_9_2489 ();
 sg13g2_decap_4 FILLER_9_2496 ();
 sg13g2_fill_1 FILLER_9_2500 ();
 sg13g2_fill_1 FILLER_9_2505 ();
 sg13g2_decap_8 FILLER_9_2516 ();
 sg13g2_decap_8 FILLER_9_2523 ();
 sg13g2_decap_8 FILLER_9_2530 ();
 sg13g2_decap_8 FILLER_9_2537 ();
 sg13g2_decap_8 FILLER_9_2544 ();
 sg13g2_decap_8 FILLER_9_2551 ();
 sg13g2_decap_8 FILLER_9_2558 ();
 sg13g2_decap_8 FILLER_9_2565 ();
 sg13g2_decap_8 FILLER_9_2572 ();
 sg13g2_decap_8 FILLER_9_2579 ();
 sg13g2_decap_8 FILLER_9_2586 ();
 sg13g2_decap_8 FILLER_9_2593 ();
 sg13g2_decap_8 FILLER_9_2600 ();
 sg13g2_decap_8 FILLER_9_2607 ();
 sg13g2_decap_8 FILLER_9_2614 ();
 sg13g2_decap_8 FILLER_9_2621 ();
 sg13g2_decap_8 FILLER_9_2628 ();
 sg13g2_decap_8 FILLER_9_2635 ();
 sg13g2_decap_8 FILLER_9_2642 ();
 sg13g2_decap_8 FILLER_9_2649 ();
 sg13g2_decap_8 FILLER_9_2656 ();
 sg13g2_decap_8 FILLER_9_2663 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_41 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_decap_4 FILLER_10_52 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_fill_1 FILLER_10_69 ();
 sg13g2_decap_4 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_decap_4 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_316 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_378 ();
 sg13g2_fill_1 FILLER_10_380 ();
 sg13g2_decap_4 FILLER_10_462 ();
 sg13g2_fill_2 FILLER_10_474 ();
 sg13g2_fill_1 FILLER_10_476 ();
 sg13g2_decap_4 FILLER_10_486 ();
 sg13g2_fill_2 FILLER_10_490 ();
 sg13g2_fill_1 FILLER_10_495 ();
 sg13g2_decap_8 FILLER_10_500 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_decap_4 FILLER_10_518 ();
 sg13g2_fill_1 FILLER_10_531 ();
 sg13g2_fill_2 FILLER_10_536 ();
 sg13g2_fill_2 FILLER_10_544 ();
 sg13g2_decap_4 FILLER_10_551 ();
 sg13g2_fill_1 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_597 ();
 sg13g2_decap_4 FILLER_10_604 ();
 sg13g2_fill_1 FILLER_10_620 ();
 sg13g2_fill_1 FILLER_10_628 ();
 sg13g2_fill_2 FILLER_10_642 ();
 sg13g2_decap_4 FILLER_10_649 ();
 sg13g2_fill_1 FILLER_10_653 ();
 sg13g2_fill_1 FILLER_10_664 ();
 sg13g2_fill_2 FILLER_10_670 ();
 sg13g2_fill_2 FILLER_10_684 ();
 sg13g2_fill_1 FILLER_10_686 ();
 sg13g2_fill_1 FILLER_10_712 ();
 sg13g2_decap_4 FILLER_10_718 ();
 sg13g2_fill_2 FILLER_10_726 ();
 sg13g2_fill_1 FILLER_10_728 ();
 sg13g2_fill_1 FILLER_10_776 ();
 sg13g2_fill_1 FILLER_10_856 ();
 sg13g2_decap_8 FILLER_10_863 ();
 sg13g2_decap_8 FILLER_10_870 ();
 sg13g2_decap_8 FILLER_10_877 ();
 sg13g2_decap_4 FILLER_10_884 ();
 sg13g2_fill_2 FILLER_10_888 ();
 sg13g2_fill_2 FILLER_10_942 ();
 sg13g2_fill_1 FILLER_10_954 ();
 sg13g2_fill_1 FILLER_10_965 ();
 sg13g2_fill_1 FILLER_10_976 ();
 sg13g2_fill_2 FILLER_10_1033 ();
 sg13g2_fill_1 FILLER_10_1049 ();
 sg13g2_fill_2 FILLER_10_1060 ();
 sg13g2_fill_1 FILLER_10_1062 ();
 sg13g2_decap_8 FILLER_10_1073 ();
 sg13g2_decap_8 FILLER_10_1080 ();
 sg13g2_decap_4 FILLER_10_1087 ();
 sg13g2_fill_2 FILLER_10_1117 ();
 sg13g2_decap_8 FILLER_10_1159 ();
 sg13g2_fill_2 FILLER_10_1166 ();
 sg13g2_fill_1 FILLER_10_1199 ();
 sg13g2_fill_1 FILLER_10_1205 ();
 sg13g2_decap_8 FILLER_10_1212 ();
 sg13g2_fill_1 FILLER_10_1223 ();
 sg13g2_fill_1 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1247 ();
 sg13g2_fill_1 FILLER_10_1254 ();
 sg13g2_decap_8 FILLER_10_1260 ();
 sg13g2_decap_4 FILLER_10_1267 ();
 sg13g2_fill_2 FILLER_10_1271 ();
 sg13g2_fill_1 FILLER_10_1306 ();
 sg13g2_decap_8 FILLER_10_1311 ();
 sg13g2_decap_4 FILLER_10_1318 ();
 sg13g2_decap_8 FILLER_10_1346 ();
 sg13g2_fill_2 FILLER_10_1366 ();
 sg13g2_fill_1 FILLER_10_1368 ();
 sg13g2_decap_4 FILLER_10_1387 ();
 sg13g2_fill_1 FILLER_10_1395 ();
 sg13g2_decap_4 FILLER_10_1414 ();
 sg13g2_fill_2 FILLER_10_1418 ();
 sg13g2_fill_2 FILLER_10_1425 ();
 sg13g2_decap_8 FILLER_10_1432 ();
 sg13g2_fill_1 FILLER_10_1439 ();
 sg13g2_fill_1 FILLER_10_1445 ();
 sg13g2_fill_1 FILLER_10_1449 ();
 sg13g2_fill_1 FILLER_10_1466 ();
 sg13g2_decap_4 FILLER_10_1503 ();
 sg13g2_fill_2 FILLER_10_1559 ();
 sg13g2_decap_8 FILLER_10_1601 ();
 sg13g2_decap_8 FILLER_10_1608 ();
 sg13g2_decap_4 FILLER_10_1615 ();
 sg13g2_decap_8 FILLER_10_1623 ();
 sg13g2_decap_8 FILLER_10_1630 ();
 sg13g2_decap_8 FILLER_10_1637 ();
 sg13g2_fill_2 FILLER_10_1644 ();
 sg13g2_decap_8 FILLER_10_1662 ();
 sg13g2_fill_1 FILLER_10_1681 ();
 sg13g2_fill_2 FILLER_10_1708 ();
 sg13g2_fill_1 FILLER_10_1710 ();
 sg13g2_decap_4 FILLER_10_1751 ();
 sg13g2_fill_2 FILLER_10_1755 ();
 sg13g2_fill_2 FILLER_10_1764 ();
 sg13g2_fill_2 FILLER_10_1784 ();
 sg13g2_fill_2 FILLER_10_1835 ();
 sg13g2_decap_4 FILLER_10_1847 ();
 sg13g2_decap_4 FILLER_10_1859 ();
 sg13g2_fill_2 FILLER_10_1863 ();
 sg13g2_decap_4 FILLER_10_1890 ();
 sg13g2_fill_1 FILLER_10_1904 ();
 sg13g2_fill_1 FILLER_10_1908 ();
 sg13g2_decap_8 FILLER_10_1977 ();
 sg13g2_decap_8 FILLER_10_1984 ();
 sg13g2_fill_1 FILLER_10_1991 ();
 sg13g2_decap_8 FILLER_10_2048 ();
 sg13g2_decap_8 FILLER_10_2055 ();
 sg13g2_decap_8 FILLER_10_2062 ();
 sg13g2_decap_8 FILLER_10_2069 ();
 sg13g2_decap_8 FILLER_10_2076 ();
 sg13g2_decap_8 FILLER_10_2083 ();
 sg13g2_decap_8 FILLER_10_2090 ();
 sg13g2_decap_8 FILLER_10_2097 ();
 sg13g2_decap_8 FILLER_10_2104 ();
 sg13g2_decap_4 FILLER_10_2111 ();
 sg13g2_fill_2 FILLER_10_2115 ();
 sg13g2_decap_8 FILLER_10_2143 ();
 sg13g2_fill_2 FILLER_10_2150 ();
 sg13g2_decap_8 FILLER_10_2209 ();
 sg13g2_fill_2 FILLER_10_2216 ();
 sg13g2_fill_1 FILLER_10_2223 ();
 sg13g2_fill_2 FILLER_10_2228 ();
 sg13g2_fill_1 FILLER_10_2230 ();
 sg13g2_decap_8 FILLER_10_2235 ();
 sg13g2_decap_8 FILLER_10_2242 ();
 sg13g2_fill_2 FILLER_10_2249 ();
 sg13g2_fill_1 FILLER_10_2251 ();
 sg13g2_fill_2 FILLER_10_2273 ();
 sg13g2_decap_4 FILLER_10_2279 ();
 sg13g2_fill_2 FILLER_10_2283 ();
 sg13g2_fill_2 FILLER_10_2295 ();
 sg13g2_fill_2 FILLER_10_2347 ();
 sg13g2_fill_1 FILLER_10_2353 ();
 sg13g2_fill_2 FILLER_10_2438 ();
 sg13g2_fill_1 FILLER_10_2471 ();
 sg13g2_decap_8 FILLER_10_2476 ();
 sg13g2_decap_8 FILLER_10_2483 ();
 sg13g2_decap_4 FILLER_10_2490 ();
 sg13g2_fill_1 FILLER_10_2494 ();
 sg13g2_decap_8 FILLER_10_2525 ();
 sg13g2_decap_8 FILLER_10_2532 ();
 sg13g2_fill_2 FILLER_10_2539 ();
 sg13g2_fill_1 FILLER_10_2541 ();
 sg13g2_fill_2 FILLER_10_2546 ();
 sg13g2_fill_1 FILLER_10_2548 ();
 sg13g2_fill_1 FILLER_10_2559 ();
 sg13g2_decap_8 FILLER_10_2586 ();
 sg13g2_decap_4 FILLER_10_2593 ();
 sg13g2_fill_2 FILLER_10_2597 ();
 sg13g2_decap_8 FILLER_10_2603 ();
 sg13g2_fill_1 FILLER_10_2610 ();
 sg13g2_decap_8 FILLER_10_2621 ();
 sg13g2_decap_8 FILLER_10_2628 ();
 sg13g2_decap_8 FILLER_10_2635 ();
 sg13g2_decap_8 FILLER_10_2642 ();
 sg13g2_decap_8 FILLER_10_2649 ();
 sg13g2_decap_8 FILLER_10_2656 ();
 sg13g2_decap_8 FILLER_10_2663 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_107 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_124 ();
 sg13g2_decap_4 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_170 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_decap_4 FILLER_11_192 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_decap_4 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_fill_1 FILLER_11_361 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_2 FILLER_11_397 ();
 sg13g2_fill_1 FILLER_11_460 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_fill_1 FILLER_11_483 ();
 sg13g2_fill_2 FILLER_11_487 ();
 sg13g2_fill_1 FILLER_11_489 ();
 sg13g2_decap_8 FILLER_11_496 ();
 sg13g2_fill_1 FILLER_11_503 ();
 sg13g2_decap_4 FILLER_11_508 ();
 sg13g2_fill_2 FILLER_11_512 ();
 sg13g2_fill_2 FILLER_11_528 ();
 sg13g2_decap_8 FILLER_11_535 ();
 sg13g2_fill_2 FILLER_11_542 ();
 sg13g2_decap_8 FILLER_11_554 ();
 sg13g2_decap_4 FILLER_11_561 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_593 ();
 sg13g2_fill_1 FILLER_11_598 ();
 sg13g2_fill_2 FILLER_11_605 ();
 sg13g2_fill_2 FILLER_11_628 ();
 sg13g2_fill_2 FILLER_11_639 ();
 sg13g2_fill_2 FILLER_11_687 ();
 sg13g2_fill_2 FILLER_11_740 ();
 sg13g2_fill_1 FILLER_11_742 ();
 sg13g2_fill_2 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_fill_1 FILLER_11_830 ();
 sg13g2_fill_2 FILLER_11_871 ();
 sg13g2_fill_1 FILLER_11_909 ();
 sg13g2_fill_2 FILLER_11_944 ();
 sg13g2_fill_1 FILLER_11_946 ();
 sg13g2_fill_2 FILLER_11_957 ();
 sg13g2_fill_1 FILLER_11_959 ();
 sg13g2_fill_2 FILLER_11_966 ();
 sg13g2_fill_2 FILLER_11_1001 ();
 sg13g2_fill_1 FILLER_11_1003 ();
 sg13g2_fill_2 FILLER_11_1040 ();
 sg13g2_fill_1 FILLER_11_1042 ();
 sg13g2_decap_4 FILLER_11_1049 ();
 sg13g2_fill_2 FILLER_11_1053 ();
 sg13g2_decap_8 FILLER_11_1059 ();
 sg13g2_fill_2 FILLER_11_1066 ();
 sg13g2_fill_1 FILLER_11_1068 ();
 sg13g2_fill_1 FILLER_11_1079 ();
 sg13g2_fill_2 FILLER_11_1084 ();
 sg13g2_fill_1 FILLER_11_1086 ();
 sg13g2_decap_4 FILLER_11_1091 ();
 sg13g2_fill_1 FILLER_11_1121 ();
 sg13g2_decap_8 FILLER_11_1148 ();
 sg13g2_decap_8 FILLER_11_1155 ();
 sg13g2_decap_8 FILLER_11_1162 ();
 sg13g2_decap_8 FILLER_11_1169 ();
 sg13g2_fill_2 FILLER_11_1176 ();
 sg13g2_fill_1 FILLER_11_1214 ();
 sg13g2_fill_2 FILLER_11_1220 ();
 sg13g2_decap_8 FILLER_11_1236 ();
 sg13g2_fill_1 FILLER_11_1251 ();
 sg13g2_decap_8 FILLER_11_1300 ();
 sg13g2_decap_8 FILLER_11_1307 ();
 sg13g2_decap_8 FILLER_11_1314 ();
 sg13g2_fill_1 FILLER_11_1321 ();
 sg13g2_decap_4 FILLER_11_1344 ();
 sg13g2_fill_2 FILLER_11_1348 ();
 sg13g2_decap_8 FILLER_11_1354 ();
 sg13g2_fill_1 FILLER_11_1361 ();
 sg13g2_fill_2 FILLER_11_1366 ();
 sg13g2_fill_1 FILLER_11_1368 ();
 sg13g2_decap_4 FILLER_11_1379 ();
 sg13g2_fill_2 FILLER_11_1383 ();
 sg13g2_fill_2 FILLER_11_1389 ();
 sg13g2_fill_1 FILLER_11_1391 ();
 sg13g2_fill_2 FILLER_11_1414 ();
 sg13g2_decap_4 FILLER_11_1424 ();
 sg13g2_fill_1 FILLER_11_1428 ();
 sg13g2_fill_2 FILLER_11_1434 ();
 sg13g2_fill_1 FILLER_11_1436 ();
 sg13g2_fill_2 FILLER_11_1457 ();
 sg13g2_decap_4 FILLER_11_1481 ();
 sg13g2_decap_8 FILLER_11_1489 ();
 sg13g2_decap_8 FILLER_11_1496 ();
 sg13g2_decap_8 FILLER_11_1503 ();
 sg13g2_fill_2 FILLER_11_1510 ();
 sg13g2_fill_1 FILLER_11_1512 ();
 sg13g2_fill_2 FILLER_11_1527 ();
 sg13g2_fill_1 FILLER_11_1539 ();
 sg13g2_fill_1 FILLER_11_1571 ();
 sg13g2_decap_8 FILLER_11_1576 ();
 sg13g2_decap_8 FILLER_11_1583 ();
 sg13g2_decap_4 FILLER_11_1590 ();
 sg13g2_decap_4 FILLER_11_1598 ();
 sg13g2_decap_8 FILLER_11_1652 ();
 sg13g2_decap_4 FILLER_11_1659 ();
 sg13g2_fill_1 FILLER_11_1663 ();
 sg13g2_decap_4 FILLER_11_1668 ();
 sg13g2_decap_4 FILLER_11_1685 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_fill_2 FILLER_11_1764 ();
 sg13g2_decap_8 FILLER_11_1846 ();
 sg13g2_fill_1 FILLER_11_1853 ();
 sg13g2_fill_2 FILLER_11_1858 ();
 sg13g2_fill_1 FILLER_11_1896 ();
 sg13g2_decap_8 FILLER_11_1958 ();
 sg13g2_fill_2 FILLER_11_1965 ();
 sg13g2_decap_8 FILLER_11_1980 ();
 sg13g2_fill_1 FILLER_11_2000 ();
 sg13g2_fill_1 FILLER_11_2036 ();
 sg13g2_fill_1 FILLER_11_2047 ();
 sg13g2_decap_8 FILLER_11_2082 ();
 sg13g2_decap_8 FILLER_11_2089 ();
 sg13g2_fill_1 FILLER_11_2096 ();
 sg13g2_decap_8 FILLER_11_2101 ();
 sg13g2_fill_2 FILLER_11_2108 ();
 sg13g2_decap_4 FILLER_11_2120 ();
 sg13g2_fill_1 FILLER_11_2124 ();
 sg13g2_decap_8 FILLER_11_2129 ();
 sg13g2_fill_1 FILLER_11_2136 ();
 sg13g2_decap_4 FILLER_11_2158 ();
 sg13g2_fill_1 FILLER_11_2162 ();
 sg13g2_decap_8 FILLER_11_2203 ();
 sg13g2_decap_8 FILLER_11_2210 ();
 sg13g2_decap_8 FILLER_11_2217 ();
 sg13g2_fill_1 FILLER_11_2224 ();
 sg13g2_decap_8 FILLER_11_2246 ();
 sg13g2_decap_8 FILLER_11_2253 ();
 sg13g2_decap_8 FILLER_11_2260 ();
 sg13g2_decap_8 FILLER_11_2267 ();
 sg13g2_decap_4 FILLER_11_2274 ();
 sg13g2_decap_8 FILLER_11_2334 ();
 sg13g2_decap_4 FILLER_11_2341 ();
 sg13g2_fill_2 FILLER_11_2345 ();
 sg13g2_decap_8 FILLER_11_2352 ();
 sg13g2_decap_4 FILLER_11_2359 ();
 sg13g2_fill_2 FILLER_11_2363 ();
 sg13g2_fill_2 FILLER_11_2369 ();
 sg13g2_fill_2 FILLER_11_2375 ();
 sg13g2_fill_1 FILLER_11_2377 ();
 sg13g2_decap_8 FILLER_11_2447 ();
 sg13g2_fill_2 FILLER_11_2454 ();
 sg13g2_fill_2 FILLER_11_2482 ();
 sg13g2_fill_2 FILLER_11_2510 ();
 sg13g2_fill_1 FILLER_11_2512 ();
 sg13g2_decap_8 FILLER_11_2539 ();
 sg13g2_decap_8 FILLER_11_2575 ();
 sg13g2_decap_4 FILLER_11_2618 ();
 sg13g2_fill_1 FILLER_11_2622 ();
 sg13g2_decap_8 FILLER_11_2649 ();
 sg13g2_decap_8 FILLER_11_2656 ();
 sg13g2_decap_8 FILLER_11_2663 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_24 ();
 sg13g2_fill_1 FILLER_12_51 ();
 sg13g2_fill_2 FILLER_12_85 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_decap_4 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_4 FILLER_12_308 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_343 ();
 sg13g2_decap_4 FILLER_12_355 ();
 sg13g2_fill_2 FILLER_12_453 ();
 sg13g2_fill_1 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_479 ();
 sg13g2_decap_4 FILLER_12_486 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_fill_1 FILLER_12_497 ();
 sg13g2_fill_2 FILLER_12_524 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_fill_2 FILLER_12_557 ();
 sg13g2_fill_2 FILLER_12_585 ();
 sg13g2_fill_2 FILLER_12_593 ();
 sg13g2_fill_1 FILLER_12_595 ();
 sg13g2_fill_2 FILLER_12_622 ();
 sg13g2_fill_2 FILLER_12_669 ();
 sg13g2_fill_2 FILLER_12_707 ();
 sg13g2_fill_1 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_4 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_4 FILLER_12_742 ();
 sg13g2_fill_2 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_752 ();
 sg13g2_fill_1 FILLER_12_769 ();
 sg13g2_fill_1 FILLER_12_774 ();
 sg13g2_fill_2 FILLER_12_780 ();
 sg13g2_fill_2 FILLER_12_788 ();
 sg13g2_fill_1 FILLER_12_790 ();
 sg13g2_fill_2 FILLER_12_799 ();
 sg13g2_fill_1 FILLER_12_801 ();
 sg13g2_fill_2 FILLER_12_828 ();
 sg13g2_fill_1 FILLER_12_830 ();
 sg13g2_decap_4 FILLER_12_915 ();
 sg13g2_fill_2 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_fill_1 FILLER_12_954 ();
 sg13g2_fill_1 FILLER_12_1084 ();
 sg13g2_decap_8 FILLER_12_1095 ();
 sg13g2_fill_2 FILLER_12_1102 ();
 sg13g2_fill_1 FILLER_12_1104 ();
 sg13g2_decap_8 FILLER_12_1120 ();
 sg13g2_decap_4 FILLER_12_1127 ();
 sg13g2_fill_2 FILLER_12_1131 ();
 sg13g2_fill_1 FILLER_12_1136 ();
 sg13g2_decap_8 FILLER_12_1141 ();
 sg13g2_fill_2 FILLER_12_1148 ();
 sg13g2_fill_1 FILLER_12_1176 ();
 sg13g2_fill_1 FILLER_12_1187 ();
 sg13g2_fill_2 FILLER_12_1194 ();
 sg13g2_fill_1 FILLER_12_1202 ();
 sg13g2_decap_4 FILLER_12_1210 ();
 sg13g2_decap_8 FILLER_12_1220 ();
 sg13g2_decap_8 FILLER_12_1233 ();
 sg13g2_decap_4 FILLER_12_1240 ();
 sg13g2_fill_1 FILLER_12_1244 ();
 sg13g2_decap_8 FILLER_12_1251 ();
 sg13g2_decap_8 FILLER_12_1258 ();
 sg13g2_fill_2 FILLER_12_1265 ();
 sg13g2_fill_1 FILLER_12_1282 ();
 sg13g2_fill_1 FILLER_12_1288 ();
 sg13g2_fill_1 FILLER_12_1294 ();
 sg13g2_fill_1 FILLER_12_1300 ();
 sg13g2_fill_1 FILLER_12_1306 ();
 sg13g2_fill_1 FILLER_12_1310 ();
 sg13g2_fill_1 FILLER_12_1340 ();
 sg13g2_fill_1 FILLER_12_1346 ();
 sg13g2_fill_1 FILLER_12_1357 ();
 sg13g2_decap_4 FILLER_12_1363 ();
 sg13g2_fill_1 FILLER_12_1367 ();
 sg13g2_fill_2 FILLER_12_1393 ();
 sg13g2_decap_4 FILLER_12_1403 ();
 sg13g2_fill_1 FILLER_12_1407 ();
 sg13g2_decap_4 FILLER_12_1431 ();
 sg13g2_fill_1 FILLER_12_1435 ();
 sg13g2_fill_1 FILLER_12_1446 ();
 sg13g2_fill_1 FILLER_12_1452 ();
 sg13g2_decap_8 FILLER_12_1479 ();
 sg13g2_decap_4 FILLER_12_1486 ();
 sg13g2_fill_2 FILLER_12_1490 ();
 sg13g2_decap_8 FILLER_12_1502 ();
 sg13g2_decap_8 FILLER_12_1509 ();
 sg13g2_decap_4 FILLER_12_1516 ();
 sg13g2_fill_2 FILLER_12_1520 ();
 sg13g2_decap_4 FILLER_12_1532 ();
 sg13g2_fill_2 FILLER_12_1536 ();
 sg13g2_fill_1 FILLER_12_1546 ();
 sg13g2_decap_8 FILLER_12_1570 ();
 sg13g2_decap_4 FILLER_12_1577 ();
 sg13g2_fill_1 FILLER_12_1581 ();
 sg13g2_decap_8 FILLER_12_1592 ();
 sg13g2_decap_8 FILLER_12_1599 ();
 sg13g2_decap_4 FILLER_12_1606 ();
 sg13g2_fill_2 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_4 FILLER_12_1666 ();
 sg13g2_fill_1 FILLER_12_1670 ();
 sg13g2_fill_1 FILLER_12_1688 ();
 sg13g2_fill_2 FILLER_12_1703 ();
 sg13g2_fill_1 FILLER_12_1731 ();
 sg13g2_fill_2 FILLER_12_1753 ();
 sg13g2_fill_1 FILLER_12_1765 ();
 sg13g2_fill_1 FILLER_12_1813 ();
 sg13g2_fill_1 FILLER_12_1835 ();
 sg13g2_decap_4 FILLER_12_1846 ();
 sg13g2_fill_1 FILLER_12_1850 ();
 sg13g2_decap_8 FILLER_12_1855 ();
 sg13g2_decap_8 FILLER_12_1862 ();
 sg13g2_decap_4 FILLER_12_1874 ();
 sg13g2_fill_1 FILLER_12_1878 ();
 sg13g2_decap_8 FILLER_12_1883 ();
 sg13g2_fill_1 FILLER_12_1903 ();
 sg13g2_decap_8 FILLER_12_1943 ();
 sg13g2_decap_8 FILLER_12_1950 ();
 sg13g2_decap_4 FILLER_12_1957 ();
 sg13g2_decap_8 FILLER_12_1987 ();
 sg13g2_fill_2 FILLER_12_1994 ();
 sg13g2_fill_2 FILLER_12_2027 ();
 sg13g2_decap_4 FILLER_12_2038 ();
 sg13g2_fill_1 FILLER_12_2042 ();
 sg13g2_fill_2 FILLER_12_2078 ();
 sg13g2_fill_1 FILLER_12_2080 ();
 sg13g2_decap_4 FILLER_12_2125 ();
 sg13g2_decap_8 FILLER_12_2159 ();
 sg13g2_decap_8 FILLER_12_2166 ();
 sg13g2_decap_8 FILLER_12_2173 ();
 sg13g2_decap_8 FILLER_12_2184 ();
 sg13g2_decap_8 FILLER_12_2191 ();
 sg13g2_decap_8 FILLER_12_2198 ();
 sg13g2_decap_8 FILLER_12_2205 ();
 sg13g2_fill_2 FILLER_12_2212 ();
 sg13g2_decap_4 FILLER_12_2264 ();
 sg13g2_fill_1 FILLER_12_2268 ();
 sg13g2_decap_4 FILLER_12_2299 ();
 sg13g2_fill_2 FILLER_12_2303 ();
 sg13g2_decap_4 FILLER_12_2326 ();
 sg13g2_decap_8 FILLER_12_2344 ();
 sg13g2_decap_8 FILLER_12_2351 ();
 sg13g2_decap_8 FILLER_12_2358 ();
 sg13g2_fill_2 FILLER_12_2365 ();
 sg13g2_fill_1 FILLER_12_2367 ();
 sg13g2_fill_1 FILLER_12_2392 ();
 sg13g2_decap_4 FILLER_12_2419 ();
 sg13g2_fill_2 FILLER_12_2423 ();
 sg13g2_decap_8 FILLER_12_2435 ();
 sg13g2_fill_2 FILLER_12_2442 ();
 sg13g2_fill_1 FILLER_12_2454 ();
 sg13g2_decap_8 FILLER_12_2499 ();
 sg13g2_fill_1 FILLER_12_2506 ();
 sg13g2_fill_1 FILLER_12_2537 ();
 sg13g2_fill_1 FILLER_12_2590 ();
 sg13g2_decap_8 FILLER_12_2643 ();
 sg13g2_decap_8 FILLER_12_2650 ();
 sg13g2_decap_8 FILLER_12_2657 ();
 sg13g2_decap_4 FILLER_12_2664 ();
 sg13g2_fill_2 FILLER_12_2668 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_8 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_118 ();
 sg13g2_fill_2 FILLER_13_124 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_333 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_decap_4 FILLER_13_400 ();
 sg13g2_fill_1 FILLER_13_404 ();
 sg13g2_fill_2 FILLER_13_409 ();
 sg13g2_fill_1 FILLER_13_411 ();
 sg13g2_fill_1 FILLER_13_416 ();
 sg13g2_decap_4 FILLER_13_438 ();
 sg13g2_fill_2 FILLER_13_456 ();
 sg13g2_fill_2 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_498 ();
 sg13g2_decap_8 FILLER_13_505 ();
 sg13g2_decap_4 FILLER_13_512 ();
 sg13g2_fill_2 FILLER_13_516 ();
 sg13g2_fill_2 FILLER_13_542 ();
 sg13g2_decap_8 FILLER_13_554 ();
 sg13g2_fill_2 FILLER_13_561 ();
 sg13g2_fill_1 FILLER_13_563 ();
 sg13g2_decap_4 FILLER_13_585 ();
 sg13g2_fill_1 FILLER_13_589 ();
 sg13g2_fill_2 FILLER_13_613 ();
 sg13g2_fill_1 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_655 ();
 sg13g2_fill_1 FILLER_13_667 ();
 sg13g2_decap_4 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_4 FILLER_13_747 ();
 sg13g2_fill_2 FILLER_13_751 ();
 sg13g2_fill_1 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_fill_2 FILLER_13_831 ();
 sg13g2_fill_1 FILLER_13_869 ();
 sg13g2_decap_8 FILLER_13_884 ();
 sg13g2_decap_8 FILLER_13_891 ();
 sg13g2_decap_4 FILLER_13_898 ();
 sg13g2_fill_2 FILLER_13_925 ();
 sg13g2_fill_1 FILLER_13_927 ();
 sg13g2_fill_2 FILLER_13_1046 ();
 sg13g2_decap_8 FILLER_13_1084 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_fill_1 FILLER_13_1098 ();
 sg13g2_fill_2 FILLER_13_1123 ();
 sg13g2_fill_1 FILLER_13_1125 ();
 sg13g2_fill_2 FILLER_13_1130 ();
 sg13g2_fill_1 FILLER_13_1132 ();
 sg13g2_fill_2 FILLER_13_1143 ();
 sg13g2_fill_1 FILLER_13_1145 ();
 sg13g2_decap_8 FILLER_13_1176 ();
 sg13g2_decap_4 FILLER_13_1251 ();
 sg13g2_fill_1 FILLER_13_1255 ();
 sg13g2_fill_2 FILLER_13_1261 ();
 sg13g2_fill_2 FILLER_13_1274 ();
 sg13g2_fill_2 FILLER_13_1282 ();
 sg13g2_fill_1 FILLER_13_1284 ();
 sg13g2_decap_4 FILLER_13_1318 ();
 sg13g2_fill_2 FILLER_13_1322 ();
 sg13g2_fill_2 FILLER_13_1328 ();
 sg13g2_fill_1 FILLER_13_1330 ();
 sg13g2_fill_1 FILLER_13_1336 ();
 sg13g2_decap_4 FILLER_13_1342 ();
 sg13g2_fill_1 FILLER_13_1346 ();
 sg13g2_fill_1 FILLER_13_1351 ();
 sg13g2_fill_2 FILLER_13_1362 ();
 sg13g2_decap_8 FILLER_13_1378 ();
 sg13g2_fill_2 FILLER_13_1416 ();
 sg13g2_fill_2 FILLER_13_1428 ();
 sg13g2_fill_1 FILLER_13_1430 ();
 sg13g2_fill_2 FILLER_13_1444 ();
 sg13g2_fill_2 FILLER_13_1451 ();
 sg13g2_fill_1 FILLER_13_1468 ();
 sg13g2_fill_2 FILLER_13_1527 ();
 sg13g2_fill_2 FILLER_13_1555 ();
 sg13g2_fill_2 FILLER_13_1561 ();
 sg13g2_fill_1 FILLER_13_1563 ();
 sg13g2_fill_2 FILLER_13_1616 ();
 sg13g2_fill_1 FILLER_13_1618 ();
 sg13g2_decap_4 FILLER_13_1666 ();
 sg13g2_decap_8 FILLER_13_1696 ();
 sg13g2_fill_2 FILLER_13_1703 ();
 sg13g2_fill_1 FILLER_13_1705 ();
 sg13g2_fill_1 FILLER_13_1716 ();
 sg13g2_fill_1 FILLER_13_1727 ();
 sg13g2_fill_2 FILLER_13_1732 ();
 sg13g2_decap_8 FILLER_13_1748 ();
 sg13g2_decap_4 FILLER_13_1755 ();
 sg13g2_decap_8 FILLER_13_1788 ();
 sg13g2_decap_4 FILLER_13_1795 ();
 sg13g2_fill_1 FILLER_13_1799 ();
 sg13g2_fill_1 FILLER_13_1833 ();
 sg13g2_decap_4 FILLER_13_1838 ();
 sg13g2_fill_2 FILLER_13_1842 ();
 sg13g2_fill_2 FILLER_13_1870 ();
 sg13g2_fill_1 FILLER_13_1872 ();
 sg13g2_decap_8 FILLER_13_1877 ();
 sg13g2_fill_1 FILLER_13_1884 ();
 sg13g2_decap_8 FILLER_13_1890 ();
 sg13g2_fill_2 FILLER_13_1897 ();
 sg13g2_fill_1 FILLER_13_1899 ();
 sg13g2_decap_8 FILLER_13_1907 ();
 sg13g2_fill_2 FILLER_13_1922 ();
 sg13g2_fill_1 FILLER_13_1924 ();
 sg13g2_decap_4 FILLER_13_1942 ();
 sg13g2_fill_1 FILLER_13_1946 ();
 sg13g2_fill_2 FILLER_13_2007 ();
 sg13g2_decap_8 FILLER_13_2013 ();
 sg13g2_fill_2 FILLER_13_2020 ();
 sg13g2_fill_1 FILLER_13_2022 ();
 sg13g2_fill_2 FILLER_13_2027 ();
 sg13g2_fill_1 FILLER_13_2029 ();
 sg13g2_fill_1 FILLER_13_2091 ();
 sg13g2_decap_8 FILLER_13_2178 ();
 sg13g2_fill_1 FILLER_13_2185 ();
 sg13g2_decap_8 FILLER_13_2190 ();
 sg13g2_decap_8 FILLER_13_2197 ();
 sg13g2_decap_8 FILLER_13_2204 ();
 sg13g2_fill_1 FILLER_13_2278 ();
 sg13g2_decap_8 FILLER_13_2289 ();
 sg13g2_decap_8 FILLER_13_2296 ();
 sg13g2_fill_1 FILLER_13_2307 ();
 sg13g2_decap_8 FILLER_13_2360 ();
 sg13g2_decap_8 FILLER_13_2367 ();
 sg13g2_decap_8 FILLER_13_2374 ();
 sg13g2_decap_8 FILLER_13_2381 ();
 sg13g2_fill_2 FILLER_13_2388 ();
 sg13g2_fill_2 FILLER_13_2400 ();
 sg13g2_decap_8 FILLER_13_2406 ();
 sg13g2_decap_8 FILLER_13_2413 ();
 sg13g2_decap_4 FILLER_13_2420 ();
 sg13g2_fill_1 FILLER_13_2424 ();
 sg13g2_decap_8 FILLER_13_2473 ();
 sg13g2_fill_1 FILLER_13_2480 ();
 sg13g2_decap_8 FILLER_13_2491 ();
 sg13g2_fill_2 FILLER_13_2498 ();
 sg13g2_fill_1 FILLER_13_2500 ();
 sg13g2_decap_8 FILLER_13_2545 ();
 sg13g2_fill_1 FILLER_13_2552 ();
 sg13g2_fill_2 FILLER_13_2557 ();
 sg13g2_fill_1 FILLER_13_2585 ();
 sg13g2_fill_2 FILLER_13_2596 ();
 sg13g2_fill_2 FILLER_13_2602 ();
 sg13g2_fill_2 FILLER_13_2625 ();
 sg13g2_decap_4 FILLER_13_2631 ();
 sg13g2_decap_8 FILLER_13_2639 ();
 sg13g2_decap_8 FILLER_13_2646 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_fill_2 FILLER_13_2667 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_48 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_decap_4 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_113 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_4 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_176 ();
 sg13g2_decap_4 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_4 FILLER_14_242 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_fill_2 FILLER_14_422 ();
 sg13g2_decap_8 FILLER_14_436 ();
 sg13g2_decap_4 FILLER_14_443 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_2 FILLER_14_472 ();
 sg13g2_fill_2 FILLER_14_480 ();
 sg13g2_fill_2 FILLER_14_487 ();
 sg13g2_decap_4 FILLER_14_510 ();
 sg13g2_fill_1 FILLER_14_519 ();
 sg13g2_fill_1 FILLER_14_530 ();
 sg13g2_fill_1 FILLER_14_537 ();
 sg13g2_fill_2 FILLER_14_544 ();
 sg13g2_fill_2 FILLER_14_556 ();
 sg13g2_fill_1 FILLER_14_558 ();
 sg13g2_fill_2 FILLER_14_563 ();
 sg13g2_fill_1 FILLER_14_583 ();
 sg13g2_fill_1 FILLER_14_624 ();
 sg13g2_fill_1 FILLER_14_632 ();
 sg13g2_fill_2 FILLER_14_644 ();
 sg13g2_fill_2 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_685 ();
 sg13g2_fill_2 FILLER_14_691 ();
 sg13g2_fill_2 FILLER_14_712 ();
 sg13g2_fill_2 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_fill_1 FILLER_14_845 ();
 sg13g2_fill_2 FILLER_14_850 ();
 sg13g2_decap_8 FILLER_14_866 ();
 sg13g2_decap_8 FILLER_14_873 ();
 sg13g2_decap_8 FILLER_14_880 ();
 sg13g2_decap_8 FILLER_14_887 ();
 sg13g2_fill_2 FILLER_14_894 ();
 sg13g2_fill_1 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_908 ();
 sg13g2_decap_8 FILLER_14_915 ();
 sg13g2_decap_8 FILLER_14_922 ();
 sg13g2_fill_2 FILLER_14_929 ();
 sg13g2_fill_1 FILLER_14_931 ();
 sg13g2_fill_2 FILLER_14_940 ();
 sg13g2_fill_2 FILLER_14_948 ();
 sg13g2_fill_2 FILLER_14_954 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_decap_8 FILLER_14_967 ();
 sg13g2_fill_1 FILLER_14_984 ();
 sg13g2_fill_1 FILLER_14_988 ();
 sg13g2_fill_2 FILLER_14_1033 ();
 sg13g2_fill_2 FILLER_14_1050 ();
 sg13g2_fill_1 FILLER_14_1052 ();
 sg13g2_fill_1 FILLER_14_1066 ();
 sg13g2_decap_8 FILLER_14_1093 ();
 sg13g2_decap_4 FILLER_14_1100 ();
 sg13g2_fill_2 FILLER_14_1137 ();
 sg13g2_decap_4 FILLER_14_1149 ();
 sg13g2_fill_1 FILLER_14_1157 ();
 sg13g2_decap_4 FILLER_14_1168 ();
 sg13g2_decap_4 FILLER_14_1199 ();
 sg13g2_fill_2 FILLER_14_1209 ();
 sg13g2_fill_2 FILLER_14_1250 ();
 sg13g2_decap_4 FILLER_14_1271 ();
 sg13g2_fill_1 FILLER_14_1275 ();
 sg13g2_fill_2 FILLER_14_1312 ();
 sg13g2_decap_4 FILLER_14_1318 ();
 sg13g2_fill_1 FILLER_14_1322 ();
 sg13g2_fill_1 FILLER_14_1336 ();
 sg13g2_fill_1 FILLER_14_1344 ();
 sg13g2_fill_2 FILLER_14_1350 ();
 sg13g2_fill_1 FILLER_14_1362 ();
 sg13g2_fill_1 FILLER_14_1383 ();
 sg13g2_fill_1 FILLER_14_1396 ();
 sg13g2_fill_1 FILLER_14_1401 ();
 sg13g2_fill_1 FILLER_14_1407 ();
 sg13g2_fill_1 FILLER_14_1420 ();
 sg13g2_decap_4 FILLER_14_1434 ();
 sg13g2_fill_1 FILLER_14_1438 ();
 sg13g2_fill_2 FILLER_14_1479 ();
 sg13g2_fill_1 FILLER_14_1481 ();
 sg13g2_decap_4 FILLER_14_1486 ();
 sg13g2_fill_2 FILLER_14_1490 ();
 sg13g2_decap_4 FILLER_14_1522 ();
 sg13g2_fill_1 FILLER_14_1526 ();
 sg13g2_decap_8 FILLER_14_1563 ();
 sg13g2_fill_2 FILLER_14_1570 ();
 sg13g2_decap_8 FILLER_14_1606 ();
 sg13g2_fill_1 FILLER_14_1613 ();
 sg13g2_decap_4 FILLER_14_1618 ();
 sg13g2_fill_2 FILLER_14_1710 ();
 sg13g2_decap_8 FILLER_14_1716 ();
 sg13g2_fill_2 FILLER_14_1723 ();
 sg13g2_decap_8 FILLER_14_1730 ();
 sg13g2_fill_1 FILLER_14_1737 ();
 sg13g2_decap_8 FILLER_14_1797 ();
 sg13g2_decap_8 FILLER_14_1804 ();
 sg13g2_fill_1 FILLER_14_1811 ();
 sg13g2_fill_1 FILLER_14_1822 ();
 sg13g2_fill_1 FILLER_14_1849 ();
 sg13g2_fill_2 FILLER_14_1886 ();
 sg13g2_fill_2 FILLER_14_1893 ();
 sg13g2_fill_1 FILLER_14_1895 ();
 sg13g2_fill_2 FILLER_14_1909 ();
 sg13g2_fill_2 FILLER_14_1916 ();
 sg13g2_fill_1 FILLER_14_1918 ();
 sg13g2_decap_8 FILLER_14_1949 ();
 sg13g2_fill_1 FILLER_14_1966 ();
 sg13g2_decap_4 FILLER_14_1996 ();
 sg13g2_fill_1 FILLER_14_2000 ();
 sg13g2_decap_4 FILLER_14_2006 ();
 sg13g2_fill_1 FILLER_14_2010 ();
 sg13g2_fill_1 FILLER_14_2019 ();
 sg13g2_fill_2 FILLER_14_2025 ();
 sg13g2_fill_1 FILLER_14_2027 ();
 sg13g2_fill_1 FILLER_14_2037 ();
 sg13g2_fill_2 FILLER_14_2047 ();
 sg13g2_fill_1 FILLER_14_2049 ();
 sg13g2_fill_1 FILLER_14_2063 ();
 sg13g2_fill_2 FILLER_14_2107 ();
 sg13g2_fill_2 FILLER_14_2147 ();
 sg13g2_decap_4 FILLER_14_2205 ();
 sg13g2_decap_8 FILLER_14_2214 ();
 sg13g2_fill_1 FILLER_14_2221 ();
 sg13g2_fill_2 FILLER_14_2273 ();
 sg13g2_fill_1 FILLER_14_2275 ();
 sg13g2_decap_8 FILLER_14_2280 ();
 sg13g2_decap_8 FILLER_14_2287 ();
 sg13g2_decap_4 FILLER_14_2294 ();
 sg13g2_fill_1 FILLER_14_2298 ();
 sg13g2_decap_4 FILLER_14_2351 ();
 sg13g2_fill_2 FILLER_14_2355 ();
 sg13g2_decap_8 FILLER_14_2397 ();
 sg13g2_decap_4 FILLER_14_2404 ();
 sg13g2_fill_1 FILLER_14_2408 ();
 sg13g2_fill_2 FILLER_14_2444 ();
 sg13g2_fill_2 FILLER_14_2458 ();
 sg13g2_decap_8 FILLER_14_2486 ();
 sg13g2_fill_1 FILLER_14_2493 ();
 sg13g2_decap_8 FILLER_14_2514 ();
 sg13g2_decap_4 FILLER_14_2521 ();
 sg13g2_fill_1 FILLER_14_2525 ();
 sg13g2_decap_8 FILLER_14_2572 ();
 sg13g2_decap_4 FILLER_14_2579 ();
 sg13g2_fill_1 FILLER_14_2583 ();
 sg13g2_decap_4 FILLER_14_2611 ();
 sg13g2_fill_2 FILLER_14_2615 ();
 sg13g2_decap_8 FILLER_14_2627 ();
 sg13g2_decap_8 FILLER_14_2634 ();
 sg13g2_decap_8 FILLER_14_2641 ();
 sg13g2_decap_8 FILLER_14_2648 ();
 sg13g2_decap_8 FILLER_14_2655 ();
 sg13g2_decap_8 FILLER_14_2662 ();
 sg13g2_fill_1 FILLER_14_2669 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_125 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_4 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_360 ();
 sg13g2_fill_2 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_decap_4 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_435 ();
 sg13g2_fill_1 FILLER_15_439 ();
 sg13g2_fill_1 FILLER_15_470 ();
 sg13g2_fill_2 FILLER_15_477 ();
 sg13g2_decap_4 FILLER_15_491 ();
 sg13g2_fill_1 FILLER_15_551 ();
 sg13g2_fill_1 FILLER_15_583 ();
 sg13g2_fill_1 FILLER_15_588 ();
 sg13g2_fill_2 FILLER_15_602 ();
 sg13g2_fill_2 FILLER_15_608 ();
 sg13g2_fill_1 FILLER_15_617 ();
 sg13g2_fill_2 FILLER_15_630 ();
 sg13g2_fill_2 FILLER_15_662 ();
 sg13g2_fill_1 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_702 ();
 sg13g2_fill_2 FILLER_15_710 ();
 sg13g2_fill_1 FILLER_15_716 ();
 sg13g2_fill_2 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_fill_2 FILLER_15_773 ();
 sg13g2_fill_1 FILLER_15_775 ();
 sg13g2_fill_1 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_4 FILLER_15_835 ();
 sg13g2_decap_4 FILLER_15_875 ();
 sg13g2_fill_2 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_911 ();
 sg13g2_fill_1 FILLER_15_918 ();
 sg13g2_fill_2 FILLER_15_980 ();
 sg13g2_fill_1 FILLER_15_982 ();
 sg13g2_decap_4 FILLER_15_1000 ();
 sg13g2_fill_2 FILLER_15_1014 ();
 sg13g2_fill_2 FILLER_15_1022 ();
 sg13g2_fill_2 FILLER_15_1029 ();
 sg13g2_decap_4 FILLER_15_1057 ();
 sg13g2_fill_2 FILLER_15_1061 ();
 sg13g2_fill_2 FILLER_15_1067 ();
 sg13g2_fill_1 FILLER_15_1082 ();
 sg13g2_fill_2 FILLER_15_1112 ();
 sg13g2_decap_8 FILLER_15_1150 ();
 sg13g2_decap_8 FILLER_15_1170 ();
 sg13g2_decap_8 FILLER_15_1177 ();
 sg13g2_fill_1 FILLER_15_1207 ();
 sg13g2_fill_2 FILLER_15_1212 ();
 sg13g2_decap_4 FILLER_15_1220 ();
 sg13g2_decap_4 FILLER_15_1234 ();
 sg13g2_decap_8 FILLER_15_1243 ();
 sg13g2_decap_8 FILLER_15_1250 ();
 sg13g2_fill_2 FILLER_15_1257 ();
 sg13g2_fill_2 FILLER_15_1264 ();
 sg13g2_fill_1 FILLER_15_1266 ();
 sg13g2_fill_2 FILLER_15_1288 ();
 sg13g2_fill_1 FILLER_15_1290 ();
 sg13g2_decap_4 FILLER_15_1311 ();
 sg13g2_fill_1 FILLER_15_1315 ();
 sg13g2_decap_4 FILLER_15_1330 ();
 sg13g2_fill_2 FILLER_15_1339 ();
 sg13g2_fill_2 FILLER_15_1346 ();
 sg13g2_fill_1 FILLER_15_1348 ();
 sg13g2_fill_2 FILLER_15_1354 ();
 sg13g2_fill_1 FILLER_15_1356 ();
 sg13g2_fill_2 FILLER_15_1361 ();
 sg13g2_fill_1 FILLER_15_1368 ();
 sg13g2_decap_4 FILLER_15_1374 ();
 sg13g2_fill_2 FILLER_15_1378 ();
 sg13g2_fill_1 FILLER_15_1394 ();
 sg13g2_fill_2 FILLER_15_1401 ();
 sg13g2_decap_8 FILLER_15_1408 ();
 sg13g2_fill_1 FILLER_15_1415 ();
 sg13g2_decap_8 FILLER_15_1442 ();
 sg13g2_decap_8 FILLER_15_1473 ();
 sg13g2_decap_8 FILLER_15_1480 ();
 sg13g2_decap_8 FILLER_15_1487 ();
 sg13g2_fill_2 FILLER_15_1494 ();
 sg13g2_fill_1 FILLER_15_1496 ();
 sg13g2_decap_4 FILLER_15_1514 ();
 sg13g2_fill_1 FILLER_15_1518 ();
 sg13g2_fill_2 FILLER_15_1577 ();
 sg13g2_decap_8 FILLER_15_1610 ();
 sg13g2_decap_8 FILLER_15_1617 ();
 sg13g2_decap_4 FILLER_15_1634 ();
 sg13g2_fill_2 FILLER_15_1638 ();
 sg13g2_decap_8 FILLER_15_1644 ();
 sg13g2_fill_2 FILLER_15_1651 ();
 sg13g2_fill_1 FILLER_15_1653 ();
 sg13g2_fill_1 FILLER_15_1664 ();
 sg13g2_fill_1 FILLER_15_1669 ();
 sg13g2_fill_1 FILLER_15_1694 ();
 sg13g2_decap_8 FILLER_15_1716 ();
 sg13g2_decap_8 FILLER_15_1723 ();
 sg13g2_fill_2 FILLER_15_1730 ();
 sg13g2_decap_8 FILLER_15_1786 ();
 sg13g2_fill_2 FILLER_15_1793 ();
 sg13g2_fill_1 FILLER_15_1805 ();
 sg13g2_decap_8 FILLER_15_1832 ();
 sg13g2_decap_8 FILLER_15_1839 ();
 sg13g2_decap_4 FILLER_15_1846 ();
 sg13g2_decap_4 FILLER_15_1854 ();
 sg13g2_fill_2 FILLER_15_1858 ();
 sg13g2_fill_1 FILLER_15_1894 ();
 sg13g2_fill_1 FILLER_15_1921 ();
 sg13g2_fill_1 FILLER_15_1927 ();
 sg13g2_fill_1 FILLER_15_1937 ();
 sg13g2_fill_2 FILLER_15_1942 ();
 sg13g2_decap_8 FILLER_15_1948 ();
 sg13g2_decap_8 FILLER_15_1955 ();
 sg13g2_decap_4 FILLER_15_1962 ();
 sg13g2_fill_1 FILLER_15_1971 ();
 sg13g2_decap_4 FILLER_15_1976 ();
 sg13g2_fill_2 FILLER_15_1984 ();
 sg13g2_fill_2 FILLER_15_1990 ();
 sg13g2_fill_1 FILLER_15_1992 ();
 sg13g2_fill_1 FILLER_15_2019 ();
 sg13g2_fill_1 FILLER_15_2029 ();
 sg13g2_fill_1 FILLER_15_2083 ();
 sg13g2_fill_1 FILLER_15_2156 ();
 sg13g2_fill_2 FILLER_15_2165 ();
 sg13g2_fill_2 FILLER_15_2177 ();
 sg13g2_fill_2 FILLER_15_2205 ();
 sg13g2_fill_1 FILLER_15_2207 ();
 sg13g2_decap_8 FILLER_15_2212 ();
 sg13g2_decap_8 FILLER_15_2219 ();
 sg13g2_decap_8 FILLER_15_2226 ();
 sg13g2_decap_4 FILLER_15_2233 ();
 sg13g2_decap_8 FILLER_15_2247 ();
 sg13g2_fill_2 FILLER_15_2258 ();
 sg13g2_decap_4 FILLER_15_2264 ();
 sg13g2_fill_2 FILLER_15_2268 ();
 sg13g2_fill_1 FILLER_15_2360 ();
 sg13g2_fill_2 FILLER_15_2387 ();
 sg13g2_fill_2 FILLER_15_2482 ();
 sg13g2_fill_1 FILLER_15_2484 ();
 sg13g2_fill_1 FILLER_15_2506 ();
 sg13g2_fill_2 FILLER_15_2533 ();
 sg13g2_decap_8 FILLER_15_2555 ();
 sg13g2_decap_8 FILLER_15_2562 ();
 sg13g2_decap_8 FILLER_15_2569 ();
 sg13g2_fill_2 FILLER_15_2576 ();
 sg13g2_fill_1 FILLER_15_2578 ();
 sg13g2_decap_8 FILLER_15_2626 ();
 sg13g2_decap_8 FILLER_15_2633 ();
 sg13g2_decap_8 FILLER_15_2640 ();
 sg13g2_decap_8 FILLER_15_2647 ();
 sg13g2_decap_8 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2661 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_4 FILLER_16_133 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_decap_4 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_373 ();
 sg13g2_fill_1 FILLER_16_375 ();
 sg13g2_fill_2 FILLER_16_399 ();
 sg13g2_decap_4 FILLER_16_427 ();
 sg13g2_decap_4 FILLER_16_447 ();
 sg13g2_decap_8 FILLER_16_481 ();
 sg13g2_decap_8 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_495 ();
 sg13g2_fill_2 FILLER_16_502 ();
 sg13g2_fill_1 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_509 ();
 sg13g2_fill_2 FILLER_16_516 ();
 sg13g2_decap_4 FILLER_16_536 ();
 sg13g2_fill_1 FILLER_16_540 ();
 sg13g2_fill_2 FILLER_16_549 ();
 sg13g2_fill_1 FILLER_16_551 ();
 sg13g2_fill_1 FILLER_16_556 ();
 sg13g2_fill_2 FILLER_16_598 ();
 sg13g2_fill_1 FILLER_16_606 ();
 sg13g2_fill_2 FILLER_16_620 ();
 sg13g2_fill_2 FILLER_16_635 ();
 sg13g2_fill_2 FILLER_16_681 ();
 sg13g2_fill_2 FILLER_16_709 ();
 sg13g2_fill_2 FILLER_16_724 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_4 FILLER_16_739 ();
 sg13g2_decap_4 FILLER_16_757 ();
 sg13g2_fill_1 FILLER_16_761 ();
 sg13g2_fill_1 FILLER_16_767 ();
 sg13g2_fill_2 FILLER_16_782 ();
 sg13g2_fill_2 FILLER_16_788 ();
 sg13g2_fill_1 FILLER_16_790 ();
 sg13g2_fill_2 FILLER_16_799 ();
 sg13g2_fill_1 FILLER_16_801 ();
 sg13g2_fill_2 FILLER_16_806 ();
 sg13g2_fill_2 FILLER_16_838 ();
 sg13g2_fill_1 FILLER_16_840 ();
 sg13g2_fill_2 FILLER_16_857 ();
 sg13g2_fill_2 FILLER_16_865 ();
 sg13g2_fill_2 FILLER_16_873 ();
 sg13g2_fill_1 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_fill_1 FILLER_16_917 ();
 sg13g2_fill_1 FILLER_16_952 ();
 sg13g2_fill_2 FILLER_16_957 ();
 sg13g2_fill_2 FILLER_16_989 ();
 sg13g2_fill_1 FILLER_16_991 ();
 sg13g2_decap_8 FILLER_16_1058 ();
 sg13g2_fill_2 FILLER_16_1065 ();
 sg13g2_fill_1 FILLER_16_1077 ();
 sg13g2_fill_2 FILLER_16_1093 ();
 sg13g2_fill_1 FILLER_16_1105 ();
 sg13g2_fill_2 FILLER_16_1120 ();
 sg13g2_fill_2 FILLER_16_1135 ();
 sg13g2_fill_1 FILLER_16_1141 ();
 sg13g2_decap_8 FILLER_16_1168 ();
 sg13g2_decap_8 FILLER_16_1175 ();
 sg13g2_decap_4 FILLER_16_1182 ();
 sg13g2_fill_1 FILLER_16_1200 ();
 sg13g2_fill_1 FILLER_16_1230 ();
 sg13g2_decap_4 FILLER_16_1252 ();
 sg13g2_fill_1 FILLER_16_1256 ();
 sg13g2_decap_8 FILLER_16_1262 ();
 sg13g2_fill_2 FILLER_16_1269 ();
 sg13g2_fill_1 FILLER_16_1271 ();
 sg13g2_decap_4 FILLER_16_1311 ();
 sg13g2_fill_1 FILLER_16_1333 ();
 sg13g2_fill_1 FILLER_16_1344 ();
 sg13g2_fill_1 FILLER_16_1348 ();
 sg13g2_decap_4 FILLER_16_1353 ();
 sg13g2_fill_1 FILLER_16_1357 ();
 sg13g2_decap_4 FILLER_16_1363 ();
 sg13g2_fill_2 FILLER_16_1367 ();
 sg13g2_fill_1 FILLER_16_1382 ();
 sg13g2_fill_2 FILLER_16_1392 ();
 sg13g2_decap_8 FILLER_16_1408 ();
 sg13g2_fill_1 FILLER_16_1420 ();
 sg13g2_decap_4 FILLER_16_1426 ();
 sg13g2_fill_1 FILLER_16_1430 ();
 sg13g2_decap_8 FILLER_16_1435 ();
 sg13g2_fill_2 FILLER_16_1442 ();
 sg13g2_fill_1 FILLER_16_1444 ();
 sg13g2_decap_4 FILLER_16_1471 ();
 sg13g2_fill_2 FILLER_16_1475 ();
 sg13g2_decap_4 FILLER_16_1481 ();
 sg13g2_decap_8 FILLER_16_1489 ();
 sg13g2_decap_8 FILLER_16_1496 ();
 sg13g2_decap_8 FILLER_16_1503 ();
 sg13g2_fill_1 FILLER_16_1510 ();
 sg13g2_fill_1 FILLER_16_1541 ();
 sg13g2_decap_8 FILLER_16_1604 ();
 sg13g2_fill_2 FILLER_16_1611 ();
 sg13g2_decap_8 FILLER_16_1627 ();
 sg13g2_decap_8 FILLER_16_1634 ();
 sg13g2_decap_4 FILLER_16_1641 ();
 sg13g2_fill_2 FILLER_16_1645 ();
 sg13g2_decap_8 FILLER_16_1651 ();
 sg13g2_decap_8 FILLER_16_1658 ();
 sg13g2_decap_8 FILLER_16_1665 ();
 sg13g2_decap_8 FILLER_16_1672 ();
 sg13g2_fill_1 FILLER_16_1679 ();
 sg13g2_decap_8 FILLER_16_1710 ();
 sg13g2_decap_8 FILLER_16_1717 ();
 sg13g2_decap_8 FILLER_16_1724 ();
 sg13g2_decap_8 FILLER_16_1735 ();
 sg13g2_decap_8 FILLER_16_1759 ();
 sg13g2_fill_2 FILLER_16_1766 ();
 sg13g2_decap_8 FILLER_16_1777 ();
 sg13g2_decap_8 FILLER_16_1784 ();
 sg13g2_fill_2 FILLER_16_1791 ();
 sg13g2_fill_1 FILLER_16_1793 ();
 sg13g2_decap_8 FILLER_16_1819 ();
 sg13g2_decap_4 FILLER_16_1826 ();
 sg13g2_fill_1 FILLER_16_1840 ();
 sg13g2_decap_4 FILLER_16_1867 ();
 sg13g2_decap_4 FILLER_16_1915 ();
 sg13g2_fill_2 FILLER_16_1924 ();
 sg13g2_fill_1 FILLER_16_1926 ();
 sg13g2_fill_1 FILLER_16_1932 ();
 sg13g2_decap_4 FILLER_16_1959 ();
 sg13g2_fill_1 FILLER_16_1963 ();
 sg13g2_decap_8 FILLER_16_1982 ();
 sg13g2_fill_2 FILLER_16_1998 ();
 sg13g2_fill_1 FILLER_16_2030 ();
 sg13g2_fill_2 FILLER_16_2057 ();
 sg13g2_fill_1 FILLER_16_2059 ();
 sg13g2_decap_4 FILLER_16_2085 ();
 sg13g2_fill_1 FILLER_16_2089 ();
 sg13g2_fill_2 FILLER_16_2108 ();
 sg13g2_fill_1 FILLER_16_2144 ();
 sg13g2_fill_2 FILLER_16_2161 ();
 sg13g2_fill_1 FILLER_16_2176 ();
 sg13g2_fill_2 FILLER_16_2221 ();
 sg13g2_decap_4 FILLER_16_2233 ();
 sg13g2_fill_2 FILLER_16_2237 ();
 sg13g2_decap_4 FILLER_16_2269 ();
 sg13g2_fill_1 FILLER_16_2273 ();
 sg13g2_fill_2 FILLER_16_2324 ();
 sg13g2_fill_1 FILLER_16_2352 ();
 sg13g2_fill_2 FILLER_16_2437 ();
 sg13g2_fill_1 FILLER_16_2439 ();
 sg13g2_fill_2 FILLER_16_2468 ();
 sg13g2_decap_4 FILLER_16_2511 ();
 sg13g2_fill_1 FILLER_16_2541 ();
 sg13g2_fill_1 FILLER_16_2568 ();
 sg13g2_fill_1 FILLER_16_2590 ();
 sg13g2_fill_1 FILLER_16_2612 ();
 sg13g2_fill_1 FILLER_16_2623 ();
 sg13g2_fill_2 FILLER_16_2628 ();
 sg13g2_decap_8 FILLER_16_2634 ();
 sg13g2_decap_8 FILLER_16_2641 ();
 sg13g2_decap_8 FILLER_16_2648 ();
 sg13g2_decap_8 FILLER_16_2655 ();
 sg13g2_decap_8 FILLER_16_2662 ();
 sg13g2_fill_1 FILLER_16_2669 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_12 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_decap_4 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_270 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_fill_2 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_1 FILLER_17_399 ();
 sg13g2_fill_1 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_decap_8 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_17_436 ();
 sg13g2_fill_1 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_444 ();
 sg13g2_decap_8 FILLER_17_451 ();
 sg13g2_fill_1 FILLER_17_458 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_fill_2 FILLER_17_561 ();
 sg13g2_fill_2 FILLER_17_610 ();
 sg13g2_fill_1 FILLER_17_630 ();
 sg13g2_fill_1 FILLER_17_686 ();
 sg13g2_fill_2 FILLER_17_723 ();
 sg13g2_fill_1 FILLER_17_728 ();
 sg13g2_fill_2 FILLER_17_732 ();
 sg13g2_fill_1 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_fill_2 FILLER_17_808 ();
 sg13g2_fill_1 FILLER_17_823 ();
 sg13g2_fill_2 FILLER_17_844 ();
 sg13g2_fill_1 FILLER_17_846 ();
 sg13g2_fill_1 FILLER_17_851 ();
 sg13g2_fill_1 FILLER_17_855 ();
 sg13g2_fill_2 FILLER_17_991 ();
 sg13g2_decap_4 FILLER_17_997 ();
 sg13g2_decap_4 FILLER_17_1005 ();
 sg13g2_decap_4 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1055 ();
 sg13g2_decap_8 FILLER_17_1062 ();
 sg13g2_decap_4 FILLER_17_1069 ();
 sg13g2_fill_2 FILLER_17_1073 ();
 sg13g2_fill_1 FILLER_17_1089 ();
 sg13g2_decap_4 FILLER_17_1100 ();
 sg13g2_fill_2 FILLER_17_1104 ();
 sg13g2_fill_2 FILLER_17_1110 ();
 sg13g2_fill_1 FILLER_17_1112 ();
 sg13g2_fill_1 FILLER_17_1153 ();
 sg13g2_decap_4 FILLER_17_1190 ();
 sg13g2_fill_2 FILLER_17_1200 ();
 sg13g2_fill_1 FILLER_17_1202 ();
 sg13g2_fill_1 FILLER_17_1240 ();
 sg13g2_fill_1 FILLER_17_1251 ();
 sg13g2_decap_8 FILLER_17_1261 ();
 sg13g2_fill_1 FILLER_17_1268 ();
 sg13g2_fill_1 FILLER_17_1285 ();
 sg13g2_decap_8 FILLER_17_1294 ();
 sg13g2_fill_2 FILLER_17_1301 ();
 sg13g2_fill_2 FILLER_17_1308 ();
 sg13g2_fill_1 FILLER_17_1310 ();
 sg13g2_decap_8 FILLER_17_1317 ();
 sg13g2_decap_4 FILLER_17_1324 ();
 sg13g2_decap_4 FILLER_17_1335 ();
 sg13g2_fill_2 FILLER_17_1339 ();
 sg13g2_decap_4 FILLER_17_1345 ();
 sg13g2_fill_1 FILLER_17_1349 ();
 sg13g2_fill_2 FILLER_17_1376 ();
 sg13g2_fill_1 FILLER_17_1411 ();
 sg13g2_fill_2 FILLER_17_1423 ();
 sg13g2_fill_1 FILLER_17_1425 ();
 sg13g2_fill_1 FILLER_17_1435 ();
 sg13g2_fill_2 FILLER_17_1441 ();
 sg13g2_fill_2 FILLER_17_1448 ();
 sg13g2_fill_2 FILLER_17_1455 ();
 sg13g2_fill_1 FILLER_17_1462 ();
 sg13g2_fill_1 FILLER_17_1540 ();
 sg13g2_fill_2 FILLER_17_1545 ();
 sg13g2_fill_1 FILLER_17_1547 ();
 sg13g2_fill_1 FILLER_17_1552 ();
 sg13g2_fill_2 FILLER_17_1568 ();
 sg13g2_fill_2 FILLER_17_1610 ();
 sg13g2_fill_2 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1674 ();
 sg13g2_decap_4 FILLER_17_1681 ();
 sg13g2_fill_2 FILLER_17_1685 ();
 sg13g2_fill_2 FILLER_17_1697 ();
 sg13g2_decap_4 FILLER_17_1709 ();
 sg13g2_fill_2 FILLER_17_1739 ();
 sg13g2_fill_2 FILLER_17_1762 ();
 sg13g2_fill_1 FILLER_17_1764 ();
 sg13g2_fill_1 FILLER_17_1775 ();
 sg13g2_fill_2 FILLER_17_1780 ();
 sg13g2_decap_4 FILLER_17_1816 ();
 sg13g2_fill_1 FILLER_17_1820 ();
 sg13g2_fill_2 FILLER_17_1825 ();
 sg13g2_fill_1 FILLER_17_1827 ();
 sg13g2_decap_8 FILLER_17_1833 ();
 sg13g2_decap_8 FILLER_17_1844 ();
 sg13g2_decap_8 FILLER_17_1851 ();
 sg13g2_decap_4 FILLER_17_1858 ();
 sg13g2_fill_1 FILLER_17_1862 ();
 sg13g2_fill_1 FILLER_17_1872 ();
 sg13g2_fill_1 FILLER_17_1894 ();
 sg13g2_decap_8 FILLER_17_1907 ();
 sg13g2_decap_8 FILLER_17_1914 ();
 sg13g2_fill_1 FILLER_17_1921 ();
 sg13g2_decap_4 FILLER_17_1956 ();
 sg13g2_fill_1 FILLER_17_1960 ();
 sg13g2_decap_4 FILLER_17_1995 ();
 sg13g2_decap_4 FILLER_17_2009 ();
 sg13g2_fill_2 FILLER_17_2013 ();
 sg13g2_decap_4 FILLER_17_2019 ();
 sg13g2_fill_1 FILLER_17_2023 ();
 sg13g2_fill_2 FILLER_17_2094 ();
 sg13g2_fill_1 FILLER_17_2096 ();
 sg13g2_fill_1 FILLER_17_2120 ();
 sg13g2_fill_2 FILLER_17_2152 ();
 sg13g2_fill_2 FILLER_17_2180 ();
 sg13g2_fill_1 FILLER_17_2182 ();
 sg13g2_fill_1 FILLER_17_2193 ();
 sg13g2_fill_2 FILLER_17_2220 ();
 sg13g2_fill_1 FILLER_17_2222 ();
 sg13g2_decap_4 FILLER_17_2259 ();
 sg13g2_fill_1 FILLER_17_2343 ();
 sg13g2_fill_1 FILLER_17_2348 ();
 sg13g2_fill_1 FILLER_17_2353 ();
 sg13g2_fill_1 FILLER_17_2358 ();
 sg13g2_fill_2 FILLER_17_2369 ();
 sg13g2_fill_1 FILLER_17_2396 ();
 sg13g2_fill_2 FILLER_17_2407 ();
 sg13g2_fill_1 FILLER_17_2409 ();
 sg13g2_fill_2 FILLER_17_2431 ();
 sg13g2_fill_1 FILLER_17_2463 ();
 sg13g2_decap_4 FILLER_17_2497 ();
 sg13g2_fill_1 FILLER_17_2532 ();
 sg13g2_fill_1 FILLER_17_2536 ();
 sg13g2_fill_2 FILLER_17_2543 ();
 sg13g2_decap_8 FILLER_17_2649 ();
 sg13g2_decap_8 FILLER_17_2656 ();
 sg13g2_decap_8 FILLER_17_2663 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_5 ();
 sg13g2_fill_1 FILLER_18_124 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_4 FILLER_18_406 ();
 sg13g2_fill_2 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_430 ();
 sg13g2_fill_2 FILLER_18_437 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_fill_2 FILLER_18_452 ();
 sg13g2_fill_2 FILLER_18_466 ();
 sg13g2_decap_4 FILLER_18_482 ();
 sg13g2_fill_1 FILLER_18_486 ();
 sg13g2_decap_8 FILLER_18_492 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_fill_2 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_4 FILLER_18_529 ();
 sg13g2_fill_1 FILLER_18_544 ();
 sg13g2_decap_4 FILLER_18_551 ();
 sg13g2_fill_1 FILLER_18_555 ();
 sg13g2_fill_2 FILLER_18_586 ();
 sg13g2_fill_1 FILLER_18_713 ();
 sg13g2_fill_2 FILLER_18_719 ();
 sg13g2_fill_2 FILLER_18_802 ();
 sg13g2_fill_2 FILLER_18_814 ();
 sg13g2_fill_1 FILLER_18_836 ();
 sg13g2_fill_2 FILLER_18_867 ();
 sg13g2_decap_8 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_18_884 ();
 sg13g2_fill_1 FILLER_18_919 ();
 sg13g2_fill_1 FILLER_18_951 ();
 sg13g2_fill_1 FILLER_18_1042 ();
 sg13g2_decap_8 FILLER_18_1047 ();
 sg13g2_decap_8 FILLER_18_1054 ();
 sg13g2_decap_8 FILLER_18_1061 ();
 sg13g2_decap_8 FILLER_18_1068 ();
 sg13g2_fill_2 FILLER_18_1075 ();
 sg13g2_fill_1 FILLER_18_1077 ();
 sg13g2_decap_8 FILLER_18_1104 ();
 sg13g2_fill_1 FILLER_18_1111 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_decap_4 FILLER_18_1159 ();
 sg13g2_decap_4 FILLER_18_1172 ();
 sg13g2_fill_1 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1184 ();
 sg13g2_fill_1 FILLER_18_1191 ();
 sg13g2_decap_4 FILLER_18_1207 ();
 sg13g2_fill_2 FILLER_18_1211 ();
 sg13g2_decap_4 FILLER_18_1218 ();
 sg13g2_fill_1 FILLER_18_1222 ();
 sg13g2_fill_1 FILLER_18_1230 ();
 sg13g2_fill_2 FILLER_18_1309 ();
 sg13g2_fill_1 FILLER_18_1311 ();
 sg13g2_fill_1 FILLER_18_1339 ();
 sg13g2_fill_2 FILLER_18_1344 ();
 sg13g2_fill_1 FILLER_18_1361 ();
 sg13g2_fill_1 FILLER_18_1389 ();
 sg13g2_decap_8 FILLER_18_1404 ();
 sg13g2_fill_2 FILLER_18_1411 ();
 sg13g2_fill_1 FILLER_18_1434 ();
 sg13g2_fill_2 FILLER_18_1446 ();
 sg13g2_fill_2 FILLER_18_1469 ();
 sg13g2_decap_4 FILLER_18_1476 ();
 sg13g2_fill_2 FILLER_18_1480 ();
 sg13g2_fill_2 FILLER_18_1528 ();
 sg13g2_fill_1 FILLER_18_1569 ();
 sg13g2_fill_2 FILLER_18_1580 ();
 sg13g2_fill_1 FILLER_18_1608 ();
 sg13g2_fill_2 FILLER_18_1635 ();
 sg13g2_fill_1 FILLER_18_1663 ();
 sg13g2_fill_2 FILLER_18_1690 ();
 sg13g2_fill_1 FILLER_18_1696 ();
 sg13g2_fill_1 FILLER_18_1723 ();
 sg13g2_decap_4 FILLER_18_1750 ();
 sg13g2_fill_2 FILLER_18_1754 ();
 sg13g2_fill_1 FILLER_18_1766 ();
 sg13g2_decap_8 FILLER_18_1793 ();
 sg13g2_fill_1 FILLER_18_1839 ();
 sg13g2_decap_8 FILLER_18_1896 ();
 sg13g2_decap_4 FILLER_18_1903 ();
 sg13g2_decap_4 FILLER_18_1963 ();
 sg13g2_fill_1 FILLER_18_1967 ();
 sg13g2_decap_4 FILLER_18_1972 ();
 sg13g2_fill_1 FILLER_18_1976 ();
 sg13g2_fill_2 FILLER_18_2011 ();
 sg13g2_decap_4 FILLER_18_2034 ();
 sg13g2_fill_2 FILLER_18_2038 ();
 sg13g2_decap_8 FILLER_18_2048 ();
 sg13g2_decap_8 FILLER_18_2055 ();
 sg13g2_fill_1 FILLER_18_2070 ();
 sg13g2_fill_2 FILLER_18_2101 ();
 sg13g2_fill_2 FILLER_18_2124 ();
 sg13g2_fill_1 FILLER_18_2149 ();
 sg13g2_decap_4 FILLER_18_2188 ();
 sg13g2_fill_2 FILLER_18_2192 ();
 sg13g2_decap_4 FILLER_18_2228 ();
 sg13g2_fill_1 FILLER_18_2232 ();
 sg13g2_fill_1 FILLER_18_2259 ();
 sg13g2_fill_2 FILLER_18_2310 ();
 sg13g2_fill_2 FILLER_18_2352 ();
 sg13g2_fill_1 FILLER_18_2370 ();
 sg13g2_fill_2 FILLER_18_2375 ();
 sg13g2_fill_2 FILLER_18_2385 ();
 sg13g2_fill_2 FILLER_18_2395 ();
 sg13g2_fill_1 FILLER_18_2397 ();
 sg13g2_decap_4 FILLER_18_2424 ();
 sg13g2_fill_1 FILLER_18_2428 ();
 sg13g2_fill_2 FILLER_18_2433 ();
 sg13g2_fill_1 FILLER_18_2461 ();
 sg13g2_fill_1 FILLER_18_2466 ();
 sg13g2_fill_1 FILLER_18_2523 ();
 sg13g2_fill_2 FILLER_18_2528 ();
 sg13g2_fill_1 FILLER_18_2536 ();
 sg13g2_fill_1 FILLER_18_2546 ();
 sg13g2_fill_1 FILLER_18_2583 ();
 sg13g2_fill_2 FILLER_18_2611 ();
 sg13g2_decap_8 FILLER_18_2639 ();
 sg13g2_decap_8 FILLER_18_2646 ();
 sg13g2_decap_8 FILLER_18_2653 ();
 sg13g2_decap_8 FILLER_18_2660 ();
 sg13g2_fill_2 FILLER_18_2667 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_61 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_fill_2 FILLER_19_251 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_357 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_421 ();
 sg13g2_fill_1 FILLER_19_458 ();
 sg13g2_fill_2 FILLER_19_472 ();
 sg13g2_fill_2 FILLER_19_479 ();
 sg13g2_fill_2 FILLER_19_487 ();
 sg13g2_fill_2 FILLER_19_525 ();
 sg13g2_fill_1 FILLER_19_579 ();
 sg13g2_fill_1 FILLER_19_606 ();
 sg13g2_fill_1 FILLER_19_611 ();
 sg13g2_fill_2 FILLER_19_638 ();
 sg13g2_fill_1 FILLER_19_654 ();
 sg13g2_fill_2 FILLER_19_796 ();
 sg13g2_fill_2 FILLER_19_830 ();
 sg13g2_fill_1 FILLER_19_841 ();
 sg13g2_fill_1 FILLER_19_846 ();
 sg13g2_decap_4 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_19_881 ();
 sg13g2_fill_1 FILLER_19_905 ();
 sg13g2_decap_4 FILLER_19_925 ();
 sg13g2_decap_4 FILLER_19_943 ();
 sg13g2_fill_1 FILLER_19_960 ();
 sg13g2_fill_2 FILLER_19_972 ();
 sg13g2_fill_1 FILLER_19_974 ();
 sg13g2_fill_1 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1031 ();
 sg13g2_decap_8 FILLER_19_1038 ();
 sg13g2_fill_2 FILLER_19_1045 ();
 sg13g2_fill_1 FILLER_19_1047 ();
 sg13g2_decap_8 FILLER_19_1058 ();
 sg13g2_decap_8 FILLER_19_1065 ();
 sg13g2_decap_8 FILLER_19_1072 ();
 sg13g2_fill_2 FILLER_19_1079 ();
 sg13g2_decap_4 FILLER_19_1108 ();
 sg13g2_fill_1 FILLER_19_1112 ();
 sg13g2_decap_8 FILLER_19_1143 ();
 sg13g2_fill_2 FILLER_19_1150 ();
 sg13g2_fill_1 FILLER_19_1152 ();
 sg13g2_fill_2 FILLER_19_1189 ();
 sg13g2_fill_1 FILLER_19_1201 ();
 sg13g2_fill_2 FILLER_19_1208 ();
 sg13g2_fill_1 FILLER_19_1216 ();
 sg13g2_fill_1 FILLER_19_1227 ();
 sg13g2_fill_2 FILLER_19_1243 ();
 sg13g2_decap_8 FILLER_19_1250 ();
 sg13g2_decap_4 FILLER_19_1257 ();
 sg13g2_fill_2 FILLER_19_1267 ();
 sg13g2_fill_1 FILLER_19_1269 ();
 sg13g2_fill_2 FILLER_19_1280 ();
 sg13g2_fill_1 FILLER_19_1282 ();
 sg13g2_decap_8 FILLER_19_1293 ();
 sg13g2_decap_4 FILLER_19_1300 ();
 sg13g2_fill_2 FILLER_19_1317 ();
 sg13g2_decap_4 FILLER_19_1324 ();
 sg13g2_fill_1 FILLER_19_1333 ();
 sg13g2_decap_8 FILLER_19_1339 ();
 sg13g2_decap_8 FILLER_19_1346 ();
 sg13g2_fill_2 FILLER_19_1357 ();
 sg13g2_fill_2 FILLER_19_1363 ();
 sg13g2_fill_1 FILLER_19_1365 ();
 sg13g2_fill_1 FILLER_19_1375 ();
 sg13g2_fill_2 FILLER_19_1381 ();
 sg13g2_fill_2 FILLER_19_1389 ();
 sg13g2_fill_2 FILLER_19_1404 ();
 sg13g2_fill_1 FILLER_19_1406 ();
 sg13g2_fill_1 FILLER_19_1420 ();
 sg13g2_fill_2 FILLER_19_1440 ();
 sg13g2_fill_1 FILLER_19_1466 ();
 sg13g2_fill_1 FILLER_19_1471 ();
 sg13g2_fill_1 FILLER_19_1479 ();
 sg13g2_fill_1 FILLER_19_1516 ();
 sg13g2_fill_2 FILLER_19_1521 ();
 sg13g2_fill_1 FILLER_19_1533 ();
 sg13g2_fill_2 FILLER_19_1560 ();
 sg13g2_fill_2 FILLER_19_1599 ();
 sg13g2_fill_1 FILLER_19_1607 ();
 sg13g2_decap_4 FILLER_19_1639 ();
 sg13g2_fill_2 FILLER_19_1643 ();
 sg13g2_fill_1 FILLER_19_1649 ();
 sg13g2_fill_1 FILLER_19_1655 ();
 sg13g2_fill_2 FILLER_19_1682 ();
 sg13g2_fill_2 FILLER_19_1688 ();
 sg13g2_fill_1 FILLER_19_1690 ();
 sg13g2_fill_2 FILLER_19_1700 ();
 sg13g2_fill_1 FILLER_19_1702 ();
 sg13g2_fill_1 FILLER_19_1707 ();
 sg13g2_fill_2 FILLER_19_1718 ();
 sg13g2_fill_1 FILLER_19_1720 ();
 sg13g2_decap_4 FILLER_19_1725 ();
 sg13g2_decap_8 FILLER_19_1759 ();
 sg13g2_decap_4 FILLER_19_1792 ();
 sg13g2_fill_2 FILLER_19_1796 ();
 sg13g2_decap_8 FILLER_19_1810 ();
 sg13g2_decap_8 FILLER_19_1817 ();
 sg13g2_fill_2 FILLER_19_1824 ();
 sg13g2_fill_1 FILLER_19_1856 ();
 sg13g2_fill_1 FILLER_19_1862 ();
 sg13g2_fill_1 FILLER_19_1889 ();
 sg13g2_fill_1 FILLER_19_1894 ();
 sg13g2_fill_2 FILLER_19_1939 ();
 sg13g2_fill_2 FILLER_19_1962 ();
 sg13g2_fill_1 FILLER_19_1964 ();
 sg13g2_decap_8 FILLER_19_2004 ();
 sg13g2_decap_8 FILLER_19_2011 ();
 sg13g2_decap_8 FILLER_19_2018 ();
 sg13g2_decap_8 FILLER_19_2025 ();
 sg13g2_decap_8 FILLER_19_2032 ();
 sg13g2_decap_8 FILLER_19_2039 ();
 sg13g2_decap_4 FILLER_19_2046 ();
 sg13g2_fill_2 FILLER_19_2059 ();
 sg13g2_decap_4 FILLER_19_2065 ();
 sg13g2_fill_1 FILLER_19_2069 ();
 sg13g2_fill_1 FILLER_19_2132 ();
 sg13g2_fill_2 FILLER_19_2194 ();
 sg13g2_decap_8 FILLER_19_2217 ();
 sg13g2_fill_1 FILLER_19_2275 ();
 sg13g2_fill_2 FILLER_19_2353 ();
 sg13g2_fill_1 FILLER_19_2387 ();
 sg13g2_fill_1 FILLER_19_2430 ();
 sg13g2_fill_1 FILLER_19_2445 ();
 sg13g2_fill_2 FILLER_19_2503 ();
 sg13g2_decap_8 FILLER_19_2509 ();
 sg13g2_decap_8 FILLER_19_2516 ();
 sg13g2_fill_1 FILLER_19_2523 ();
 sg13g2_fill_1 FILLER_19_2560 ();
 sg13g2_decap_8 FILLER_19_2571 ();
 sg13g2_decap_4 FILLER_19_2578 ();
 sg13g2_fill_1 FILLER_19_2582 ();
 sg13g2_fill_2 FILLER_19_2587 ();
 sg13g2_decap_8 FILLER_19_2594 ();
 sg13g2_fill_2 FILLER_19_2601 ();
 sg13g2_fill_1 FILLER_19_2603 ();
 sg13g2_decap_8 FILLER_19_2614 ();
 sg13g2_decap_8 FILLER_19_2621 ();
 sg13g2_decap_8 FILLER_19_2628 ();
 sg13g2_decap_8 FILLER_19_2635 ();
 sg13g2_decap_8 FILLER_19_2642 ();
 sg13g2_decap_8 FILLER_19_2649 ();
 sg13g2_decap_8 FILLER_19_2656 ();
 sg13g2_decap_8 FILLER_19_2663 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_fill_2 FILLER_20_388 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_457 ();
 sg13g2_fill_1 FILLER_20_467 ();
 sg13g2_fill_1 FILLER_20_473 ();
 sg13g2_fill_2 FILLER_20_478 ();
 sg13g2_fill_2 FILLER_20_490 ();
 sg13g2_fill_1 FILLER_20_492 ();
 sg13g2_fill_2 FILLER_20_505 ();
 sg13g2_fill_1 FILLER_20_507 ();
 sg13g2_fill_2 FILLER_20_512 ();
 sg13g2_fill_1 FILLER_20_514 ();
 sg13g2_fill_2 FILLER_20_525 ();
 sg13g2_fill_1 FILLER_20_527 ();
 sg13g2_fill_1 FILLER_20_559 ();
 sg13g2_fill_1 FILLER_20_586 ();
 sg13g2_fill_1 FILLER_20_601 ();
 sg13g2_fill_1 FILLER_20_608 ();
 sg13g2_fill_1 FILLER_20_629 ();
 sg13g2_fill_1 FILLER_20_634 ();
 sg13g2_fill_2 FILLER_20_639 ();
 sg13g2_fill_1 FILLER_20_649 ();
 sg13g2_fill_2 FILLER_20_673 ();
 sg13g2_fill_1 FILLER_20_685 ();
 sg13g2_fill_2 FILLER_20_716 ();
 sg13g2_fill_2 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_fill_1 FILLER_20_782 ();
 sg13g2_fill_2 FILLER_20_789 ();
 sg13g2_fill_1 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_796 ();
 sg13g2_decap_4 FILLER_20_803 ();
 sg13g2_fill_1 FILLER_20_807 ();
 sg13g2_decap_4 FILLER_20_812 ();
 sg13g2_decap_4 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_4 FILLER_20_841 ();
 sg13g2_fill_1 FILLER_20_845 ();
 sg13g2_fill_2 FILLER_20_863 ();
 sg13g2_fill_1 FILLER_20_865 ();
 sg13g2_decap_4 FILLER_20_870 ();
 sg13g2_fill_2 FILLER_20_914 ();
 sg13g2_fill_2 FILLER_20_958 ();
 sg13g2_fill_1 FILLER_20_960 ();
 sg13g2_fill_1 FILLER_20_990 ();
 sg13g2_fill_2 FILLER_20_1000 ();
 sg13g2_fill_1 FILLER_20_1012 ();
 sg13g2_decap_4 FILLER_20_1017 ();
 sg13g2_fill_2 FILLER_20_1021 ();
 sg13g2_fill_2 FILLER_20_1085 ();
 sg13g2_decap_4 FILLER_20_1117 ();
 sg13g2_decap_4 FILLER_20_1125 ();
 sg13g2_fill_2 FILLER_20_1155 ();
 sg13g2_fill_1 FILLER_20_1165 ();
 sg13g2_fill_1 FILLER_20_1180 ();
 sg13g2_fill_2 FILLER_20_1208 ();
 sg13g2_fill_2 FILLER_20_1228 ();
 sg13g2_fill_1 FILLER_20_1230 ();
 sg13g2_decap_8 FILLER_20_1238 ();
 sg13g2_decap_8 FILLER_20_1258 ();
 sg13g2_decap_4 FILLER_20_1265 ();
 sg13g2_fill_1 FILLER_20_1269 ();
 sg13g2_decap_4 FILLER_20_1275 ();
 sg13g2_fill_1 FILLER_20_1279 ();
 sg13g2_decap_4 FILLER_20_1288 ();
 sg13g2_fill_1 FILLER_20_1292 ();
 sg13g2_decap_4 FILLER_20_1306 ();
 sg13g2_fill_1 FILLER_20_1310 ();
 sg13g2_fill_1 FILLER_20_1321 ();
 sg13g2_fill_1 FILLER_20_1327 ();
 sg13g2_fill_2 FILLER_20_1333 ();
 sg13g2_fill_1 FILLER_20_1378 ();
 sg13g2_fill_1 FILLER_20_1389 ();
 sg13g2_fill_2 FILLER_20_1396 ();
 sg13g2_fill_2 FILLER_20_1403 ();
 sg13g2_fill_1 FILLER_20_1426 ();
 sg13g2_fill_1 FILLER_20_1453 ();
 sg13g2_fill_2 FILLER_20_1467 ();
 sg13g2_fill_1 FILLER_20_1469 ();
 sg13g2_decap_8 FILLER_20_1476 ();
 sg13g2_fill_1 FILLER_20_1483 ();
 sg13g2_decap_4 FILLER_20_1494 ();
 sg13g2_decap_8 FILLER_20_1506 ();
 sg13g2_decap_4 FILLER_20_1513 ();
 sg13g2_fill_2 FILLER_20_1517 ();
 sg13g2_decap_8 FILLER_20_1550 ();
 sg13g2_decap_4 FILLER_20_1591 ();
 sg13g2_fill_2 FILLER_20_1595 ();
 sg13g2_decap_8 FILLER_20_1627 ();
 sg13g2_decap_4 FILLER_20_1634 ();
 sg13g2_fill_1 FILLER_20_1638 ();
 sg13g2_fill_2 FILLER_20_1644 ();
 sg13g2_fill_1 FILLER_20_1659 ();
 sg13g2_fill_2 FILLER_20_1690 ();
 sg13g2_fill_1 FILLER_20_1692 ();
 sg13g2_decap_8 FILLER_20_1698 ();
 sg13g2_decap_4 FILLER_20_1705 ();
 sg13g2_fill_1 FILLER_20_1718 ();
 sg13g2_fill_1 FILLER_20_1723 ();
 sg13g2_decap_4 FILLER_20_1730 ();
 sg13g2_fill_1 FILLER_20_1734 ();
 sg13g2_decap_8 FILLER_20_1745 ();
 sg13g2_decap_8 FILLER_20_1752 ();
 sg13g2_fill_2 FILLER_20_1759 ();
 sg13g2_fill_2 FILLER_20_1831 ();
 sg13g2_fill_1 FILLER_20_1833 ();
 sg13g2_fill_2 FILLER_20_1847 ();
 sg13g2_fill_2 FILLER_20_1863 ();
 sg13g2_fill_1 FILLER_20_1865 ();
 sg13g2_fill_1 FILLER_20_1870 ();
 sg13g2_fill_1 FILLER_20_1875 ();
 sg13g2_fill_1 FILLER_20_1924 ();
 sg13g2_decap_4 FILLER_20_1951 ();
 sg13g2_decap_8 FILLER_20_2013 ();
 sg13g2_decap_8 FILLER_20_2020 ();
 sg13g2_decap_8 FILLER_20_2027 ();
 sg13g2_decap_4 FILLER_20_2034 ();
 sg13g2_fill_2 FILLER_20_2069 ();
 sg13g2_fill_1 FILLER_20_2071 ();
 sg13g2_fill_2 FILLER_20_2082 ();
 sg13g2_fill_1 FILLER_20_2127 ();
 sg13g2_decap_8 FILLER_20_2157 ();
 sg13g2_decap_8 FILLER_20_2168 ();
 sg13g2_decap_4 FILLER_20_2175 ();
 sg13g2_fill_2 FILLER_20_2208 ();
 sg13g2_decap_4 FILLER_20_2214 ();
 sg13g2_fill_2 FILLER_20_2226 ();
 sg13g2_fill_1 FILLER_20_2228 ();
 sg13g2_fill_2 FILLER_20_2244 ();
 sg13g2_fill_1 FILLER_20_2246 ();
 sg13g2_fill_1 FILLER_20_2255 ();
 sg13g2_decap_8 FILLER_20_2260 ();
 sg13g2_decap_4 FILLER_20_2267 ();
 sg13g2_fill_1 FILLER_20_2271 ();
 sg13g2_fill_1 FILLER_20_2301 ();
 sg13g2_fill_1 FILLER_20_2308 ();
 sg13g2_fill_1 FILLER_20_2330 ();
 sg13g2_fill_2 FILLER_20_2378 ();
 sg13g2_decap_4 FILLER_20_2384 ();
 sg13g2_decap_4 FILLER_20_2403 ();
 sg13g2_fill_2 FILLER_20_2417 ();
 sg13g2_fill_1 FILLER_20_2419 ();
 sg13g2_decap_8 FILLER_20_2428 ();
 sg13g2_decap_8 FILLER_20_2435 ();
 sg13g2_decap_8 FILLER_20_2442 ();
 sg13g2_decap_8 FILLER_20_2449 ();
 sg13g2_decap_4 FILLER_20_2456 ();
 sg13g2_fill_1 FILLER_20_2470 ();
 sg13g2_fill_1 FILLER_20_2476 ();
 sg13g2_decap_8 FILLER_20_2481 ();
 sg13g2_decap_8 FILLER_20_2488 ();
 sg13g2_fill_1 FILLER_20_2495 ();
 sg13g2_fill_1 FILLER_20_2505 ();
 sg13g2_decap_8 FILLER_20_2516 ();
 sg13g2_fill_2 FILLER_20_2523 ();
 sg13g2_fill_1 FILLER_20_2536 ();
 sg13g2_fill_1 FILLER_20_2546 ();
 sg13g2_decap_4 FILLER_20_2567 ();
 sg13g2_fill_1 FILLER_20_2571 ();
 sg13g2_decap_8 FILLER_20_2593 ();
 sg13g2_fill_2 FILLER_20_2600 ();
 sg13g2_fill_1 FILLER_20_2602 ();
 sg13g2_decap_8 FILLER_20_2613 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_4 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_111 ();
 sg13g2_fill_1 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_4 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_4 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_decap_4 FILLER_21_382 ();
 sg13g2_fill_2 FILLER_21_386 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_413 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_21_440 ();
 sg13g2_fill_1 FILLER_21_455 ();
 sg13g2_fill_2 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_fill_2 FILLER_21_508 ();
 sg13g2_fill_2 FILLER_21_530 ();
 sg13g2_fill_2 FILLER_21_542 ();
 sg13g2_fill_2 FILLER_21_562 ();
 sg13g2_fill_2 FILLER_21_573 ();
 sg13g2_decap_8 FILLER_21_579 ();
 sg13g2_fill_1 FILLER_21_586 ();
 sg13g2_fill_1 FILLER_21_640 ();
 sg13g2_fill_2 FILLER_21_680 ();
 sg13g2_fill_1 FILLER_21_686 ();
 sg13g2_fill_2 FILLER_21_691 ();
 sg13g2_fill_1 FILLER_21_709 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_fill_1 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_811 ();
 sg13g2_fill_2 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_4 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_fill_2 FILLER_21_869 ();
 sg13g2_fill_1 FILLER_21_907 ();
 sg13g2_fill_2 FILLER_21_952 ();
 sg13g2_fill_2 FILLER_21_979 ();
 sg13g2_fill_1 FILLER_21_990 ();
 sg13g2_fill_2 FILLER_21_1005 ();
 sg13g2_fill_1 FILLER_21_1007 ();
 sg13g2_decap_4 FILLER_21_1018 ();
 sg13g2_fill_2 FILLER_21_1040 ();
 sg13g2_fill_1 FILLER_21_1042 ();
 sg13g2_fill_1 FILLER_21_1072 ();
 sg13g2_fill_2 FILLER_21_1086 ();
 sg13g2_fill_1 FILLER_21_1088 ();
 sg13g2_fill_2 FILLER_21_1093 ();
 sg13g2_fill_1 FILLER_21_1095 ();
 sg13g2_fill_1 FILLER_21_1106 ();
 sg13g2_fill_2 FILLER_21_1133 ();
 sg13g2_fill_1 FILLER_21_1135 ();
 sg13g2_decap_4 FILLER_21_1140 ();
 sg13g2_fill_2 FILLER_21_1144 ();
 sg13g2_fill_2 FILLER_21_1233 ();
 sg13g2_decap_8 FILLER_21_1251 ();
 sg13g2_decap_8 FILLER_21_1258 ();
 sg13g2_decap_8 FILLER_21_1265 ();
 sg13g2_decap_8 FILLER_21_1272 ();
 sg13g2_decap_8 FILLER_21_1279 ();
 sg13g2_fill_2 FILLER_21_1286 ();
 sg13g2_decap_4 FILLER_21_1305 ();
 sg13g2_fill_2 FILLER_21_1320 ();
 sg13g2_fill_1 FILLER_21_1335 ();
 sg13g2_fill_1 FILLER_21_1345 ();
 sg13g2_fill_1 FILLER_21_1355 ();
 sg13g2_fill_2 FILLER_21_1361 ();
 sg13g2_fill_1 FILLER_21_1369 ();
 sg13g2_fill_2 FILLER_21_1373 ();
 sg13g2_fill_1 FILLER_21_1375 ();
 sg13g2_fill_2 FILLER_21_1391 ();
 sg13g2_fill_2 FILLER_21_1398 ();
 sg13g2_fill_1 FILLER_21_1441 ();
 sg13g2_fill_2 FILLER_21_1447 ();
 sg13g2_fill_2 FILLER_21_1479 ();
 sg13g2_fill_1 FILLER_21_1481 ();
 sg13g2_decap_8 FILLER_21_1492 ();
 sg13g2_decap_8 FILLER_21_1499 ();
 sg13g2_decap_8 FILLER_21_1506 ();
 sg13g2_decap_8 FILLER_21_1513 ();
 sg13g2_decap_8 FILLER_21_1520 ();
 sg13g2_fill_2 FILLER_21_1527 ();
 sg13g2_fill_1 FILLER_21_1529 ();
 sg13g2_fill_1 FILLER_21_1605 ();
 sg13g2_decap_8 FILLER_21_1632 ();
 sg13g2_fill_1 FILLER_21_1639 ();
 sg13g2_decap_4 FILLER_21_1650 ();
 sg13g2_fill_1 FILLER_21_1654 ();
 sg13g2_fill_2 FILLER_21_1664 ();
 sg13g2_fill_1 FILLER_21_1666 ();
 sg13g2_fill_2 FILLER_21_1689 ();
 sg13g2_fill_1 FILLER_21_1691 ();
 sg13g2_fill_2 FILLER_21_1743 ();
 sg13g2_fill_1 FILLER_21_1745 ();
 sg13g2_fill_1 FILLER_21_1772 ();
 sg13g2_fill_1 FILLER_21_1777 ();
 sg13g2_fill_1 FILLER_21_1842 ();
 sg13g2_decap_8 FILLER_21_1847 ();
 sg13g2_decap_4 FILLER_21_1854 ();
 sg13g2_fill_1 FILLER_21_1884 ();
 sg13g2_fill_1 FILLER_21_1941 ();
 sg13g2_decap_8 FILLER_21_1956 ();
 sg13g2_fill_2 FILLER_21_1963 ();
 sg13g2_fill_1 FILLER_21_1965 ();
 sg13g2_decap_4 FILLER_21_1970 ();
 sg13g2_decap_8 FILLER_21_1978 ();
 sg13g2_fill_2 FILLER_21_1985 ();
 sg13g2_fill_2 FILLER_21_2091 ();
 sg13g2_fill_1 FILLER_21_2093 ();
 sg13g2_decap_8 FILLER_21_2122 ();
 sg13g2_decap_4 FILLER_21_2129 ();
 sg13g2_fill_1 FILLER_21_2133 ();
 sg13g2_decap_8 FILLER_21_2143 ();
 sg13g2_fill_1 FILLER_21_2150 ();
 sg13g2_fill_1 FILLER_21_2187 ();
 sg13g2_fill_1 FILLER_21_2196 ();
 sg13g2_fill_1 FILLER_21_2201 ();
 sg13g2_fill_2 FILLER_21_2236 ();
 sg13g2_decap_8 FILLER_21_2248 ();
 sg13g2_decap_4 FILLER_21_2255 ();
 sg13g2_fill_2 FILLER_21_2259 ();
 sg13g2_fill_1 FILLER_21_2270 ();
 sg13g2_fill_1 FILLER_21_2318 ();
 sg13g2_fill_1 FILLER_21_2345 ();
 sg13g2_fill_1 FILLER_21_2356 ();
 sg13g2_fill_2 FILLER_21_2361 ();
 sg13g2_decap_8 FILLER_21_2367 ();
 sg13g2_decap_8 FILLER_21_2374 ();
 sg13g2_fill_2 FILLER_21_2381 ();
 sg13g2_fill_1 FILLER_21_2383 ();
 sg13g2_fill_2 FILLER_21_2424 ();
 sg13g2_fill_1 FILLER_21_2426 ();
 sg13g2_decap_8 FILLER_21_2437 ();
 sg13g2_decap_8 FILLER_21_2444 ();
 sg13g2_fill_1 FILLER_21_2451 ();
 sg13g2_decap_4 FILLER_21_2465 ();
 sg13g2_fill_1 FILLER_21_2469 ();
 sg13g2_fill_2 FILLER_21_2499 ();
 sg13g2_fill_1 FILLER_21_2505 ();
 sg13g2_fill_1 FILLER_21_2568 ();
 sg13g2_decap_4 FILLER_21_2579 ();
 sg13g2_fill_1 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2588 ();
 sg13g2_decap_4 FILLER_21_2621 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_decap_4 FILLER_21_2665 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_fill_2 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_decap_8 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_229 ();
 sg13g2_decap_4 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_decap_4 FILLER_22_281 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_4 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_decap_4 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_22_436 ();
 sg13g2_decap_4 FILLER_22_443 ();
 sg13g2_fill_1 FILLER_22_447 ();
 sg13g2_fill_1 FILLER_22_458 ();
 sg13g2_decap_4 FILLER_22_463 ();
 sg13g2_decap_8 FILLER_22_498 ();
 sg13g2_fill_2 FILLER_22_535 ();
 sg13g2_fill_2 FILLER_22_549 ();
 sg13g2_fill_1 FILLER_22_556 ();
 sg13g2_fill_2 FILLER_22_578 ();
 sg13g2_fill_1 FILLER_22_621 ();
 sg13g2_fill_2 FILLER_22_648 ();
 sg13g2_fill_1 FILLER_22_670 ();
 sg13g2_fill_2 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_771 ();
 sg13g2_fill_1 FILLER_22_834 ();
 sg13g2_fill_1 FILLER_22_841 ();
 sg13g2_fill_2 FILLER_22_858 ();
 sg13g2_fill_2 FILLER_22_866 ();
 sg13g2_fill_1 FILLER_22_878 ();
 sg13g2_decap_4 FILLER_22_945 ();
 sg13g2_fill_1 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_960 ();
 sg13g2_decap_8 FILLER_22_967 ();
 sg13g2_fill_2 FILLER_22_978 ();
 sg13g2_fill_2 FILLER_22_1011 ();
 sg13g2_fill_2 FILLER_22_1039 ();
 sg13g2_fill_2 FILLER_22_1064 ();
 sg13g2_fill_1 FILLER_22_1072 ();
 sg13g2_decap_4 FILLER_22_1092 ();
 sg13g2_fill_2 FILLER_22_1096 ();
 sg13g2_fill_2 FILLER_22_1103 ();
 sg13g2_fill_1 FILLER_22_1105 ();
 sg13g2_fill_1 FILLER_22_1168 ();
 sg13g2_decap_8 FILLER_22_1250 ();
 sg13g2_fill_1 FILLER_22_1257 ();
 sg13g2_fill_2 FILLER_22_1264 ();
 sg13g2_fill_1 FILLER_22_1266 ();
 sg13g2_decap_4 FILLER_22_1274 ();
 sg13g2_decap_4 FILLER_22_1283 ();
 sg13g2_fill_1 FILLER_22_1287 ();
 sg13g2_decap_4 FILLER_22_1304 ();
 sg13g2_decap_8 FILLER_22_1316 ();
 sg13g2_fill_1 FILLER_22_1323 ();
 sg13g2_fill_1 FILLER_22_1409 ();
 sg13g2_fill_2 FILLER_22_1439 ();
 sg13g2_fill_2 FILLER_22_1447 ();
 sg13g2_fill_2 FILLER_22_1465 ();
 sg13g2_fill_1 FILLER_22_1472 ();
 sg13g2_fill_2 FILLER_22_1488 ();
 sg13g2_fill_2 FILLER_22_1516 ();
 sg13g2_fill_2 FILLER_22_1522 ();
 sg13g2_decap_8 FILLER_22_1589 ();
 sg13g2_fill_1 FILLER_22_1596 ();
 sg13g2_fill_2 FILLER_22_1601 ();
 sg13g2_fill_1 FILLER_22_1603 ();
 sg13g2_decap_4 FILLER_22_1653 ();
 sg13g2_fill_2 FILLER_22_1739 ();
 sg13g2_decap_8 FILLER_22_1817 ();
 sg13g2_fill_2 FILLER_22_1824 ();
 sg13g2_fill_1 FILLER_22_1826 ();
 sg13g2_decap_8 FILLER_22_1840 ();
 sg13g2_decap_8 FILLER_22_1847 ();
 sg13g2_decap_8 FILLER_22_1854 ();
 sg13g2_decap_8 FILLER_22_1861 ();
 sg13g2_decap_4 FILLER_22_1868 ();
 sg13g2_fill_1 FILLER_22_1881 ();
 sg13g2_decap_4 FILLER_22_1886 ();
 sg13g2_decap_4 FILLER_22_1899 ();
 sg13g2_fill_1 FILLER_22_1903 ();
 sg13g2_fill_2 FILLER_22_1921 ();
 sg13g2_decap_4 FILLER_22_1936 ();
 sg13g2_decap_8 FILLER_22_1944 ();
 sg13g2_decap_8 FILLER_22_1951 ();
 sg13g2_decap_8 FILLER_22_1958 ();
 sg13g2_decap_8 FILLER_22_1965 ();
 sg13g2_fill_1 FILLER_22_2010 ();
 sg13g2_decap_4 FILLER_22_2015 ();
 sg13g2_fill_1 FILLER_22_2019 ();
 sg13g2_decap_8 FILLER_22_2024 ();
 sg13g2_decap_4 FILLER_22_2031 ();
 sg13g2_fill_1 FILLER_22_2035 ();
 sg13g2_fill_1 FILLER_22_2091 ();
 sg13g2_decap_8 FILLER_22_2126 ();
 sg13g2_decap_8 FILLER_22_2133 ();
 sg13g2_decap_8 FILLER_22_2140 ();
 sg13g2_fill_2 FILLER_22_2147 ();
 sg13g2_decap_4 FILLER_22_2225 ();
 sg13g2_fill_2 FILLER_22_2229 ();
 sg13g2_fill_1 FILLER_22_2270 ();
 sg13g2_fill_1 FILLER_22_2274 ();
 sg13g2_fill_2 FILLER_22_2303 ();
 sg13g2_fill_2 FILLER_22_2324 ();
 sg13g2_decap_8 FILLER_22_2347 ();
 sg13g2_decap_8 FILLER_22_2354 ();
 sg13g2_fill_2 FILLER_22_2361 ();
 sg13g2_fill_1 FILLER_22_2363 ();
 sg13g2_decap_4 FILLER_22_2374 ();
 sg13g2_decap_8 FILLER_22_2388 ();
 sg13g2_fill_2 FILLER_22_2395 ();
 sg13g2_fill_1 FILLER_22_2397 ();
 sg13g2_fill_2 FILLER_22_2402 ();
 sg13g2_fill_2 FILLER_22_2430 ();
 sg13g2_fill_1 FILLER_22_2432 ();
 sg13g2_fill_2 FILLER_22_2459 ();
 sg13g2_fill_1 FILLER_22_2461 ();
 sg13g2_fill_1 FILLER_22_2490 ();
 sg13g2_fill_2 FILLER_22_2547 ();
 sg13g2_decap_8 FILLER_22_2661 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_decap_4 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_248 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_23_422 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_fill_1 FILLER_23_441 ();
 sg13g2_fill_1 FILLER_23_448 ();
 sg13g2_fill_1 FILLER_23_525 ();
 sg13g2_fill_2 FILLER_23_540 ();
 sg13g2_decap_8 FILLER_23_562 ();
 sg13g2_fill_2 FILLER_23_569 ();
 sg13g2_fill_1 FILLER_23_571 ();
 sg13g2_fill_2 FILLER_23_581 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_fill_2 FILLER_23_602 ();
 sg13g2_fill_1 FILLER_23_604 ();
 sg13g2_fill_1 FILLER_23_630 ();
 sg13g2_fill_2 FILLER_23_648 ();
 sg13g2_fill_2 FILLER_23_796 ();
 sg13g2_fill_1 FILLER_23_798 ();
 sg13g2_fill_1 FILLER_23_887 ();
 sg13g2_fill_1 FILLER_23_910 ();
 sg13g2_fill_1 FILLER_23_923 ();
 sg13g2_fill_1 FILLER_23_939 ();
 sg13g2_decap_8 FILLER_23_979 ();
 sg13g2_fill_1 FILLER_23_986 ();
 sg13g2_decap_4 FILLER_23_992 ();
 sg13g2_fill_2 FILLER_23_996 ();
 sg13g2_decap_8 FILLER_23_1002 ();
 sg13g2_decap_8 FILLER_23_1009 ();
 sg13g2_decap_8 FILLER_23_1016 ();
 sg13g2_decap_8 FILLER_23_1023 ();
 sg13g2_decap_8 FILLER_23_1030 ();
 sg13g2_decap_8 FILLER_23_1037 ();
 sg13g2_decap_4 FILLER_23_1044 ();
 sg13g2_fill_2 FILLER_23_1061 ();
 sg13g2_fill_1 FILLER_23_1087 ();
 sg13g2_fill_2 FILLER_23_1101 ();
 sg13g2_fill_1 FILLER_23_1103 ();
 sg13g2_decap_8 FILLER_23_1118 ();
 sg13g2_fill_1 FILLER_23_1125 ();
 sg13g2_decap_4 FILLER_23_1156 ();
 sg13g2_fill_2 FILLER_23_1160 ();
 sg13g2_fill_2 FILLER_23_1183 ();
 sg13g2_fill_1 FILLER_23_1231 ();
 sg13g2_fill_2 FILLER_23_1237 ();
 sg13g2_fill_2 FILLER_23_1250 ();
 sg13g2_decap_8 FILLER_23_1257 ();
 sg13g2_fill_2 FILLER_23_1264 ();
 sg13g2_fill_1 FILLER_23_1266 ();
 sg13g2_decap_8 FILLER_23_1284 ();
 sg13g2_decap_4 FILLER_23_1296 ();
 sg13g2_fill_1 FILLER_23_1305 ();
 sg13g2_fill_2 FILLER_23_1310 ();
 sg13g2_fill_1 FILLER_23_1312 ();
 sg13g2_fill_2 FILLER_23_1319 ();
 sg13g2_fill_1 FILLER_23_1326 ();
 sg13g2_fill_2 FILLER_23_1336 ();
 sg13g2_fill_1 FILLER_23_1343 ();
 sg13g2_fill_1 FILLER_23_1361 ();
 sg13g2_fill_1 FILLER_23_1367 ();
 sg13g2_fill_2 FILLER_23_1373 ();
 sg13g2_fill_1 FILLER_23_1391 ();
 sg13g2_fill_1 FILLER_23_1396 ();
 sg13g2_fill_1 FILLER_23_1410 ();
 sg13g2_fill_2 FILLER_23_1424 ();
 sg13g2_fill_2 FILLER_23_1441 ();
 sg13g2_fill_2 FILLER_23_1471 ();
 sg13g2_fill_1 FILLER_23_1483 ();
 sg13g2_fill_2 FILLER_23_1494 ();
 sg13g2_fill_1 FILLER_23_1496 ();
 sg13g2_decap_4 FILLER_23_1501 ();
 sg13g2_fill_1 FILLER_23_1515 ();
 sg13g2_fill_2 FILLER_23_1542 ();
 sg13g2_fill_1 FILLER_23_1577 ();
 sg13g2_fill_2 FILLER_23_1609 ();
 sg13g2_fill_1 FILLER_23_1611 ();
 sg13g2_fill_2 FILLER_23_1630 ();
 sg13g2_fill_1 FILLER_23_1666 ();
 sg13g2_fill_1 FILLER_23_1688 ();
 sg13g2_fill_2 FILLER_23_1727 ();
 sg13g2_fill_1 FILLER_23_1755 ();
 sg13g2_decap_8 FILLER_23_1825 ();
 sg13g2_fill_1 FILLER_23_1832 ();
 sg13g2_fill_1 FILLER_23_1863 ();
 sg13g2_fill_1 FILLER_23_1885 ();
 sg13g2_decap_8 FILLER_23_1892 ();
 sg13g2_decap_8 FILLER_23_1911 ();
 sg13g2_decap_8 FILLER_23_1918 ();
 sg13g2_fill_1 FILLER_23_1925 ();
 sg13g2_decap_8 FILLER_23_1934 ();
 sg13g2_decap_4 FILLER_23_1941 ();
 sg13g2_fill_2 FILLER_23_1945 ();
 sg13g2_fill_1 FILLER_23_1990 ();
 sg13g2_fill_1 FILLER_23_1999 ();
 sg13g2_decap_8 FILLER_23_2007 ();
 sg13g2_decap_4 FILLER_23_2014 ();
 sg13g2_fill_2 FILLER_23_2018 ();
 sg13g2_decap_8 FILLER_23_2028 ();
 sg13g2_fill_2 FILLER_23_2035 ();
 sg13g2_fill_2 FILLER_23_2042 ();
 sg13g2_fill_2 FILLER_23_2052 ();
 sg13g2_fill_1 FILLER_23_2054 ();
 sg13g2_fill_2 FILLER_23_2091 ();
 sg13g2_fill_1 FILLER_23_2093 ();
 sg13g2_fill_2 FILLER_23_2098 ();
 sg13g2_fill_1 FILLER_23_2100 ();
 sg13g2_fill_2 FILLER_23_2127 ();
 sg13g2_fill_2 FILLER_23_2155 ();
 sg13g2_fill_1 FILLER_23_2161 ();
 sg13g2_fill_1 FILLER_23_2170 ();
 sg13g2_decap_4 FILLER_23_2192 ();
 sg13g2_fill_1 FILLER_23_2196 ();
 sg13g2_decap_8 FILLER_23_2233 ();
 sg13g2_fill_1 FILLER_23_2240 ();
 sg13g2_fill_2 FILLER_23_2276 ();
 sg13g2_fill_1 FILLER_23_2304 ();
 sg13g2_decap_8 FILLER_23_2367 ();
 sg13g2_fill_2 FILLER_23_2400 ();
 sg13g2_fill_2 FILLER_23_2412 ();
 sg13g2_fill_1 FILLER_23_2414 ();
 sg13g2_fill_1 FILLER_23_2425 ();
 sg13g2_fill_2 FILLER_23_2430 ();
 sg13g2_fill_1 FILLER_23_2432 ();
 sg13g2_decap_4 FILLER_23_2570 ();
 sg13g2_fill_1 FILLER_23_2574 ();
 sg13g2_fill_2 FILLER_23_2601 ();
 sg13g2_fill_2 FILLER_23_2607 ();
 sg13g2_fill_2 FILLER_23_2619 ();
 sg13g2_fill_2 FILLER_23_2631 ();
 sg13g2_fill_1 FILLER_23_2633 ();
 sg13g2_fill_1 FILLER_23_2648 ();
 sg13g2_decap_8 FILLER_23_2653 ();
 sg13g2_decap_8 FILLER_23_2660 ();
 sg13g2_fill_2 FILLER_23_2667 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_37 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_decap_4 FILLER_24_222 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_decap_4 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_446 ();
 sg13g2_fill_2 FILLER_24_450 ();
 sg13g2_fill_2 FILLER_24_455 ();
 sg13g2_fill_1 FILLER_24_457 ();
 sg13g2_decap_8 FILLER_24_461 ();
 sg13g2_decap_4 FILLER_24_468 ();
 sg13g2_fill_2 FILLER_24_472 ();
 sg13g2_decap_4 FILLER_24_482 ();
 sg13g2_fill_1 FILLER_24_486 ();
 sg13g2_decap_8 FILLER_24_491 ();
 sg13g2_fill_2 FILLER_24_498 ();
 sg13g2_fill_1 FILLER_24_536 ();
 sg13g2_fill_1 FILLER_24_563 ();
 sg13g2_fill_1 FILLER_24_570 ();
 sg13g2_fill_1 FILLER_24_625 ();
 sg13g2_fill_1 FILLER_24_689 ();
 sg13g2_fill_1 FILLER_24_737 ();
 sg13g2_fill_1 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_775 ();
 sg13g2_decap_4 FILLER_24_780 ();
 sg13g2_fill_2 FILLER_24_784 ();
 sg13g2_fill_2 FILLER_24_796 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_fill_1 FILLER_24_841 ();
 sg13g2_fill_2 FILLER_24_880 ();
 sg13g2_fill_2 FILLER_24_906 ();
 sg13g2_fill_1 FILLER_24_950 ();
 sg13g2_fill_2 FILLER_24_961 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_fill_1 FILLER_24_1007 ();
 sg13g2_decap_8 FILLER_24_1026 ();
 sg13g2_decap_8 FILLER_24_1033 ();
 sg13g2_fill_2 FILLER_24_1040 ();
 sg13g2_fill_1 FILLER_24_1042 ();
 sg13g2_fill_1 FILLER_24_1075 ();
 sg13g2_decap_8 FILLER_24_1109 ();
 sg13g2_fill_1 FILLER_24_1116 ();
 sg13g2_fill_2 FILLER_24_1140 ();
 sg13g2_fill_1 FILLER_24_1146 ();
 sg13g2_fill_1 FILLER_24_1161 ();
 sg13g2_fill_2 FILLER_24_1215 ();
 sg13g2_fill_1 FILLER_24_1222 ();
 sg13g2_fill_2 FILLER_24_1228 ();
 sg13g2_decap_4 FILLER_24_1241 ();
 sg13g2_fill_1 FILLER_24_1245 ();
 sg13g2_fill_2 FILLER_24_1251 ();
 sg13g2_fill_1 FILLER_24_1253 ();
 sg13g2_fill_2 FILLER_24_1272 ();
 sg13g2_decap_4 FILLER_24_1288 ();
 sg13g2_fill_1 FILLER_24_1296 ();
 sg13g2_decap_4 FILLER_24_1304 ();
 sg13g2_fill_2 FILLER_24_1316 ();
 sg13g2_fill_1 FILLER_24_1330 ();
 sg13g2_fill_1 FILLER_24_1342 ();
 sg13g2_fill_1 FILLER_24_1361 ();
 sg13g2_fill_1 FILLER_24_1379 ();
 sg13g2_fill_2 FILLER_24_1403 ();
 sg13g2_fill_1 FILLER_24_1434 ();
 sg13g2_fill_1 FILLER_24_1461 ();
 sg13g2_fill_1 FILLER_24_1469 ();
 sg13g2_fill_2 FILLER_24_1491 ();
 sg13g2_decap_4 FILLER_24_1503 ();
 sg13g2_fill_1 FILLER_24_1507 ();
 sg13g2_fill_1 FILLER_24_1534 ();
 sg13g2_fill_1 FILLER_24_1561 ();
 sg13g2_fill_2 FILLER_24_1566 ();
 sg13g2_fill_2 FILLER_24_1604 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_fill_2 FILLER_24_1624 ();
 sg13g2_fill_1 FILLER_24_1626 ();
 sg13g2_fill_1 FILLER_24_1635 ();
 sg13g2_fill_2 FILLER_24_1662 ();
 sg13g2_fill_1 FILLER_24_1664 ();
 sg13g2_decap_4 FILLER_24_1687 ();
 sg13g2_decap_8 FILLER_24_1695 ();
 sg13g2_fill_1 FILLER_24_1702 ();
 sg13g2_fill_2 FILLER_24_1707 ();
 sg13g2_fill_1 FILLER_24_1709 ();
 sg13g2_fill_1 FILLER_24_1732 ();
 sg13g2_fill_1 FILLER_24_1799 ();
 sg13g2_fill_1 FILLER_24_1821 ();
 sg13g2_fill_1 FILLER_24_1848 ();
 sg13g2_fill_1 FILLER_24_1854 ();
 sg13g2_decap_8 FILLER_24_1876 ();
 sg13g2_fill_2 FILLER_24_1883 ();
 sg13g2_fill_1 FILLER_24_1885 ();
 sg13g2_fill_2 FILLER_24_1890 ();
 sg13g2_fill_1 FILLER_24_1892 ();
 sg13g2_fill_2 FILLER_24_1928 ();
 sg13g2_fill_2 FILLER_24_1951 ();
 sg13g2_fill_1 FILLER_24_1953 ();
 sg13g2_fill_1 FILLER_24_1963 ();
 sg13g2_fill_2 FILLER_24_1990 ();
 sg13g2_fill_2 FILLER_24_2013 ();
 sg13g2_fill_1 FILLER_24_2015 ();
 sg13g2_fill_2 FILLER_24_2042 ();
 sg13g2_fill_1 FILLER_24_2044 ();
 sg13g2_decap_4 FILLER_24_2080 ();
 sg13g2_fill_1 FILLER_24_2084 ();
 sg13g2_decap_4 FILLER_24_2150 ();
 sg13g2_fill_1 FILLER_24_2154 ();
 sg13g2_decap_8 FILLER_24_2189 ();
 sg13g2_decap_8 FILLER_24_2196 ();
 sg13g2_decap_8 FILLER_24_2207 ();
 sg13g2_decap_8 FILLER_24_2214 ();
 sg13g2_fill_2 FILLER_24_2246 ();
 sg13g2_decap_4 FILLER_24_2274 ();
 sg13g2_fill_1 FILLER_24_2278 ();
 sg13g2_fill_2 FILLER_24_2345 ();
 sg13g2_decap_8 FILLER_24_2351 ();
 sg13g2_fill_2 FILLER_24_2384 ();
 sg13g2_fill_2 FILLER_24_2412 ();
 sg13g2_fill_1 FILLER_24_2414 ();
 sg13g2_fill_2 FILLER_24_2448 ();
 sg13g2_fill_1 FILLER_24_2454 ();
 sg13g2_fill_2 FILLER_24_2504 ();
 sg13g2_decap_4 FILLER_24_2526 ();
 sg13g2_fill_1 FILLER_24_2530 ();
 sg13g2_fill_2 FILLER_24_2541 ();
 sg13g2_decap_8 FILLER_24_2547 ();
 sg13g2_decap_8 FILLER_24_2554 ();
 sg13g2_decap_8 FILLER_24_2561 ();
 sg13g2_decap_4 FILLER_24_2568 ();
 sg13g2_fill_2 FILLER_24_2582 ();
 sg13g2_fill_1 FILLER_24_2584 ();
 sg13g2_decap_8 FILLER_24_2602 ();
 sg13g2_decap_8 FILLER_24_2609 ();
 sg13g2_decap_8 FILLER_24_2616 ();
 sg13g2_decap_8 FILLER_24_2623 ();
 sg13g2_fill_1 FILLER_24_2630 ();
 sg13g2_fill_2 FILLER_24_2667 ();
 sg13g2_fill_1 FILLER_24_2669 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_4 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_decap_4 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_4 FILLER_25_434 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_1 FILLER_25_457 ();
 sg13g2_fill_2 FILLER_25_463 ();
 sg13g2_decap_8 FILLER_25_491 ();
 sg13g2_decap_4 FILLER_25_554 ();
 sg13g2_fill_1 FILLER_25_599 ();
 sg13g2_fill_2 FILLER_25_625 ();
 sg13g2_fill_2 FILLER_25_642 ();
 sg13g2_fill_1 FILLER_25_698 ();
 sg13g2_fill_2 FILLER_25_712 ();
 sg13g2_fill_2 FILLER_25_729 ();
 sg13g2_fill_1 FILLER_25_743 ();
 sg13g2_fill_1 FILLER_25_748 ();
 sg13g2_fill_2 FILLER_25_754 ();
 sg13g2_fill_1 FILLER_25_792 ();
 sg13g2_fill_1 FILLER_25_830 ();
 sg13g2_fill_1 FILLER_25_841 ();
 sg13g2_fill_1 FILLER_25_874 ();
 sg13g2_fill_2 FILLER_25_888 ();
 sg13g2_fill_1 FILLER_25_930 ();
 sg13g2_decap_8 FILLER_25_957 ();
 sg13g2_decap_4 FILLER_25_964 ();
 sg13g2_fill_1 FILLER_25_968 ();
 sg13g2_fill_2 FILLER_25_998 ();
 sg13g2_fill_1 FILLER_25_1005 ();
 sg13g2_fill_2 FILLER_25_1010 ();
 sg13g2_fill_2 FILLER_25_1022 ();
 sg13g2_fill_2 FILLER_25_1044 ();
 sg13g2_fill_1 FILLER_25_1046 ();
 sg13g2_decap_8 FILLER_25_1054 ();
 sg13g2_fill_1 FILLER_25_1178 ();
 sg13g2_fill_2 FILLER_25_1235 ();
 sg13g2_fill_1 FILLER_25_1247 ();
 sg13g2_fill_2 FILLER_25_1262 ();
 sg13g2_decap_4 FILLER_25_1272 ();
 sg13g2_fill_1 FILLER_25_1301 ();
 sg13g2_fill_2 FILLER_25_1321 ();
 sg13g2_fill_2 FILLER_25_1353 ();
 sg13g2_fill_1 FILLER_25_1370 ();
 sg13g2_fill_1 FILLER_25_1378 ();
 sg13g2_fill_2 FILLER_25_1387 ();
 sg13g2_fill_2 FILLER_25_1397 ();
 sg13g2_fill_2 FILLER_25_1421 ();
 sg13g2_fill_1 FILLER_25_1440 ();
 sg13g2_fill_1 FILLER_25_1461 ();
 sg13g2_fill_1 FILLER_25_1472 ();
 sg13g2_fill_2 FILLER_25_1482 ();
 sg13g2_fill_1 FILLER_25_1487 ();
 sg13g2_decap_8 FILLER_25_1514 ();
 sg13g2_decap_4 FILLER_25_1521 ();
 sg13g2_fill_2 FILLER_25_1525 ();
 sg13g2_fill_1 FILLER_25_1537 ();
 sg13g2_fill_2 FILLER_25_1548 ();
 sg13g2_decap_8 FILLER_25_1558 ();
 sg13g2_decap_4 FILLER_25_1565 ();
 sg13g2_decap_8 FILLER_25_1579 ();
 sg13g2_fill_2 FILLER_25_1594 ();
 sg13g2_fill_2 FILLER_25_1632 ();
 sg13g2_fill_1 FILLER_25_1638 ();
 sg13g2_fill_1 FILLER_25_1648 ();
 sg13g2_fill_1 FILLER_25_1701 ();
 sg13g2_decap_8 FILLER_25_1706 ();
 sg13g2_fill_2 FILLER_25_1713 ();
 sg13g2_fill_2 FILLER_25_1727 ();
 sg13g2_fill_1 FILLER_25_1745 ();
 sg13g2_fill_2 FILLER_25_1818 ();
 sg13g2_decap_4 FILLER_25_1881 ();
 sg13g2_fill_1 FILLER_25_1966 ();
 sg13g2_fill_1 FILLER_25_1997 ();
 sg13g2_fill_1 FILLER_25_2050 ();
 sg13g2_fill_1 FILLER_25_2102 ();
 sg13g2_fill_1 FILLER_25_2108 ();
 sg13g2_fill_1 FILLER_25_2113 ();
 sg13g2_fill_2 FILLER_25_2211 ();
 sg13g2_fill_1 FILLER_25_2213 ();
 sg13g2_fill_1 FILLER_25_2239 ();
 sg13g2_fill_1 FILLER_25_2250 ();
 sg13g2_fill_2 FILLER_25_2259 ();
 sg13g2_fill_1 FILLER_25_2261 ();
 sg13g2_fill_2 FILLER_25_2266 ();
 sg13g2_fill_2 FILLER_25_2339 ();
 sg13g2_fill_1 FILLER_25_2351 ();
 sg13g2_decap_8 FILLER_25_2356 ();
 sg13g2_fill_2 FILLER_25_2363 ();
 sg13g2_fill_2 FILLER_25_2377 ();
 sg13g2_fill_2 FILLER_25_2432 ();
 sg13g2_fill_1 FILLER_25_2458 ();
 sg13g2_fill_1 FILLER_25_2499 ();
 sg13g2_fill_1 FILLER_25_2526 ();
 sg13g2_decap_8 FILLER_25_2558 ();
 sg13g2_decap_8 FILLER_25_2565 ();
 sg13g2_decap_8 FILLER_25_2572 ();
 sg13g2_fill_2 FILLER_25_2579 ();
 sg13g2_decap_8 FILLER_25_2622 ();
 sg13g2_fill_2 FILLER_25_2629 ();
 sg13g2_fill_2 FILLER_25_2667 ();
 sg13g2_fill_1 FILLER_25_2669 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_13 ();
 sg13g2_decap_4 FILLER_26_19 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_131 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_157 ();
 sg13g2_decap_4 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_368 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_decap_4 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_26_432 ();
 sg13g2_decap_4 FILLER_26_479 ();
 sg13g2_fill_2 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_495 ();
 sg13g2_decap_8 FILLER_26_502 ();
 sg13g2_decap_4 FILLER_26_509 ();
 sg13g2_fill_1 FILLER_26_513 ();
 sg13g2_fill_1 FILLER_26_518 ();
 sg13g2_fill_1 FILLER_26_533 ();
 sg13g2_decap_4 FILLER_26_554 ();
 sg13g2_fill_1 FILLER_26_576 ();
 sg13g2_fill_2 FILLER_26_638 ();
 sg13g2_fill_1 FILLER_26_661 ();
 sg13g2_fill_2 FILLER_26_674 ();
 sg13g2_fill_2 FILLER_26_746 ();
 sg13g2_fill_2 FILLER_26_771 ();
 sg13g2_fill_2 FILLER_26_777 ();
 sg13g2_fill_2 FILLER_26_783 ();
 sg13g2_fill_1 FILLER_26_785 ();
 sg13g2_fill_2 FILLER_26_791 ();
 sg13g2_fill_1 FILLER_26_793 ();
 sg13g2_fill_2 FILLER_26_818 ();
 sg13g2_fill_1 FILLER_26_834 ();
 sg13g2_fill_1 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_936 ();
 sg13g2_decap_8 FILLER_26_942 ();
 sg13g2_decap_8 FILLER_26_949 ();
 sg13g2_fill_1 FILLER_26_956 ();
 sg13g2_fill_2 FILLER_26_965 ();
 sg13g2_fill_1 FILLER_26_967 ();
 sg13g2_fill_1 FILLER_26_1022 ();
 sg13g2_fill_1 FILLER_26_1031 ();
 sg13g2_fill_1 FILLER_26_1047 ();
 sg13g2_fill_2 FILLER_26_1069 ();
 sg13g2_fill_2 FILLER_26_1080 ();
 sg13g2_fill_1 FILLER_26_1086 ();
 sg13g2_fill_2 FILLER_26_1113 ();
 sg13g2_fill_2 FILLER_26_1131 ();
 sg13g2_fill_2 FILLER_26_1153 ();
 sg13g2_fill_1 FILLER_26_1216 ();
 sg13g2_decap_4 FILLER_26_1235 ();
 sg13g2_fill_1 FILLER_26_1258 ();
 sg13g2_fill_1 FILLER_26_1264 ();
 sg13g2_fill_1 FILLER_26_1269 ();
 sg13g2_fill_1 FILLER_26_1276 ();
 sg13g2_fill_1 FILLER_26_1285 ();
 sg13g2_decap_4 FILLER_26_1327 ();
 sg13g2_fill_2 FILLER_26_1344 ();
 sg13g2_fill_2 FILLER_26_1380 ();
 sg13g2_decap_4 FILLER_26_1395 ();
 sg13g2_fill_1 FILLER_26_1416 ();
 sg13g2_fill_2 FILLER_26_1460 ();
 sg13g2_fill_1 FILLER_26_1493 ();
 sg13g2_decap_4 FILLER_26_1501 ();
 sg13g2_decap_8 FILLER_26_1541 ();
 sg13g2_decap_8 FILLER_26_1548 ();
 sg13g2_decap_8 FILLER_26_1555 ();
 sg13g2_decap_8 FILLER_26_1562 ();
 sg13g2_decap_8 FILLER_26_1569 ();
 sg13g2_decap_8 FILLER_26_1576 ();
 sg13g2_fill_2 FILLER_26_1583 ();
 sg13g2_fill_1 FILLER_26_1585 ();
 sg13g2_decap_8 FILLER_26_1590 ();
 sg13g2_decap_8 FILLER_26_1597 ();
 sg13g2_fill_2 FILLER_26_1604 ();
 sg13g2_fill_1 FILLER_26_1606 ();
 sg13g2_decap_8 FILLER_26_1624 ();
 sg13g2_decap_8 FILLER_26_1631 ();
 sg13g2_decap_8 FILLER_26_1638 ();
 sg13g2_fill_2 FILLER_26_1645 ();
 sg13g2_decap_4 FILLER_26_1651 ();
 sg13g2_decap_8 FILLER_26_1659 ();
 sg13g2_decap_8 FILLER_26_1666 ();
 sg13g2_fill_2 FILLER_26_1673 ();
 sg13g2_fill_1 FILLER_26_1675 ();
 sg13g2_fill_1 FILLER_26_1690 ();
 sg13g2_fill_2 FILLER_26_1722 ();
 sg13g2_fill_1 FILLER_26_1770 ();
 sg13g2_fill_2 FILLER_26_1795 ();
 sg13g2_decap_4 FILLER_26_1808 ();
 sg13g2_fill_1 FILLER_26_1812 ();
 sg13g2_fill_2 FILLER_26_1826 ();
 sg13g2_fill_2 FILLER_26_1832 ();
 sg13g2_fill_1 FILLER_26_1834 ();
 sg13g2_fill_2 FILLER_26_1897 ();
 sg13g2_fill_1 FILLER_26_1899 ();
 sg13g2_fill_2 FILLER_26_1978 ();
 sg13g2_fill_2 FILLER_26_2015 ();
 sg13g2_fill_1 FILLER_26_2056 ();
 sg13g2_decap_8 FILLER_26_2069 ();
 sg13g2_decap_8 FILLER_26_2076 ();
 sg13g2_decap_8 FILLER_26_2083 ();
 sg13g2_decap_8 FILLER_26_2090 ();
 sg13g2_decap_8 FILLER_26_2097 ();
 sg13g2_decap_8 FILLER_26_2104 ();
 sg13g2_decap_8 FILLER_26_2111 ();
 sg13g2_fill_2 FILLER_26_2118 ();
 sg13g2_fill_1 FILLER_26_2120 ();
 sg13g2_fill_1 FILLER_26_2130 ();
 sg13g2_decap_8 FILLER_26_2135 ();
 sg13g2_decap_8 FILLER_26_2142 ();
 sg13g2_decap_4 FILLER_26_2149 ();
 sg13g2_decap_8 FILLER_26_2249 ();
 sg13g2_decap_4 FILLER_26_2256 ();
 sg13g2_decap_8 FILLER_26_2270 ();
 sg13g2_fill_2 FILLER_26_2287 ();
 sg13g2_decap_4 FILLER_26_2302 ();
 sg13g2_fill_2 FILLER_26_2306 ();
 sg13g2_fill_2 FILLER_26_2334 ();
 sg13g2_decap_4 FILLER_26_2380 ();
 sg13g2_fill_1 FILLER_26_2405 ();
 sg13g2_fill_2 FILLER_26_2432 ();
 sg13g2_fill_2 FILLER_26_2553 ();
 sg13g2_fill_2 FILLER_26_2576 ();
 sg13g2_fill_2 FILLER_26_2604 ();
 sg13g2_fill_1 FILLER_26_2606 ();
 sg13g2_fill_2 FILLER_26_2633 ();
 sg13g2_fill_1 FILLER_26_2635 ();
 sg13g2_fill_2 FILLER_26_2662 ();
 sg13g2_fill_1 FILLER_26_2664 ();
 sg13g2_fill_1 FILLER_26_2669 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_decap_4 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_4 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_4 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_fill_2 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_fill_2 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_445 ();
 sg13g2_fill_2 FILLER_27_450 ();
 sg13g2_fill_1 FILLER_27_452 ();
 sg13g2_fill_1 FILLER_27_457 ();
 sg13g2_fill_1 FILLER_27_475 ();
 sg13g2_fill_2 FILLER_27_481 ();
 sg13g2_fill_1 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_493 ();
 sg13g2_decap_8 FILLER_27_500 ();
 sg13g2_decap_4 FILLER_27_507 ();
 sg13g2_fill_1 FILLER_27_511 ();
 sg13g2_fill_1 FILLER_27_531 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_fill_2 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_551 ();
 sg13g2_decap_8 FILLER_27_558 ();
 sg13g2_fill_2 FILLER_27_565 ();
 sg13g2_fill_2 FILLER_27_586 ();
 sg13g2_fill_2 FILLER_27_620 ();
 sg13g2_fill_1 FILLER_27_635 ();
 sg13g2_fill_2 FILLER_27_656 ();
 sg13g2_fill_1 FILLER_27_667 ();
 sg13g2_fill_2 FILLER_27_690 ();
 sg13g2_fill_1 FILLER_27_702 ();
 sg13g2_fill_1 FILLER_27_706 ();
 sg13g2_fill_1 FILLER_27_711 ();
 sg13g2_fill_1 FILLER_27_716 ();
 sg13g2_fill_2 FILLER_27_747 ();
 sg13g2_fill_1 FILLER_27_765 ();
 sg13g2_fill_2 FILLER_27_784 ();
 sg13g2_fill_1 FILLER_27_786 ();
 sg13g2_fill_2 FILLER_27_823 ();
 sg13g2_fill_2 FILLER_27_836 ();
 sg13g2_fill_1 FILLER_27_902 ();
 sg13g2_decap_8 FILLER_27_913 ();
 sg13g2_decap_8 FILLER_27_920 ();
 sg13g2_decap_8 FILLER_27_927 ();
 sg13g2_decap_8 FILLER_27_934 ();
 sg13g2_decap_8 FILLER_27_941 ();
 sg13g2_fill_1 FILLER_27_958 ();
 sg13g2_fill_1 FILLER_27_964 ();
 sg13g2_decap_4 FILLER_27_970 ();
 sg13g2_fill_1 FILLER_27_982 ();
 sg13g2_fill_1 FILLER_27_990 ();
 sg13g2_fill_2 FILLER_27_996 ();
 sg13g2_fill_1 FILLER_27_998 ();
 sg13g2_fill_1 FILLER_27_1008 ();
 sg13g2_fill_2 FILLER_27_1031 ();
 sg13g2_fill_1 FILLER_27_1045 ();
 sg13g2_fill_1 FILLER_27_1053 ();
 sg13g2_fill_2 FILLER_27_1072 ();
 sg13g2_fill_2 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1092 ();
 sg13g2_fill_2 FILLER_27_1098 ();
 sg13g2_fill_1 FILLER_27_1110 ();
 sg13g2_fill_2 FILLER_27_1145 ();
 sg13g2_fill_2 FILLER_27_1245 ();
 sg13g2_fill_1 FILLER_27_1251 ();
 sg13g2_fill_1 FILLER_27_1262 ();
 sg13g2_fill_2 FILLER_27_1289 ();
 sg13g2_fill_2 FILLER_27_1299 ();
 sg13g2_fill_2 FILLER_27_1320 ();
 sg13g2_fill_1 FILLER_27_1322 ();
 sg13g2_decap_8 FILLER_27_1336 ();
 sg13g2_fill_1 FILLER_27_1372 ();
 sg13g2_fill_1 FILLER_27_1377 ();
 sg13g2_fill_1 FILLER_27_1382 ();
 sg13g2_fill_1 FILLER_27_1393 ();
 sg13g2_fill_1 FILLER_27_1399 ();
 sg13g2_decap_4 FILLER_27_1404 ();
 sg13g2_fill_2 FILLER_27_1469 ();
 sg13g2_fill_1 FILLER_27_1485 ();
 sg13g2_decap_8 FILLER_27_1512 ();
 sg13g2_decap_4 FILLER_27_1519 ();
 sg13g2_decap_4 FILLER_27_1527 ();
 sg13g2_fill_1 FILLER_27_1531 ();
 sg13g2_fill_2 FILLER_27_1537 ();
 sg13g2_fill_2 FILLER_27_1604 ();
 sg13g2_fill_1 FILLER_27_1606 ();
 sg13g2_fill_1 FILLER_27_1637 ();
 sg13g2_fill_2 FILLER_27_1642 ();
 sg13g2_fill_2 FILLER_27_1675 ();
 sg13g2_decap_8 FILLER_27_1736 ();
 sg13g2_fill_2 FILLER_27_1743 ();
 sg13g2_fill_2 FILLER_27_1780 ();
 sg13g2_fill_1 FILLER_27_1789 ();
 sg13g2_fill_1 FILLER_27_1808 ();
 sg13g2_fill_2 FILLER_27_1814 ();
 sg13g2_fill_1 FILLER_27_1816 ();
 sg13g2_decap_8 FILLER_27_1821 ();
 sg13g2_decap_4 FILLER_27_1828 ();
 sg13g2_fill_1 FILLER_27_1832 ();
 sg13g2_decap_4 FILLER_27_1886 ();
 sg13g2_fill_1 FILLER_27_1890 ();
 sg13g2_fill_2 FILLER_27_1912 ();
 sg13g2_fill_1 FILLER_27_1914 ();
 sg13g2_fill_2 FILLER_27_1920 ();
 sg13g2_fill_2 FILLER_27_1939 ();
 sg13g2_fill_1 FILLER_27_1962 ();
 sg13g2_fill_2 FILLER_27_1993 ();
 sg13g2_fill_2 FILLER_27_2016 ();
 sg13g2_fill_1 FILLER_27_2018 ();
 sg13g2_fill_2 FILLER_27_2066 ();
 sg13g2_decap_4 FILLER_27_2072 ();
 sg13g2_decap_8 FILLER_27_2080 ();
 sg13g2_fill_2 FILLER_27_2087 ();
 sg13g2_fill_2 FILLER_27_2093 ();
 sg13g2_decap_8 FILLER_27_2100 ();
 sg13g2_fill_2 FILLER_27_2107 ();
 sg13g2_fill_1 FILLER_27_2113 ();
 sg13g2_fill_1 FILLER_27_2135 ();
 sg13g2_fill_1 FILLER_27_2140 ();
 sg13g2_decap_8 FILLER_27_2145 ();
 sg13g2_decap_8 FILLER_27_2152 ();
 sg13g2_fill_2 FILLER_27_2159 ();
 sg13g2_fill_1 FILLER_27_2161 ();
 sg13g2_fill_1 FILLER_27_2171 ();
 sg13g2_fill_2 FILLER_27_2202 ();
 sg13g2_fill_1 FILLER_27_2204 ();
 sg13g2_fill_1 FILLER_27_2210 ();
 sg13g2_fill_1 FILLER_27_2215 ();
 sg13g2_fill_2 FILLER_27_2242 ();
 sg13g2_decap_4 FILLER_27_2249 ();
 sg13g2_fill_1 FILLER_27_2352 ();
 sg13g2_fill_1 FILLER_27_2357 ();
 sg13g2_fill_2 FILLER_27_2387 ();
 sg13g2_fill_2 FILLER_27_2421 ();
 sg13g2_fill_1 FILLER_27_2423 ();
 sg13g2_fill_1 FILLER_27_2455 ();
 sg13g2_decap_8 FILLER_27_2464 ();
 sg13g2_decap_4 FILLER_27_2471 ();
 sg13g2_decap_8 FILLER_27_2515 ();
 sg13g2_fill_1 FILLER_27_2522 ();
 sg13g2_fill_2 FILLER_27_2589 ();
 sg13g2_fill_1 FILLER_27_2591 ();
 sg13g2_fill_2 FILLER_27_2668 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_120 ();
 sg13g2_decap_4 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_decap_4 FILLER_28_364 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_decap_4 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_415 ();
 sg13g2_fill_2 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_435 ();
 sg13g2_decap_4 FILLER_28_445 ();
 sg13g2_decap_4 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_481 ();
 sg13g2_fill_1 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_492 ();
 sg13g2_fill_1 FILLER_28_499 ();
 sg13g2_fill_2 FILLER_28_536 ();
 sg13g2_fill_1 FILLER_28_538 ();
 sg13g2_fill_1 FILLER_28_585 ();
 sg13g2_decap_4 FILLER_28_596 ();
 sg13g2_fill_2 FILLER_28_600 ();
 sg13g2_fill_2 FILLER_28_607 ();
 sg13g2_fill_1 FILLER_28_639 ();
 sg13g2_fill_1 FILLER_28_647 ();
 sg13g2_fill_2 FILLER_28_708 ();
 sg13g2_fill_2 FILLER_28_741 ();
 sg13g2_fill_1 FILLER_28_746 ();
 sg13g2_fill_2 FILLER_28_768 ();
 sg13g2_fill_2 FILLER_28_796 ();
 sg13g2_fill_1 FILLER_28_798 ();
 sg13g2_fill_2 FILLER_28_829 ();
 sg13g2_fill_2 FILLER_28_854 ();
 sg13g2_fill_2 FILLER_28_875 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_decap_8 FILLER_28_924 ();
 sg13g2_decap_8 FILLER_28_931 ();
 sg13g2_fill_2 FILLER_28_938 ();
 sg13g2_fill_1 FILLER_28_940 ();
 sg13g2_fill_2 FILLER_28_961 ();
 sg13g2_fill_2 FILLER_28_973 ();
 sg13g2_fill_2 FILLER_28_980 ();
 sg13g2_fill_2 FILLER_28_987 ();
 sg13g2_fill_1 FILLER_28_989 ();
 sg13g2_fill_2 FILLER_28_995 ();
 sg13g2_fill_1 FILLER_28_997 ();
 sg13g2_fill_1 FILLER_28_1023 ();
 sg13g2_fill_1 FILLER_28_1051 ();
 sg13g2_fill_1 FILLER_28_1057 ();
 sg13g2_fill_1 FILLER_28_1063 ();
 sg13g2_fill_1 FILLER_28_1073 ();
 sg13g2_fill_1 FILLER_28_1090 ();
 sg13g2_fill_2 FILLER_28_1119 ();
 sg13g2_fill_1 FILLER_28_1130 ();
 sg13g2_fill_1 FILLER_28_1236 ();
 sg13g2_fill_2 FILLER_28_1245 ();
 sg13g2_fill_2 FILLER_28_1261 ();
 sg13g2_fill_1 FILLER_28_1282 ();
 sg13g2_fill_1 FILLER_28_1301 ();
 sg13g2_fill_1 FILLER_28_1306 ();
 sg13g2_fill_1 FILLER_28_1312 ();
 sg13g2_decap_4 FILLER_28_1360 ();
 sg13g2_fill_2 FILLER_28_1368 ();
 sg13g2_fill_1 FILLER_28_1370 ();
 sg13g2_decap_4 FILLER_28_1400 ();
 sg13g2_fill_2 FILLER_28_1404 ();
 sg13g2_decap_8 FILLER_28_1411 ();
 sg13g2_fill_1 FILLER_28_1432 ();
 sg13g2_fill_2 FILLER_28_1447 ();
 sg13g2_decap_8 FILLER_28_1509 ();
 sg13g2_decap_8 FILLER_28_1516 ();
 sg13g2_fill_2 FILLER_28_1523 ();
 sg13g2_fill_1 FILLER_28_1659 ();
 sg13g2_fill_2 FILLER_28_1694 ();
 sg13g2_fill_1 FILLER_28_1696 ();
 sg13g2_fill_1 FILLER_28_1724 ();
 sg13g2_fill_2 FILLER_28_1784 ();
 sg13g2_decap_8 FILLER_28_1833 ();
 sg13g2_fill_2 FILLER_28_1840 ();
 sg13g2_fill_1 FILLER_28_1865 ();
 sg13g2_decap_8 FILLER_28_1893 ();
 sg13g2_decap_4 FILLER_28_1904 ();
 sg13g2_fill_1 FILLER_28_1908 ();
 sg13g2_fill_1 FILLER_28_1999 ();
 sg13g2_decap_4 FILLER_28_2030 ();
 sg13g2_fill_1 FILLER_28_2060 ();
 sg13g2_fill_1 FILLER_28_2087 ();
 sg13g2_fill_1 FILLER_28_2093 ();
 sg13g2_fill_2 FILLER_28_2154 ();
 sg13g2_fill_2 FILLER_28_2177 ();
 sg13g2_fill_1 FILLER_28_2188 ();
 sg13g2_fill_1 FILLER_28_2193 ();
 sg13g2_decap_4 FILLER_28_2198 ();
 sg13g2_fill_2 FILLER_28_2207 ();
 sg13g2_fill_1 FILLER_28_2209 ();
 sg13g2_fill_2 FILLER_28_2330 ();
 sg13g2_fill_1 FILLER_28_2359 ();
 sg13g2_fill_2 FILLER_28_2412 ();
 sg13g2_fill_1 FILLER_28_2482 ();
 sg13g2_fill_1 FILLER_28_2515 ();
 sg13g2_decap_8 FILLER_28_2524 ();
 sg13g2_fill_2 FILLER_28_2531 ();
 sg13g2_fill_2 FILLER_28_2537 ();
 sg13g2_fill_1 FILLER_28_2539 ();
 sg13g2_decap_4 FILLER_28_2544 ();
 sg13g2_fill_2 FILLER_28_2585 ();
 sg13g2_fill_1 FILLER_28_2587 ();
 sg13g2_decap_8 FILLER_28_2657 ();
 sg13g2_decap_4 FILLER_28_2664 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_13 ();
 sg13g2_fill_1 FILLER_29_17 ();
 sg13g2_decap_8 FILLER_29_22 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_2 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_424 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_29_456 ();
 sg13g2_fill_2 FILLER_29_484 ();
 sg13g2_fill_1 FILLER_29_486 ();
 sg13g2_decap_8 FILLER_29_531 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_decap_4 FILLER_29_598 ();
 sg13g2_decap_4 FILLER_29_607 ();
 sg13g2_fill_1 FILLER_29_664 ();
 sg13g2_fill_2 FILLER_29_674 ();
 sg13g2_fill_1 FILLER_29_696 ();
 sg13g2_fill_1 FILLER_29_717 ();
 sg13g2_fill_1 FILLER_29_739 ();
 sg13g2_fill_1 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_788 ();
 sg13g2_fill_1 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_fill_2 FILLER_29_821 ();
 sg13g2_fill_1 FILLER_29_823 ();
 sg13g2_fill_1 FILLER_29_836 ();
 sg13g2_fill_1 FILLER_29_844 ();
 sg13g2_fill_1 FILLER_29_849 ();
 sg13g2_fill_2 FILLER_29_867 ();
 sg13g2_decap_8 FILLER_29_914 ();
 sg13g2_decap_8 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_928 ();
 sg13g2_fill_2 FILLER_29_977 ();
 sg13g2_fill_1 FILLER_29_979 ();
 sg13g2_decap_8 FILLER_29_985 ();
 sg13g2_fill_2 FILLER_29_997 ();
 sg13g2_fill_1 FILLER_29_1030 ();
 sg13g2_fill_2 FILLER_29_1036 ();
 sg13g2_fill_2 FILLER_29_1074 ();
 sg13g2_fill_2 FILLER_29_1095 ();
 sg13g2_fill_2 FILLER_29_1122 ();
 sg13g2_fill_2 FILLER_29_1231 ();
 sg13g2_fill_2 FILLER_29_1242 ();
 sg13g2_fill_2 FILLER_29_1248 ();
 sg13g2_fill_1 FILLER_29_1264 ();
 sg13g2_fill_1 FILLER_29_1274 ();
 sg13g2_fill_2 FILLER_29_1286 ();
 sg13g2_fill_1 FILLER_29_1295 ();
 sg13g2_fill_2 FILLER_29_1335 ();
 sg13g2_fill_1 FILLER_29_1350 ();
 sg13g2_fill_2 FILLER_29_1356 ();
 sg13g2_fill_1 FILLER_29_1358 ();
 sg13g2_decap_4 FILLER_29_1416 ();
 sg13g2_fill_1 FILLER_29_1430 ();
 sg13g2_fill_2 FILLER_29_1448 ();
 sg13g2_fill_2 FILLER_29_1456 ();
 sg13g2_fill_2 FILLER_29_1484 ();
 sg13g2_fill_2 FILLER_29_1567 ();
 sg13g2_fill_1 FILLER_29_1609 ();
 sg13g2_decap_4 FILLER_29_1623 ();
 sg13g2_fill_1 FILLER_29_1632 ();
 sg13g2_decap_8 FILLER_29_1662 ();
 sg13g2_decap_8 FILLER_29_1690 ();
 sg13g2_decap_4 FILLER_29_1697 ();
 sg13g2_fill_1 FILLER_29_1701 ();
 sg13g2_decap_8 FILLER_29_1706 ();
 sg13g2_fill_1 FILLER_29_1720 ();
 sg13g2_fill_1 FILLER_29_1779 ();
 sg13g2_decap_8 FILLER_29_1806 ();
 sg13g2_decap_8 FILLER_29_1839 ();
 sg13g2_fill_2 FILLER_29_1846 ();
 sg13g2_fill_1 FILLER_29_1848 ();
 sg13g2_decap_4 FILLER_29_1944 ();
 sg13g2_decap_4 FILLER_29_1952 ();
 sg13g2_fill_2 FILLER_29_1956 ();
 sg13g2_fill_1 FILLER_29_2031 ();
 sg13g2_fill_1 FILLER_29_2037 ();
 sg13g2_fill_1 FILLER_29_2043 ();
 sg13g2_fill_1 FILLER_29_2106 ();
 sg13g2_fill_1 FILLER_29_2158 ();
 sg13g2_fill_2 FILLER_29_2167 ();
 sg13g2_decap_8 FILLER_29_2195 ();
 sg13g2_decap_8 FILLER_29_2202 ();
 sg13g2_decap_8 FILLER_29_2209 ();
 sg13g2_fill_2 FILLER_29_2216 ();
 sg13g2_fill_2 FILLER_29_2230 ();
 sg13g2_fill_2 FILLER_29_2248 ();
 sg13g2_fill_1 FILLER_29_2311 ();
 sg13g2_fill_2 FILLER_29_2323 ();
 sg13g2_decap_4 FILLER_29_2371 ();
 sg13g2_fill_2 FILLER_29_2401 ();
 sg13g2_fill_2 FILLER_29_2440 ();
 sg13g2_fill_1 FILLER_29_2468 ();
 sg13g2_fill_1 FILLER_29_2495 ();
 sg13g2_fill_1 FILLER_29_2517 ();
 sg13g2_decap_8 FILLER_29_2544 ();
 sg13g2_decap_8 FILLER_29_2551 ();
 sg13g2_decap_8 FILLER_29_2558 ();
 sg13g2_decap_4 FILLER_29_2565 ();
 sg13g2_fill_1 FILLER_29_2569 ();
 sg13g2_decap_8 FILLER_29_2580 ();
 sg13g2_decap_8 FILLER_29_2587 ();
 sg13g2_decap_8 FILLER_29_2619 ();
 sg13g2_decap_8 FILLER_29_2626 ();
 sg13g2_decap_8 FILLER_29_2633 ();
 sg13g2_decap_8 FILLER_29_2640 ();
 sg13g2_decap_8 FILLER_29_2647 ();
 sg13g2_decap_8 FILLER_29_2654 ();
 sg13g2_decap_8 FILLER_29_2661 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_decap_8 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_43 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_decap_4 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_decap_4 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_fill_1 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_460 ();
 sg13g2_fill_2 FILLER_30_471 ();
 sg13g2_fill_2 FILLER_30_512 ();
 sg13g2_fill_1 FILLER_30_514 ();
 sg13g2_fill_1 FILLER_30_531 ();
 sg13g2_decap_8 FILLER_30_552 ();
 sg13g2_fill_2 FILLER_30_559 ();
 sg13g2_decap_4 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_605 ();
 sg13g2_decap_4 FILLER_30_617 ();
 sg13g2_fill_1 FILLER_30_621 ();
 sg13g2_decap_4 FILLER_30_625 ();
 sg13g2_fill_2 FILLER_30_629 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_fill_2 FILLER_30_658 ();
 sg13g2_fill_1 FILLER_30_660 ();
 sg13g2_fill_1 FILLER_30_676 ();
 sg13g2_fill_2 FILLER_30_685 ();
 sg13g2_fill_2 FILLER_30_692 ();
 sg13g2_fill_1 FILLER_30_707 ();
 sg13g2_fill_2 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_fill_1 FILLER_30_771 ();
 sg13g2_decap_8 FILLER_30_782 ();
 sg13g2_decap_8 FILLER_30_789 ();
 sg13g2_decap_4 FILLER_30_796 ();
 sg13g2_fill_2 FILLER_30_821 ();
 sg13g2_decap_4 FILLER_30_877 ();
 sg13g2_fill_2 FILLER_30_881 ();
 sg13g2_decap_8 FILLER_30_886 ();
 sg13g2_fill_2 FILLER_30_893 ();
 sg13g2_decap_8 FILLER_30_911 ();
 sg13g2_fill_2 FILLER_30_918 ();
 sg13g2_decap_4 FILLER_30_924 ();
 sg13g2_fill_1 FILLER_30_942 ();
 sg13g2_fill_2 FILLER_30_952 ();
 sg13g2_fill_1 FILLER_30_972 ();
 sg13g2_fill_1 FILLER_30_989 ();
 sg13g2_fill_2 FILLER_30_1011 ();
 sg13g2_fill_1 FILLER_30_1036 ();
 sg13g2_fill_2 FILLER_30_1054 ();
 sg13g2_fill_1 FILLER_30_1067 ();
 sg13g2_fill_2 FILLER_30_1076 ();
 sg13g2_fill_1 FILLER_30_1088 ();
 sg13g2_fill_1 FILLER_30_1115 ();
 sg13g2_fill_2 FILLER_30_1146 ();
 sg13g2_fill_1 FILLER_30_1181 ();
 sg13g2_fill_2 FILLER_30_1215 ();
 sg13g2_fill_1 FILLER_30_1220 ();
 sg13g2_fill_2 FILLER_30_1225 ();
 sg13g2_fill_2 FILLER_30_1239 ();
 sg13g2_fill_2 FILLER_30_1288 ();
 sg13g2_fill_1 FILLER_30_1290 ();
 sg13g2_fill_1 FILLER_30_1323 ();
 sg13g2_decap_4 FILLER_30_1346 ();
 sg13g2_fill_1 FILLER_30_1350 ();
 sg13g2_fill_2 FILLER_30_1356 ();
 sg13g2_decap_4 FILLER_30_1362 ();
 sg13g2_fill_2 FILLER_30_1374 ();
 sg13g2_fill_2 FILLER_30_1389 ();
 sg13g2_fill_1 FILLER_30_1395 ();
 sg13g2_fill_1 FILLER_30_1400 ();
 sg13g2_fill_1 FILLER_30_1405 ();
 sg13g2_fill_2 FILLER_30_1411 ();
 sg13g2_fill_2 FILLER_30_1423 ();
 sg13g2_fill_2 FILLER_30_1437 ();
 sg13g2_fill_2 FILLER_30_1488 ();
 sg13g2_fill_2 FILLER_30_1498 ();
 sg13g2_fill_2 FILLER_30_1526 ();
 sg13g2_fill_1 FILLER_30_1590 ();
 sg13g2_fill_1 FILLER_30_1604 ();
 sg13g2_fill_1 FILLER_30_1631 ();
 sg13g2_decap_8 FILLER_30_1664 ();
 sg13g2_fill_2 FILLER_30_1685 ();
 sg13g2_decap_8 FILLER_30_1691 ();
 sg13g2_fill_2 FILLER_30_1698 ();
 sg13g2_fill_1 FILLER_30_1700 ();
 sg13g2_fill_2 FILLER_30_1709 ();
 sg13g2_fill_1 FILLER_30_1734 ();
 sg13g2_fill_2 FILLER_30_1743 ();
 sg13g2_fill_2 FILLER_30_1765 ();
 sg13g2_fill_1 FILLER_30_1767 ();
 sg13g2_decap_4 FILLER_30_1823 ();
 sg13g2_fill_2 FILLER_30_1827 ();
 sg13g2_decap_8 FILLER_30_1859 ();
 sg13g2_fill_2 FILLER_30_1869 ();
 sg13g2_decap_4 FILLER_30_1969 ();
 sg13g2_fill_1 FILLER_30_1973 ();
 sg13g2_fill_1 FILLER_30_1978 ();
 sg13g2_fill_1 FILLER_30_2010 ();
 sg13g2_fill_2 FILLER_30_2032 ();
 sg13g2_fill_1 FILLER_30_2039 ();
 sg13g2_fill_1 FILLER_30_2044 ();
 sg13g2_fill_1 FILLER_30_2049 ();
 sg13g2_decap_8 FILLER_30_2080 ();
 sg13g2_fill_1 FILLER_30_2087 ();
 sg13g2_fill_1 FILLER_30_2092 ();
 sg13g2_fill_2 FILLER_30_2136 ();
 sg13g2_fill_1 FILLER_30_2164 ();
 sg13g2_fill_1 FILLER_30_2169 ();
 sg13g2_fill_1 FILLER_30_2196 ();
 sg13g2_decap_8 FILLER_30_2232 ();
 sg13g2_decap_4 FILLER_30_2239 ();
 sg13g2_fill_2 FILLER_30_2243 ();
 sg13g2_fill_2 FILLER_30_2270 ();
 sg13g2_fill_1 FILLER_30_2291 ();
 sg13g2_fill_2 FILLER_30_2315 ();
 sg13g2_decap_4 FILLER_30_2335 ();
 sg13g2_fill_1 FILLER_30_2344 ();
 sg13g2_fill_2 FILLER_30_2351 ();
 sg13g2_fill_1 FILLER_30_2436 ();
 sg13g2_fill_2 FILLER_30_2461 ();
 sg13g2_fill_1 FILLER_30_2473 ();
 sg13g2_fill_2 FILLER_30_2490 ();
 sg13g2_fill_1 FILLER_30_2518 ();
 sg13g2_fill_2 FILLER_30_2540 ();
 sg13g2_fill_1 FILLER_30_2542 ();
 sg13g2_fill_2 FILLER_30_2547 ();
 sg13g2_decap_8 FILLER_30_2563 ();
 sg13g2_fill_1 FILLER_30_2570 ();
 sg13g2_fill_2 FILLER_30_2592 ();
 sg13g2_fill_1 FILLER_30_2594 ();
 sg13g2_fill_1 FILLER_30_2599 ();
 sg13g2_fill_2 FILLER_30_2624 ();
 sg13g2_fill_1 FILLER_30_2626 ();
 sg13g2_decap_8 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2644 ();
 sg13g2_decap_8 FILLER_30_2651 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_4 FILLER_30_2665 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_78 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_decap_4 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_decap_4 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_31_421 ();
 sg13g2_fill_2 FILLER_31_429 ();
 sg13g2_decap_4 FILLER_31_452 ();
 sg13g2_fill_2 FILLER_31_508 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_decap_4 FILLER_31_554 ();
 sg13g2_fill_1 FILLER_31_558 ();
 sg13g2_fill_2 FILLER_31_569 ();
 sg13g2_fill_1 FILLER_31_575 ();
 sg13g2_fill_2 FILLER_31_596 ();
 sg13g2_fill_1 FILLER_31_615 ();
 sg13g2_decap_8 FILLER_31_628 ();
 sg13g2_decap_4 FILLER_31_635 ();
 sg13g2_fill_1 FILLER_31_642 ();
 sg13g2_fill_1 FILLER_31_672 ();
 sg13g2_fill_1 FILLER_31_679 ();
 sg13g2_fill_2 FILLER_31_698 ();
 sg13g2_fill_1 FILLER_31_705 ();
 sg13g2_fill_1 FILLER_31_713 ();
 sg13g2_fill_1 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_4 FILLER_31_764 ();
 sg13g2_fill_1 FILLER_31_768 ();
 sg13g2_fill_2 FILLER_31_785 ();
 sg13g2_fill_2 FILLER_31_803 ();
 sg13g2_fill_1 FILLER_31_819 ();
 sg13g2_fill_1 FILLER_31_828 ();
 sg13g2_fill_1 FILLER_31_836 ();
 sg13g2_fill_2 FILLER_31_848 ();
 sg13g2_fill_2 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_fill_1 FILLER_31_882 ();
 sg13g2_fill_1 FILLER_31_893 ();
 sg13g2_decap_8 FILLER_31_914 ();
 sg13g2_fill_2 FILLER_31_921 ();
 sg13g2_decap_4 FILLER_31_931 ();
 sg13g2_fill_2 FILLER_31_935 ();
 sg13g2_fill_2 FILLER_31_958 ();
 sg13g2_fill_1 FILLER_31_988 ();
 sg13g2_fill_1 FILLER_31_999 ();
 sg13g2_decap_8 FILLER_31_1004 ();
 sg13g2_decap_4 FILLER_31_1015 ();
 sg13g2_fill_1 FILLER_31_1019 ();
 sg13g2_fill_2 FILLER_31_1037 ();
 sg13g2_fill_1 FILLER_31_1044 ();
 sg13g2_fill_1 FILLER_31_1072 ();
 sg13g2_fill_1 FILLER_31_1110 ();
 sg13g2_fill_2 FILLER_31_1119 ();
 sg13g2_fill_1 FILLER_31_1191 ();
 sg13g2_fill_1 FILLER_31_1195 ();
 sg13g2_fill_2 FILLER_31_1243 ();
 sg13g2_fill_2 FILLER_31_1269 ();
 sg13g2_fill_1 FILLER_31_1280 ();
 sg13g2_fill_1 FILLER_31_1326 ();
 sg13g2_decap_8 FILLER_31_1333 ();
 sg13g2_decap_8 FILLER_31_1340 ();
 sg13g2_decap_8 FILLER_31_1351 ();
 sg13g2_fill_2 FILLER_31_1358 ();
 sg13g2_fill_1 FILLER_31_1360 ();
 sg13g2_fill_2 FILLER_31_1371 ();
 sg13g2_fill_2 FILLER_31_1382 ();
 sg13g2_decap_8 FILLER_31_1394 ();
 sg13g2_decap_4 FILLER_31_1401 ();
 sg13g2_fill_2 FILLER_31_1405 ();
 sg13g2_fill_1 FILLER_31_1412 ();
 sg13g2_decap_8 FILLER_31_1416 ();
 sg13g2_fill_1 FILLER_31_1423 ();
 sg13g2_fill_2 FILLER_31_1456 ();
 sg13g2_fill_2 FILLER_31_1490 ();
 sg13g2_decap_4 FILLER_31_1525 ();
 sg13g2_fill_2 FILLER_31_1534 ();
 sg13g2_fill_2 FILLER_31_1545 ();
 sg13g2_fill_1 FILLER_31_1630 ();
 sg13g2_fill_2 FILLER_31_1635 ();
 sg13g2_fill_1 FILLER_31_1663 ();
 sg13g2_fill_2 FILLER_31_1667 ();
 sg13g2_fill_1 FILLER_31_1669 ();
 sg13g2_fill_1 FILLER_31_1706 ();
 sg13g2_decap_8 FILLER_31_1761 ();
 sg13g2_decap_8 FILLER_31_1768 ();
 sg13g2_decap_4 FILLER_31_1775 ();
 sg13g2_fill_1 FILLER_31_1779 ();
 sg13g2_decap_8 FILLER_31_1815 ();
 sg13g2_decap_8 FILLER_31_1822 ();
 sg13g2_decap_4 FILLER_31_1829 ();
 sg13g2_fill_1 FILLER_31_1833 ();
 sg13g2_decap_4 FILLER_31_1839 ();
 sg13g2_fill_2 FILLER_31_1843 ();
 sg13g2_fill_1 FILLER_31_1875 ();
 sg13g2_fill_2 FILLER_31_1887 ();
 sg13g2_fill_2 FILLER_31_1910 ();
 sg13g2_fill_1 FILLER_31_1912 ();
 sg13g2_fill_2 FILLER_31_1918 ();
 sg13g2_decap_4 FILLER_31_1946 ();
 sg13g2_fill_2 FILLER_31_1950 ();
 sg13g2_decap_8 FILLER_31_1977 ();
 sg13g2_fill_2 FILLER_31_2062 ();
 sg13g2_decap_8 FILLER_31_2085 ();
 sg13g2_fill_1 FILLER_31_2092 ();
 sg13g2_decap_4 FILLER_31_2097 ();
 sg13g2_fill_1 FILLER_31_2101 ();
 sg13g2_fill_1 FILLER_31_2106 ();
 sg13g2_fill_1 FILLER_31_2112 ();
 sg13g2_fill_1 FILLER_31_2125 ();
 sg13g2_fill_2 FILLER_31_2131 ();
 sg13g2_fill_2 FILLER_31_2155 ();
 sg13g2_decap_4 FILLER_31_2182 ();
 sg13g2_fill_2 FILLER_31_2186 ();
 sg13g2_fill_2 FILLER_31_2235 ();
 sg13g2_fill_2 FILLER_31_2241 ();
 sg13g2_fill_1 FILLER_31_2263 ();
 sg13g2_fill_2 FILLER_31_2271 ();
 sg13g2_fill_2 FILLER_31_2286 ();
 sg13g2_fill_2 FILLER_31_2331 ();
 sg13g2_fill_2 FILLER_31_2353 ();
 sg13g2_fill_1 FILLER_31_2365 ();
 sg13g2_decap_8 FILLER_31_2382 ();
 sg13g2_fill_2 FILLER_31_2393 ();
 sg13g2_fill_1 FILLER_31_2395 ();
 sg13g2_fill_2 FILLER_31_2468 ();
 sg13g2_fill_1 FILLER_31_2498 ();
 sg13g2_fill_1 FILLER_31_2610 ();
 sg13g2_fill_1 FILLER_31_2637 ();
 sg13g2_decap_4 FILLER_31_2664 ();
 sg13g2_fill_2 FILLER_31_2668 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_decap_8 FILLER_32_268 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_4 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_decap_4 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_decap_4 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_394 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_418 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_32_430 ();
 sg13g2_decap_8 FILLER_32_466 ();
 sg13g2_fill_2 FILLER_32_473 ();
 sg13g2_fill_1 FILLER_32_475 ();
 sg13g2_fill_2 FILLER_32_496 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_1 FILLER_32_513 ();
 sg13g2_decap_4 FILLER_32_522 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_fill_1 FILLER_32_532 ();
 sg13g2_decap_4 FILLER_32_537 ();
 sg13g2_fill_1 FILLER_32_541 ();
 sg13g2_fill_2 FILLER_32_573 ();
 sg13g2_fill_1 FILLER_32_575 ();
 sg13g2_decap_4 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_712 ();
 sg13g2_fill_1 FILLER_32_723 ();
 sg13g2_fill_1 FILLER_32_732 ();
 sg13g2_fill_1 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_786 ();
 sg13g2_fill_1 FILLER_32_793 ();
 sg13g2_fill_1 FILLER_32_820 ();
 sg13g2_decap_4 FILLER_32_849 ();
 sg13g2_fill_2 FILLER_32_853 ();
 sg13g2_fill_1 FILLER_32_866 ();
 sg13g2_fill_1 FILLER_32_893 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_fill_2 FILLER_32_931 ();
 sg13g2_fill_1 FILLER_32_933 ();
 sg13g2_fill_1 FILLER_32_947 ();
 sg13g2_fill_1 FILLER_32_961 ();
 sg13g2_fill_1 FILLER_32_970 ();
 sg13g2_fill_1 FILLER_32_992 ();
 sg13g2_fill_2 FILLER_32_1008 ();
 sg13g2_fill_1 FILLER_32_1010 ();
 sg13g2_fill_1 FILLER_32_1016 ();
 sg13g2_fill_2 FILLER_32_1033 ();
 sg13g2_fill_2 FILLER_32_1062 ();
 sg13g2_fill_2 FILLER_32_1146 ();
 sg13g2_fill_2 FILLER_32_1151 ();
 sg13g2_fill_1 FILLER_32_1191 ();
 sg13g2_fill_1 FILLER_32_1221 ();
 sg13g2_fill_1 FILLER_32_1233 ();
 sg13g2_fill_2 FILLER_32_1289 ();
 sg13g2_fill_2 FILLER_32_1339 ();
 sg13g2_decap_4 FILLER_32_1367 ();
 sg13g2_fill_2 FILLER_32_1371 ();
 sg13g2_decap_4 FILLER_32_1377 ();
 sg13g2_decap_8 FILLER_32_1411 ();
 sg13g2_fill_1 FILLER_32_1418 ();
 sg13g2_fill_2 FILLER_32_1428 ();
 sg13g2_fill_1 FILLER_32_1430 ();
 sg13g2_fill_1 FILLER_32_1456 ();
 sg13g2_decap_4 FILLER_32_1483 ();
 sg13g2_fill_1 FILLER_32_1487 ();
 sg13g2_decap_4 FILLER_32_1518 ();
 sg13g2_fill_2 FILLER_32_1531 ();
 sg13g2_fill_1 FILLER_32_1545 ();
 sg13g2_fill_1 FILLER_32_1571 ();
 sg13g2_fill_2 FILLER_32_1578 ();
 sg13g2_decap_8 FILLER_32_1611 ();
 sg13g2_decap_4 FILLER_32_1618 ();
 sg13g2_decap_4 FILLER_32_1652 ();
 sg13g2_fill_2 FILLER_32_1661 ();
 sg13g2_fill_1 FILLER_32_1663 ();
 sg13g2_fill_2 FILLER_32_1703 ();
 sg13g2_fill_1 FILLER_32_1705 ();
 sg13g2_decap_8 FILLER_32_1743 ();
 sg13g2_fill_1 FILLER_32_1750 ();
 sg13g2_decap_8 FILLER_32_1761 ();
 sg13g2_fill_2 FILLER_32_1768 ();
 sg13g2_fill_1 FILLER_32_1780 ();
 sg13g2_decap_8 FILLER_32_1807 ();
 sg13g2_decap_8 FILLER_32_1814 ();
 sg13g2_decap_8 FILLER_32_1844 ();
 sg13g2_decap_4 FILLER_32_1851 ();
 sg13g2_fill_1 FILLER_32_1855 ();
 sg13g2_decap_8 FILLER_32_1860 ();
 sg13g2_decap_8 FILLER_32_1867 ();
 sg13g2_fill_1 FILLER_32_1874 ();
 sg13g2_fill_2 FILLER_32_1904 ();
 sg13g2_fill_1 FILLER_32_1906 ();
 sg13g2_decap_8 FILLER_32_1941 ();
 sg13g2_decap_8 FILLER_32_1948 ();
 sg13g2_fill_2 FILLER_32_1955 ();
 sg13g2_decap_8 FILLER_32_1978 ();
 sg13g2_fill_2 FILLER_32_2041 ();
 sg13g2_decap_8 FILLER_32_2047 ();
 sg13g2_decap_8 FILLER_32_2054 ();
 sg13g2_decap_4 FILLER_32_2097 ();
 sg13g2_fill_1 FILLER_32_2101 ();
 sg13g2_decap_4 FILLER_32_2128 ();
 sg13g2_fill_1 FILLER_32_2132 ();
 sg13g2_decap_4 FILLER_32_2172 ();
 sg13g2_fill_1 FILLER_32_2176 ();
 sg13g2_decap_4 FILLER_32_2181 ();
 sg13g2_decap_8 FILLER_32_2199 ();
 sg13g2_fill_2 FILLER_32_2206 ();
 sg13g2_fill_1 FILLER_32_2208 ();
 sg13g2_fill_2 FILLER_32_2349 ();
 sg13g2_fill_1 FILLER_32_2361 ();
 sg13g2_fill_2 FILLER_32_2422 ();
 sg13g2_fill_1 FILLER_32_2440 ();
 sg13g2_fill_2 FILLER_32_2475 ();
 sg13g2_fill_2 FILLER_32_2523 ();
 sg13g2_fill_1 FILLER_32_2525 ();
 sg13g2_fill_1 FILLER_32_2560 ();
 sg13g2_decap_8 FILLER_32_2662 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_2 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_439 ();
 sg13g2_decap_4 FILLER_33_489 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_decap_4 FILLER_33_530 ();
 sg13g2_fill_2 FILLER_33_534 ();
 sg13g2_fill_2 FILLER_33_559 ();
 sg13g2_fill_2 FILLER_33_571 ();
 sg13g2_fill_2 FILLER_33_582 ();
 sg13g2_fill_1 FILLER_33_584 ();
 sg13g2_fill_1 FILLER_33_617 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_decap_4 FILLER_33_637 ();
 sg13g2_fill_2 FILLER_33_655 ();
 sg13g2_fill_1 FILLER_33_657 ();
 sg13g2_fill_1 FILLER_33_662 ();
 sg13g2_fill_1 FILLER_33_673 ();
 sg13g2_fill_2 FILLER_33_680 ();
 sg13g2_fill_1 FILLER_33_697 ();
 sg13g2_fill_1 FILLER_33_703 ();
 sg13g2_fill_1 FILLER_33_710 ();
 sg13g2_fill_2 FILLER_33_785 ();
 sg13g2_fill_2 FILLER_33_816 ();
 sg13g2_fill_1 FILLER_33_828 ();
 sg13g2_fill_2 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_860 ();
 sg13g2_decap_4 FILLER_33_867 ();
 sg13g2_fill_2 FILLER_33_871 ();
 sg13g2_fill_1 FILLER_33_885 ();
 sg13g2_fill_2 FILLER_33_905 ();
 sg13g2_decap_8 FILLER_33_915 ();
 sg13g2_fill_2 FILLER_33_927 ();
 sg13g2_fill_1 FILLER_33_929 ();
 sg13g2_decap_8 FILLER_33_934 ();
 sg13g2_fill_1 FILLER_33_941 ();
 sg13g2_decap_4 FILLER_33_954 ();
 sg13g2_fill_2 FILLER_33_958 ();
 sg13g2_decap_8 FILLER_33_964 ();
 sg13g2_decap_8 FILLER_33_971 ();
 sg13g2_fill_2 FILLER_33_978 ();
 sg13g2_fill_1 FILLER_33_980 ();
 sg13g2_fill_2 FILLER_33_1012 ();
 sg13g2_fill_1 FILLER_33_1024 ();
 sg13g2_fill_1 FILLER_33_1041 ();
 sg13g2_decap_4 FILLER_33_1045 ();
 sg13g2_fill_1 FILLER_33_1049 ();
 sg13g2_fill_1 FILLER_33_1076 ();
 sg13g2_fill_2 FILLER_33_1081 ();
 sg13g2_fill_1 FILLER_33_1095 ();
 sg13g2_fill_1 FILLER_33_1100 ();
 sg13g2_fill_2 FILLER_33_1151 ();
 sg13g2_fill_1 FILLER_33_1203 ();
 sg13g2_fill_1 FILLER_33_1207 ();
 sg13g2_fill_2 FILLER_33_1237 ();
 sg13g2_fill_1 FILLER_33_1283 ();
 sg13g2_decap_4 FILLER_33_1292 ();
 sg13g2_fill_2 FILLER_33_1296 ();
 sg13g2_fill_1 FILLER_33_1308 ();
 sg13g2_fill_1 FILLER_33_1316 ();
 sg13g2_decap_8 FILLER_33_1333 ();
 sg13g2_decap_8 FILLER_33_1340 ();
 sg13g2_decap_8 FILLER_33_1347 ();
 sg13g2_decap_8 FILLER_33_1354 ();
 sg13g2_fill_1 FILLER_33_1361 ();
 sg13g2_fill_1 FILLER_33_1372 ();
 sg13g2_decap_8 FILLER_33_1377 ();
 sg13g2_fill_2 FILLER_33_1394 ();
 sg13g2_fill_1 FILLER_33_1430 ();
 sg13g2_fill_1 FILLER_33_1463 ();
 sg13g2_decap_4 FILLER_33_1468 ();
 sg13g2_fill_1 FILLER_33_1472 ();
 sg13g2_decap_4 FILLER_33_1486 ();
 sg13g2_decap_4 FILLER_33_1493 ();
 sg13g2_decap_4 FILLER_33_1514 ();
 sg13g2_fill_2 FILLER_33_1518 ();
 sg13g2_fill_2 FILLER_33_1556 ();
 sg13g2_fill_1 FILLER_33_1562 ();
 sg13g2_fill_2 FILLER_33_1576 ();
 sg13g2_fill_1 FILLER_33_1585 ();
 sg13g2_fill_1 FILLER_33_1612 ();
 sg13g2_fill_1 FILLER_33_1619 ();
 sg13g2_fill_1 FILLER_33_1625 ();
 sg13g2_fill_1 FILLER_33_1630 ();
 sg13g2_fill_2 FILLER_33_1651 ();
 sg13g2_decap_8 FILLER_33_1669 ();
 sg13g2_fill_1 FILLER_33_1676 ();
 sg13g2_decap_8 FILLER_33_1721 ();
 sg13g2_decap_8 FILLER_33_1728 ();
 sg13g2_decap_8 FILLER_33_1735 ();
 sg13g2_fill_2 FILLER_33_1742 ();
 sg13g2_fill_1 FILLER_33_1821 ();
 sg13g2_fill_1 FILLER_33_1826 ();
 sg13g2_fill_1 FILLER_33_1874 ();
 sg13g2_fill_2 FILLER_33_1897 ();
 sg13g2_decap_8 FILLER_33_1924 ();
 sg13g2_decap_8 FILLER_33_1931 ();
 sg13g2_decap_4 FILLER_33_1942 ();
 sg13g2_decap_4 FILLER_33_1972 ();
 sg13g2_decap_4 FILLER_33_2006 ();
 sg13g2_decap_4 FILLER_33_2018 ();
 sg13g2_fill_2 FILLER_33_2022 ();
 sg13g2_decap_8 FILLER_33_2028 ();
 sg13g2_decap_8 FILLER_33_2035 ();
 sg13g2_fill_2 FILLER_33_2042 ();
 sg13g2_decap_4 FILLER_33_2054 ();
 sg13g2_decap_8 FILLER_33_2088 ();
 sg13g2_decap_4 FILLER_33_2095 ();
 sg13g2_fill_2 FILLER_33_2099 ();
 sg13g2_decap_8 FILLER_33_2174 ();
 sg13g2_decap_8 FILLER_33_2181 ();
 sg13g2_decap_8 FILLER_33_2188 ();
 sg13g2_decap_8 FILLER_33_2195 ();
 sg13g2_fill_1 FILLER_33_2202 ();
 sg13g2_decap_8 FILLER_33_2239 ();
 sg13g2_fill_2 FILLER_33_2246 ();
 sg13g2_decap_4 FILLER_33_2297 ();
 sg13g2_fill_1 FILLER_33_2309 ();
 sg13g2_decap_4 FILLER_33_2335 ();
 sg13g2_decap_4 FILLER_33_2365 ();
 sg13g2_fill_2 FILLER_33_2369 ();
 sg13g2_fill_2 FILLER_33_2405 ();
 sg13g2_fill_1 FILLER_33_2411 ();
 sg13g2_fill_1 FILLER_33_2464 ();
 sg13g2_decap_8 FILLER_33_2486 ();
 sg13g2_decap_8 FILLER_33_2493 ();
 sg13g2_decap_8 FILLER_33_2556 ();
 sg13g2_decap_4 FILLER_33_2563 ();
 sg13g2_fill_2 FILLER_33_2567 ();
 sg13g2_fill_1 FILLER_33_2579 ();
 sg13g2_fill_1 FILLER_33_2606 ();
 sg13g2_decap_8 FILLER_33_2638 ();
 sg13g2_decap_8 FILLER_33_2653 ();
 sg13g2_decap_8 FILLER_33_2660 ();
 sg13g2_fill_2 FILLER_33_2667 ();
 sg13g2_fill_1 FILLER_33_2669 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_16 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_32 ();
 sg13g2_decap_4 FILLER_34_39 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_4 FILLER_34_374 ();
 sg13g2_fill_1 FILLER_34_383 ();
 sg13g2_fill_2 FILLER_34_410 ();
 sg13g2_fill_1 FILLER_34_412 ();
 sg13g2_fill_1 FILLER_34_439 ();
 sg13g2_decap_4 FILLER_34_444 ();
 sg13g2_fill_2 FILLER_34_452 ();
 sg13g2_decap_4 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_477 ();
 sg13g2_fill_2 FILLER_34_496 ();
 sg13g2_decap_8 FILLER_34_528 ();
 sg13g2_decap_4 FILLER_34_535 ();
 sg13g2_fill_2 FILLER_34_557 ();
 sg13g2_fill_2 FILLER_34_565 ();
 sg13g2_fill_1 FILLER_34_597 ();
 sg13g2_fill_2 FILLER_34_609 ();
 sg13g2_decap_4 FILLER_34_624 ();
 sg13g2_fill_1 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_634 ();
 sg13g2_decap_8 FILLER_34_641 ();
 sg13g2_decap_8 FILLER_34_648 ();
 sg13g2_decap_8 FILLER_34_655 ();
 sg13g2_fill_2 FILLER_34_662 ();
 sg13g2_decap_4 FILLER_34_674 ();
 sg13g2_decap_4 FILLER_34_708 ();
 sg13g2_fill_2 FILLER_34_736 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_4 FILLER_34_756 ();
 sg13g2_fill_1 FILLER_34_764 ();
 sg13g2_fill_1 FILLER_34_769 ();
 sg13g2_fill_1 FILLER_34_774 ();
 sg13g2_fill_1 FILLER_34_785 ();
 sg13g2_decap_4 FILLER_34_794 ();
 sg13g2_fill_1 FILLER_34_808 ();
 sg13g2_fill_1 FILLER_34_819 ();
 sg13g2_fill_1 FILLER_34_824 ();
 sg13g2_fill_1 FILLER_34_848 ();
 sg13g2_fill_1 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_decap_8 FILLER_34_870 ();
 sg13g2_decap_4 FILLER_34_877 ();
 sg13g2_fill_2 FILLER_34_881 ();
 sg13g2_fill_2 FILLER_34_892 ();
 sg13g2_fill_1 FILLER_34_897 ();
 sg13g2_fill_2 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_930 ();
 sg13g2_decap_8 FILLER_34_937 ();
 sg13g2_decap_8 FILLER_34_944 ();
 sg13g2_decap_8 FILLER_34_951 ();
 sg13g2_decap_8 FILLER_34_958 ();
 sg13g2_decap_8 FILLER_34_965 ();
 sg13g2_decap_8 FILLER_34_972 ();
 sg13g2_fill_2 FILLER_34_979 ();
 sg13g2_fill_1 FILLER_34_996 ();
 sg13g2_fill_1 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1018 ();
 sg13g2_fill_2 FILLER_34_1034 ();
 sg13g2_fill_1 FILLER_34_1036 ();
 sg13g2_decap_8 FILLER_34_1042 ();
 sg13g2_fill_1 FILLER_34_1049 ();
 sg13g2_fill_1 FILLER_34_1076 ();
 sg13g2_fill_1 FILLER_34_1091 ();
 sg13g2_fill_1 FILLER_34_1132 ();
 sg13g2_fill_1 FILLER_34_1143 ();
 sg13g2_fill_2 FILLER_34_1170 ();
 sg13g2_fill_2 FILLER_34_1196 ();
 sg13g2_decap_4 FILLER_34_1294 ();
 sg13g2_fill_1 FILLER_34_1322 ();
 sg13g2_fill_2 FILLER_34_1358 ();
 sg13g2_fill_1 FILLER_34_1416 ();
 sg13g2_decap_4 FILLER_34_1450 ();
 sg13g2_fill_2 FILLER_34_1454 ();
 sg13g2_fill_1 FILLER_34_1486 ();
 sg13g2_fill_2 FILLER_34_1500 ();
 sg13g2_fill_1 FILLER_34_1502 ();
 sg13g2_fill_1 FILLER_34_1529 ();
 sg13g2_fill_2 FILLER_34_1534 ();
 sg13g2_fill_1 FILLER_34_1544 ();
 sg13g2_fill_1 FILLER_34_1563 ();
 sg13g2_decap_8 FILLER_34_1567 ();
 sg13g2_decap_4 FILLER_34_1574 ();
 sg13g2_fill_1 FILLER_34_1578 ();
 sg13g2_fill_2 FILLER_34_1587 ();
 sg13g2_decap_8 FILLER_34_1603 ();
 sg13g2_decap_4 FILLER_34_1610 ();
 sg13g2_fill_1 FILLER_34_1614 ();
 sg13g2_decap_4 FILLER_34_1620 ();
 sg13g2_decap_4 FILLER_34_1628 ();
 sg13g2_fill_2 FILLER_34_1632 ();
 sg13g2_decap_4 FILLER_34_1639 ();
 sg13g2_fill_2 FILLER_34_1643 ();
 sg13g2_decap_8 FILLER_34_1724 ();
 sg13g2_fill_1 FILLER_34_1731 ();
 sg13g2_fill_2 FILLER_34_1750 ();
 sg13g2_fill_1 FILLER_34_1752 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_8 FILLER_34_1764 ();
 sg13g2_fill_2 FILLER_34_1771 ();
 sg13g2_fill_1 FILLER_34_1787 ();
 sg13g2_fill_2 FILLER_34_1819 ();
 sg13g2_fill_1 FILLER_34_1873 ();
 sg13g2_fill_2 FILLER_34_1939 ();
 sg13g2_fill_1 FILLER_34_1941 ();
 sg13g2_decap_4 FILLER_34_1986 ();
 sg13g2_fill_2 FILLER_34_1990 ();
 sg13g2_decap_4 FILLER_34_2002 ();
 sg13g2_fill_2 FILLER_34_2006 ();
 sg13g2_decap_8 FILLER_34_2021 ();
 sg13g2_fill_2 FILLER_34_2028 ();
 sg13g2_fill_1 FILLER_34_2030 ();
 sg13g2_fill_1 FILLER_34_2041 ();
 sg13g2_decap_8 FILLER_34_2078 ();
 sg13g2_fill_2 FILLER_34_2085 ();
 sg13g2_fill_2 FILLER_34_2113 ();
 sg13g2_fill_2 FILLER_34_2141 ();
 sg13g2_fill_1 FILLER_34_2143 ();
 sg13g2_fill_1 FILLER_34_2149 ();
 sg13g2_fill_2 FILLER_34_2176 ();
 sg13g2_fill_1 FILLER_34_2178 ();
 sg13g2_fill_1 FILLER_34_2205 ();
 sg13g2_decap_8 FILLER_34_2214 ();
 sg13g2_decap_4 FILLER_34_2221 ();
 sg13g2_fill_1 FILLER_34_2225 ();
 sg13g2_decap_4 FILLER_34_2236 ();
 sg13g2_fill_1 FILLER_34_2240 ();
 sg13g2_decap_8 FILLER_34_2298 ();
 sg13g2_decap_8 FILLER_34_2305 ();
 sg13g2_fill_2 FILLER_34_2312 ();
 sg13g2_decap_8 FILLER_34_2324 ();
 sg13g2_decap_4 FILLER_34_2331 ();
 sg13g2_decap_8 FILLER_34_2340 ();
 sg13g2_decap_8 FILLER_34_2347 ();
 sg13g2_fill_2 FILLER_34_2354 ();
 sg13g2_fill_1 FILLER_34_2356 ();
 sg13g2_fill_1 FILLER_34_2378 ();
 sg13g2_fill_2 FILLER_34_2405 ();
 sg13g2_fill_1 FILLER_34_2433 ();
 sg13g2_fill_2 FILLER_34_2455 ();
 sg13g2_fill_2 FILLER_34_2467 ();
 sg13g2_fill_1 FILLER_34_2495 ();
 sg13g2_fill_2 FILLER_34_2511 ();
 sg13g2_decap_8 FILLER_34_2564 ();
 sg13g2_decap_4 FILLER_34_2571 ();
 sg13g2_fill_1 FILLER_34_2575 ();
 sg13g2_decap_8 FILLER_34_2605 ();
 sg13g2_decap_8 FILLER_34_2612 ();
 sg13g2_decap_8 FILLER_34_2623 ();
 sg13g2_decap_8 FILLER_34_2630 ();
 sg13g2_decap_8 FILLER_34_2637 ();
 sg13g2_decap_8 FILLER_34_2644 ();
 sg13g2_decap_8 FILLER_34_2651 ();
 sg13g2_decap_8 FILLER_34_2658 ();
 sg13g2_decap_4 FILLER_34_2665 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_102 ();
 sg13g2_decap_4 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_decap_4 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_4 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_372 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_4 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_2 FILLER_35_409 ();
 sg13g2_fill_1 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_439 ();
 sg13g2_fill_1 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_447 ();
 sg13g2_decap_8 FILLER_35_454 ();
 sg13g2_fill_2 FILLER_35_461 ();
 sg13g2_decap_4 FILLER_35_493 ();
 sg13g2_fill_2 FILLER_35_504 ();
 sg13g2_fill_1 FILLER_35_533 ();
 sg13g2_fill_2 FILLER_35_560 ();
 sg13g2_fill_1 FILLER_35_567 ();
 sg13g2_fill_1 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_592 ();
 sg13g2_fill_2 FILLER_35_599 ();
 sg13g2_fill_1 FILLER_35_611 ();
 sg13g2_fill_1 FILLER_35_638 ();
 sg13g2_decap_4 FILLER_35_670 ();
 sg13g2_fill_2 FILLER_35_674 ();
 sg13g2_fill_1 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_727 ();
 sg13g2_decap_4 FILLER_35_740 ();
 sg13g2_fill_1 FILLER_35_744 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_fill_1 FILLER_35_815 ();
 sg13g2_decap_4 FILLER_35_820 ();
 sg13g2_fill_2 FILLER_35_837 ();
 sg13g2_fill_1 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_866 ();
 sg13g2_decap_8 FILLER_35_873 ();
 sg13g2_decap_4 FILLER_35_880 ();
 sg13g2_fill_2 FILLER_35_884 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_decap_8 FILLER_35_897 ();
 sg13g2_fill_2 FILLER_35_904 ();
 sg13g2_decap_8 FILLER_35_950 ();
 sg13g2_decap_4 FILLER_35_957 ();
 sg13g2_decap_8 FILLER_35_965 ();
 sg13g2_decap_8 FILLER_35_972 ();
 sg13g2_fill_2 FILLER_35_979 ();
 sg13g2_fill_1 FILLER_35_984 ();
 sg13g2_fill_1 FILLER_35_1020 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_decap_4 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1047 ();
 sg13g2_fill_1 FILLER_35_1054 ();
 sg13g2_fill_1 FILLER_35_1077 ();
 sg13g2_fill_1 FILLER_35_1085 ();
 sg13g2_fill_2 FILLER_35_1117 ();
 sg13g2_fill_2 FILLER_35_1184 ();
 sg13g2_fill_1 FILLER_35_1214 ();
 sg13g2_fill_1 FILLER_35_1241 ();
 sg13g2_fill_2 FILLER_35_1273 ();
 sg13g2_fill_2 FILLER_35_1280 ();
 sg13g2_fill_1 FILLER_35_1282 ();
 sg13g2_fill_2 FILLER_35_1314 ();
 sg13g2_decap_8 FILLER_35_1346 ();
 sg13g2_fill_1 FILLER_35_1353 ();
 sg13g2_fill_2 FILLER_35_1359 ();
 sg13g2_fill_2 FILLER_35_1365 ();
 sg13g2_decap_8 FILLER_35_1371 ();
 sg13g2_decap_4 FILLER_35_1378 ();
 sg13g2_fill_1 FILLER_35_1400 ();
 sg13g2_fill_1 FILLER_35_1439 ();
 sg13g2_decap_4 FILLER_35_1456 ();
 sg13g2_decap_4 FILLER_35_1486 ();
 sg13g2_fill_1 FILLER_35_1490 ();
 sg13g2_fill_1 FILLER_35_1525 ();
 sg13g2_fill_2 FILLER_35_1634 ();
 sg13g2_fill_1 FILLER_35_1636 ();
 sg13g2_decap_4 FILLER_35_1643 ();
 sg13g2_fill_2 FILLER_35_1647 ();
 sg13g2_fill_1 FILLER_35_1712 ();
 sg13g2_decap_8 FILLER_35_1763 ();
 sg13g2_decap_8 FILLER_35_1770 ();
 sg13g2_decap_8 FILLER_35_1777 ();
 sg13g2_decap_4 FILLER_35_1784 ();
 sg13g2_fill_1 FILLER_35_1788 ();
 sg13g2_decap_8 FILLER_35_1807 ();
 sg13g2_fill_1 FILLER_35_1814 ();
 sg13g2_fill_1 FILLER_35_1829 ();
 sg13g2_fill_1 FILLER_35_1865 ();
 sg13g2_fill_1 FILLER_35_1890 ();
 sg13g2_fill_1 FILLER_35_1901 ();
 sg13g2_fill_2 FILLER_35_1932 ();
 sg13g2_fill_1 FILLER_35_1938 ();
 sg13g2_decap_8 FILLER_35_1994 ();
 sg13g2_decap_8 FILLER_35_2001 ();
 sg13g2_decap_8 FILLER_35_2008 ();
 sg13g2_decap_8 FILLER_35_2015 ();
 sg13g2_fill_2 FILLER_35_2022 ();
 sg13g2_fill_1 FILLER_35_2024 ();
 sg13g2_decap_8 FILLER_35_2059 ();
 sg13g2_fill_1 FILLER_35_2066 ();
 sg13g2_fill_1 FILLER_35_2094 ();
 sg13g2_decap_4 FILLER_35_2099 ();
 sg13g2_fill_1 FILLER_35_2103 ();
 sg13g2_fill_2 FILLER_35_2119 ();
 sg13g2_fill_2 FILLER_35_2173 ();
 sg13g2_fill_2 FILLER_35_2179 ();
 sg13g2_fill_1 FILLER_35_2181 ();
 sg13g2_decap_4 FILLER_35_2208 ();
 sg13g2_fill_1 FILLER_35_2212 ();
 sg13g2_fill_2 FILLER_35_2369 ();
 sg13g2_fill_1 FILLER_35_2371 ();
 sg13g2_fill_2 FILLER_35_2431 ();
 sg13g2_decap_4 FILLER_35_2469 ();
 sg13g2_fill_2 FILLER_35_2473 ();
 sg13g2_decap_8 FILLER_35_2479 ();
 sg13g2_fill_2 FILLER_35_2486 ();
 sg13g2_fill_1 FILLER_35_2488 ();
 sg13g2_decap_4 FILLER_35_2499 ();
 sg13g2_fill_1 FILLER_35_2532 ();
 sg13g2_decap_8 FILLER_35_2580 ();
 sg13g2_fill_2 FILLER_35_2587 ();
 sg13g2_decap_4 FILLER_35_2599 ();
 sg13g2_fill_2 FILLER_35_2603 ();
 sg13g2_decap_8 FILLER_35_2626 ();
 sg13g2_decap_8 FILLER_35_2633 ();
 sg13g2_decap_8 FILLER_35_2640 ();
 sg13g2_decap_8 FILLER_35_2647 ();
 sg13g2_decap_8 FILLER_35_2654 ();
 sg13g2_decap_8 FILLER_35_2661 ();
 sg13g2_fill_2 FILLER_35_2668 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_8 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_decap_4 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_369 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_decap_4 FILLER_36_420 ();
 sg13g2_decap_4 FILLER_36_465 ();
 sg13g2_fill_1 FILLER_36_473 ();
 sg13g2_fill_2 FILLER_36_478 ();
 sg13g2_fill_1 FILLER_36_480 ();
 sg13g2_fill_1 FILLER_36_489 ();
 sg13g2_fill_1 FILLER_36_516 ();
 sg13g2_fill_2 FILLER_36_537 ();
 sg13g2_decap_4 FILLER_36_544 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_2 FILLER_36_570 ();
 sg13g2_fill_1 FILLER_36_598 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_fill_1 FILLER_36_644 ();
 sg13g2_fill_1 FILLER_36_649 ();
 sg13g2_decap_4 FILLER_36_681 ();
 sg13g2_fill_2 FILLER_36_704 ();
 sg13g2_fill_2 FILLER_36_749 ();
 sg13g2_fill_1 FILLER_36_751 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_772 ();
 sg13g2_fill_2 FILLER_36_787 ();
 sg13g2_fill_1 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_4 FILLER_36_828 ();
 sg13g2_fill_1 FILLER_36_849 ();
 sg13g2_fill_1 FILLER_36_855 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_1 FILLER_36_867 ();
 sg13g2_decap_8 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_36_884 ();
 sg13g2_decap_8 FILLER_36_891 ();
 sg13g2_fill_1 FILLER_36_939 ();
 sg13g2_decap_4 FILLER_36_949 ();
 sg13g2_fill_2 FILLER_36_953 ();
 sg13g2_fill_1 FILLER_36_981 ();
 sg13g2_decap_8 FILLER_36_988 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_fill_1 FILLER_36_1008 ();
 sg13g2_fill_1 FILLER_36_1014 ();
 sg13g2_fill_2 FILLER_36_1020 ();
 sg13g2_decap_8 FILLER_36_1030 ();
 sg13g2_fill_2 FILLER_36_1037 ();
 sg13g2_fill_1 FILLER_36_1039 ();
 sg13g2_fill_1 FILLER_36_1050 ();
 sg13g2_fill_1 FILLER_36_1059 ();
 sg13g2_fill_1 FILLER_36_1065 ();
 sg13g2_fill_2 FILLER_36_1081 ();
 sg13g2_decap_8 FILLER_36_1092 ();
 sg13g2_fill_2 FILLER_36_1099 ();
 sg13g2_fill_2 FILLER_36_1113 ();
 sg13g2_fill_2 FILLER_36_1140 ();
 sg13g2_fill_2 FILLER_36_1147 ();
 sg13g2_fill_2 FILLER_36_1196 ();
 sg13g2_fill_2 FILLER_36_1201 ();
 sg13g2_fill_1 FILLER_36_1231 ();
 sg13g2_fill_1 FILLER_36_1246 ();
 sg13g2_fill_1 FILLER_36_1264 ();
 sg13g2_fill_2 FILLER_36_1278 ();
 sg13g2_fill_1 FILLER_36_1280 ();
 sg13g2_fill_1 FILLER_36_1284 ();
 sg13g2_fill_1 FILLER_36_1290 ();
 sg13g2_fill_1 FILLER_36_1305 ();
 sg13g2_decap_8 FILLER_36_1332 ();
 sg13g2_decap_8 FILLER_36_1339 ();
 sg13g2_decap_8 FILLER_36_1346 ();
 sg13g2_fill_2 FILLER_36_1353 ();
 sg13g2_fill_1 FILLER_36_1355 ();
 sg13g2_decap_8 FILLER_36_1382 ();
 sg13g2_fill_2 FILLER_36_1389 ();
 sg13g2_fill_2 FILLER_36_1404 ();
 sg13g2_decap_8 FILLER_36_1415 ();
 sg13g2_decap_8 FILLER_36_1422 ();
 sg13g2_decap_8 FILLER_36_1429 ();
 sg13g2_decap_8 FILLER_36_1436 ();
 sg13g2_decap_4 FILLER_36_1446 ();
 sg13g2_decap_8 FILLER_36_1489 ();
 sg13g2_fill_2 FILLER_36_1496 ();
 sg13g2_fill_1 FILLER_36_1498 ();
 sg13g2_decap_8 FILLER_36_1508 ();
 sg13g2_fill_2 FILLER_36_1524 ();
 sg13g2_fill_2 FILLER_36_1541 ();
 sg13g2_fill_1 FILLER_36_1543 ();
 sg13g2_fill_2 FILLER_36_1548 ();
 sg13g2_fill_1 FILLER_36_1550 ();
 sg13g2_decap_4 FILLER_36_1556 ();
 sg13g2_fill_2 FILLER_36_1560 ();
 sg13g2_decap_4 FILLER_36_1574 ();
 sg13g2_fill_1 FILLER_36_1578 ();
 sg13g2_fill_1 FILLER_36_1584 ();
 sg13g2_decap_8 FILLER_36_1594 ();
 sg13g2_decap_8 FILLER_36_1601 ();
 sg13g2_fill_2 FILLER_36_1608 ();
 sg13g2_fill_1 FILLER_36_1610 ();
 sg13g2_fill_1 FILLER_36_1653 ();
 sg13g2_fill_2 FILLER_36_1690 ();
 sg13g2_fill_2 FILLER_36_1700 ();
 sg13g2_fill_1 FILLER_36_1732 ();
 sg13g2_decap_8 FILLER_36_1775 ();
 sg13g2_decap_8 FILLER_36_1782 ();
 sg13g2_decap_8 FILLER_36_1789 ();
 sg13g2_decap_8 FILLER_36_1796 ();
 sg13g2_decap_8 FILLER_36_1803 ();
 sg13g2_decap_8 FILLER_36_1810 ();
 sg13g2_decap_8 FILLER_36_1817 ();
 sg13g2_decap_8 FILLER_36_1824 ();
 sg13g2_fill_1 FILLER_36_1831 ();
 sg13g2_fill_2 FILLER_36_1842 ();
 sg13g2_fill_1 FILLER_36_1852 ();
 sg13g2_decap_8 FILLER_36_1863 ();
 sg13g2_decap_8 FILLER_36_1870 ();
 sg13g2_fill_2 FILLER_36_1877 ();
 sg13g2_fill_2 FILLER_36_1895 ();
 sg13g2_fill_2 FILLER_36_1913 ();
 sg13g2_decap_8 FILLER_36_1941 ();
 sg13g2_fill_1 FILLER_36_1948 ();
 sg13g2_decap_8 FILLER_36_1986 ();
 sg13g2_fill_1 FILLER_36_1993 ();
 sg13g2_decap_8 FILLER_36_2008 ();
 sg13g2_decap_4 FILLER_36_2015 ();
 sg13g2_fill_1 FILLER_36_2019 ();
 sg13g2_decap_4 FILLER_36_2024 ();
 sg13g2_fill_1 FILLER_36_2028 ();
 sg13g2_decap_8 FILLER_36_2033 ();
 sg13g2_decap_8 FILLER_36_2040 ();
 sg13g2_decap_8 FILLER_36_2047 ();
 sg13g2_decap_4 FILLER_36_2054 ();
 sg13g2_fill_2 FILLER_36_2058 ();
 sg13g2_decap_8 FILLER_36_2065 ();
 sg13g2_decap_8 FILLER_36_2072 ();
 sg13g2_fill_1 FILLER_36_2079 ();
 sg13g2_decap_8 FILLER_36_2090 ();
 sg13g2_decap_8 FILLER_36_2097 ();
 sg13g2_decap_8 FILLER_36_2104 ();
 sg13g2_decap_8 FILLER_36_2111 ();
 sg13g2_fill_2 FILLER_36_2136 ();
 sg13g2_fill_1 FILLER_36_2138 ();
 sg13g2_decap_4 FILLER_36_2149 ();
 sg13g2_fill_2 FILLER_36_2153 ();
 sg13g2_decap_4 FILLER_36_2163 ();
 sg13g2_fill_2 FILLER_36_2177 ();
 sg13g2_decap_8 FILLER_36_2193 ();
 sg13g2_fill_1 FILLER_36_2200 ();
 sg13g2_fill_1 FILLER_36_2205 ();
 sg13g2_fill_2 FILLER_36_2246 ();
 sg13g2_decap_4 FILLER_36_2262 ();
 sg13g2_fill_2 FILLER_36_2266 ();
 sg13g2_fill_2 FILLER_36_2319 ();
 sg13g2_decap_8 FILLER_36_2351 ();
 sg13g2_fill_1 FILLER_36_2358 ();
 sg13g2_fill_2 FILLER_36_2377 ();
 sg13g2_fill_2 FILLER_36_2387 ();
 sg13g2_fill_1 FILLER_36_2389 ();
 sg13g2_fill_1 FILLER_36_2394 ();
 sg13g2_fill_2 FILLER_36_2400 ();
 sg13g2_fill_2 FILLER_36_2415 ();
 sg13g2_fill_2 FILLER_36_2421 ();
 sg13g2_fill_1 FILLER_36_2449 ();
 sg13g2_fill_2 FILLER_36_2454 ();
 sg13g2_decap_4 FILLER_36_2486 ();
 sg13g2_fill_1 FILLER_36_2490 ();
 sg13g2_fill_1 FILLER_36_2504 ();
 sg13g2_fill_2 FILLER_36_2509 ();
 sg13g2_fill_1 FILLER_36_2511 ();
 sg13g2_fill_1 FILLER_36_2539 ();
 sg13g2_fill_2 FILLER_36_2622 ();
 sg13g2_decap_8 FILLER_36_2654 ();
 sg13g2_decap_8 FILLER_36_2661 ();
 sg13g2_fill_2 FILLER_36_2668 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_38 ();
 sg13g2_decap_8 FILLER_37_43 ();
 sg13g2_decap_8 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_57 ();
 sg13g2_fill_1 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_decap_4 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_4 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_2 FILLER_37_383 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_2 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_fill_2 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_461 ();
 sg13g2_decap_4 FILLER_37_468 ();
 sg13g2_fill_2 FILLER_37_472 ();
 sg13g2_decap_4 FILLER_37_480 ();
 sg13g2_fill_1 FILLER_37_484 ();
 sg13g2_fill_1 FILLER_37_489 ();
 sg13g2_decap_8 FILLER_37_535 ();
 sg13g2_decap_8 FILLER_37_552 ();
 sg13g2_fill_1 FILLER_37_559 ();
 sg13g2_decap_4 FILLER_37_568 ();
 sg13g2_fill_2 FILLER_37_572 ();
 sg13g2_fill_2 FILLER_37_586 ();
 sg13g2_fill_1 FILLER_37_598 ();
 sg13g2_fill_2 FILLER_37_635 ();
 sg13g2_decap_4 FILLER_37_657 ();
 sg13g2_fill_1 FILLER_37_661 ();
 sg13g2_fill_2 FILLER_37_666 ();
 sg13g2_fill_1 FILLER_37_668 ();
 sg13g2_decap_4 FILLER_37_674 ();
 sg13g2_fill_1 FILLER_37_684 ();
 sg13g2_decap_4 FILLER_37_689 ();
 sg13g2_fill_2 FILLER_37_754 ();
 sg13g2_fill_1 FILLER_37_756 ();
 sg13g2_fill_2 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_824 ();
 sg13g2_fill_1 FILLER_37_837 ();
 sg13g2_decap_4 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_855 ();
 sg13g2_decap_8 FILLER_37_862 ();
 sg13g2_decap_8 FILLER_37_877 ();
 sg13g2_decap_8 FILLER_37_884 ();
 sg13g2_fill_2 FILLER_37_891 ();
 sg13g2_fill_2 FILLER_37_904 ();
 sg13g2_fill_1 FILLER_37_921 ();
 sg13g2_fill_1 FILLER_37_926 ();
 sg13g2_fill_1 FILLER_37_932 ();
 sg13g2_fill_1 FILLER_37_938 ();
 sg13g2_decap_4 FILLER_37_944 ();
 sg13g2_fill_1 FILLER_37_948 ();
 sg13g2_fill_1 FILLER_37_983 ();
 sg13g2_fill_1 FILLER_37_1034 ();
 sg13g2_fill_1 FILLER_37_1039 ();
 sg13g2_fill_2 FILLER_37_1053 ();
 sg13g2_fill_1 FILLER_37_1055 ();
 sg13g2_fill_1 FILLER_37_1103 ();
 sg13g2_fill_1 FILLER_37_1118 ();
 sg13g2_fill_1 FILLER_37_1125 ();
 sg13g2_fill_2 FILLER_37_1179 ();
 sg13g2_fill_2 FILLER_37_1193 ();
 sg13g2_fill_2 FILLER_37_1207 ();
 sg13g2_fill_2 FILLER_37_1219 ();
 sg13g2_fill_2 FILLER_37_1246 ();
 sg13g2_fill_1 FILLER_37_1248 ();
 sg13g2_fill_2 FILLER_37_1257 ();
 sg13g2_fill_1 FILLER_37_1259 ();
 sg13g2_fill_2 FILLER_37_1279 ();
 sg13g2_fill_2 FILLER_37_1284 ();
 sg13g2_fill_1 FILLER_37_1286 ();
 sg13g2_fill_1 FILLER_37_1321 ();
 sg13g2_decap_8 FILLER_37_1338 ();
 sg13g2_decap_4 FILLER_37_1345 ();
 sg13g2_fill_1 FILLER_37_1349 ();
 sg13g2_decap_8 FILLER_37_1368 ();
 sg13g2_decap_8 FILLER_37_1375 ();
 sg13g2_decap_8 FILLER_37_1382 ();
 sg13g2_decap_8 FILLER_37_1389 ();
 sg13g2_decap_4 FILLER_37_1396 ();
 sg13g2_decap_8 FILLER_37_1404 ();
 sg13g2_decap_8 FILLER_37_1411 ();
 sg13g2_decap_8 FILLER_37_1418 ();
 sg13g2_decap_8 FILLER_37_1425 ();
 sg13g2_decap_8 FILLER_37_1432 ();
 sg13g2_decap_8 FILLER_37_1439 ();
 sg13g2_decap_4 FILLER_37_1446 ();
 sg13g2_fill_1 FILLER_37_1450 ();
 sg13g2_fill_1 FILLER_37_1477 ();
 sg13g2_fill_2 FILLER_37_1487 ();
 sg13g2_fill_2 FILLER_37_1493 ();
 sg13g2_fill_2 FILLER_37_1525 ();
 sg13g2_fill_1 FILLER_37_1589 ();
 sg13g2_fill_2 FILLER_37_1598 ();
 sg13g2_fill_2 FILLER_37_1605 ();
 sg13g2_fill_1 FILLER_37_1672 ();
 sg13g2_fill_2 FILLER_37_1685 ();
 sg13g2_fill_2 FILLER_37_1696 ();
 sg13g2_fill_1 FILLER_37_1732 ();
 sg13g2_fill_1 FILLER_37_1746 ();
 sg13g2_fill_2 FILLER_37_1773 ();
 sg13g2_fill_2 FILLER_37_1805 ();
 sg13g2_fill_1 FILLER_37_1813 ();
 sg13g2_fill_2 FILLER_37_1817 ();
 sg13g2_decap_8 FILLER_37_1845 ();
 sg13g2_decap_8 FILLER_37_1852 ();
 sg13g2_decap_8 FILLER_37_1859 ();
 sg13g2_decap_8 FILLER_37_1866 ();
 sg13g2_decap_4 FILLER_37_1883 ();
 sg13g2_fill_1 FILLER_37_1891 ();
 sg13g2_decap_4 FILLER_37_1935 ();
 sg13g2_fill_2 FILLER_37_1943 ();
 sg13g2_fill_1 FILLER_37_1969 ();
 sg13g2_decap_4 FILLER_37_1980 ();
 sg13g2_fill_2 FILLER_37_2010 ();
 sg13g2_fill_1 FILLER_37_2012 ();
 sg13g2_decap_8 FILLER_37_2039 ();
 sg13g2_decap_8 FILLER_37_2046 ();
 sg13g2_decap_8 FILLER_37_2053 ();
 sg13g2_fill_2 FILLER_37_2074 ();
 sg13g2_fill_1 FILLER_37_2076 ();
 sg13g2_decap_8 FILLER_37_2103 ();
 sg13g2_decap_8 FILLER_37_2110 ();
 sg13g2_decap_8 FILLER_37_2117 ();
 sg13g2_decap_8 FILLER_37_2124 ();
 sg13g2_decap_8 FILLER_37_2131 ();
 sg13g2_decap_4 FILLER_37_2138 ();
 sg13g2_fill_1 FILLER_37_2142 ();
 sg13g2_decap_4 FILLER_37_2153 ();
 sg13g2_decap_8 FILLER_37_2181 ();
 sg13g2_decap_8 FILLER_37_2188 ();
 sg13g2_decap_8 FILLER_37_2195 ();
 sg13g2_decap_8 FILLER_37_2202 ();
 sg13g2_fill_2 FILLER_37_2213 ();
 sg13g2_fill_2 FILLER_37_2230 ();
 sg13g2_fill_1 FILLER_37_2232 ();
 sg13g2_decap_8 FILLER_37_2243 ();
 sg13g2_decap_8 FILLER_37_2250 ();
 sg13g2_decap_4 FILLER_37_2257 ();
 sg13g2_fill_1 FILLER_37_2261 ();
 sg13g2_decap_8 FILLER_37_2314 ();
 sg13g2_decap_4 FILLER_37_2335 ();
 sg13g2_fill_2 FILLER_37_2339 ();
 sg13g2_fill_2 FILLER_37_2398 ();
 sg13g2_fill_2 FILLER_37_2413 ();
 sg13g2_fill_1 FILLER_37_2415 ();
 sg13g2_fill_1 FILLER_37_2424 ();
 sg13g2_fill_2 FILLER_37_2435 ();
 sg13g2_fill_1 FILLER_37_2437 ();
 sg13g2_decap_8 FILLER_37_2442 ();
 sg13g2_decap_8 FILLER_37_2449 ();
 sg13g2_decap_4 FILLER_37_2456 ();
 sg13g2_fill_1 FILLER_37_2460 ();
 sg13g2_decap_4 FILLER_37_2471 ();
 sg13g2_decap_4 FILLER_37_2511 ();
 sg13g2_fill_2 FILLER_37_2515 ();
 sg13g2_fill_1 FILLER_37_2540 ();
 sg13g2_decap_8 FILLER_37_2553 ();
 sg13g2_fill_2 FILLER_37_2560 ();
 sg13g2_fill_2 FILLER_37_2572 ();
 sg13g2_decap_8 FILLER_37_2578 ();
 sg13g2_fill_1 FILLER_37_2585 ();
 sg13g2_decap_8 FILLER_37_2612 ();
 sg13g2_fill_1 FILLER_37_2619 ();
 sg13g2_decap_8 FILLER_37_2630 ();
 sg13g2_decap_8 FILLER_37_2637 ();
 sg13g2_decap_8 FILLER_37_2644 ();
 sg13g2_decap_8 FILLER_37_2651 ();
 sg13g2_decap_8 FILLER_37_2658 ();
 sg13g2_decap_4 FILLER_37_2665 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_fill_2 FILLER_38_31 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_decap_4 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_4 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_318 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_decap_4 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_4 FILLER_38_378 ();
 sg13g2_fill_2 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_411 ();
 sg13g2_fill_2 FILLER_38_418 ();
 sg13g2_fill_2 FILLER_38_424 ();
 sg13g2_fill_1 FILLER_38_431 ();
 sg13g2_fill_1 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_454 ();
 sg13g2_fill_1 FILLER_38_493 ();
 sg13g2_fill_1 FILLER_38_542 ();
 sg13g2_decap_4 FILLER_38_553 ();
 sg13g2_fill_1 FILLER_38_557 ();
 sg13g2_fill_2 FILLER_38_561 ();
 sg13g2_fill_1 FILLER_38_563 ();
 sg13g2_decap_4 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_572 ();
 sg13g2_decap_4 FILLER_38_580 ();
 sg13g2_fill_2 FILLER_38_588 ();
 sg13g2_fill_1 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_632 ();
 sg13g2_fill_2 FILLER_38_664 ();
 sg13g2_fill_1 FILLER_38_666 ();
 sg13g2_decap_4 FILLER_38_672 ();
 sg13g2_fill_1 FILLER_38_676 ();
 sg13g2_fill_2 FILLER_38_695 ();
 sg13g2_fill_2 FILLER_38_711 ();
 sg13g2_fill_1 FILLER_38_713 ();
 sg13g2_fill_1 FILLER_38_724 ();
 sg13g2_fill_1 FILLER_38_733 ();
 sg13g2_fill_2 FILLER_38_752 ();
 sg13g2_fill_2 FILLER_38_855 ();
 sg13g2_fill_2 FILLER_38_870 ();
 sg13g2_fill_1 FILLER_38_872 ();
 sg13g2_fill_2 FILLER_38_887 ();
 sg13g2_fill_1 FILLER_38_889 ();
 sg13g2_fill_1 FILLER_38_899 ();
 sg13g2_fill_1 FILLER_38_908 ();
 sg13g2_fill_1 FILLER_38_916 ();
 sg13g2_fill_1 FILLER_38_921 ();
 sg13g2_decap_4 FILLER_38_928 ();
 sg13g2_fill_2 FILLER_38_937 ();
 sg13g2_fill_1 FILLER_38_944 ();
 sg13g2_fill_1 FILLER_38_954 ();
 sg13g2_fill_1 FILLER_38_959 ();
 sg13g2_decap_4 FILLER_38_988 ();
 sg13g2_fill_2 FILLER_38_992 ();
 sg13g2_fill_2 FILLER_38_998 ();
 sg13g2_fill_2 FILLER_38_1010 ();
 sg13g2_decap_8 FILLER_38_1030 ();
 sg13g2_decap_8 FILLER_38_1037 ();
 sg13g2_decap_8 FILLER_38_1044 ();
 sg13g2_fill_2 FILLER_38_1051 ();
 sg13g2_fill_1 FILLER_38_1057 ();
 sg13g2_fill_2 FILLER_38_1118 ();
 sg13g2_decap_8 FILLER_38_1130 ();
 sg13g2_fill_1 FILLER_38_1137 ();
 sg13g2_fill_2 FILLER_38_1142 ();
 sg13g2_fill_1 FILLER_38_1155 ();
 sg13g2_fill_2 FILLER_38_1176 ();
 sg13g2_fill_2 FILLER_38_1186 ();
 sg13g2_fill_2 FILLER_38_1196 ();
 sg13g2_fill_1 FILLER_38_1212 ();
 sg13g2_fill_1 FILLER_38_1245 ();
 sg13g2_fill_2 FILLER_38_1251 ();
 sg13g2_fill_1 FILLER_38_1262 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1304 ();
 sg13g2_decap_8 FILLER_38_1311 ();
 sg13g2_fill_1 FILLER_38_1346 ();
 sg13g2_decap_4 FILLER_38_1377 ();
 sg13g2_fill_1 FILLER_38_1385 ();
 sg13g2_fill_2 FILLER_38_1412 ();
 sg13g2_decap_8 FILLER_38_1419 ();
 sg13g2_fill_2 FILLER_38_1426 ();
 sg13g2_fill_1 FILLER_38_1428 ();
 sg13g2_decap_8 FILLER_38_1437 ();
 sg13g2_decap_8 FILLER_38_1444 ();
 sg13g2_decap_8 FILLER_38_1451 ();
 sg13g2_fill_1 FILLER_38_1458 ();
 sg13g2_decap_4 FILLER_38_1463 ();
 sg13g2_fill_1 FILLER_38_1467 ();
 sg13g2_fill_1 FILLER_38_1472 ();
 sg13g2_fill_1 FILLER_38_1483 ();
 sg13g2_decap_4 FILLER_38_1527 ();
 sg13g2_decap_8 FILLER_38_1535 ();
 sg13g2_fill_2 FILLER_38_1542 ();
 sg13g2_decap_4 FILLER_38_1574 ();
 sg13g2_fill_1 FILLER_38_1578 ();
 sg13g2_fill_2 FILLER_38_1622 ();
 sg13g2_fill_1 FILLER_38_1640 ();
 sg13g2_fill_1 FILLER_38_1645 ();
 sg13g2_fill_1 FILLER_38_1693 ();
 sg13g2_fill_2 FILLER_38_1707 ();
 sg13g2_fill_2 FILLER_38_1724 ();
 sg13g2_fill_1 FILLER_38_1797 ();
 sg13g2_decap_8 FILLER_38_1844 ();
 sg13g2_decap_8 FILLER_38_1851 ();
 sg13g2_decap_8 FILLER_38_1858 ();
 sg13g2_decap_4 FILLER_38_1865 ();
 sg13g2_fill_2 FILLER_38_1869 ();
 sg13g2_fill_2 FILLER_38_1897 ();
 sg13g2_fill_1 FILLER_38_1899 ();
 sg13g2_fill_1 FILLER_38_1929 ();
 sg13g2_decap_4 FILLER_38_2020 ();
 sg13g2_fill_1 FILLER_38_2024 ();
 sg13g2_fill_1 FILLER_38_2035 ();
 sg13g2_fill_1 FILLER_38_2041 ();
 sg13g2_fill_2 FILLER_38_2146 ();
 sg13g2_fill_1 FILLER_38_2148 ();
 sg13g2_decap_8 FILLER_38_2196 ();
 sg13g2_decap_4 FILLER_38_2203 ();
 sg13g2_fill_2 FILLER_38_2211 ();
 sg13g2_fill_1 FILLER_38_2213 ();
 sg13g2_decap_8 FILLER_38_2224 ();
 sg13g2_decap_8 FILLER_38_2252 ();
 sg13g2_decap_8 FILLER_38_2259 ();
 sg13g2_fill_2 FILLER_38_2266 ();
 sg13g2_decap_8 FILLER_38_2293 ();
 sg13g2_decap_8 FILLER_38_2300 ();
 sg13g2_decap_4 FILLER_38_2307 ();
 sg13g2_fill_1 FILLER_38_2311 ();
 sg13g2_decap_4 FILLER_38_2338 ();
 sg13g2_fill_1 FILLER_38_2342 ();
 sg13g2_decap_8 FILLER_38_2347 ();
 sg13g2_decap_4 FILLER_38_2354 ();
 sg13g2_decap_4 FILLER_38_2362 ();
 sg13g2_fill_2 FILLER_38_2366 ();
 sg13g2_decap_8 FILLER_38_2410 ();
 sg13g2_fill_2 FILLER_38_2417 ();
 sg13g2_decap_8 FILLER_38_2424 ();
 sg13g2_decap_8 FILLER_38_2431 ();
 sg13g2_decap_8 FILLER_38_2438 ();
 sg13g2_decap_8 FILLER_38_2445 ();
 sg13g2_decap_8 FILLER_38_2452 ();
 sg13g2_fill_2 FILLER_38_2459 ();
 sg13g2_decap_4 FILLER_38_2487 ();
 sg13g2_decap_8 FILLER_38_2512 ();
 sg13g2_fill_1 FILLER_38_2519 ();
 sg13g2_fill_2 FILLER_38_2523 ();
 sg13g2_fill_2 FILLER_38_2549 ();
 sg13g2_decap_8 FILLER_38_2555 ();
 sg13g2_fill_2 FILLER_38_2562 ();
 sg13g2_decap_8 FILLER_38_2574 ();
 sg13g2_fill_2 FILLER_38_2581 ();
 sg13g2_fill_1 FILLER_38_2583 ();
 sg13g2_fill_2 FILLER_38_2611 ();
 sg13g2_decap_4 FILLER_38_2623 ();
 sg13g2_decap_8 FILLER_38_2653 ();
 sg13g2_decap_8 FILLER_38_2660 ();
 sg13g2_fill_2 FILLER_38_2667 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_24 ();
 sg13g2_decap_8 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_44 ();
 sg13g2_fill_1 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_174 ();
 sg13g2_decap_4 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_185 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_decap_4 FILLER_39_196 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_decap_4 FILLER_39_306 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_fill_2 FILLER_39_414 ();
 sg13g2_fill_2 FILLER_39_485 ();
 sg13g2_fill_1 FILLER_39_519 ();
 sg13g2_fill_2 FILLER_39_568 ();
 sg13g2_fill_1 FILLER_39_585 ();
 sg13g2_fill_2 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_fill_2 FILLER_39_735 ();
 sg13g2_fill_2 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_818 ();
 sg13g2_decap_4 FILLER_39_825 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_1 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_39_884 ();
 sg13g2_fill_1 FILLER_39_886 ();
 sg13g2_fill_1 FILLER_39_894 ();
 sg13g2_fill_2 FILLER_39_905 ();
 sg13g2_fill_1 FILLER_39_934 ();
 sg13g2_fill_1 FILLER_39_943 ();
 sg13g2_fill_1 FILLER_39_949 ();
 sg13g2_fill_1 FILLER_39_982 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_fill_1 FILLER_39_1001 ();
 sg13g2_fill_2 FILLER_39_1029 ();
 sg13g2_decap_8 FILLER_39_1035 ();
 sg13g2_decap_4 FILLER_39_1042 ();
 sg13g2_fill_1 FILLER_39_1053 ();
 sg13g2_fill_2 FILLER_39_1059 ();
 sg13g2_fill_1 FILLER_39_1079 ();
 sg13g2_decap_4 FILLER_39_1086 ();
 sg13g2_fill_1 FILLER_39_1116 ();
 sg13g2_decap_8 FILLER_39_1121 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_4 FILLER_39_1135 ();
 sg13g2_fill_1 FILLER_39_1139 ();
 sg13g2_fill_2 FILLER_39_1148 ();
 sg13g2_fill_1 FILLER_39_1153 ();
 sg13g2_fill_1 FILLER_39_1177 ();
 sg13g2_fill_1 FILLER_39_1201 ();
 sg13g2_fill_2 FILLER_39_1212 ();
 sg13g2_fill_2 FILLER_39_1231 ();
 sg13g2_fill_1 FILLER_39_1233 ();
 sg13g2_fill_2 FILLER_39_1238 ();
 sg13g2_fill_1 FILLER_39_1267 ();
 sg13g2_fill_2 FILLER_39_1273 ();
 sg13g2_decap_8 FILLER_39_1295 ();
 sg13g2_decap_8 FILLER_39_1302 ();
 sg13g2_decap_8 FILLER_39_1309 ();
 sg13g2_decap_4 FILLER_39_1316 ();
 sg13g2_fill_1 FILLER_39_1320 ();
 sg13g2_decap_4 FILLER_39_1351 ();
 sg13g2_fill_2 FILLER_39_1359 ();
 sg13g2_fill_1 FILLER_39_1361 ();
 sg13g2_fill_2 FILLER_39_1424 ();
 sg13g2_fill_2 FILLER_39_1465 ();
 sg13g2_fill_2 FILLER_39_1472 ();
 sg13g2_fill_2 FILLER_39_1478 ();
 sg13g2_decap_4 FILLER_39_1485 ();
 sg13g2_fill_2 FILLER_39_1489 ();
 sg13g2_decap_8 FILLER_39_1530 ();
 sg13g2_fill_2 FILLER_39_1537 ();
 sg13g2_fill_1 FILLER_39_1539 ();
 sg13g2_fill_2 FILLER_39_1579 ();
 sg13g2_decap_8 FILLER_39_1598 ();
 sg13g2_decap_8 FILLER_39_1605 ();
 sg13g2_decap_4 FILLER_39_1612 ();
 sg13g2_fill_1 FILLER_39_1647 ();
 sg13g2_fill_2 FILLER_39_1777 ();
 sg13g2_fill_2 FILLER_39_1805 ();
 sg13g2_decap_8 FILLER_39_1843 ();
 sg13g2_decap_4 FILLER_39_1850 ();
 sg13g2_decap_8 FILLER_39_1858 ();
 sg13g2_fill_1 FILLER_39_1931 ();
 sg13g2_fill_2 FILLER_39_1968 ();
 sg13g2_fill_1 FILLER_39_1995 ();
 sg13g2_fill_2 FILLER_39_2022 ();
 sg13g2_fill_1 FILLER_39_2024 ();
 sg13g2_decap_4 FILLER_39_2035 ();
 sg13g2_fill_2 FILLER_39_2039 ();
 sg13g2_fill_2 FILLER_39_2080 ();
 sg13g2_fill_1 FILLER_39_2112 ();
 sg13g2_fill_2 FILLER_39_2173 ();
 sg13g2_decap_4 FILLER_39_2201 ();
 sg13g2_fill_1 FILLER_39_2205 ();
 sg13g2_fill_2 FILLER_39_2232 ();
 sg13g2_fill_1 FILLER_39_2234 ();
 sg13g2_fill_2 FILLER_39_2280 ();
 sg13g2_decap_4 FILLER_39_2312 ();
 sg13g2_fill_1 FILLER_39_2316 ();
 sg13g2_fill_2 FILLER_39_2331 ();
 sg13g2_fill_1 FILLER_39_2333 ();
 sg13g2_fill_2 FILLER_39_2355 ();
 sg13g2_fill_1 FILLER_39_2357 ();
 sg13g2_decap_8 FILLER_39_2443 ();
 sg13g2_fill_2 FILLER_39_2450 ();
 sg13g2_fill_1 FILLER_39_2462 ();
 sg13g2_decap_8 FILLER_39_2489 ();
 sg13g2_fill_2 FILLER_39_2496 ();
 sg13g2_fill_2 FILLER_39_2541 ();
 sg13g2_decap_8 FILLER_39_2595 ();
 sg13g2_decap_4 FILLER_39_2602 ();
 sg13g2_fill_2 FILLER_39_2606 ();
 sg13g2_decap_8 FILLER_39_2612 ();
 sg13g2_decap_8 FILLER_39_2619 ();
 sg13g2_decap_8 FILLER_39_2626 ();
 sg13g2_fill_2 FILLER_39_2633 ();
 sg13g2_decap_8 FILLER_39_2639 ();
 sg13g2_decap_8 FILLER_39_2646 ();
 sg13g2_decap_8 FILLER_39_2653 ();
 sg13g2_decap_8 FILLER_39_2660 ();
 sg13g2_fill_2 FILLER_39_2667 ();
 sg13g2_fill_1 FILLER_39_2669 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_11 ();
 sg13g2_decap_4 FILLER_40_16 ();
 sg13g2_fill_1 FILLER_40_20 ();
 sg13g2_decap_4 FILLER_40_33 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_77 ();
 sg13g2_fill_2 FILLER_40_86 ();
 sg13g2_fill_1 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_97 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_134 ();
 sg13g2_fill_1 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_179 ();
 sg13g2_decap_8 FILLER_40_185 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_230 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_decap_4 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_fill_2 FILLER_40_295 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_fill_1 FILLER_40_351 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_454 ();
 sg13g2_fill_1 FILLER_40_525 ();
 sg13g2_fill_2 FILLER_40_552 ();
 sg13g2_fill_2 FILLER_40_566 ();
 sg13g2_fill_2 FILLER_40_573 ();
 sg13g2_decap_8 FILLER_40_584 ();
 sg13g2_decap_8 FILLER_40_591 ();
 sg13g2_decap_8 FILLER_40_598 ();
 sg13g2_fill_1 FILLER_40_605 ();
 sg13g2_decap_4 FILLER_40_614 ();
 sg13g2_decap_8 FILLER_40_622 ();
 sg13g2_decap_8 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_636 ();
 sg13g2_decap_4 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_652 ();
 sg13g2_fill_2 FILLER_40_688 ();
 sg13g2_decap_4 FILLER_40_730 ();
 sg13g2_fill_1 FILLER_40_734 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_fill_1 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_fill_2 FILLER_40_859 ();
 sg13g2_fill_1 FILLER_40_921 ();
 sg13g2_fill_1 FILLER_40_927 ();
 sg13g2_fill_1 FILLER_40_935 ();
 sg13g2_fill_1 FILLER_40_940 ();
 sg13g2_fill_2 FILLER_40_982 ();
 sg13g2_fill_1 FILLER_40_993 ();
 sg13g2_fill_2 FILLER_40_999 ();
 sg13g2_fill_1 FILLER_40_1008 ();
 sg13g2_fill_2 FILLER_40_1014 ();
 sg13g2_fill_1 FILLER_40_1016 ();
 sg13g2_fill_2 FILLER_40_1021 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_fill_2 FILLER_40_1037 ();
 sg13g2_fill_1 FILLER_40_1043 ();
 sg13g2_fill_2 FILLER_40_1049 ();
 sg13g2_fill_1 FILLER_40_1074 ();
 sg13g2_decap_8 FILLER_40_1080 ();
 sg13g2_fill_2 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1089 ();
 sg13g2_fill_2 FILLER_40_1094 ();
 sg13g2_fill_2 FILLER_40_1100 ();
 sg13g2_fill_2 FILLER_40_1107 ();
 sg13g2_fill_1 FILLER_40_1127 ();
 sg13g2_fill_2 FILLER_40_1160 ();
 sg13g2_fill_1 FILLER_40_1167 ();
 sg13g2_fill_1 FILLER_40_1185 ();
 sg13g2_decap_8 FILLER_40_1231 ();
 sg13g2_decap_8 FILLER_40_1238 ();
 sg13g2_decap_4 FILLER_40_1245 ();
 sg13g2_fill_2 FILLER_40_1257 ();
 sg13g2_fill_1 FILLER_40_1259 ();
 sg13g2_fill_1 FILLER_40_1287 ();
 sg13g2_fill_1 FILLER_40_1293 ();
 sg13g2_fill_2 FILLER_40_1332 ();
 sg13g2_decap_8 FILLER_40_1360 ();
 sg13g2_decap_8 FILLER_40_1367 ();
 sg13g2_decap_8 FILLER_40_1374 ();
 sg13g2_decap_4 FILLER_40_1381 ();
 sg13g2_decap_8 FILLER_40_1399 ();
 sg13g2_fill_1 FILLER_40_1406 ();
 sg13g2_decap_4 FILLER_40_1411 ();
 sg13g2_fill_2 FILLER_40_1415 ();
 sg13g2_fill_1 FILLER_40_1448 ();
 sg13g2_decap_8 FILLER_40_1459 ();
 sg13g2_decap_8 FILLER_40_1466 ();
 sg13g2_fill_2 FILLER_40_1473 ();
 sg13g2_fill_2 FILLER_40_1483 ();
 sg13g2_decap_8 FILLER_40_1511 ();
 sg13g2_decap_8 FILLER_40_1518 ();
 sg13g2_decap_8 FILLER_40_1525 ();
 sg13g2_fill_2 FILLER_40_1543 ();
 sg13g2_fill_1 FILLER_40_1545 ();
 sg13g2_fill_1 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1556 ();
 sg13g2_decap_8 FILLER_40_1563 ();
 sg13g2_fill_2 FILLER_40_1570 ();
 sg13g2_fill_2 FILLER_40_1602 ();
 sg13g2_fill_1 FILLER_40_1604 ();
 sg13g2_decap_4 FILLER_40_1609 ();
 sg13g2_fill_1 FILLER_40_1622 ();
 sg13g2_fill_1 FILLER_40_1649 ();
 sg13g2_fill_2 FILLER_40_1659 ();
 sg13g2_fill_1 FILLER_40_1661 ();
 sg13g2_fill_1 FILLER_40_1666 ();
 sg13g2_fill_1 FILLER_40_1671 ();
 sg13g2_fill_2 FILLER_40_1676 ();
 sg13g2_fill_1 FILLER_40_1823 ();
 sg13g2_fill_1 FILLER_40_1828 ();
 sg13g2_fill_1 FILLER_40_1833 ();
 sg13g2_fill_1 FILLER_40_1844 ();
 sg13g2_fill_2 FILLER_40_1893 ();
 sg13g2_decap_4 FILLER_40_1920 ();
 sg13g2_fill_1 FILLER_40_1950 ();
 sg13g2_fill_2 FILLER_40_1954 ();
 sg13g2_fill_1 FILLER_40_2006 ();
 sg13g2_fill_2 FILLER_40_2021 ();
 sg13g2_fill_1 FILLER_40_2028 ();
 sg13g2_fill_1 FILLER_40_2037 ();
 sg13g2_fill_2 FILLER_40_2048 ();
 sg13g2_fill_1 FILLER_40_2050 ();
 sg13g2_fill_1 FILLER_40_2060 ();
 sg13g2_fill_1 FILLER_40_2075 ();
 sg13g2_fill_1 FILLER_40_2081 ();
 sg13g2_decap_4 FILLER_40_2139 ();
 sg13g2_fill_2 FILLER_40_2153 ();
 sg13g2_fill_1 FILLER_40_2155 ();
 sg13g2_decap_8 FILLER_40_2192 ();
 sg13g2_decap_4 FILLER_40_2199 ();
 sg13g2_fill_2 FILLER_40_2207 ();
 sg13g2_fill_2 FILLER_40_2235 ();
 sg13g2_fill_1 FILLER_40_2237 ();
 sg13g2_decap_4 FILLER_40_2268 ();
 sg13g2_fill_1 FILLER_40_2272 ();
 sg13g2_decap_8 FILLER_40_2313 ();
 sg13g2_decap_8 FILLER_40_2320 ();
 sg13g2_fill_1 FILLER_40_2345 ();
 sg13g2_decap_8 FILLER_40_2350 ();
 sg13g2_fill_2 FILLER_40_2374 ();
 sg13g2_fill_1 FILLER_40_2406 ();
 sg13g2_fill_1 FILLER_40_2433 ();
 sg13g2_fill_1 FILLER_40_2455 ();
 sg13g2_fill_1 FILLER_40_2466 ();
 sg13g2_fill_2 FILLER_40_2479 ();
 sg13g2_fill_2 FILLER_40_2558 ();
 sg13g2_decap_8 FILLER_40_2564 ();
 sg13g2_decap_4 FILLER_40_2571 ();
 sg13g2_fill_1 FILLER_40_2575 ();
 sg13g2_decap_8 FILLER_40_2610 ();
 sg13g2_decap_8 FILLER_40_2627 ();
 sg13g2_decap_8 FILLER_40_2634 ();
 sg13g2_decap_8 FILLER_40_2641 ();
 sg13g2_decap_8 FILLER_40_2648 ();
 sg13g2_decap_8 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2662 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_fill_2 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_89 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_fill_2 FILLER_41_205 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_232 ();
 sg13g2_fill_1 FILLER_41_237 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_311 ();
 sg13g2_fill_2 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_323 ();
 sg13g2_fill_1 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_1 FILLER_41_379 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_fill_1 FILLER_41_506 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_521 ();
 sg13g2_decap_4 FILLER_41_526 ();
 sg13g2_fill_1 FILLER_41_530 ();
 sg13g2_fill_2 FILLER_41_535 ();
 sg13g2_decap_4 FILLER_41_541 ();
 sg13g2_fill_1 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_569 ();
 sg13g2_decap_8 FILLER_41_582 ();
 sg13g2_decap_8 FILLER_41_589 ();
 sg13g2_decap_4 FILLER_41_596 ();
 sg13g2_fill_2 FILLER_41_600 ();
 sg13g2_decap_8 FILLER_41_606 ();
 sg13g2_decap_8 FILLER_41_613 ();
 sg13g2_decap_4 FILLER_41_624 ();
 sg13g2_fill_2 FILLER_41_628 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_fill_1 FILLER_41_652 ();
 sg13g2_decap_4 FILLER_41_658 ();
 sg13g2_fill_2 FILLER_41_692 ();
 sg13g2_decap_4 FILLER_41_705 ();
 sg13g2_fill_2 FILLER_41_709 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_4 FILLER_41_721 ();
 sg13g2_fill_1 FILLER_41_725 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_decap_4 FILLER_41_745 ();
 sg13g2_fill_2 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_755 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_decap_8 FILLER_41_767 ();
 sg13g2_decap_8 FILLER_41_774 ();
 sg13g2_decap_8 FILLER_41_781 ();
 sg13g2_fill_2 FILLER_41_788 ();
 sg13g2_fill_1 FILLER_41_799 ();
 sg13g2_decap_4 FILLER_41_804 ();
 sg13g2_fill_1 FILLER_41_813 ();
 sg13g2_fill_2 FILLER_41_829 ();
 sg13g2_fill_1 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_841 ();
 sg13g2_decap_8 FILLER_41_848 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_decap_4 FILLER_41_862 ();
 sg13g2_fill_2 FILLER_41_878 ();
 sg13g2_fill_1 FILLER_41_880 ();
 sg13g2_fill_1 FILLER_41_886 ();
 sg13g2_fill_1 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_897 ();
 sg13g2_fill_1 FILLER_41_904 ();
 sg13g2_decap_4 FILLER_41_931 ();
 sg13g2_fill_1 FILLER_41_935 ();
 sg13g2_fill_1 FILLER_41_971 ();
 sg13g2_fill_1 FILLER_41_976 ();
 sg13g2_fill_1 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_985 ();
 sg13g2_fill_1 FILLER_41_992 ();
 sg13g2_decap_8 FILLER_41_998 ();
 sg13g2_fill_2 FILLER_41_1005 ();
 sg13g2_fill_1 FILLER_41_1007 ();
 sg13g2_fill_1 FILLER_41_1017 ();
 sg13g2_fill_1 FILLER_41_1040 ();
 sg13g2_fill_2 FILLER_41_1075 ();
 sg13g2_fill_1 FILLER_41_1110 ();
 sg13g2_fill_1 FILLER_41_1125 ();
 sg13g2_fill_1 FILLER_41_1143 ();
 sg13g2_fill_2 FILLER_41_1165 ();
 sg13g2_fill_1 FILLER_41_1172 ();
 sg13g2_fill_2 FILLER_41_1189 ();
 sg13g2_decap_8 FILLER_41_1244 ();
 sg13g2_decap_4 FILLER_41_1251 ();
 sg13g2_fill_1 FILLER_41_1255 ();
 sg13g2_fill_2 FILLER_41_1282 ();
 sg13g2_fill_1 FILLER_41_1294 ();
 sg13g2_fill_1 FILLER_41_1321 ();
 sg13g2_fill_1 FILLER_41_1346 ();
 sg13g2_decap_8 FILLER_41_1386 ();
 sg13g2_decap_8 FILLER_41_1393 ();
 sg13g2_decap_4 FILLER_41_1400 ();
 sg13g2_fill_2 FILLER_41_1404 ();
 sg13g2_decap_4 FILLER_41_1445 ();
 sg13g2_decap_8 FILLER_41_1455 ();
 sg13g2_decap_4 FILLER_41_1462 ();
 sg13g2_decap_4 FILLER_41_1500 ();
 sg13g2_fill_2 FILLER_41_1504 ();
 sg13g2_fill_2 FILLER_41_1545 ();
 sg13g2_fill_1 FILLER_41_1547 ();
 sg13g2_decap_8 FILLER_41_1558 ();
 sg13g2_fill_2 FILLER_41_1565 ();
 sg13g2_fill_1 FILLER_41_1567 ();
 sg13g2_fill_2 FILLER_41_1607 ();
 sg13g2_fill_1 FILLER_41_1609 ();
 sg13g2_fill_2 FILLER_41_1650 ();
 sg13g2_fill_1 FILLER_41_1676 ();
 sg13g2_fill_2 FILLER_41_1717 ();
 sg13g2_fill_1 FILLER_41_1744 ();
 sg13g2_fill_2 FILLER_41_1751 ();
 sg13g2_fill_2 FILLER_41_1761 ();
 sg13g2_fill_2 FILLER_41_1837 ();
 sg13g2_fill_1 FILLER_41_1839 ();
 sg13g2_decap_8 FILLER_41_1854 ();
 sg13g2_decap_4 FILLER_41_1861 ();
 sg13g2_decap_4 FILLER_41_1874 ();
 sg13g2_decap_8 FILLER_41_1904 ();
 sg13g2_fill_1 FILLER_41_1911 ();
 sg13g2_decap_4 FILLER_41_1916 ();
 sg13g2_fill_2 FILLER_41_1930 ();
 sg13g2_fill_2 FILLER_41_1941 ();
 sg13g2_fill_2 FILLER_41_1960 ();
 sg13g2_fill_1 FILLER_41_1972 ();
 sg13g2_decap_8 FILLER_41_2010 ();
 sg13g2_decap_8 FILLER_41_2017 ();
 sg13g2_fill_1 FILLER_41_2024 ();
 sg13g2_fill_2 FILLER_41_2047 ();
 sg13g2_fill_1 FILLER_41_2059 ();
 sg13g2_decap_4 FILLER_41_2106 ();
 sg13g2_fill_1 FILLER_41_2120 ();
 sg13g2_decap_4 FILLER_41_2142 ();
 sg13g2_fill_1 FILLER_41_2146 ();
 sg13g2_decap_8 FILLER_41_2157 ();
 sg13g2_decap_8 FILLER_41_2164 ();
 sg13g2_fill_2 FILLER_41_2171 ();
 sg13g2_fill_1 FILLER_41_2173 ();
 sg13g2_decap_4 FILLER_41_2178 ();
 sg13g2_fill_2 FILLER_41_2182 ();
 sg13g2_decap_8 FILLER_41_2188 ();
 sg13g2_fill_2 FILLER_41_2195 ();
 sg13g2_decap_4 FILLER_41_2201 ();
 sg13g2_fill_2 FILLER_41_2205 ();
 sg13g2_decap_4 FILLER_41_2259 ();
 sg13g2_fill_1 FILLER_41_2263 ();
 sg13g2_fill_1 FILLER_41_2274 ();
 sg13g2_fill_1 FILLER_41_2301 ();
 sg13g2_fill_2 FILLER_41_2332 ();
 sg13g2_fill_1 FILLER_41_2334 ();
 sg13g2_fill_2 FILLER_41_2361 ();
 sg13g2_decap_4 FILLER_41_2379 ();
 sg13g2_fill_2 FILLER_41_2422 ();
 sg13g2_fill_2 FILLER_41_2464 ();
 sg13g2_decap_4 FILLER_41_2474 ();
 sg13g2_decap_8 FILLER_41_2488 ();
 sg13g2_fill_2 FILLER_41_2495 ();
 sg13g2_fill_1 FILLER_41_2497 ();
 sg13g2_decap_8 FILLER_41_2523 ();
 sg13g2_decap_4 FILLER_41_2530 ();
 sg13g2_fill_1 FILLER_41_2534 ();
 sg13g2_fill_2 FILLER_41_2585 ();
 sg13g2_fill_1 FILLER_41_2587 ();
 sg13g2_fill_1 FILLER_41_2609 ();
 sg13g2_decap_8 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2653 ();
 sg13g2_decap_8 FILLER_41_2660 ();
 sg13g2_fill_2 FILLER_41_2667 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_43 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_55 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_fill_2 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_105 ();
 sg13g2_decap_4 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_158 ();
 sg13g2_fill_2 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_decap_4 FILLER_42_226 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_decap_4 FILLER_42_258 ();
 sg13g2_fill_2 FILLER_42_262 ();
 sg13g2_decap_4 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_272 ();
 sg13g2_fill_1 FILLER_42_316 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_fill_1 FILLER_42_348 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_372 ();
 sg13g2_fill_1 FILLER_42_379 ();
 sg13g2_fill_2 FILLER_42_392 ();
 sg13g2_fill_1 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_2 FILLER_42_424 ();
 sg13g2_fill_1 FILLER_42_426 ();
 sg13g2_decap_4 FILLER_42_434 ();
 sg13g2_fill_2 FILLER_42_449 ();
 sg13g2_fill_1 FILLER_42_459 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_518 ();
 sg13g2_decap_4 FILLER_42_536 ();
 sg13g2_decap_8 FILLER_42_544 ();
 sg13g2_fill_1 FILLER_42_551 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_fill_1 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_591 ();
 sg13g2_decap_8 FILLER_42_598 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_fill_2 FILLER_42_616 ();
 sg13g2_fill_1 FILLER_42_618 ();
 sg13g2_decap_4 FILLER_42_629 ();
 sg13g2_fill_2 FILLER_42_661 ();
 sg13g2_decap_8 FILLER_42_667 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_fill_2 FILLER_42_740 ();
 sg13g2_fill_1 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_4 FILLER_42_784 ();
 sg13g2_decap_4 FILLER_42_844 ();
 sg13g2_fill_1 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_fill_1 FILLER_42_863 ();
 sg13g2_fill_1 FILLER_42_869 ();
 sg13g2_fill_2 FILLER_42_900 ();
 sg13g2_fill_1 FILLER_42_902 ();
 sg13g2_fill_2 FILLER_42_917 ();
 sg13g2_decap_4 FILLER_42_923 ();
 sg13g2_fill_1 FILLER_42_927 ();
 sg13g2_fill_2 FILLER_42_938 ();
 sg13g2_fill_1 FILLER_42_974 ();
 sg13g2_decap_4 FILLER_42_980 ();
 sg13g2_fill_1 FILLER_42_984 ();
 sg13g2_decap_4 FILLER_42_989 ();
 sg13g2_fill_1 FILLER_42_993 ();
 sg13g2_fill_1 FILLER_42_999 ();
 sg13g2_decap_4 FILLER_42_1004 ();
 sg13g2_decap_4 FILLER_42_1016 ();
 sg13g2_decap_4 FILLER_42_1037 ();
 sg13g2_fill_1 FILLER_42_1041 ();
 sg13g2_decap_4 FILLER_42_1059 ();
 sg13g2_fill_2 FILLER_42_1063 ();
 sg13g2_fill_1 FILLER_42_1069 ();
 sg13g2_fill_2 FILLER_42_1080 ();
 sg13g2_fill_2 FILLER_42_1087 ();
 sg13g2_fill_1 FILLER_42_1100 ();
 sg13g2_fill_1 FILLER_42_1118 ();
 sg13g2_fill_1 FILLER_42_1127 ();
 sg13g2_fill_2 FILLER_42_1135 ();
 sg13g2_fill_1 FILLER_42_1159 ();
 sg13g2_fill_1 FILLER_42_1185 ();
 sg13g2_fill_1 FILLER_42_1193 ();
 sg13g2_fill_2 FILLER_42_1207 ();
 sg13g2_fill_1 FILLER_42_1217 ();
 sg13g2_fill_2 FILLER_42_1228 ();
 sg13g2_decap_8 FILLER_42_1239 ();
 sg13g2_fill_1 FILLER_42_1283 ();
 sg13g2_fill_2 FILLER_42_1289 ();
 sg13g2_fill_1 FILLER_42_1291 ();
 sg13g2_fill_2 FILLER_42_1306 ();
 sg13g2_decap_4 FILLER_42_1330 ();
 sg13g2_decap_8 FILLER_42_1339 ();
 sg13g2_fill_1 FILLER_42_1346 ();
 sg13g2_fill_1 FILLER_42_1354 ();
 sg13g2_decap_8 FILLER_42_1359 ();
 sg13g2_decap_8 FILLER_42_1396 ();
 sg13g2_decap_4 FILLER_42_1403 ();
 sg13g2_fill_1 FILLER_42_1437 ();
 sg13g2_fill_2 FILLER_42_1469 ();
 sg13g2_fill_1 FILLER_42_1471 ();
 sg13g2_fill_2 FILLER_42_1495 ();
 sg13g2_fill_2 FILLER_42_1518 ();
 sg13g2_fill_2 FILLER_42_1537 ();
 sg13g2_decap_8 FILLER_42_1570 ();
 sg13g2_decap_8 FILLER_42_1577 ();
 sg13g2_fill_1 FILLER_42_1584 ();
 sg13g2_fill_2 FILLER_42_1604 ();
 sg13g2_decap_8 FILLER_42_1636 ();
 sg13g2_fill_1 FILLER_42_1643 ();
 sg13g2_fill_2 FILLER_42_1674 ();
 sg13g2_fill_1 FILLER_42_1685 ();
 sg13g2_fill_2 FILLER_42_1703 ();
 sg13g2_fill_1 FILLER_42_1734 ();
 sg13g2_fill_1 FILLER_42_1745 ();
 sg13g2_fill_1 FILLER_42_1804 ();
 sg13g2_decap_8 FILLER_42_1831 ();
 sg13g2_fill_1 FILLER_42_1838 ();
 sg13g2_fill_1 FILLER_42_1869 ();
 sg13g2_fill_2 FILLER_42_1880 ();
 sg13g2_fill_1 FILLER_42_1882 ();
 sg13g2_decap_8 FILLER_42_1909 ();
 sg13g2_fill_1 FILLER_42_1916 ();
 sg13g2_fill_1 FILLER_42_1926 ();
 sg13g2_fill_2 FILLER_42_1931 ();
 sg13g2_fill_2 FILLER_42_1942 ();
 sg13g2_fill_1 FILLER_42_1944 ();
 sg13g2_fill_2 FILLER_42_2009 ();
 sg13g2_decap_8 FILLER_42_2016 ();
 sg13g2_decap_4 FILLER_42_2023 ();
 sg13g2_fill_2 FILLER_42_2027 ();
 sg13g2_fill_2 FILLER_42_2052 ();
 sg13g2_fill_2 FILLER_42_2059 ();
 sg13g2_fill_2 FILLER_42_2084 ();
 sg13g2_fill_1 FILLER_42_2086 ();
 sg13g2_decap_4 FILLER_42_2131 ();
 sg13g2_fill_2 FILLER_42_2139 ();
 sg13g2_fill_1 FILLER_42_2141 ();
 sg13g2_fill_1 FILLER_42_2156 ();
 sg13g2_decap_8 FILLER_42_2183 ();
 sg13g2_decap_4 FILLER_42_2190 ();
 sg13g2_fill_2 FILLER_42_2194 ();
 sg13g2_fill_1 FILLER_42_2234 ();
 sg13g2_decap_8 FILLER_42_2262 ();
 sg13g2_decap_8 FILLER_42_2269 ();
 sg13g2_fill_1 FILLER_42_2276 ();
 sg13g2_fill_1 FILLER_42_2281 ();
 sg13g2_fill_1 FILLER_42_2296 ();
 sg13g2_decap_8 FILLER_42_2318 ();
 sg13g2_decap_8 FILLER_42_2325 ();
 sg13g2_fill_2 FILLER_42_2332 ();
 sg13g2_fill_1 FILLER_42_2334 ();
 sg13g2_fill_1 FILLER_42_2339 ();
 sg13g2_decap_8 FILLER_42_2344 ();
 sg13g2_decap_8 FILLER_42_2351 ();
 sg13g2_fill_1 FILLER_42_2358 ();
 sg13g2_decap_4 FILLER_42_2363 ();
 sg13g2_fill_2 FILLER_42_2367 ();
 sg13g2_fill_1 FILLER_42_2390 ();
 sg13g2_decap_4 FILLER_42_2396 ();
 sg13g2_fill_2 FILLER_42_2400 ();
 sg13g2_fill_2 FILLER_42_2406 ();
 sg13g2_decap_8 FILLER_42_2413 ();
 sg13g2_decap_8 FILLER_42_2420 ();
 sg13g2_fill_2 FILLER_42_2427 ();
 sg13g2_fill_2 FILLER_42_2439 ();
 sg13g2_fill_2 FILLER_42_2445 ();
 sg13g2_decap_8 FILLER_42_2451 ();
 sg13g2_decap_8 FILLER_42_2458 ();
 sg13g2_decap_8 FILLER_42_2465 ();
 sg13g2_decap_8 FILLER_42_2472 ();
 sg13g2_fill_2 FILLER_42_2479 ();
 sg13g2_fill_1 FILLER_42_2481 ();
 sg13g2_decap_4 FILLER_42_2518 ();
 sg13g2_fill_1 FILLER_42_2522 ();
 sg13g2_fill_1 FILLER_42_2532 ();
 sg13g2_decap_8 FILLER_42_2554 ();
 sg13g2_decap_4 FILLER_42_2561 ();
 sg13g2_fill_2 FILLER_42_2565 ();
 sg13g2_fill_2 FILLER_42_2624 ();
 sg13g2_decap_8 FILLER_42_2652 ();
 sg13g2_decap_8 FILLER_42_2659 ();
 sg13g2_decap_4 FILLER_42_2666 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_fill_2 FILLER_43_94 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_126 ();
 sg13g2_decap_4 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_175 ();
 sg13g2_fill_1 FILLER_43_177 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_fill_1 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_275 ();
 sg13g2_decap_4 FILLER_43_282 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_decap_4 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_304 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_decap_8 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_decap_8 FILLER_43_341 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_fill_2 FILLER_43_355 ();
 sg13g2_fill_1 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_fill_1 FILLER_43_489 ();
 sg13g2_fill_2 FILLER_43_496 ();
 sg13g2_fill_2 FILLER_43_522 ();
 sg13g2_fill_2 FILLER_43_559 ();
 sg13g2_fill_2 FILLER_43_584 ();
 sg13g2_decap_8 FILLER_43_591 ();
 sg13g2_fill_1 FILLER_43_598 ();
 sg13g2_decap_4 FILLER_43_603 ();
 sg13g2_fill_1 FILLER_43_612 ();
 sg13g2_decap_8 FILLER_43_635 ();
 sg13g2_fill_2 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_fill_1 FILLER_43_670 ();
 sg13g2_fill_1 FILLER_43_678 ();
 sg13g2_fill_2 FILLER_43_686 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_fill_2 FILLER_43_746 ();
 sg13g2_fill_2 FILLER_43_753 ();
 sg13g2_fill_1 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_4 FILLER_43_845 ();
 sg13g2_fill_2 FILLER_43_853 ();
 sg13g2_fill_1 FILLER_43_889 ();
 sg13g2_fill_1 FILLER_43_894 ();
 sg13g2_decap_4 FILLER_43_900 ();
 sg13g2_fill_2 FILLER_43_904 ();
 sg13g2_fill_2 FILLER_43_930 ();
 sg13g2_fill_1 FILLER_43_945 ();
 sg13g2_fill_1 FILLER_43_952 ();
 sg13g2_decap_4 FILLER_43_975 ();
 sg13g2_fill_2 FILLER_43_979 ();
 sg13g2_fill_1 FILLER_43_986 ();
 sg13g2_fill_1 FILLER_43_991 ();
 sg13g2_fill_2 FILLER_43_997 ();
 sg13g2_fill_1 FILLER_43_1007 ();
 sg13g2_fill_1 FILLER_43_1013 ();
 sg13g2_fill_2 FILLER_43_1034 ();
 sg13g2_fill_1 FILLER_43_1036 ();
 sg13g2_fill_1 FILLER_43_1062 ();
 sg13g2_fill_1 FILLER_43_1084 ();
 sg13g2_fill_1 FILLER_43_1106 ();
 sg13g2_fill_2 FILLER_43_1115 ();
 sg13g2_fill_1 FILLER_43_1157 ();
 sg13g2_fill_1 FILLER_43_1165 ();
 sg13g2_fill_1 FILLER_43_1181 ();
 sg13g2_fill_2 FILLER_43_1185 ();
 sg13g2_fill_2 FILLER_43_1192 ();
 sg13g2_fill_2 FILLER_43_1209 ();
 sg13g2_fill_2 FILLER_43_1217 ();
 sg13g2_fill_1 FILLER_43_1222 ();
 sg13g2_fill_1 FILLER_43_1229 ();
 sg13g2_fill_2 FILLER_43_1245 ();
 sg13g2_decap_4 FILLER_43_1251 ();
 sg13g2_fill_1 FILLER_43_1259 ();
 sg13g2_decap_4 FILLER_43_1263 ();
 sg13g2_fill_1 FILLER_43_1312 ();
 sg13g2_decap_8 FILLER_43_1339 ();
 sg13g2_fill_2 FILLER_43_1346 ();
 sg13g2_decap_8 FILLER_43_1373 ();
 sg13g2_decap_4 FILLER_43_1380 ();
 sg13g2_fill_1 FILLER_43_1384 ();
 sg13g2_decap_8 FILLER_43_1401 ();
 sg13g2_decap_4 FILLER_43_1408 ();
 sg13g2_fill_2 FILLER_43_1412 ();
 sg13g2_fill_1 FILLER_43_1423 ();
 sg13g2_fill_2 FILLER_43_1433 ();
 sg13g2_fill_1 FILLER_43_1435 ();
 sg13g2_decap_4 FILLER_43_1445 ();
 sg13g2_fill_1 FILLER_43_1449 ();
 sg13g2_fill_1 FILLER_43_1484 ();
 sg13g2_fill_1 FILLER_43_1501 ();
 sg13g2_fill_1 FILLER_43_1507 ();
 sg13g2_fill_1 FILLER_43_1512 ();
 sg13g2_fill_2 FILLER_43_1563 ();
 sg13g2_decap_4 FILLER_43_1569 ();
 sg13g2_decap_4 FILLER_43_1579 ();
 sg13g2_fill_2 FILLER_43_1583 ();
 sg13g2_fill_1 FILLER_43_1603 ();
 sg13g2_fill_2 FILLER_43_1609 ();
 sg13g2_decap_4 FILLER_43_1624 ();
 sg13g2_fill_1 FILLER_43_1628 ();
 sg13g2_decap_8 FILLER_43_1635 ();
 sg13g2_fill_2 FILLER_43_1642 ();
 sg13g2_fill_1 FILLER_43_1644 ();
 sg13g2_decap_8 FILLER_43_1655 ();
 sg13g2_decap_4 FILLER_43_1662 ();
 sg13g2_fill_2 FILLER_43_1720 ();
 sg13g2_fill_2 FILLER_43_1757 ();
 sg13g2_fill_1 FILLER_43_1790 ();
 sg13g2_fill_1 FILLER_43_1821 ();
 sg13g2_fill_2 FILLER_43_1832 ();
 sg13g2_decap_4 FILLER_43_1880 ();
 sg13g2_fill_1 FILLER_43_1888 ();
 sg13g2_fill_1 FILLER_43_1893 ();
 sg13g2_fill_2 FILLER_43_1941 ();
 sg13g2_fill_1 FILLER_43_1959 ();
 sg13g2_fill_2 FILLER_43_1968 ();
 sg13g2_decap_4 FILLER_43_1996 ();
 sg13g2_fill_2 FILLER_43_2000 ();
 sg13g2_decap_4 FILLER_43_2028 ();
 sg13g2_fill_1 FILLER_43_2032 ();
 sg13g2_decap_8 FILLER_43_2038 ();
 sg13g2_fill_1 FILLER_43_2045 ();
 sg13g2_fill_1 FILLER_43_2060 ();
 sg13g2_fill_1 FILLER_43_2073 ();
 sg13g2_fill_1 FILLER_43_2110 ();
 sg13g2_decap_8 FILLER_43_2142 ();
 sg13g2_decap_8 FILLER_43_2179 ();
 sg13g2_decap_8 FILLER_43_2186 ();
 sg13g2_fill_1 FILLER_43_2193 ();
 sg13g2_fill_2 FILLER_43_2234 ();
 sg13g2_decap_8 FILLER_43_2261 ();
 sg13g2_decap_8 FILLER_43_2268 ();
 sg13g2_decap_8 FILLER_43_2275 ();
 sg13g2_decap_8 FILLER_43_2282 ();
 sg13g2_decap_8 FILLER_43_2289 ();
 sg13g2_fill_2 FILLER_43_2296 ();
 sg13g2_decap_8 FILLER_43_2308 ();
 sg13g2_decap_4 FILLER_43_2315 ();
 sg13g2_fill_2 FILLER_43_2319 ();
 sg13g2_decap_8 FILLER_43_2408 ();
 sg13g2_decap_8 FILLER_43_2415 ();
 sg13g2_fill_2 FILLER_43_2422 ();
 sg13g2_fill_2 FILLER_43_2437 ();
 sg13g2_fill_1 FILLER_43_2439 ();
 sg13g2_decap_8 FILLER_43_2470 ();
 sg13g2_decap_4 FILLER_43_2487 ();
 sg13g2_decap_8 FILLER_43_2562 ();
 sg13g2_fill_2 FILLER_43_2569 ();
 sg13g2_decap_4 FILLER_43_2581 ();
 sg13g2_decap_8 FILLER_43_2657 ();
 sg13g2_decap_4 FILLER_43_2664 ();
 sg13g2_fill_2 FILLER_43_2668 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_9 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_64 ();
 sg13g2_fill_1 FILLER_44_87 ();
 sg13g2_fill_1 FILLER_44_97 ();
 sg13g2_fill_2 FILLER_44_129 ();
 sg13g2_fill_2 FILLER_44_137 ();
 sg13g2_fill_1 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_159 ();
 sg13g2_decap_8 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_181 ();
 sg13g2_fill_2 FILLER_44_192 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_decap_8 FILLER_44_233 ();
 sg13g2_decap_4 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_258 ();
 sg13g2_decap_8 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_fill_2 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_fill_1 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_fill_1 FILLER_44_470 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_fill_1 FILLER_44_509 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_fill_2 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_611 ();
 sg13g2_fill_1 FILLER_44_621 ();
 sg13g2_fill_1 FILLER_44_626 ();
 sg13g2_decap_8 FILLER_44_632 ();
 sg13g2_decap_8 FILLER_44_639 ();
 sg13g2_decap_4 FILLER_44_646 ();
 sg13g2_decap_4 FILLER_44_656 ();
 sg13g2_fill_2 FILLER_44_660 ();
 sg13g2_fill_2 FILLER_44_694 ();
 sg13g2_fill_1 FILLER_44_710 ();
 sg13g2_fill_2 FILLER_44_757 ();
 sg13g2_fill_2 FILLER_44_780 ();
 sg13g2_fill_1 FILLER_44_782 ();
 sg13g2_decap_4 FILLER_44_787 ();
 sg13g2_decap_4 FILLER_44_817 ();
 sg13g2_decap_4 FILLER_44_825 ();
 sg13g2_fill_1 FILLER_44_829 ();
 sg13g2_fill_1 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_fill_1 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_942 ();
 sg13g2_fill_2 FILLER_44_949 ();
 sg13g2_fill_1 FILLER_44_951 ();
 sg13g2_fill_1 FILLER_44_958 ();
 sg13g2_fill_2 FILLER_44_975 ();
 sg13g2_fill_1 FILLER_44_977 ();
 sg13g2_decap_4 FILLER_44_1004 ();
 sg13g2_fill_2 FILLER_44_1008 ();
 sg13g2_decap_8 FILLER_44_1014 ();
 sg13g2_fill_2 FILLER_44_1021 ();
 sg13g2_fill_1 FILLER_44_1062 ();
 sg13g2_fill_1 FILLER_44_1098 ();
 sg13g2_fill_1 FILLER_44_1121 ();
 sg13g2_fill_1 FILLER_44_1156 ();
 sg13g2_fill_2 FILLER_44_1195 ();
 sg13g2_fill_1 FILLER_44_1204 ();
 sg13g2_fill_2 FILLER_44_1239 ();
 sg13g2_fill_1 FILLER_44_1267 ();
 sg13g2_fill_1 FILLER_44_1299 ();
 sg13g2_decap_8 FILLER_44_1330 ();
 sg13g2_decap_8 FILLER_44_1337 ();
 sg13g2_decap_8 FILLER_44_1344 ();
 sg13g2_decap_8 FILLER_44_1356 ();
 sg13g2_decap_8 FILLER_44_1363 ();
 sg13g2_fill_1 FILLER_44_1375 ();
 sg13g2_decap_4 FILLER_44_1380 ();
 sg13g2_fill_1 FILLER_44_1384 ();
 sg13g2_decap_8 FILLER_44_1389 ();
 sg13g2_decap_4 FILLER_44_1396 ();
 sg13g2_fill_2 FILLER_44_1400 ();
 sg13g2_fill_2 FILLER_44_1486 ();
 sg13g2_fill_1 FILLER_44_1488 ();
 sg13g2_fill_1 FILLER_44_1493 ();
 sg13g2_fill_1 FILLER_44_1520 ();
 sg13g2_fill_1 FILLER_44_1547 ();
 sg13g2_fill_1 FILLER_44_1574 ();
 sg13g2_fill_1 FILLER_44_1579 ();
 sg13g2_fill_1 FILLER_44_1606 ();
 sg13g2_fill_2 FILLER_44_1613 ();
 sg13g2_fill_1 FILLER_44_1615 ();
 sg13g2_decap_4 FILLER_44_1664 ();
 sg13g2_fill_1 FILLER_44_1668 ();
 sg13g2_fill_2 FILLER_44_1734 ();
 sg13g2_fill_1 FILLER_44_1798 ();
 sg13g2_fill_2 FILLER_44_1809 ();
 sg13g2_decap_4 FILLER_44_1855 ();
 sg13g2_fill_1 FILLER_44_1859 ();
 sg13g2_fill_2 FILLER_44_1912 ();
 sg13g2_fill_1 FILLER_44_1964 ();
 sg13g2_fill_1 FILLER_44_1973 ();
 sg13g2_fill_2 FILLER_44_1988 ();
 sg13g2_fill_1 FILLER_44_2000 ();
 sg13g2_fill_1 FILLER_44_2005 ();
 sg13g2_fill_1 FILLER_44_2040 ();
 sg13g2_fill_1 FILLER_44_2048 ();
 sg13g2_fill_1 FILLER_44_2064 ();
 sg13g2_fill_1 FILLER_44_2068 ();
 sg13g2_fill_2 FILLER_44_2117 ();
 sg13g2_decap_8 FILLER_44_2145 ();
 sg13g2_decap_4 FILLER_44_2152 ();
 sg13g2_decap_8 FILLER_44_2160 ();
 sg13g2_decap_8 FILLER_44_2167 ();
 sg13g2_decap_8 FILLER_44_2174 ();
 sg13g2_decap_8 FILLER_44_2181 ();
 sg13g2_fill_2 FILLER_44_2188 ();
 sg13g2_fill_1 FILLER_44_2190 ();
 sg13g2_fill_1 FILLER_44_2196 ();
 sg13g2_fill_1 FILLER_44_2202 ();
 sg13g2_fill_1 FILLER_44_2207 ();
 sg13g2_fill_2 FILLER_44_2212 ();
 sg13g2_fill_1 FILLER_44_2224 ();
 sg13g2_fill_2 FILLER_44_2229 ();
 sg13g2_decap_4 FILLER_44_2252 ();
 sg13g2_fill_1 FILLER_44_2256 ();
 sg13g2_decap_4 FILLER_44_2317 ();
 sg13g2_fill_2 FILLER_44_2321 ();
 sg13g2_decap_8 FILLER_44_2333 ();
 sg13g2_fill_2 FILLER_44_2340 ();
 sg13g2_decap_8 FILLER_44_2347 ();
 sg13g2_fill_1 FILLER_44_2354 ();
 sg13g2_fill_1 FILLER_44_2419 ();
 sg13g2_fill_1 FILLER_44_2450 ();
 sg13g2_decap_4 FILLER_44_2492 ();
 sg13g2_decap_4 FILLER_44_2504 ();
 sg13g2_decap_4 FILLER_44_2565 ();
 sg13g2_fill_2 FILLER_44_2569 ();
 sg13g2_decap_4 FILLER_44_2581 ();
 sg13g2_decap_8 FILLER_44_2611 ();
 sg13g2_fill_2 FILLER_44_2628 ();
 sg13g2_fill_1 FILLER_44_2630 ();
 sg13g2_fill_2 FILLER_44_2635 ();
 sg13g2_fill_1 FILLER_44_2637 ();
 sg13g2_decap_8 FILLER_44_2642 ();
 sg13g2_decap_8 FILLER_44_2649 ();
 sg13g2_decap_8 FILLER_44_2656 ();
 sg13g2_decap_8 FILLER_44_2663 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_31 ();
 sg13g2_decap_8 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_45 ();
 sg13g2_fill_1 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_57 ();
 sg13g2_decap_4 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_76 ();
 sg13g2_decap_8 FILLER_45_83 ();
 sg13g2_decap_4 FILLER_45_90 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_decap_8 FILLER_45_101 ();
 sg13g2_fill_2 FILLER_45_108 ();
 sg13g2_decap_8 FILLER_45_114 ();
 sg13g2_decap_4 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_fill_2 FILLER_45_146 ();
 sg13g2_decap_4 FILLER_45_152 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_fill_2 FILLER_45_209 ();
 sg13g2_fill_1 FILLER_45_211 ();
 sg13g2_fill_2 FILLER_45_240 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_fill_1 FILLER_45_248 ();
 sg13g2_decap_8 FILLER_45_253 ();
 sg13g2_fill_1 FILLER_45_260 ();
 sg13g2_decap_4 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_fill_2 FILLER_45_455 ();
 sg13g2_fill_1 FILLER_45_505 ();
 sg13g2_fill_1 FILLER_45_519 ();
 sg13g2_fill_2 FILLER_45_548 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_fill_2 FILLER_45_579 ();
 sg13g2_fill_1 FILLER_45_622 ();
 sg13g2_fill_1 FILLER_45_631 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_fill_2 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_671 ();
 sg13g2_fill_1 FILLER_45_699 ();
 sg13g2_fill_1 FILLER_45_710 ();
 sg13g2_fill_1 FILLER_45_720 ();
 sg13g2_fill_1 FILLER_45_729 ();
 sg13g2_fill_1 FILLER_45_735 ();
 sg13g2_fill_1 FILLER_45_740 ();
 sg13g2_fill_1 FILLER_45_746 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_fill_2 FILLER_45_847 ();
 sg13g2_fill_1 FILLER_45_857 ();
 sg13g2_fill_1 FILLER_45_909 ();
 sg13g2_fill_2 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_924 ();
 sg13g2_fill_2 FILLER_45_934 ();
 sg13g2_fill_1 FILLER_45_936 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_fill_2 FILLER_45_952 ();
 sg13g2_fill_1 FILLER_45_954 ();
 sg13g2_decap_4 FILLER_45_970 ();
 sg13g2_fill_1 FILLER_45_979 ();
 sg13g2_fill_1 FILLER_45_986 ();
 sg13g2_fill_2 FILLER_45_991 ();
 sg13g2_fill_1 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1003 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_fill_1 FILLER_45_1022 ();
 sg13g2_fill_2 FILLER_45_1033 ();
 sg13g2_fill_2 FILLER_45_1074 ();
 sg13g2_fill_2 FILLER_45_1079 ();
 sg13g2_fill_1 FILLER_45_1112 ();
 sg13g2_fill_1 FILLER_45_1121 ();
 sg13g2_fill_2 FILLER_45_1125 ();
 sg13g2_fill_1 FILLER_45_1158 ();
 sg13g2_fill_1 FILLER_45_1185 ();
 sg13g2_fill_1 FILLER_45_1191 ();
 sg13g2_fill_1 FILLER_45_1197 ();
 sg13g2_fill_1 FILLER_45_1213 ();
 sg13g2_fill_2 FILLER_45_1217 ();
 sg13g2_fill_2 FILLER_45_1227 ();
 sg13g2_fill_1 FILLER_45_1246 ();
 sg13g2_fill_1 FILLER_45_1281 ();
 sg13g2_fill_1 FILLER_45_1318 ();
 sg13g2_decap_4 FILLER_45_1379 ();
 sg13g2_fill_2 FILLER_45_1383 ();
 sg13g2_fill_2 FILLER_45_1395 ();
 sg13g2_fill_1 FILLER_45_1397 ();
 sg13g2_fill_2 FILLER_45_1504 ();
 sg13g2_fill_2 FILLER_45_1516 ();
 sg13g2_fill_2 FILLER_45_1530 ();
 sg13g2_fill_2 FILLER_45_1536 ();
 sg13g2_fill_1 FILLER_45_1538 ();
 sg13g2_fill_1 FILLER_45_1544 ();
 sg13g2_fill_2 FILLER_45_1549 ();
 sg13g2_fill_1 FILLER_45_1556 ();
 sg13g2_fill_2 FILLER_45_1561 ();
 sg13g2_fill_2 FILLER_45_1567 ();
 sg13g2_fill_1 FILLER_45_1569 ();
 sg13g2_fill_2 FILLER_45_1576 ();
 sg13g2_fill_1 FILLER_45_1578 ();
 sg13g2_fill_2 FILLER_45_1592 ();
 sg13g2_fill_2 FILLER_45_1604 ();
 sg13g2_fill_1 FILLER_45_1606 ();
 sg13g2_fill_1 FILLER_45_1650 ();
 sg13g2_fill_1 FILLER_45_1681 ();
 sg13g2_fill_1 FILLER_45_1802 ();
 sg13g2_fill_2 FILLER_45_1815 ();
 sg13g2_fill_2 FILLER_45_1830 ();
 sg13g2_fill_1 FILLER_45_1832 ();
 sg13g2_decap_4 FILLER_45_1843 ();
 sg13g2_fill_1 FILLER_45_1847 ();
 sg13g2_decap_8 FILLER_45_1862 ();
 sg13g2_decap_8 FILLER_45_1869 ();
 sg13g2_decap_8 FILLER_45_1876 ();
 sg13g2_decap_4 FILLER_45_1883 ();
 sg13g2_fill_1 FILLER_45_1887 ();
 sg13g2_fill_2 FILLER_45_1950 ();
 sg13g2_fill_2 FILLER_45_1962 ();
 sg13g2_fill_1 FILLER_45_1974 ();
 sg13g2_decap_8 FILLER_45_1985 ();
 sg13g2_decap_8 FILLER_45_1992 ();
 sg13g2_fill_2 FILLER_45_1999 ();
 sg13g2_fill_2 FILLER_45_2011 ();
 sg13g2_fill_2 FILLER_45_2020 ();
 sg13g2_fill_1 FILLER_45_2027 ();
 sg13g2_fill_2 FILLER_45_2034 ();
 sg13g2_fill_2 FILLER_45_2041 ();
 sg13g2_fill_2 FILLER_45_2060 ();
 sg13g2_fill_1 FILLER_45_2127 ();
 sg13g2_decap_8 FILLER_45_2140 ();
 sg13g2_fill_1 FILLER_45_2147 ();
 sg13g2_decap_8 FILLER_45_2174 ();
 sg13g2_decap_8 FILLER_45_2181 ();
 sg13g2_fill_2 FILLER_45_2188 ();
 sg13g2_fill_1 FILLER_45_2190 ();
 sg13g2_fill_1 FILLER_45_2219 ();
 sg13g2_fill_2 FILLER_45_2224 ();
 sg13g2_fill_2 FILLER_45_2240 ();
 sg13g2_fill_1 FILLER_45_2242 ();
 sg13g2_fill_1 FILLER_45_2279 ();
 sg13g2_decap_4 FILLER_45_2327 ();
 sg13g2_fill_1 FILLER_45_2331 ();
 sg13g2_decap_4 FILLER_45_2358 ();
 sg13g2_fill_1 FILLER_45_2454 ();
 sg13g2_decap_8 FILLER_45_2487 ();
 sg13g2_decap_4 FILLER_45_2494 ();
 sg13g2_fill_2 FILLER_45_2501 ();
 sg13g2_fill_2 FILLER_45_2557 ();
 sg13g2_decap_4 FILLER_45_2585 ();
 sg13g2_fill_2 FILLER_45_2613 ();
 sg13g2_decap_8 FILLER_45_2619 ();
 sg13g2_decap_8 FILLER_45_2626 ();
 sg13g2_decap_8 FILLER_45_2633 ();
 sg13g2_decap_8 FILLER_45_2640 ();
 sg13g2_decap_8 FILLER_45_2647 ();
 sg13g2_decap_8 FILLER_45_2654 ();
 sg13g2_decap_8 FILLER_45_2661 ();
 sg13g2_fill_2 FILLER_45_2668 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_11 ();
 sg13g2_decap_4 FILLER_46_16 ();
 sg13g2_fill_1 FILLER_46_20 ();
 sg13g2_decap_8 FILLER_46_47 ();
 sg13g2_decap_8 FILLER_46_54 ();
 sg13g2_decap_8 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_68 ();
 sg13g2_decap_4 FILLER_46_75 ();
 sg13g2_fill_1 FILLER_46_79 ();
 sg13g2_decap_8 FILLER_46_93 ();
 sg13g2_decap_8 FILLER_46_100 ();
 sg13g2_decap_8 FILLER_46_107 ();
 sg13g2_decap_4 FILLER_46_123 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_decap_4 FILLER_46_181 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_decap_8 FILLER_46_227 ();
 sg13g2_decap_8 FILLER_46_265 ();
 sg13g2_decap_4 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_1 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_fill_2 FILLER_46_350 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_409 ();
 sg13g2_fill_2 FILLER_46_451 ();
 sg13g2_fill_1 FILLER_46_484 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_1 FILLER_46_494 ();
 sg13g2_fill_2 FILLER_46_514 ();
 sg13g2_fill_1 FILLER_46_526 ();
 sg13g2_fill_2 FILLER_46_540 ();
 sg13g2_fill_1 FILLER_46_639 ();
 sg13g2_fill_1 FILLER_46_644 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_1 FILLER_46_691 ();
 sg13g2_decap_4 FILLER_46_726 ();
 sg13g2_fill_1 FILLER_46_749 ();
 sg13g2_fill_2 FILLER_46_758 ();
 sg13g2_fill_1 FILLER_46_760 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_fill_2 FILLER_46_779 ();
 sg13g2_fill_1 FILLER_46_781 ();
 sg13g2_decap_4 FILLER_46_786 ();
 sg13g2_fill_2 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_4 FILLER_46_821 ();
 sg13g2_fill_1 FILLER_46_825 ();
 sg13g2_decap_4 FILLER_46_858 ();
 sg13g2_fill_2 FILLER_46_862 ();
 sg13g2_fill_1 FILLER_46_868 ();
 sg13g2_fill_2 FILLER_46_874 ();
 sg13g2_fill_2 FILLER_46_884 ();
 sg13g2_fill_2 FILLER_46_889 ();
 sg13g2_fill_1 FILLER_46_903 ();
 sg13g2_fill_1 FILLER_46_913 ();
 sg13g2_decap_8 FILLER_46_951 ();
 sg13g2_decap_8 FILLER_46_958 ();
 sg13g2_fill_1 FILLER_46_965 ();
 sg13g2_fill_1 FILLER_46_977 ();
 sg13g2_fill_1 FILLER_46_994 ();
 sg13g2_decap_4 FILLER_46_1000 ();
 sg13g2_fill_1 FILLER_46_1004 ();
 sg13g2_decap_8 FILLER_46_1009 ();
 sg13g2_decap_4 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1030 ();
 sg13g2_fill_1 FILLER_46_1081 ();
 sg13g2_fill_1 FILLER_46_1118 ();
 sg13g2_fill_2 FILLER_46_1132 ();
 sg13g2_fill_2 FILLER_46_1177 ();
 sg13g2_fill_1 FILLER_46_1186 ();
 sg13g2_fill_1 FILLER_46_1259 ();
 sg13g2_fill_2 FILLER_46_1271 ();
 sg13g2_fill_1 FILLER_46_1307 ();
 sg13g2_fill_2 FILLER_46_1311 ();
 sg13g2_fill_1 FILLER_46_1327 ();
 sg13g2_fill_1 FILLER_46_1338 ();
 sg13g2_fill_2 FILLER_46_1346 ();
 sg13g2_fill_2 FILLER_46_1351 ();
 sg13g2_decap_8 FILLER_46_1357 ();
 sg13g2_decap_4 FILLER_46_1364 ();
 sg13g2_fill_2 FILLER_46_1433 ();
 sg13g2_fill_2 FILLER_46_1447 ();
 sg13g2_fill_2 FILLER_46_1458 ();
 sg13g2_fill_2 FILLER_46_1465 ();
 sg13g2_fill_2 FILLER_46_1471 ();
 sg13g2_fill_1 FILLER_46_1477 ();
 sg13g2_fill_1 FILLER_46_1483 ();
 sg13g2_decap_8 FILLER_46_1492 ();
 sg13g2_fill_2 FILLER_46_1499 ();
 sg13g2_fill_1 FILLER_46_1512 ();
 sg13g2_decap_4 FILLER_46_1519 ();
 sg13g2_fill_1 FILLER_46_1527 ();
 sg13g2_fill_1 FILLER_46_1533 ();
 sg13g2_fill_2 FILLER_46_1543 ();
 sg13g2_fill_1 FILLER_46_1545 ();
 sg13g2_fill_1 FILLER_46_1606 ();
 sg13g2_fill_2 FILLER_46_1612 ();
 sg13g2_fill_1 FILLER_46_1614 ();
 sg13g2_fill_1 FILLER_46_1664 ();
 sg13g2_fill_1 FILLER_46_1698 ();
 sg13g2_fill_2 FILLER_46_1712 ();
 sg13g2_fill_1 FILLER_46_1728 ();
 sg13g2_fill_1 FILLER_46_1766 ();
 sg13g2_fill_1 FILLER_46_1800 ();
 sg13g2_decap_4 FILLER_46_1837 ();
 sg13g2_fill_1 FILLER_46_1841 ();
 sg13g2_fill_1 FILLER_46_1874 ();
 sg13g2_fill_1 FILLER_46_1933 ();
 sg13g2_fill_1 FILLER_46_1955 ();
 sg13g2_decap_8 FILLER_46_1986 ();
 sg13g2_decap_8 FILLER_46_1993 ();
 sg13g2_fill_2 FILLER_46_2000 ();
 sg13g2_fill_1 FILLER_46_2002 ();
 sg13g2_fill_2 FILLER_46_2046 ();
 sg13g2_fill_1 FILLER_46_2055 ();
 sg13g2_fill_1 FILLER_46_2065 ();
 sg13g2_fill_1 FILLER_46_2084 ();
 sg13g2_fill_2 FILLER_46_2130 ();
 sg13g2_decap_8 FILLER_46_2136 ();
 sg13g2_decap_4 FILLER_46_2153 ();
 sg13g2_fill_1 FILLER_46_2157 ();
 sg13g2_decap_8 FILLER_46_2167 ();
 sg13g2_decap_8 FILLER_46_2174 ();
 sg13g2_fill_2 FILLER_46_2181 ();
 sg13g2_fill_1 FILLER_46_2183 ();
 sg13g2_fill_1 FILLER_46_2208 ();
 sg13g2_fill_2 FILLER_46_2213 ();
 sg13g2_fill_1 FILLER_46_2240 ();
 sg13g2_decap_4 FILLER_46_2245 ();
 sg13g2_fill_1 FILLER_46_2249 ();
 sg13g2_fill_2 FILLER_46_2260 ();
 sg13g2_fill_1 FILLER_46_2266 ();
 sg13g2_fill_1 FILLER_46_2271 ();
 sg13g2_fill_1 FILLER_46_2276 ();
 sg13g2_fill_1 FILLER_46_2287 ();
 sg13g2_fill_1 FILLER_46_2298 ();
 sg13g2_fill_2 FILLER_46_2303 ();
 sg13g2_fill_2 FILLER_46_2331 ();
 sg13g2_fill_1 FILLER_46_2333 ();
 sg13g2_decap_8 FILLER_46_2342 ();
 sg13g2_fill_2 FILLER_46_2349 ();
 sg13g2_fill_1 FILLER_46_2361 ();
 sg13g2_decap_8 FILLER_46_2366 ();
 sg13g2_decap_8 FILLER_46_2373 ();
 sg13g2_fill_1 FILLER_46_2390 ();
 sg13g2_fill_2 FILLER_46_2403 ();
 sg13g2_fill_1 FILLER_46_2405 ();
 sg13g2_decap_8 FILLER_46_2553 ();
 sg13g2_decap_4 FILLER_46_2560 ();
 sg13g2_fill_1 FILLER_46_2564 ();
 sg13g2_decap_8 FILLER_46_2634 ();
 sg13g2_decap_8 FILLER_46_2641 ();
 sg13g2_decap_8 FILLER_46_2648 ();
 sg13g2_decap_8 FILLER_46_2655 ();
 sg13g2_decap_8 FILLER_46_2662 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_61 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_116 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_143 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_205 ();
 sg13g2_decap_8 FILLER_47_214 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_fill_1 FILLER_47_232 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_260 ();
 sg13g2_fill_2 FILLER_47_266 ();
 sg13g2_fill_2 FILLER_47_273 ();
 sg13g2_fill_1 FILLER_47_275 ();
 sg13g2_fill_2 FILLER_47_312 ();
 sg13g2_decap_8 FILLER_47_318 ();
 sg13g2_decap_4 FILLER_47_325 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_decap_8 FILLER_47_341 ();
 sg13g2_decap_8 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_412 ();
 sg13g2_fill_1 FILLER_47_418 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_fill_2 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_440 ();
 sg13g2_fill_2 FILLER_47_517 ();
 sg13g2_fill_2 FILLER_47_586 ();
 sg13g2_fill_1 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_626 ();
 sg13g2_fill_2 FILLER_47_641 ();
 sg13g2_fill_2 FILLER_47_658 ();
 sg13g2_fill_1 FILLER_47_660 ();
 sg13g2_fill_1 FILLER_47_688 ();
 sg13g2_fill_1 FILLER_47_722 ();
 sg13g2_fill_1 FILLER_47_766 ();
 sg13g2_fill_1 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_fill_2 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_decap_4 FILLER_47_870 ();
 sg13g2_decap_4 FILLER_47_888 ();
 sg13g2_fill_2 FILLER_47_892 ();
 sg13g2_decap_4 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_908 ();
 sg13g2_fill_2 FILLER_47_915 ();
 sg13g2_fill_1 FILLER_47_925 ();
 sg13g2_fill_2 FILLER_47_943 ();
 sg13g2_fill_1 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_fill_2 FILLER_47_976 ();
 sg13g2_fill_2 FILLER_47_985 ();
 sg13g2_fill_2 FILLER_47_1038 ();
 sg13g2_fill_2 FILLER_47_1065 ();
 sg13g2_fill_1 FILLER_47_1114 ();
 sg13g2_fill_1 FILLER_47_1149 ();
 sg13g2_fill_1 FILLER_47_1160 ();
 sg13g2_fill_1 FILLER_47_1166 ();
 sg13g2_fill_1 FILLER_47_1171 ();
 sg13g2_fill_1 FILLER_47_1179 ();
 sg13g2_fill_2 FILLER_47_1255 ();
 sg13g2_fill_1 FILLER_47_1318 ();
 sg13g2_fill_2 FILLER_47_1355 ();
 sg13g2_fill_2 FILLER_47_1383 ();
 sg13g2_decap_4 FILLER_47_1389 ();
 sg13g2_fill_1 FILLER_47_1397 ();
 sg13g2_fill_2 FILLER_47_1402 ();
 sg13g2_fill_2 FILLER_47_1408 ();
 sg13g2_decap_4 FILLER_47_1414 ();
 sg13g2_fill_2 FILLER_47_1418 ();
 sg13g2_decap_8 FILLER_47_1440 ();
 sg13g2_fill_1 FILLER_47_1447 ();
 sg13g2_decap_8 FILLER_47_1480 ();
 sg13g2_fill_2 FILLER_47_1487 ();
 sg13g2_decap_8 FILLER_47_1493 ();
 sg13g2_decap_4 FILLER_47_1500 ();
 sg13g2_fill_2 FILLER_47_1560 ();
 sg13g2_fill_2 FILLER_47_1576 ();
 sg13g2_fill_2 FILLER_47_1591 ();
 sg13g2_decap_8 FILLER_47_1606 ();
 sg13g2_fill_2 FILLER_47_1617 ();
 sg13g2_fill_1 FILLER_47_1619 ();
 sg13g2_fill_1 FILLER_47_1756 ();
 sg13g2_fill_1 FILLER_47_1796 ();
 sg13g2_decap_8 FILLER_47_1823 ();
 sg13g2_fill_2 FILLER_47_1830 ();
 sg13g2_decap_8 FILLER_47_1849 ();
 sg13g2_decap_4 FILLER_47_1856 ();
 sg13g2_fill_1 FILLER_47_1860 ();
 sg13g2_fill_2 FILLER_47_1867 ();
 sg13g2_fill_1 FILLER_47_1869 ();
 sg13g2_fill_1 FILLER_47_1891 ();
 sg13g2_fill_1 FILLER_47_1925 ();
 sg13g2_fill_1 FILLER_47_1936 ();
 sg13g2_fill_1 FILLER_47_1967 ();
 sg13g2_decap_4 FILLER_47_1994 ();
 sg13g2_fill_1 FILLER_47_2020 ();
 sg13g2_fill_2 FILLER_47_2027 ();
 sg13g2_fill_2 FILLER_47_2032 ();
 sg13g2_fill_1 FILLER_47_2044 ();
 sg13g2_fill_1 FILLER_47_2142 ();
 sg13g2_decap_8 FILLER_47_2147 ();
 sg13g2_fill_1 FILLER_47_2163 ();
 sg13g2_fill_2 FILLER_47_2177 ();
 sg13g2_fill_1 FILLER_47_2187 ();
 sg13g2_fill_1 FILLER_47_2193 ();
 sg13g2_fill_2 FILLER_47_2199 ();
 sg13g2_fill_1 FILLER_47_2201 ();
 sg13g2_decap_8 FILLER_47_2257 ();
 sg13g2_decap_4 FILLER_47_2264 ();
 sg13g2_fill_1 FILLER_47_2268 ();
 sg13g2_fill_2 FILLER_47_2299 ();
 sg13g2_fill_1 FILLER_47_2301 ();
 sg13g2_decap_4 FILLER_47_2337 ();
 sg13g2_fill_2 FILLER_47_2341 ();
 sg13g2_fill_2 FILLER_47_2384 ();
 sg13g2_fill_1 FILLER_47_2386 ();
 sg13g2_fill_1 FILLER_47_2444 ();
 sg13g2_fill_1 FILLER_47_2510 ();
 sg13g2_fill_2 FILLER_47_2517 ();
 sg13g2_fill_1 FILLER_47_2523 ();
 sg13g2_decap_8 FILLER_47_2550 ();
 sg13g2_decap_8 FILLER_47_2557 ();
 sg13g2_decap_8 FILLER_47_2564 ();
 sg13g2_decap_4 FILLER_47_2571 ();
 sg13g2_fill_1 FILLER_47_2575 ();
 sg13g2_fill_1 FILLER_47_2580 ();
 sg13g2_fill_1 FILLER_47_2606 ();
 sg13g2_fill_1 FILLER_47_2633 ();
 sg13g2_decap_8 FILLER_47_2660 ();
 sg13g2_fill_2 FILLER_47_2667 ();
 sg13g2_fill_1 FILLER_47_2669 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_fill_1 FILLER_48_103 ();
 sg13g2_fill_1 FILLER_48_134 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_174 ();
 sg13g2_decap_8 FILLER_48_180 ();
 sg13g2_decap_4 FILLER_48_187 ();
 sg13g2_fill_1 FILLER_48_208 ();
 sg13g2_fill_2 FILLER_48_213 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_decap_4 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_229 ();
 sg13g2_decap_4 FILLER_48_234 ();
 sg13g2_fill_2 FILLER_48_246 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_fill_1 FILLER_48_255 ();
 sg13g2_decap_8 FILLER_48_260 ();
 sg13g2_decap_4 FILLER_48_267 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_fill_2 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_410 ();
 sg13g2_fill_1 FILLER_48_417 ();
 sg13g2_decap_8 FILLER_48_433 ();
 sg13g2_fill_2 FILLER_48_444 ();
 sg13g2_fill_1 FILLER_48_451 ();
 sg13g2_fill_2 FILLER_48_526 ();
 sg13g2_fill_1 FILLER_48_542 ();
 sg13g2_fill_2 FILLER_48_548 ();
 sg13g2_fill_2 FILLER_48_622 ();
 sg13g2_fill_2 FILLER_48_664 ();
 sg13g2_fill_1 FILLER_48_666 ();
 sg13g2_fill_1 FILLER_48_677 ();
 sg13g2_fill_1 FILLER_48_695 ();
 sg13g2_fill_1 FILLER_48_713 ();
 sg13g2_fill_2 FILLER_48_727 ();
 sg13g2_fill_2 FILLER_48_744 ();
 sg13g2_fill_2 FILLER_48_755 ();
 sg13g2_fill_1 FILLER_48_757 ();
 sg13g2_decap_4 FILLER_48_777 ();
 sg13g2_fill_1 FILLER_48_781 ();
 sg13g2_fill_2 FILLER_48_839 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_fill_2 FILLER_48_887 ();
 sg13g2_fill_1 FILLER_48_894 ();
 sg13g2_fill_1 FILLER_48_899 ();
 sg13g2_fill_2 FILLER_48_905 ();
 sg13g2_fill_2 FILLER_48_912 ();
 sg13g2_fill_2 FILLER_48_921 ();
 sg13g2_fill_1 FILLER_48_923 ();
 sg13g2_decap_8 FILLER_48_933 ();
 sg13g2_decap_8 FILLER_48_940 ();
 sg13g2_decap_8 FILLER_48_947 ();
 sg13g2_decap_8 FILLER_48_954 ();
 sg13g2_fill_2 FILLER_48_961 ();
 sg13g2_decap_8 FILLER_48_971 ();
 sg13g2_decap_8 FILLER_48_978 ();
 sg13g2_decap_4 FILLER_48_985 ();
 sg13g2_fill_1 FILLER_48_989 ();
 sg13g2_decap_4 FILLER_48_1000 ();
 sg13g2_fill_2 FILLER_48_1008 ();
 sg13g2_fill_2 FILLER_48_1019 ();
 sg13g2_fill_2 FILLER_48_1036 ();
 sg13g2_fill_1 FILLER_48_1056 ();
 sg13g2_fill_1 FILLER_48_1157 ();
 sg13g2_fill_1 FILLER_48_1198 ();
 sg13g2_fill_1 FILLER_48_1248 ();
 sg13g2_fill_2 FILLER_48_1326 ();
 sg13g2_decap_4 FILLER_48_1335 ();
 sg13g2_decap_8 FILLER_48_1382 ();
 sg13g2_decap_8 FILLER_48_1389 ();
 sg13g2_fill_2 FILLER_48_1396 ();
 sg13g2_decap_4 FILLER_48_1402 ();
 sg13g2_fill_2 FILLER_48_1429 ();
 sg13g2_fill_1 FILLER_48_1431 ();
 sg13g2_fill_2 FILLER_48_1441 ();
 sg13g2_fill_1 FILLER_48_1443 ();
 sg13g2_fill_2 FILLER_48_1449 ();
 sg13g2_fill_1 FILLER_48_1451 ();
 sg13g2_decap_4 FILLER_48_1456 ();
 sg13g2_decap_8 FILLER_48_1464 ();
 sg13g2_fill_2 FILLER_48_1471 ();
 sg13g2_fill_1 FILLER_48_1473 ();
 sg13g2_fill_1 FILLER_48_1508 ();
 sg13g2_fill_1 FILLER_48_1515 ();
 sg13g2_fill_2 FILLER_48_1527 ();
 sg13g2_decap_8 FILLER_48_1551 ();
 sg13g2_decap_4 FILLER_48_1558 ();
 sg13g2_fill_2 FILLER_48_1562 ();
 sg13g2_fill_1 FILLER_48_1593 ();
 sg13g2_decap_4 FILLER_48_1612 ();
 sg13g2_fill_1 FILLER_48_1633 ();
 sg13g2_fill_1 FILLER_48_1664 ();
 sg13g2_fill_1 FILLER_48_1726 ();
 sg13g2_fill_2 FILLER_48_1747 ();
 sg13g2_fill_2 FILLER_48_1803 ();
 sg13g2_fill_1 FILLER_48_1825 ();
 sg13g2_fill_1 FILLER_48_1952 ();
 sg13g2_decap_4 FILLER_48_1966 ();
 sg13g2_fill_1 FILLER_48_2015 ();
 sg13g2_fill_1 FILLER_48_2033 ();
 sg13g2_fill_2 FILLER_48_2063 ();
 sg13g2_fill_2 FILLER_48_2070 ();
 sg13g2_fill_2 FILLER_48_2077 ();
 sg13g2_fill_2 FILLER_48_2105 ();
 sg13g2_fill_1 FILLER_48_2137 ();
 sg13g2_decap_4 FILLER_48_2148 ();
 sg13g2_decap_4 FILLER_48_2221 ();
 sg13g2_fill_2 FILLER_48_2251 ();
 sg13g2_fill_2 FILLER_48_2351 ();
 sg13g2_fill_1 FILLER_48_2404 ();
 sg13g2_fill_2 FILLER_48_2423 ();
 sg13g2_fill_1 FILLER_48_2483 ();
 sg13g2_fill_1 FILLER_48_2510 ();
 sg13g2_decap_8 FILLER_48_2558 ();
 sg13g2_decap_8 FILLER_48_2565 ();
 sg13g2_decap_8 FILLER_48_2572 ();
 sg13g2_decap_8 FILLER_48_2579 ();
 sg13g2_fill_1 FILLER_48_2586 ();
 sg13g2_fill_2 FILLER_48_2623 ();
 sg13g2_fill_2 FILLER_48_2629 ();
 sg13g2_fill_1 FILLER_48_2641 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_13 ();
 sg13g2_decap_4 FILLER_49_52 ();
 sg13g2_fill_2 FILLER_49_56 ();
 sg13g2_fill_1 FILLER_49_66 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_fill_1 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_143 ();
 sg13g2_fill_2 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_fill_2 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_fill_1 FILLER_49_326 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_379 ();
 sg13g2_fill_2 FILLER_49_384 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_decap_4 FILLER_49_407 ();
 sg13g2_fill_2 FILLER_49_411 ();
 sg13g2_fill_1 FILLER_49_428 ();
 sg13g2_decap_4 FILLER_49_455 ();
 sg13g2_fill_1 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_464 ();
 sg13g2_fill_2 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_521 ();
 sg13g2_fill_1 FILLER_49_532 ();
 sg13g2_fill_2 FILLER_49_546 ();
 sg13g2_fill_1 FILLER_49_629 ();
 sg13g2_fill_1 FILLER_49_654 ();
 sg13g2_fill_1 FILLER_49_660 ();
 sg13g2_fill_1 FILLER_49_666 ();
 sg13g2_decap_4 FILLER_49_672 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_fill_2 FILLER_49_717 ();
 sg13g2_decap_4 FILLER_49_724 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_fill_1 FILLER_49_739 ();
 sg13g2_fill_2 FILLER_49_744 ();
 sg13g2_fill_2 FILLER_49_760 ();
 sg13g2_fill_1 FILLER_49_762 ();
 sg13g2_decap_4 FILLER_49_777 ();
 sg13g2_fill_1 FILLER_49_787 ();
 sg13g2_fill_1 FILLER_49_793 ();
 sg13g2_fill_1 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_872 ();
 sg13g2_fill_1 FILLER_49_879 ();
 sg13g2_decap_4 FILLER_49_898 ();
 sg13g2_decap_8 FILLER_49_906 ();
 sg13g2_decap_4 FILLER_49_918 ();
 sg13g2_fill_2 FILLER_49_922 ();
 sg13g2_fill_2 FILLER_49_972 ();
 sg13g2_fill_2 FILLER_49_979 ();
 sg13g2_decap_4 FILLER_49_987 ();
 sg13g2_fill_2 FILLER_49_991 ();
 sg13g2_decap_4 FILLER_49_1001 ();
 sg13g2_fill_2 FILLER_49_1010 ();
 sg13g2_fill_1 FILLER_49_1012 ();
 sg13g2_fill_2 FILLER_49_1032 ();
 sg13g2_fill_1 FILLER_49_1041 ();
 sg13g2_fill_1 FILLER_49_1052 ();
 sg13g2_fill_1 FILLER_49_1092 ();
 sg13g2_fill_1 FILLER_49_1146 ();
 sg13g2_fill_2 FILLER_49_1152 ();
 sg13g2_fill_2 FILLER_49_1159 ();
 sg13g2_fill_1 FILLER_49_1192 ();
 sg13g2_fill_2 FILLER_49_1201 ();
 sg13g2_fill_1 FILLER_49_1234 ();
 sg13g2_fill_1 FILLER_49_1263 ();
 sg13g2_fill_2 FILLER_49_1281 ();
 sg13g2_decap_4 FILLER_49_1325 ();
 sg13g2_fill_2 FILLER_49_1329 ();
 sg13g2_decap_8 FILLER_49_1374 ();
 sg13g2_decap_4 FILLER_49_1381 ();
 sg13g2_fill_1 FILLER_49_1385 ();
 sg13g2_fill_1 FILLER_49_1396 ();
 sg13g2_fill_1 FILLER_49_1437 ();
 sg13g2_decap_4 FILLER_49_1498 ();
 sg13g2_fill_1 FILLER_49_1526 ();
 sg13g2_fill_2 FILLER_49_1553 ();
 sg13g2_fill_1 FILLER_49_1555 ();
 sg13g2_fill_2 FILLER_49_1560 ();
 sg13g2_fill_1 FILLER_49_1562 ();
 sg13g2_fill_2 FILLER_49_1571 ();
 sg13g2_fill_1 FILLER_49_1573 ();
 sg13g2_fill_1 FILLER_49_1608 ();
 sg13g2_fill_2 FILLER_49_1650 ();
 sg13g2_fill_1 FILLER_49_1683 ();
 sg13g2_fill_1 FILLER_49_1720 ();
 sg13g2_fill_2 FILLER_49_1753 ();
 sg13g2_fill_1 FILLER_49_1765 ();
 sg13g2_fill_2 FILLER_49_1829 ();
 sg13g2_fill_1 FILLER_49_1837 ();
 sg13g2_fill_2 FILLER_49_1846 ();
 sg13g2_fill_2 FILLER_49_1861 ();
 sg13g2_fill_1 FILLER_49_1873 ();
 sg13g2_fill_2 FILLER_49_1950 ();
 sg13g2_fill_2 FILLER_49_1972 ();
 sg13g2_fill_2 FILLER_49_2009 ();
 sg13g2_fill_1 FILLER_49_2022 ();
 sg13g2_fill_2 FILLER_49_2100 ();
 sg13g2_fill_2 FILLER_49_2130 ();
 sg13g2_fill_2 FILLER_49_2163 ();
 sg13g2_fill_1 FILLER_49_2165 ();
 sg13g2_decap_4 FILLER_49_2171 ();
 sg13g2_fill_1 FILLER_49_2175 ();
 sg13g2_fill_1 FILLER_49_2185 ();
 sg13g2_fill_1 FILLER_49_2190 ();
 sg13g2_fill_2 FILLER_49_2195 ();
 sg13g2_decap_8 FILLER_49_2253 ();
 sg13g2_fill_1 FILLER_49_2260 ();
 sg13g2_decap_4 FILLER_49_2265 ();
 sg13g2_fill_1 FILLER_49_2269 ();
 sg13g2_fill_1 FILLER_49_2278 ();
 sg13g2_fill_1 FILLER_49_2287 ();
 sg13g2_fill_1 FILLER_49_2334 ();
 sg13g2_fill_2 FILLER_49_2347 ();
 sg13g2_decap_8 FILLER_49_2364 ();
 sg13g2_decap_4 FILLER_49_2371 ();
 sg13g2_fill_2 FILLER_49_2375 ();
 sg13g2_fill_2 FILLER_49_2407 ();
 sg13g2_decap_4 FILLER_49_2417 ();
 sg13g2_fill_2 FILLER_49_2469 ();
 sg13g2_fill_1 FILLER_49_2507 ();
 sg13g2_decap_8 FILLER_49_2553 ();
 sg13g2_decap_8 FILLER_49_2560 ();
 sg13g2_decap_4 FILLER_49_2593 ();
 sg13g2_fill_1 FILLER_49_2597 ();
 sg13g2_fill_2 FILLER_49_2612 ();
 sg13g2_fill_1 FILLER_49_2614 ();
 sg13g2_decap_4 FILLER_49_2623 ();
 sg13g2_fill_1 FILLER_49_2627 ();
 sg13g2_decap_4 FILLER_49_2638 ();
 sg13g2_fill_1 FILLER_49_2642 ();
 sg13g2_fill_2 FILLER_49_2647 ();
 sg13g2_fill_1 FILLER_49_2649 ();
 sg13g2_decap_8 FILLER_49_2654 ();
 sg13g2_decap_8 FILLER_49_2661 ();
 sg13g2_fill_2 FILLER_49_2668 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_51 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_fill_2 FILLER_50_100 ();
 sg13g2_fill_2 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_117 ();
 sg13g2_fill_2 FILLER_50_136 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_200 ();
 sg13g2_fill_2 FILLER_50_207 ();
 sg13g2_decap_8 FILLER_50_214 ();
 sg13g2_fill_1 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_227 ();
 sg13g2_fill_2 FILLER_50_253 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_decap_4 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_fill_2 FILLER_50_299 ();
 sg13g2_fill_1 FILLER_50_301 ();
 sg13g2_fill_1 FILLER_50_327 ();
 sg13g2_fill_2 FILLER_50_348 ();
 sg13g2_decap_8 FILLER_50_355 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_393 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_409 ();
 sg13g2_fill_1 FILLER_50_414 ();
 sg13g2_fill_2 FILLER_50_420 ();
 sg13g2_fill_1 FILLER_50_483 ();
 sg13g2_fill_2 FILLER_50_533 ();
 sg13g2_fill_2 FILLER_50_549 ();
 sg13g2_fill_2 FILLER_50_570 ();
 sg13g2_fill_1 FILLER_50_575 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_fill_2 FILLER_50_606 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_fill_1 FILLER_50_624 ();
 sg13g2_fill_1 FILLER_50_635 ();
 sg13g2_fill_1 FILLER_50_646 ();
 sg13g2_fill_2 FILLER_50_656 ();
 sg13g2_fill_1 FILLER_50_702 ();
 sg13g2_fill_1 FILLER_50_718 ();
 sg13g2_fill_2 FILLER_50_728 ();
 sg13g2_fill_1 FILLER_50_740 ();
 sg13g2_fill_1 FILLER_50_765 ();
 sg13g2_fill_2 FILLER_50_771 ();
 sg13g2_fill_2 FILLER_50_804 ();
 sg13g2_fill_1 FILLER_50_806 ();
 sg13g2_fill_2 FILLER_50_839 ();
 sg13g2_fill_1 FILLER_50_867 ();
 sg13g2_fill_1 FILLER_50_872 ();
 sg13g2_fill_2 FILLER_50_883 ();
 sg13g2_fill_2 FILLER_50_896 ();
 sg13g2_fill_2 FILLER_50_912 ();
 sg13g2_fill_1 FILLER_50_914 ();
 sg13g2_fill_2 FILLER_50_919 ();
 sg13g2_decap_4 FILLER_50_926 ();
 sg13g2_fill_1 FILLER_50_930 ();
 sg13g2_fill_2 FILLER_50_935 ();
 sg13g2_fill_2 FILLER_50_942 ();
 sg13g2_fill_1 FILLER_50_944 ();
 sg13g2_decap_8 FILLER_50_949 ();
 sg13g2_decap_4 FILLER_50_956 ();
 sg13g2_fill_2 FILLER_50_960 ();
 sg13g2_decap_8 FILLER_50_975 ();
 sg13g2_decap_8 FILLER_50_982 ();
 sg13g2_decap_8 FILLER_50_989 ();
 sg13g2_fill_1 FILLER_50_996 ();
 sg13g2_fill_1 FILLER_50_1036 ();
 sg13g2_fill_1 FILLER_50_1051 ();
 sg13g2_fill_1 FILLER_50_1068 ();
 sg13g2_fill_1 FILLER_50_1074 ();
 sg13g2_fill_2 FILLER_50_1111 ();
 sg13g2_fill_2 FILLER_50_1118 ();
 sg13g2_fill_2 FILLER_50_1132 ();
 sg13g2_fill_1 FILLER_50_1138 ();
 sg13g2_fill_2 FILLER_50_1156 ();
 sg13g2_fill_2 FILLER_50_1174 ();
 sg13g2_fill_2 FILLER_50_1241 ();
 sg13g2_fill_1 FILLER_50_1247 ();
 sg13g2_fill_1 FILLER_50_1274 ();
 sg13g2_fill_1 FILLER_50_1288 ();
 sg13g2_fill_2 FILLER_50_1308 ();
 sg13g2_decap_8 FILLER_50_1318 ();
 sg13g2_decap_8 FILLER_50_1374 ();
 sg13g2_decap_8 FILLER_50_1381 ();
 sg13g2_decap_8 FILLER_50_1388 ();
 sg13g2_decap_4 FILLER_50_1395 ();
 sg13g2_decap_4 FILLER_50_1409 ();
 sg13g2_fill_1 FILLER_50_1413 ();
 sg13g2_fill_1 FILLER_50_1444 ();
 sg13g2_fill_1 FILLER_50_1471 ();
 sg13g2_fill_1 FILLER_50_1483 ();
 sg13g2_fill_1 FILLER_50_1494 ();
 sg13g2_fill_2 FILLER_50_1509 ();
 sg13g2_fill_1 FILLER_50_1545 ();
 sg13g2_decap_4 FILLER_50_1561 ();
 sg13g2_fill_2 FILLER_50_1602 ();
 sg13g2_decap_4 FILLER_50_1669 ();
 sg13g2_fill_1 FILLER_50_1673 ();
 sg13g2_fill_1 FILLER_50_1688 ();
 sg13g2_fill_1 FILLER_50_1693 ();
 sg13g2_fill_2 FILLER_50_1702 ();
 sg13g2_fill_2 FILLER_50_1799 ();
 sg13g2_fill_1 FILLER_50_1818 ();
 sg13g2_fill_1 FILLER_50_1832 ();
 sg13g2_fill_1 FILLER_50_1848 ();
 sg13g2_fill_2 FILLER_50_1854 ();
 sg13g2_fill_2 FILLER_50_1860 ();
 sg13g2_fill_1 FILLER_50_1898 ();
 sg13g2_fill_2 FILLER_50_1977 ();
 sg13g2_fill_1 FILLER_50_1979 ();
 sg13g2_decap_8 FILLER_50_1984 ();
 sg13g2_decap_8 FILLER_50_1991 ();
 sg13g2_fill_2 FILLER_50_1998 ();
 sg13g2_fill_1 FILLER_50_2000 ();
 sg13g2_fill_1 FILLER_50_2012 ();
 sg13g2_fill_1 FILLER_50_2052 ();
 sg13g2_fill_2 FILLER_50_2106 ();
 sg13g2_fill_1 FILLER_50_2119 ();
 sg13g2_fill_1 FILLER_50_2126 ();
 sg13g2_fill_2 FILLER_50_2159 ();
 sg13g2_decap_8 FILLER_50_2165 ();
 sg13g2_fill_2 FILLER_50_2172 ();
 sg13g2_fill_1 FILLER_50_2174 ();
 sg13g2_decap_8 FILLER_50_2180 ();
 sg13g2_fill_2 FILLER_50_2187 ();
 sg13g2_decap_8 FILLER_50_2194 ();
 sg13g2_fill_1 FILLER_50_2232 ();
 sg13g2_decap_4 FILLER_50_2237 ();
 sg13g2_fill_2 FILLER_50_2251 ();
 sg13g2_fill_1 FILLER_50_2282 ();
 sg13g2_decap_4 FILLER_50_2303 ();
 sg13g2_fill_1 FILLER_50_2339 ();
 sg13g2_fill_1 FILLER_50_2348 ();
 sg13g2_fill_1 FILLER_50_2356 ();
 sg13g2_fill_1 FILLER_50_2402 ();
 sg13g2_decap_4 FILLER_50_2412 ();
 sg13g2_fill_2 FILLER_50_2416 ();
 sg13g2_fill_2 FILLER_50_2449 ();
 sg13g2_fill_2 FILLER_50_2518 ();
 sg13g2_decap_4 FILLER_50_2559 ();
 sg13g2_decap_8 FILLER_50_2588 ();
 sg13g2_fill_1 FILLER_50_2595 ();
 sg13g2_decap_8 FILLER_50_2606 ();
 sg13g2_decap_8 FILLER_50_2613 ();
 sg13g2_fill_2 FILLER_50_2620 ();
 sg13g2_decap_8 FILLER_50_2643 ();
 sg13g2_decap_8 FILLER_50_2650 ();
 sg13g2_decap_8 FILLER_50_2657 ();
 sg13g2_decap_4 FILLER_50_2664 ();
 sg13g2_fill_2 FILLER_50_2668 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_13 ();
 sg13g2_decap_4 FILLER_51_20 ();
 sg13g2_decap_4 FILLER_51_37 ();
 sg13g2_decap_4 FILLER_51_45 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_fill_2 FILLER_51_130 ();
 sg13g2_decap_8 FILLER_51_136 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_fill_1 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_2 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_322 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_342 ();
 sg13g2_fill_2 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_fill_2 FILLER_51_373 ();
 sg13g2_fill_1 FILLER_51_375 ();
 sg13g2_fill_2 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_fill_1 FILLER_51_389 ();
 sg13g2_fill_2 FILLER_51_419 ();
 sg13g2_fill_1 FILLER_51_441 ();
 sg13g2_fill_2 FILLER_51_484 ();
 sg13g2_fill_2 FILLER_51_522 ();
 sg13g2_fill_1 FILLER_51_529 ();
 sg13g2_fill_1 FILLER_51_560 ();
 sg13g2_fill_1 FILLER_51_566 ();
 sg13g2_fill_2 FILLER_51_593 ();
 sg13g2_fill_1 FILLER_51_623 ();
 sg13g2_fill_1 FILLER_51_629 ();
 sg13g2_fill_2 FILLER_51_647 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_fill_1 FILLER_51_695 ();
 sg13g2_fill_1 FILLER_51_724 ();
 sg13g2_fill_1 FILLER_51_729 ();
 sg13g2_decap_8 FILLER_51_740 ();
 sg13g2_decap_8 FILLER_51_747 ();
 sg13g2_decap_4 FILLER_51_754 ();
 sg13g2_fill_2 FILLER_51_769 ();
 sg13g2_fill_2 FILLER_51_793 ();
 sg13g2_fill_2 FILLER_51_805 ();
 sg13g2_fill_1 FILLER_51_807 ();
 sg13g2_decap_4 FILLER_51_854 ();
 sg13g2_fill_2 FILLER_51_877 ();
 sg13g2_decap_4 FILLER_51_921 ();
 sg13g2_fill_1 FILLER_51_967 ();
 sg13g2_fill_1 FILLER_51_973 ();
 sg13g2_decap_8 FILLER_51_983 ();
 sg13g2_fill_2 FILLER_51_994 ();
 sg13g2_decap_4 FILLER_51_1010 ();
 sg13g2_fill_1 FILLER_51_1014 ();
 sg13g2_decap_4 FILLER_51_1019 ();
 sg13g2_fill_1 FILLER_51_1023 ();
 sg13g2_fill_2 FILLER_51_1029 ();
 sg13g2_fill_1 FILLER_51_1031 ();
 sg13g2_fill_1 FILLER_51_1062 ();
 sg13g2_fill_2 FILLER_51_1163 ();
 sg13g2_fill_2 FILLER_51_1214 ();
 sg13g2_fill_2 FILLER_51_1236 ();
 sg13g2_fill_1 FILLER_51_1284 ();
 sg13g2_fill_1 FILLER_51_1295 ();
 sg13g2_fill_1 FILLER_51_1307 ();
 sg13g2_decap_8 FILLER_51_1316 ();
 sg13g2_decap_8 FILLER_51_1323 ();
 sg13g2_fill_1 FILLER_51_1330 ();
 sg13g2_decap_4 FILLER_51_1337 ();
 sg13g2_fill_1 FILLER_51_1341 ();
 sg13g2_fill_2 FILLER_51_1346 ();
 sg13g2_fill_1 FILLER_51_1348 ();
 sg13g2_fill_1 FILLER_51_1436 ();
 sg13g2_fill_1 FILLER_51_1462 ();
 sg13g2_fill_2 FILLER_51_1548 ();
 sg13g2_fill_1 FILLER_51_1550 ();
 sg13g2_decap_8 FILLER_51_1580 ();
 sg13g2_fill_1 FILLER_51_1621 ();
 sg13g2_decap_8 FILLER_51_1632 ();
 sg13g2_fill_2 FILLER_51_1639 ();
 sg13g2_fill_1 FILLER_51_1641 ();
 sg13g2_fill_2 FILLER_51_1652 ();
 sg13g2_fill_2 FILLER_51_1663 ();
 sg13g2_fill_2 FILLER_51_1678 ();
 sg13g2_fill_1 FILLER_51_1770 ();
 sg13g2_fill_2 FILLER_51_1817 ();
 sg13g2_fill_1 FILLER_51_1844 ();
 sg13g2_fill_2 FILLER_51_1875 ();
 sg13g2_fill_2 FILLER_51_1888 ();
 sg13g2_fill_2 FILLER_51_1919 ();
 sg13g2_fill_2 FILLER_51_1950 ();
 sg13g2_decap_8 FILLER_51_1998 ();
 sg13g2_fill_2 FILLER_51_2005 ();
 sg13g2_fill_1 FILLER_51_2007 ();
 sg13g2_fill_1 FILLER_51_2030 ();
 sg13g2_fill_1 FILLER_51_2035 ();
 sg13g2_fill_1 FILLER_51_2040 ();
 sg13g2_fill_2 FILLER_51_2061 ();
 sg13g2_fill_2 FILLER_51_2143 ();
 sg13g2_decap_8 FILLER_51_2164 ();
 sg13g2_decap_8 FILLER_51_2171 ();
 sg13g2_decap_8 FILLER_51_2178 ();
 sg13g2_fill_2 FILLER_51_2185 ();
 sg13g2_fill_1 FILLER_51_2187 ();
 sg13g2_fill_1 FILLER_51_2195 ();
 sg13g2_decap_8 FILLER_51_2210 ();
 sg13g2_fill_2 FILLER_51_2217 ();
 sg13g2_fill_1 FILLER_51_2249 ();
 sg13g2_fill_1 FILLER_51_2254 ();
 sg13g2_fill_1 FILLER_51_2259 ();
 sg13g2_fill_1 FILLER_51_2286 ();
 sg13g2_fill_1 FILLER_51_2325 ();
 sg13g2_decap_4 FILLER_51_2396 ();
 sg13g2_fill_1 FILLER_51_2400 ();
 sg13g2_fill_1 FILLER_51_2440 ();
 sg13g2_fill_1 FILLER_51_2523 ();
 sg13g2_fill_2 FILLER_51_2549 ();
 sg13g2_fill_1 FILLER_51_2551 ();
 sg13g2_decap_4 FILLER_51_2562 ();
 sg13g2_decap_8 FILLER_51_2610 ();
 sg13g2_decap_8 FILLER_51_2617 ();
 sg13g2_fill_1 FILLER_51_2624 ();
 sg13g2_decap_4 FILLER_51_2635 ();
 sg13g2_decap_4 FILLER_51_2665 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_33 ();
 sg13g2_decap_4 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_57 ();
 sg13g2_fill_2 FILLER_52_90 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_decap_8 FILLER_52_123 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_1 FILLER_52_139 ();
 sg13g2_fill_1 FILLER_52_155 ();
 sg13g2_fill_2 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_179 ();
 sg13g2_decap_4 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_decap_4 FILLER_52_194 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_204 ();
 sg13g2_fill_1 FILLER_52_209 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_244 ();
 sg13g2_decap_8 FILLER_52_251 ();
 sg13g2_fill_1 FILLER_52_258 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_295 ();
 sg13g2_fill_1 FILLER_52_297 ();
 sg13g2_fill_2 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_305 ();
 sg13g2_decap_8 FILLER_52_310 ();
 sg13g2_decap_8 FILLER_52_326 ();
 sg13g2_decap_4 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_4 FILLER_52_370 ();
 sg13g2_fill_1 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_398 ();
 sg13g2_fill_1 FILLER_52_400 ();
 sg13g2_decap_4 FILLER_52_417 ();
 sg13g2_decap_8 FILLER_52_426 ();
 sg13g2_decap_8 FILLER_52_433 ();
 sg13g2_fill_2 FILLER_52_440 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_decap_4 FILLER_52_460 ();
 sg13g2_fill_2 FILLER_52_487 ();
 sg13g2_fill_2 FILLER_52_543 ();
 sg13g2_fill_1 FILLER_52_554 ();
 sg13g2_fill_1 FILLER_52_575 ();
 sg13g2_fill_2 FILLER_52_585 ();
 sg13g2_fill_2 FILLER_52_596 ();
 sg13g2_fill_1 FILLER_52_615 ();
 sg13g2_fill_2 FILLER_52_643 ();
 sg13g2_fill_2 FILLER_52_674 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_fill_2 FILLER_52_693 ();
 sg13g2_fill_1 FILLER_52_695 ();
 sg13g2_fill_2 FILLER_52_700 ();
 sg13g2_fill_2 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_708 ();
 sg13g2_decap_4 FILLER_52_717 ();
 sg13g2_fill_2 FILLER_52_731 ();
 sg13g2_fill_2 FILLER_52_737 ();
 sg13g2_fill_2 FILLER_52_743 ();
 sg13g2_fill_2 FILLER_52_759 ();
 sg13g2_fill_2 FILLER_52_776 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_fill_1 FILLER_52_817 ();
 sg13g2_decap_4 FILLER_52_851 ();
 sg13g2_fill_2 FILLER_52_855 ();
 sg13g2_decap_8 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_52_868 ();
 sg13g2_fill_2 FILLER_52_875 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_fill_1 FILLER_52_888 ();
 sg13g2_fill_1 FILLER_52_917 ();
 sg13g2_fill_1 FILLER_52_923 ();
 sg13g2_fill_1 FILLER_52_928 ();
 sg13g2_fill_1 FILLER_52_934 ();
 sg13g2_fill_2 FILLER_52_940 ();
 sg13g2_fill_1 FILLER_52_950 ();
 sg13g2_fill_2 FILLER_52_957 ();
 sg13g2_fill_1 FILLER_52_964 ();
 sg13g2_fill_2 FILLER_52_973 ();
 sg13g2_fill_2 FILLER_52_979 ();
 sg13g2_decap_4 FILLER_52_993 ();
 sg13g2_decap_8 FILLER_52_1005 ();
 sg13g2_decap_8 FILLER_52_1012 ();
 sg13g2_fill_1 FILLER_52_1019 ();
 sg13g2_fill_1 FILLER_52_1027 ();
 sg13g2_fill_2 FILLER_52_1032 ();
 sg13g2_fill_1 FILLER_52_1034 ();
 sg13g2_fill_2 FILLER_52_1039 ();
 sg13g2_fill_1 FILLER_52_1041 ();
 sg13g2_decap_4 FILLER_52_1046 ();
 sg13g2_decap_8 FILLER_52_1054 ();
 sg13g2_fill_1 FILLER_52_1064 ();
 sg13g2_fill_2 FILLER_52_1109 ();
 sg13g2_fill_2 FILLER_52_1115 ();
 sg13g2_fill_2 FILLER_52_1129 ();
 sg13g2_fill_2 FILLER_52_1140 ();
 sg13g2_fill_2 FILLER_52_1156 ();
 sg13g2_fill_1 FILLER_52_1247 ();
 sg13g2_fill_1 FILLER_52_1306 ();
 sg13g2_fill_2 FILLER_52_1312 ();
 sg13g2_decap_4 FILLER_52_1344 ();
 sg13g2_decap_4 FILLER_52_1382 ();
 sg13g2_fill_1 FILLER_52_1390 ();
 sg13g2_fill_1 FILLER_52_1395 ();
 sg13g2_fill_2 FILLER_52_1401 ();
 sg13g2_fill_2 FILLER_52_1412 ();
 sg13g2_fill_1 FILLER_52_1414 ();
 sg13g2_fill_1 FILLER_52_1419 ();
 sg13g2_fill_2 FILLER_52_1430 ();
 sg13g2_fill_1 FILLER_52_1432 ();
 sg13g2_decap_8 FILLER_52_1441 ();
 sg13g2_decap_8 FILLER_52_1448 ();
 sg13g2_decap_8 FILLER_52_1455 ();
 sg13g2_fill_2 FILLER_52_1462 ();
 sg13g2_decap_4 FILLER_52_1470 ();
 sg13g2_decap_8 FILLER_52_1525 ();
 sg13g2_decap_4 FILLER_52_1532 ();
 sg13g2_fill_1 FILLER_52_1540 ();
 sg13g2_fill_1 FILLER_52_1567 ();
 sg13g2_fill_2 FILLER_52_1572 ();
 sg13g2_fill_2 FILLER_52_1581 ();
 sg13g2_fill_2 FILLER_52_1596 ();
 sg13g2_fill_1 FILLER_52_1598 ();
 sg13g2_fill_1 FILLER_52_1608 ();
 sg13g2_fill_1 FILLER_52_1653 ();
 sg13g2_decap_8 FILLER_52_1668 ();
 sg13g2_fill_1 FILLER_52_1678 ();
 sg13g2_fill_2 FILLER_52_1687 ();
 sg13g2_fill_1 FILLER_52_1689 ();
 sg13g2_fill_1 FILLER_52_1750 ();
 sg13g2_fill_2 FILLER_52_1829 ();
 sg13g2_fill_1 FILLER_52_1870 ();
 sg13g2_fill_2 FILLER_52_1906 ();
 sg13g2_fill_2 FILLER_52_2016 ();
 sg13g2_fill_1 FILLER_52_2048 ();
 sg13g2_fill_2 FILLER_52_2073 ();
 sg13g2_fill_1 FILLER_52_2143 ();
 sg13g2_fill_1 FILLER_52_2158 ();
 sg13g2_fill_1 FILLER_52_2195 ();
 sg13g2_decap_4 FILLER_52_2223 ();
 sg13g2_fill_2 FILLER_52_2227 ();
 sg13g2_fill_2 FILLER_52_2234 ();
 sg13g2_fill_2 FILLER_52_2240 ();
 sg13g2_fill_1 FILLER_52_2242 ();
 sg13g2_decap_4 FILLER_52_2263 ();
 sg13g2_fill_2 FILLER_52_2267 ();
 sg13g2_fill_2 FILLER_52_2324 ();
 sg13g2_fill_1 FILLER_52_2388 ();
 sg13g2_fill_1 FILLER_52_2393 ();
 sg13g2_fill_1 FILLER_52_2420 ();
 sg13g2_fill_1 FILLER_52_2447 ();
 sg13g2_fill_2 FILLER_52_2458 ();
 sg13g2_fill_2 FILLER_52_2550 ();
 sg13g2_fill_1 FILLER_52_2552 ();
 sg13g2_fill_2 FILLER_52_2599 ();
 sg13g2_fill_1 FILLER_52_2601 ();
 sg13g2_decap_4 FILLER_52_2664 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_1 FILLER_53_62 ();
 sg13g2_fill_2 FILLER_53_71 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_decap_8 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_85 ();
 sg13g2_fill_2 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_125 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_decap_8 FILLER_53_132 ();
 sg13g2_decap_8 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_fill_1 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_214 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_2 FILLER_53_252 ();
 sg13g2_fill_2 FILLER_53_267 ();
 sg13g2_fill_1 FILLER_53_278 ();
 sg13g2_decap_8 FILLER_53_342 ();
 sg13g2_fill_2 FILLER_53_349 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_fill_1 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_372 ();
 sg13g2_fill_2 FILLER_53_378 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_53_436 ();
 sg13g2_fill_1 FILLER_53_443 ();
 sg13g2_decap_8 FILLER_53_447 ();
 sg13g2_decap_8 FILLER_53_454 ();
 sg13g2_fill_2 FILLER_53_461 ();
 sg13g2_fill_1 FILLER_53_463 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_2 FILLER_53_496 ();
 sg13g2_fill_2 FILLER_53_508 ();
 sg13g2_fill_2 FILLER_53_545 ();
 sg13g2_fill_1 FILLER_53_555 ();
 sg13g2_fill_2 FILLER_53_560 ();
 sg13g2_fill_1 FILLER_53_578 ();
 sg13g2_fill_2 FILLER_53_593 ();
 sg13g2_fill_1 FILLER_53_696 ();
 sg13g2_fill_1 FILLER_53_770 ();
 sg13g2_fill_2 FILLER_53_791 ();
 sg13g2_fill_2 FILLER_53_811 ();
 sg13g2_fill_2 FILLER_53_825 ();
 sg13g2_fill_2 FILLER_53_832 ();
 sg13g2_fill_2 FILLER_53_838 ();
 sg13g2_decap_8 FILLER_53_844 ();
 sg13g2_fill_1 FILLER_53_886 ();
 sg13g2_fill_2 FILLER_53_913 ();
 sg13g2_decap_4 FILLER_53_938 ();
 sg13g2_fill_1 FILLER_53_1004 ();
 sg13g2_fill_1 FILLER_53_1019 ();
 sg13g2_decap_8 FILLER_53_1024 ();
 sg13g2_decap_4 FILLER_53_1031 ();
 sg13g2_fill_1 FILLER_53_1035 ();
 sg13g2_fill_2 FILLER_53_1051 ();
 sg13g2_fill_2 FILLER_53_1066 ();
 sg13g2_fill_1 FILLER_53_1084 ();
 sg13g2_fill_2 FILLER_53_1093 ();
 sg13g2_fill_2 FILLER_53_1100 ();
 sg13g2_fill_1 FILLER_53_1133 ();
 sg13g2_fill_2 FILLER_53_1140 ();
 sg13g2_fill_2 FILLER_53_1154 ();
 sg13g2_fill_2 FILLER_53_1166 ();
 sg13g2_fill_1 FILLER_53_1194 ();
 sg13g2_fill_1 FILLER_53_1199 ();
 sg13g2_fill_2 FILLER_53_1204 ();
 sg13g2_fill_2 FILLER_53_1256 ();
 sg13g2_fill_1 FILLER_53_1281 ();
 sg13g2_fill_2 FILLER_53_1293 ();
 sg13g2_decap_8 FILLER_53_1368 ();
 sg13g2_decap_4 FILLER_53_1375 ();
 sg13g2_fill_2 FILLER_53_1379 ();
 sg13g2_fill_1 FILLER_53_1387 ();
 sg13g2_decap_8 FILLER_53_1395 ();
 sg13g2_decap_4 FILLER_53_1402 ();
 sg13g2_decap_8 FILLER_53_1416 ();
 sg13g2_fill_2 FILLER_53_1423 ();
 sg13g2_decap_8 FILLER_53_1429 ();
 sg13g2_decap_8 FILLER_53_1436 ();
 sg13g2_fill_2 FILLER_53_1443 ();
 sg13g2_fill_1 FILLER_53_1445 ();
 sg13g2_decap_4 FILLER_53_1454 ();
 sg13g2_fill_2 FILLER_53_1458 ();
 sg13g2_decap_4 FILLER_53_1499 ();
 sg13g2_fill_1 FILLER_53_1503 ();
 sg13g2_decap_8 FILLER_53_1508 ();
 sg13g2_decap_8 FILLER_53_1515 ();
 sg13g2_decap_8 FILLER_53_1522 ();
 sg13g2_decap_8 FILLER_53_1529 ();
 sg13g2_fill_2 FILLER_53_1536 ();
 sg13g2_fill_2 FILLER_53_1550 ();
 sg13g2_fill_1 FILLER_53_1552 ();
 sg13g2_decap_4 FILLER_53_1561 ();
 sg13g2_decap_4 FILLER_53_1570 ();
 sg13g2_fill_2 FILLER_53_1574 ();
 sg13g2_decap_8 FILLER_53_1586 ();
 sg13g2_fill_2 FILLER_53_1593 ();
 sg13g2_fill_1 FILLER_53_1595 ();
 sg13g2_fill_2 FILLER_53_1655 ();
 sg13g2_fill_1 FILLER_53_1699 ();
 sg13g2_fill_1 FILLER_53_1714 ();
 sg13g2_fill_2 FILLER_53_1742 ();
 sg13g2_fill_1 FILLER_53_1771 ();
 sg13g2_decap_4 FILLER_53_1851 ();
 sg13g2_fill_2 FILLER_53_1897 ();
 sg13g2_fill_1 FILLER_53_1961 ();
 sg13g2_fill_1 FILLER_53_1988 ();
 sg13g2_fill_2 FILLER_53_2002 ();
 sg13g2_fill_1 FILLER_53_2011 ();
 sg13g2_fill_1 FILLER_53_2025 ();
 sg13g2_fill_2 FILLER_53_2060 ();
 sg13g2_fill_1 FILLER_53_2078 ();
 sg13g2_fill_2 FILLER_53_2098 ();
 sg13g2_fill_1 FILLER_53_2136 ();
 sg13g2_fill_1 FILLER_53_2191 ();
 sg13g2_fill_1 FILLER_53_2203 ();
 sg13g2_fill_1 FILLER_53_2208 ();
 sg13g2_decap_8 FILLER_53_2237 ();
 sg13g2_fill_1 FILLER_53_2244 ();
 sg13g2_fill_2 FILLER_53_2249 ();
 sg13g2_decap_8 FILLER_53_2261 ();
 sg13g2_fill_1 FILLER_53_2268 ();
 sg13g2_decap_8 FILLER_53_2274 ();
 sg13g2_fill_1 FILLER_53_2281 ();
 sg13g2_fill_1 FILLER_53_2355 ();
 sg13g2_fill_1 FILLER_53_2399 ();
 sg13g2_decap_4 FILLER_53_2410 ();
 sg13g2_fill_1 FILLER_53_2414 ();
 sg13g2_fill_2 FILLER_53_2418 ();
 sg13g2_fill_1 FILLER_53_2424 ();
 sg13g2_fill_1 FILLER_53_2471 ();
 sg13g2_decap_8 FILLER_53_2489 ();
 sg13g2_decap_4 FILLER_53_2496 ();
 sg13g2_fill_2 FILLER_53_2500 ();
 sg13g2_fill_2 FILLER_53_2519 ();
 sg13g2_fill_1 FILLER_53_2547 ();
 sg13g2_fill_2 FILLER_53_2601 ();
 sg13g2_fill_1 FILLER_53_2603 ();
 sg13g2_decap_8 FILLER_53_2630 ();
 sg13g2_decap_4 FILLER_53_2637 ();
 sg13g2_decap_8 FILLER_53_2649 ();
 sg13g2_decap_8 FILLER_53_2656 ();
 sg13g2_decap_8 FILLER_53_2663 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_36 ();
 sg13g2_fill_2 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_69 ();
 sg13g2_decap_4 FILLER_54_76 ();
 sg13g2_fill_2 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_216 ();
 sg13g2_fill_2 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_fill_1 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_393 ();
 sg13g2_fill_2 FILLER_54_400 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_54_416 ();
 sg13g2_decap_8 FILLER_54_423 ();
 sg13g2_fill_2 FILLER_54_496 ();
 sg13g2_fill_1 FILLER_54_506 ();
 sg13g2_fill_2 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_597 ();
 sg13g2_fill_1 FILLER_54_606 ();
 sg13g2_fill_1 FILLER_54_612 ();
 sg13g2_fill_2 FILLER_54_639 ();
 sg13g2_fill_1 FILLER_54_696 ();
 sg13g2_fill_2 FILLER_54_723 ();
 sg13g2_fill_1 FILLER_54_725 ();
 sg13g2_fill_1 FILLER_54_772 ();
 sg13g2_fill_1 FILLER_54_806 ();
 sg13g2_fill_1 FILLER_54_811 ();
 sg13g2_fill_2 FILLER_54_816 ();
 sg13g2_fill_2 FILLER_54_823 ();
 sg13g2_decap_4 FILLER_54_832 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_decap_4 FILLER_54_846 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_decap_8 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_54_868 ();
 sg13g2_fill_1 FILLER_54_896 ();
 sg13g2_fill_1 FILLER_54_915 ();
 sg13g2_fill_2 FILLER_54_920 ();
 sg13g2_fill_2 FILLER_54_930 ();
 sg13g2_fill_2 FILLER_54_938 ();
 sg13g2_decap_8 FILLER_54_962 ();
 sg13g2_fill_1 FILLER_54_969 ();
 sg13g2_fill_2 FILLER_54_999 ();
 sg13g2_fill_2 FILLER_54_1009 ();
 sg13g2_fill_1 FILLER_54_1011 ();
 sg13g2_fill_1 FILLER_54_1027 ();
 sg13g2_fill_2 FILLER_54_1038 ();
 sg13g2_decap_8 FILLER_54_1044 ();
 sg13g2_decap_4 FILLER_54_1051 ();
 sg13g2_fill_1 FILLER_54_1055 ();
 sg13g2_fill_1 FILLER_54_1066 ();
 sg13g2_fill_2 FILLER_54_1077 ();
 sg13g2_fill_1 FILLER_54_1099 ();
 sg13g2_fill_2 FILLER_54_1116 ();
 sg13g2_fill_2 FILLER_54_1147 ();
 sg13g2_fill_1 FILLER_54_1176 ();
 sg13g2_fill_1 FILLER_54_1186 ();
 sg13g2_fill_2 FILLER_54_1231 ();
 sg13g2_fill_2 FILLER_54_1265 ();
 sg13g2_fill_1 FILLER_54_1272 ();
 sg13g2_fill_1 FILLER_54_1276 ();
 sg13g2_fill_2 FILLER_54_1287 ();
 sg13g2_fill_1 FILLER_54_1294 ();
 sg13g2_decap_4 FILLER_54_1345 ();
 sg13g2_fill_1 FILLER_54_1349 ();
 sg13g2_fill_1 FILLER_54_1374 ();
 sg13g2_fill_2 FILLER_54_1419 ();
 sg13g2_fill_1 FILLER_54_1421 ();
 sg13g2_decap_4 FILLER_54_1453 ();
 sg13g2_fill_1 FILLER_54_1457 ();
 sg13g2_fill_2 FILLER_54_1488 ();
 sg13g2_fill_1 FILLER_54_1490 ();
 sg13g2_decap_8 FILLER_54_1495 ();
 sg13g2_decap_8 FILLER_54_1502 ();
 sg13g2_decap_4 FILLER_54_1509 ();
 sg13g2_fill_2 FILLER_54_1513 ();
 sg13g2_decap_4 FILLER_54_1520 ();
 sg13g2_decap_8 FILLER_54_1567 ();
 sg13g2_decap_8 FILLER_54_1574 ();
 sg13g2_decap_8 FILLER_54_1581 ();
 sg13g2_fill_2 FILLER_54_1588 ();
 sg13g2_fill_1 FILLER_54_1590 ();
 sg13g2_fill_2 FILLER_54_1640 ();
 sg13g2_fill_2 FILLER_54_1645 ();
 sg13g2_fill_1 FILLER_54_1647 ();
 sg13g2_fill_1 FILLER_54_1661 ();
 sg13g2_fill_1 FILLER_54_1665 ();
 sg13g2_fill_1 FILLER_54_1702 ();
 sg13g2_fill_1 FILLER_54_1763 ();
 sg13g2_fill_2 FILLER_54_1802 ();
 sg13g2_fill_1 FILLER_54_1838 ();
 sg13g2_decap_4 FILLER_54_1843 ();
 sg13g2_fill_1 FILLER_54_1851 ();
 sg13g2_fill_2 FILLER_54_1856 ();
 sg13g2_fill_1 FILLER_54_1858 ();
 sg13g2_fill_2 FILLER_54_1869 ();
 sg13g2_fill_1 FILLER_54_1871 ();
 sg13g2_fill_2 FILLER_54_1893 ();
 sg13g2_fill_2 FILLER_54_1905 ();
 sg13g2_fill_1 FILLER_54_1955 ();
 sg13g2_fill_1 FILLER_54_2015 ();
 sg13g2_fill_2 FILLER_54_2020 ();
 sg13g2_fill_1 FILLER_54_2032 ();
 sg13g2_fill_2 FILLER_54_2043 ();
 sg13g2_fill_1 FILLER_54_2048 ();
 sg13g2_fill_1 FILLER_54_2057 ();
 sg13g2_fill_2 FILLER_54_2088 ();
 sg13g2_fill_1 FILLER_54_2100 ();
 sg13g2_decap_4 FILLER_54_2200 ();
 sg13g2_fill_1 FILLER_54_2230 ();
 sg13g2_fill_2 FILLER_54_2244 ();
 sg13g2_fill_1 FILLER_54_2256 ();
 sg13g2_fill_1 FILLER_54_2283 ();
 sg13g2_fill_2 FILLER_54_2310 ();
 sg13g2_fill_2 FILLER_54_2316 ();
 sg13g2_fill_1 FILLER_54_2354 ();
 sg13g2_decap_8 FILLER_54_2395 ();
 sg13g2_decap_8 FILLER_54_2402 ();
 sg13g2_decap_4 FILLER_54_2409 ();
 sg13g2_fill_2 FILLER_54_2413 ();
 sg13g2_fill_2 FILLER_54_2442 ();
 sg13g2_decap_4 FILLER_54_2450 ();
 sg13g2_fill_2 FILLER_54_2454 ();
 sg13g2_decap_4 FILLER_54_2464 ();
 sg13g2_decap_8 FILLER_54_2497 ();
 sg13g2_fill_1 FILLER_54_2504 ();
 sg13g2_fill_1 FILLER_54_2508 ();
 sg13g2_decap_8 FILLER_54_2586 ();
 sg13g2_decap_8 FILLER_54_2593 ();
 sg13g2_decap_8 FILLER_54_2600 ();
 sg13g2_fill_2 FILLER_54_2607 ();
 sg13g2_fill_2 FILLER_54_2617 ();
 sg13g2_decap_8 FILLER_54_2640 ();
 sg13g2_decap_8 FILLER_54_2647 ();
 sg13g2_decap_8 FILLER_54_2654 ();
 sg13g2_decap_8 FILLER_54_2661 ();
 sg13g2_fill_2 FILLER_54_2668 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_73 ();
 sg13g2_decap_8 FILLER_55_80 ();
 sg13g2_fill_2 FILLER_55_87 ();
 sg13g2_fill_1 FILLER_55_115 ();
 sg13g2_decap_8 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_145 ();
 sg13g2_fill_2 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_185 ();
 sg13g2_fill_2 FILLER_55_196 ();
 sg13g2_fill_1 FILLER_55_224 ();
 sg13g2_fill_2 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_278 ();
 sg13g2_fill_2 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_55_416 ();
 sg13g2_fill_1 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_436 ();
 sg13g2_fill_2 FILLER_55_509 ();
 sg13g2_fill_1 FILLER_55_525 ();
 sg13g2_fill_2 FILLER_55_531 ();
 sg13g2_fill_2 FILLER_55_603 ();
 sg13g2_fill_2 FILLER_55_610 ();
 sg13g2_fill_1 FILLER_55_620 ();
 sg13g2_fill_1 FILLER_55_625 ();
 sg13g2_fill_1 FILLER_55_631 ();
 sg13g2_decap_4 FILLER_55_639 ();
 sg13g2_fill_1 FILLER_55_698 ();
 sg13g2_fill_2 FILLER_55_771 ();
 sg13g2_fill_2 FILLER_55_790 ();
 sg13g2_fill_1 FILLER_55_817 ();
 sg13g2_fill_1 FILLER_55_841 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_890 ();
 sg13g2_fill_1 FILLER_55_892 ();
 sg13g2_decap_8 FILLER_55_924 ();
 sg13g2_decap_8 FILLER_55_931 ();
 sg13g2_decap_4 FILLER_55_938 ();
 sg13g2_fill_1 FILLER_55_942 ();
 sg13g2_decap_4 FILLER_55_957 ();
 sg13g2_fill_2 FILLER_55_961 ();
 sg13g2_fill_1 FILLER_55_967 ();
 sg13g2_fill_2 FILLER_55_972 ();
 sg13g2_fill_1 FILLER_55_978 ();
 sg13g2_fill_2 FILLER_55_1026 ();
 sg13g2_fill_2 FILLER_55_1032 ();
 sg13g2_decap_8 FILLER_55_1038 ();
 sg13g2_decap_4 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1049 ();
 sg13g2_fill_1 FILLER_55_1088 ();
 sg13g2_fill_1 FILLER_55_1102 ();
 sg13g2_fill_2 FILLER_55_1139 ();
 sg13g2_fill_2 FILLER_55_1154 ();
 sg13g2_fill_2 FILLER_55_1171 ();
 sg13g2_fill_1 FILLER_55_1185 ();
 sg13g2_fill_2 FILLER_55_1206 ();
 sg13g2_fill_1 FILLER_55_1219 ();
 sg13g2_fill_2 FILLER_55_1233 ();
 sg13g2_fill_1 FILLER_55_1260 ();
 sg13g2_fill_2 FILLER_55_1311 ();
 sg13g2_fill_2 FILLER_55_1326 ();
 sg13g2_fill_1 FILLER_55_1328 ();
 sg13g2_decap_8 FILLER_55_1335 ();
 sg13g2_decap_8 FILLER_55_1342 ();
 sg13g2_decap_4 FILLER_55_1349 ();
 sg13g2_fill_2 FILLER_55_1379 ();
 sg13g2_fill_1 FILLER_55_1393 ();
 sg13g2_fill_2 FILLER_55_1490 ();
 sg13g2_fill_1 FILLER_55_1492 ();
 sg13g2_decap_8 FILLER_55_1498 ();
 sg13g2_decap_4 FILLER_55_1505 ();
 sg13g2_fill_2 FILLER_55_1509 ();
 sg13g2_decap_4 FILLER_55_1564 ();
 sg13g2_fill_2 FILLER_55_1568 ();
 sg13g2_fill_1 FILLER_55_1614 ();
 sg13g2_fill_1 FILLER_55_1632 ();
 sg13g2_decap_8 FILLER_55_1698 ();
 sg13g2_fill_2 FILLER_55_1705 ();
 sg13g2_fill_1 FILLER_55_1707 ();
 sg13g2_fill_2 FILLER_55_1713 ();
 sg13g2_fill_2 FILLER_55_1749 ();
 sg13g2_fill_1 FILLER_55_1814 ();
 sg13g2_decap_8 FILLER_55_1859 ();
 sg13g2_decap_4 FILLER_55_1866 ();
 sg13g2_fill_1 FILLER_55_1870 ();
 sg13g2_decap_4 FILLER_55_1881 ();
 sg13g2_fill_2 FILLER_55_1885 ();
 sg13g2_fill_2 FILLER_55_1903 ();
 sg13g2_fill_2 FILLER_55_1908 ();
 sg13g2_fill_2 FILLER_55_1979 ();
 sg13g2_fill_2 FILLER_55_2007 ();
 sg13g2_fill_2 FILLER_55_2038 ();
 sg13g2_fill_1 FILLER_55_2058 ();
 sg13g2_fill_1 FILLER_55_2083 ();
 sg13g2_fill_1 FILLER_55_2102 ();
 sg13g2_fill_1 FILLER_55_2108 ();
 sg13g2_fill_2 FILLER_55_2120 ();
 sg13g2_fill_1 FILLER_55_2168 ();
 sg13g2_fill_1 FILLER_55_2201 ();
 sg13g2_decap_8 FILLER_55_2210 ();
 sg13g2_decap_4 FILLER_55_2217 ();
 sg13g2_fill_2 FILLER_55_2221 ();
 sg13g2_fill_1 FILLER_55_2231 ();
 sg13g2_fill_2 FILLER_55_2266 ();
 sg13g2_decap_4 FILLER_55_2272 ();
 sg13g2_decap_8 FILLER_55_2306 ();
 sg13g2_decap_8 FILLER_55_2313 ();
 sg13g2_decap_8 FILLER_55_2320 ();
 sg13g2_fill_2 FILLER_55_2327 ();
 sg13g2_fill_2 FILLER_55_2333 ();
 sg13g2_decap_8 FILLER_55_2343 ();
 sg13g2_decap_4 FILLER_55_2350 ();
 sg13g2_fill_1 FILLER_55_2375 ();
 sg13g2_fill_2 FILLER_55_2404 ();
 sg13g2_fill_1 FILLER_55_2411 ();
 sg13g2_fill_2 FILLER_55_2458 ();
 sg13g2_decap_8 FILLER_55_2470 ();
 sg13g2_fill_2 FILLER_55_2477 ();
 sg13g2_decap_4 FILLER_55_2509 ();
 sg13g2_fill_1 FILLER_55_2513 ();
 sg13g2_fill_1 FILLER_55_2518 ();
 sg13g2_decap_4 FILLER_55_2545 ();
 sg13g2_decap_8 FILLER_55_2612 ();
 sg13g2_decap_8 FILLER_55_2619 ();
 sg13g2_fill_1 FILLER_55_2647 ();
 sg13g2_decap_8 FILLER_55_2652 ();
 sg13g2_decap_8 FILLER_55_2659 ();
 sg13g2_decap_4 FILLER_55_2666 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_47 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_125 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_187 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_fill_2 FILLER_56_217 ();
 sg13g2_fill_2 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_279 ();
 sg13g2_fill_2 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_fill_1 FILLER_56_378 ();
 sg13g2_fill_2 FILLER_56_384 ();
 sg13g2_fill_1 FILLER_56_392 ();
 sg13g2_fill_2 FILLER_56_404 ();
 sg13g2_decap_4 FILLER_56_414 ();
 sg13g2_fill_1 FILLER_56_446 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_1 FILLER_56_511 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_553 ();
 sg13g2_fill_2 FILLER_56_570 ();
 sg13g2_fill_2 FILLER_56_588 ();
 sg13g2_fill_1 FILLER_56_595 ();
 sg13g2_fill_1 FILLER_56_611 ();
 sg13g2_fill_2 FILLER_56_615 ();
 sg13g2_fill_1 FILLER_56_627 ();
 sg13g2_decap_8 FILLER_56_638 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_fill_1 FILLER_56_765 ();
 sg13g2_fill_1 FILLER_56_791 ();
 sg13g2_fill_1 FILLER_56_818 ();
 sg13g2_fill_2 FILLER_56_825 ();
 sg13g2_fill_2 FILLER_56_836 ();
 sg13g2_decap_8 FILLER_56_847 ();
 sg13g2_decap_4 FILLER_56_854 ();
 sg13g2_fill_1 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_867 ();
 sg13g2_fill_2 FILLER_56_873 ();
 sg13g2_fill_1 FILLER_56_875 ();
 sg13g2_fill_2 FILLER_56_881 ();
 sg13g2_decap_8 FILLER_56_887 ();
 sg13g2_decap_8 FILLER_56_894 ();
 sg13g2_decap_8 FILLER_56_905 ();
 sg13g2_decap_8 FILLER_56_921 ();
 sg13g2_decap_8 FILLER_56_928 ();
 sg13g2_decap_8 FILLER_56_935 ();
 sg13g2_decap_8 FILLER_56_942 ();
 sg13g2_decap_8 FILLER_56_949 ();
 sg13g2_fill_2 FILLER_56_985 ();
 sg13g2_fill_1 FILLER_56_1050 ();
 sg13g2_fill_1 FILLER_56_1103 ();
 sg13g2_fill_1 FILLER_56_1117 ();
 sg13g2_fill_1 FILLER_56_1123 ();
 sg13g2_fill_1 FILLER_56_1129 ();
 sg13g2_fill_2 FILLER_56_1134 ();
 sg13g2_fill_1 FILLER_56_1145 ();
 sg13g2_fill_1 FILLER_56_1150 ();
 sg13g2_fill_2 FILLER_56_1158 ();
 sg13g2_fill_1 FILLER_56_1171 ();
 sg13g2_fill_2 FILLER_56_1181 ();
 sg13g2_fill_2 FILLER_56_1193 ();
 sg13g2_fill_1 FILLER_56_1219 ();
 sg13g2_fill_2 FILLER_56_1251 ();
 sg13g2_fill_2 FILLER_56_1260 ();
 sg13g2_fill_2 FILLER_56_1267 ();
 sg13g2_fill_1 FILLER_56_1277 ();
 sg13g2_fill_2 FILLER_56_1304 ();
 sg13g2_fill_1 FILLER_56_1306 ();
 sg13g2_decap_4 FILLER_56_1311 ();
 sg13g2_fill_2 FILLER_56_1368 ();
 sg13g2_fill_2 FILLER_56_1380 ();
 sg13g2_fill_2 FILLER_56_1389 ();
 sg13g2_decap_8 FILLER_56_1450 ();
 sg13g2_fill_2 FILLER_56_1457 ();
 sg13g2_fill_1 FILLER_56_1459 ();
 sg13g2_fill_2 FILLER_56_1465 ();
 sg13g2_fill_2 FILLER_56_1476 ();
 sg13g2_fill_1 FILLER_56_1486 ();
 sg13g2_decap_4 FILLER_56_1491 ();
 sg13g2_fill_1 FILLER_56_1529 ();
 sg13g2_fill_2 FILLER_56_1556 ();
 sg13g2_fill_2 FILLER_56_1563 ();
 sg13g2_fill_1 FILLER_56_1565 ();
 sg13g2_fill_2 FILLER_56_1614 ();
 sg13g2_fill_2 FILLER_56_1629 ();
 sg13g2_fill_1 FILLER_56_1638 ();
 sg13g2_fill_1 FILLER_56_1665 ();
 sg13g2_fill_2 FILLER_56_1677 ();
 sg13g2_decap_4 FILLER_56_1690 ();
 sg13g2_decap_4 FILLER_56_1763 ();
 sg13g2_fill_2 FILLER_56_1767 ();
 sg13g2_fill_2 FILLER_56_1773 ();
 sg13g2_fill_2 FILLER_56_1781 ();
 sg13g2_fill_2 FILLER_56_1787 ();
 sg13g2_decap_8 FILLER_56_1832 ();
 sg13g2_fill_1 FILLER_56_1839 ();
 sg13g2_decap_8 FILLER_56_1848 ();
 sg13g2_fill_1 FILLER_56_1855 ();
 sg13g2_fill_1 FILLER_56_1882 ();
 sg13g2_fill_1 FILLER_56_1893 ();
 sg13g2_fill_2 FILLER_56_1989 ();
 sg13g2_fill_1 FILLER_56_1991 ();
 sg13g2_fill_1 FILLER_56_2050 ();
 sg13g2_fill_1 FILLER_56_2056 ();
 sg13g2_fill_1 FILLER_56_2063 ();
 sg13g2_fill_1 FILLER_56_2069 ();
 sg13g2_fill_1 FILLER_56_2102 ();
 sg13g2_fill_1 FILLER_56_2107 ();
 sg13g2_fill_2 FILLER_56_2112 ();
 sg13g2_fill_1 FILLER_56_2134 ();
 sg13g2_fill_2 FILLER_56_2160 ();
 sg13g2_fill_1 FILLER_56_2205 ();
 sg13g2_decap_4 FILLER_56_2217 ();
 sg13g2_fill_2 FILLER_56_2221 ();
 sg13g2_fill_1 FILLER_56_2227 ();
 sg13g2_fill_1 FILLER_56_2236 ();
 sg13g2_decap_8 FILLER_56_2263 ();
 sg13g2_fill_2 FILLER_56_2313 ();
 sg13g2_fill_2 FILLER_56_2350 ();
 sg13g2_decap_4 FILLER_56_2402 ();
 sg13g2_fill_2 FILLER_56_2419 ();
 sg13g2_fill_2 FILLER_56_2424 ();
 sg13g2_fill_2 FILLER_56_2439 ();
 sg13g2_fill_2 FILLER_56_2445 ();
 sg13g2_fill_2 FILLER_56_2452 ();
 sg13g2_fill_2 FILLER_56_2459 ();
 sg13g2_fill_1 FILLER_56_2461 ();
 sg13g2_decap_8 FILLER_56_2498 ();
 sg13g2_decap_8 FILLER_56_2508 ();
 sg13g2_fill_2 FILLER_56_2519 ();
 sg13g2_fill_2 FILLER_56_2525 ();
 sg13g2_fill_2 FILLER_56_2531 ();
 sg13g2_fill_2 FILLER_56_2543 ();
 sg13g2_decap_8 FILLER_56_2559 ();
 sg13g2_fill_2 FILLER_56_2566 ();
 sg13g2_decap_8 FILLER_56_2594 ();
 sg13g2_fill_1 FILLER_56_2601 ();
 sg13g2_fill_2 FILLER_56_2628 ();
 sg13g2_fill_1 FILLER_56_2630 ();
 sg13g2_fill_2 FILLER_56_2667 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_15 ();
 sg13g2_decap_8 FILLER_57_22 ();
 sg13g2_fill_1 FILLER_57_29 ();
 sg13g2_decap_4 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_39 ();
 sg13g2_fill_2 FILLER_57_51 ();
 sg13g2_fill_1 FILLER_57_53 ();
 sg13g2_decap_4 FILLER_57_71 ();
 sg13g2_fill_2 FILLER_57_115 ();
 sg13g2_fill_1 FILLER_57_121 ();
 sg13g2_decap_8 FILLER_57_152 ();
 sg13g2_decap_4 FILLER_57_159 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_decap_4 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_202 ();
 sg13g2_decap_4 FILLER_57_209 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_4 FILLER_57_224 ();
 sg13g2_fill_2 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_333 ();
 sg13g2_decap_8 FILLER_57_340 ();
 sg13g2_decap_8 FILLER_57_347 ();
 sg13g2_decap_4 FILLER_57_354 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_4 FILLER_57_375 ();
 sg13g2_decap_4 FILLER_57_399 ();
 sg13g2_fill_1 FILLER_57_403 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_fill_1 FILLER_57_434 ();
 sg13g2_fill_2 FILLER_57_442 ();
 sg13g2_fill_1 FILLER_57_453 ();
 sg13g2_decap_4 FILLER_57_458 ();
 sg13g2_fill_2 FILLER_57_462 ();
 sg13g2_fill_1 FILLER_57_472 ();
 sg13g2_fill_2 FILLER_57_493 ();
 sg13g2_fill_1 FILLER_57_550 ();
 sg13g2_fill_1 FILLER_57_612 ();
 sg13g2_fill_2 FILLER_57_621 ();
 sg13g2_fill_2 FILLER_57_636 ();
 sg13g2_fill_1 FILLER_57_638 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_decap_8 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_fill_2 FILLER_57_700 ();
 sg13g2_fill_1 FILLER_57_702 ();
 sg13g2_fill_1 FILLER_57_721 ();
 sg13g2_fill_2 FILLER_57_761 ();
 sg13g2_fill_1 FILLER_57_767 ();
 sg13g2_fill_2 FILLER_57_781 ();
 sg13g2_fill_2 FILLER_57_789 ();
 sg13g2_fill_1 FILLER_57_800 ();
 sg13g2_fill_1 FILLER_57_805 ();
 sg13g2_fill_2 FILLER_57_812 ();
 sg13g2_fill_1 FILLER_57_814 ();
 sg13g2_decap_4 FILLER_57_830 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_8 FILLER_57_857 ();
 sg13g2_decap_4 FILLER_57_864 ();
 sg13g2_decap_8 FILLER_57_873 ();
 sg13g2_decap_8 FILLER_57_880 ();
 sg13g2_decap_8 FILLER_57_887 ();
 sg13g2_decap_8 FILLER_57_898 ();
 sg13g2_fill_2 FILLER_57_910 ();
 sg13g2_fill_1 FILLER_57_912 ();
 sg13g2_decap_8 FILLER_57_917 ();
 sg13g2_decap_8 FILLER_57_924 ();
 sg13g2_fill_2 FILLER_57_931 ();
 sg13g2_fill_1 FILLER_57_933 ();
 sg13g2_decap_8 FILLER_57_944 ();
 sg13g2_decap_8 FILLER_57_951 ();
 sg13g2_decap_8 FILLER_57_958 ();
 sg13g2_decap_8 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_972 ();
 sg13g2_decap_8 FILLER_57_979 ();
 sg13g2_decap_8 FILLER_57_986 ();
 sg13g2_decap_8 FILLER_57_993 ();
 sg13g2_decap_4 FILLER_57_1008 ();
 sg13g2_fill_1 FILLER_57_1012 ();
 sg13g2_decap_8 FILLER_57_1017 ();
 sg13g2_decap_8 FILLER_57_1024 ();
 sg13g2_fill_2 FILLER_57_1031 ();
 sg13g2_decap_8 FILLER_57_1038 ();
 sg13g2_decap_8 FILLER_57_1045 ();
 sg13g2_fill_2 FILLER_57_1052 ();
 sg13g2_fill_1 FILLER_57_1059 ();
 sg13g2_fill_2 FILLER_57_1065 ();
 sg13g2_fill_2 FILLER_57_1071 ();
 sg13g2_fill_2 FILLER_57_1079 ();
 sg13g2_fill_1 FILLER_57_1081 ();
 sg13g2_fill_1 FILLER_57_1139 ();
 sg13g2_fill_1 FILLER_57_1145 ();
 sg13g2_fill_1 FILLER_57_1151 ();
 sg13g2_fill_2 FILLER_57_1174 ();
 sg13g2_fill_1 FILLER_57_1191 ();
 sg13g2_fill_2 FILLER_57_1206 ();
 sg13g2_fill_1 FILLER_57_1230 ();
 sg13g2_fill_1 FILLER_57_1245 ();
 sg13g2_fill_1 FILLER_57_1254 ();
 sg13g2_decap_4 FILLER_57_1269 ();
 sg13g2_fill_2 FILLER_57_1273 ();
 sg13g2_fill_2 FILLER_57_1289 ();
 sg13g2_fill_1 FILLER_57_1291 ();
 sg13g2_fill_2 FILLER_57_1302 ();
 sg13g2_decap_4 FILLER_57_1340 ();
 sg13g2_fill_1 FILLER_57_1353 ();
 sg13g2_fill_1 FILLER_57_1364 ();
 sg13g2_fill_2 FILLER_57_1373 ();
 sg13g2_fill_1 FILLER_57_1389 ();
 sg13g2_fill_2 FILLER_57_1404 ();
 sg13g2_fill_2 FILLER_57_1445 ();
 sg13g2_decap_8 FILLER_57_1453 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_fill_2 FILLER_57_1467 ();
 sg13g2_fill_1 FILLER_57_1469 ();
 sg13g2_fill_2 FILLER_57_1475 ();
 sg13g2_decap_4 FILLER_57_1503 ();
 sg13g2_fill_1 FILLER_57_1516 ();
 sg13g2_fill_1 FILLER_57_1521 ();
 sg13g2_fill_2 FILLER_57_1536 ();
 sg13g2_fill_1 FILLER_57_1538 ();
 sg13g2_fill_1 FILLER_57_1543 ();
 sg13g2_fill_1 FILLER_57_1548 ();
 sg13g2_decap_4 FILLER_57_1579 ();
 sg13g2_fill_1 FILLER_57_1583 ();
 sg13g2_fill_2 FILLER_57_1590 ();
 sg13g2_fill_1 FILLER_57_1601 ();
 sg13g2_fill_1 FILLER_57_1623 ();
 sg13g2_fill_2 FILLER_57_1656 ();
 sg13g2_fill_1 FILLER_57_1658 ();
 sg13g2_fill_1 FILLER_57_1732 ();
 sg13g2_decap_8 FILLER_57_1747 ();
 sg13g2_fill_1 FILLER_57_1754 ();
 sg13g2_fill_2 FILLER_57_1797 ();
 sg13g2_fill_1 FILLER_57_1799 ();
 sg13g2_fill_2 FILLER_57_1889 ();
 sg13g2_fill_1 FILLER_57_1938 ();
 sg13g2_fill_2 FILLER_57_1999 ();
 sg13g2_fill_1 FILLER_57_2018 ();
 sg13g2_fill_2 FILLER_57_2036 ();
 sg13g2_fill_2 FILLER_57_2077 ();
 sg13g2_fill_2 FILLER_57_2084 ();
 sg13g2_fill_2 FILLER_57_2090 ();
 sg13g2_fill_2 FILLER_57_2121 ();
 sg13g2_fill_2 FILLER_57_2139 ();
 sg13g2_fill_1 FILLER_57_2171 ();
 sg13g2_fill_1 FILLER_57_2177 ();
 sg13g2_fill_1 FILLER_57_2183 ();
 sg13g2_fill_2 FILLER_57_2194 ();
 sg13g2_fill_1 FILLER_57_2201 ();
 sg13g2_fill_2 FILLER_57_2256 ();
 sg13g2_fill_1 FILLER_57_2258 ();
 sg13g2_decap_8 FILLER_57_2263 ();
 sg13g2_decap_8 FILLER_57_2270 ();
 sg13g2_fill_2 FILLER_57_2277 ();
 sg13g2_fill_1 FILLER_57_2279 ();
 sg13g2_decap_8 FILLER_57_2315 ();
 sg13g2_decap_8 FILLER_57_2322 ();
 sg13g2_decap_4 FILLER_57_2329 ();
 sg13g2_fill_2 FILLER_57_2333 ();
 sg13g2_fill_2 FILLER_57_2374 ();
 sg13g2_fill_2 FILLER_57_2388 ();
 sg13g2_fill_2 FILLER_57_2413 ();
 sg13g2_fill_1 FILLER_57_2428 ();
 sg13g2_decap_8 FILLER_57_2448 ();
 sg13g2_decap_8 FILLER_57_2455 ();
 sg13g2_decap_4 FILLER_57_2462 ();
 sg13g2_fill_1 FILLER_57_2470 ();
 sg13g2_decap_8 FILLER_57_2481 ();
 sg13g2_fill_1 FILLER_57_2488 ();
 sg13g2_decap_8 FILLER_57_2541 ();
 sg13g2_fill_2 FILLER_57_2548 ();
 sg13g2_fill_2 FILLER_57_2638 ();
 sg13g2_fill_1 FILLER_57_2640 ();
 sg13g2_fill_2 FILLER_57_2667 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_decap_8 FILLER_58_30 ();
 sg13g2_decap_8 FILLER_58_37 ();
 sg13g2_fill_1 FILLER_58_85 ();
 sg13g2_fill_2 FILLER_58_116 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_122 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_151 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_decap_8 FILLER_58_197 ();
 sg13g2_decap_8 FILLER_58_204 ();
 sg13g2_decap_8 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_fill_1 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_276 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_1 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_decap_4 FILLER_58_365 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_decap_4 FILLER_58_391 ();
 sg13g2_fill_2 FILLER_58_400 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_417 ();
 sg13g2_fill_1 FILLER_58_427 ();
 sg13g2_fill_2 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_469 ();
 sg13g2_fill_2 FILLER_58_474 ();
 sg13g2_fill_1 FILLER_58_476 ();
 sg13g2_fill_2 FILLER_58_508 ();
 sg13g2_fill_1 FILLER_58_516 ();
 sg13g2_fill_1 FILLER_58_538 ();
 sg13g2_fill_2 FILLER_58_548 ();
 sg13g2_fill_1 FILLER_58_555 ();
 sg13g2_decap_8 FILLER_58_625 ();
 sg13g2_decap_8 FILLER_58_632 ();
 sg13g2_fill_2 FILLER_58_639 ();
 sg13g2_fill_1 FILLER_58_641 ();
 sg13g2_decap_8 FILLER_58_673 ();
 sg13g2_decap_8 FILLER_58_680 ();
 sg13g2_decap_8 FILLER_58_687 ();
 sg13g2_decap_8 FILLER_58_694 ();
 sg13g2_decap_8 FILLER_58_701 ();
 sg13g2_decap_8 FILLER_58_708 ();
 sg13g2_decap_4 FILLER_58_715 ();
 sg13g2_fill_2 FILLER_58_719 ();
 sg13g2_fill_1 FILLER_58_734 ();
 sg13g2_fill_2 FILLER_58_744 ();
 sg13g2_fill_1 FILLER_58_790 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_830 ();
 sg13g2_decap_8 FILLER_58_837 ();
 sg13g2_fill_1 FILLER_58_844 ();
 sg13g2_fill_2 FILLER_58_850 ();
 sg13g2_fill_1 FILLER_58_862 ();
 sg13g2_decap_8 FILLER_58_867 ();
 sg13g2_fill_1 FILLER_58_878 ();
 sg13g2_fill_2 FILLER_58_883 ();
 sg13g2_fill_2 FILLER_58_893 ();
 sg13g2_fill_1 FILLER_58_895 ();
 sg13g2_fill_1 FILLER_58_902 ();
 sg13g2_fill_2 FILLER_58_908 ();
 sg13g2_fill_1 FILLER_58_910 ();
 sg13g2_decap_4 FILLER_58_950 ();
 sg13g2_decap_4 FILLER_58_958 ();
 sg13g2_fill_1 FILLER_58_962 ();
 sg13g2_decap_4 FILLER_58_984 ();
 sg13g2_fill_1 FILLER_58_988 ();
 sg13g2_decap_4 FILLER_58_995 ();
 sg13g2_fill_1 FILLER_58_999 ();
 sg13g2_decap_8 FILLER_58_1004 ();
 sg13g2_decap_8 FILLER_58_1011 ();
 sg13g2_decap_8 FILLER_58_1018 ();
 sg13g2_fill_1 FILLER_58_1025 ();
 sg13g2_decap_4 FILLER_58_1031 ();
 sg13g2_fill_2 FILLER_58_1035 ();
 sg13g2_fill_1 FILLER_58_1051 ();
 sg13g2_decap_8 FILLER_58_1056 ();
 sg13g2_fill_2 FILLER_58_1063 ();
 sg13g2_fill_1 FILLER_58_1065 ();
 sg13g2_decap_8 FILLER_58_1078 ();
 sg13g2_fill_1 FILLER_58_1085 ();
 sg13g2_fill_1 FILLER_58_1099 ();
 sg13g2_fill_2 FILLER_58_1103 ();
 sg13g2_fill_2 FILLER_58_1124 ();
 sg13g2_fill_2 FILLER_58_1156 ();
 sg13g2_fill_1 FILLER_58_1200 ();
 sg13g2_fill_1 FILLER_58_1206 ();
 sg13g2_fill_2 FILLER_58_1231 ();
 sg13g2_fill_2 FILLER_58_1237 ();
 sg13g2_fill_2 FILLER_58_1246 ();
 sg13g2_fill_1 FILLER_58_1267 ();
 sg13g2_decap_8 FILLER_58_1281 ();
 sg13g2_decap_8 FILLER_58_1288 ();
 sg13g2_fill_2 FILLER_58_1295 ();
 sg13g2_fill_1 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1305 ();
 sg13g2_fill_2 FILLER_58_1312 ();
 sg13g2_decap_8 FILLER_58_1331 ();
 sg13g2_fill_1 FILLER_58_1342 ();
 sg13g2_decap_4 FILLER_58_1347 ();
 sg13g2_fill_1 FILLER_58_1351 ();
 sg13g2_fill_1 FILLER_58_1357 ();
 sg13g2_fill_1 FILLER_58_1367 ();
 sg13g2_fill_2 FILLER_58_1397 ();
 sg13g2_fill_1 FILLER_58_1419 ();
 sg13g2_fill_2 FILLER_58_1446 ();
 sg13g2_decap_8 FILLER_58_1452 ();
 sg13g2_decap_4 FILLER_58_1459 ();
 sg13g2_fill_1 FILLER_58_1463 ();
 sg13g2_fill_2 FILLER_58_1483 ();
 sg13g2_decap_4 FILLER_58_1490 ();
 sg13g2_fill_2 FILLER_58_1494 ();
 sg13g2_fill_2 FILLER_58_1527 ();
 sg13g2_fill_2 FILLER_58_1538 ();
 sg13g2_fill_1 FILLER_58_1540 ();
 sg13g2_decap_8 FILLER_58_1545 ();
 sg13g2_decap_4 FILLER_58_1552 ();
 sg13g2_fill_1 FILLER_58_1556 ();
 sg13g2_fill_1 FILLER_58_1583 ();
 sg13g2_fill_1 FILLER_58_1632 ();
 sg13g2_fill_2 FILLER_58_1643 ();
 sg13g2_fill_1 FILLER_58_1645 ();
 sg13g2_decap_8 FILLER_58_1651 ();
 sg13g2_fill_1 FILLER_58_1658 ();
 sg13g2_fill_2 FILLER_58_1663 ();
 sg13g2_decap_8 FILLER_58_1669 ();
 sg13g2_fill_2 FILLER_58_1676 ();
 sg13g2_decap_4 FILLER_58_1681 ();
 sg13g2_decap_4 FILLER_58_1689 ();
 sg13g2_fill_1 FILLER_58_1697 ();
 sg13g2_decap_4 FILLER_58_1703 ();
 sg13g2_decap_8 FILLER_58_1719 ();
 sg13g2_decap_8 FILLER_58_1726 ();
 sg13g2_decap_8 FILLER_58_1733 ();
 sg13g2_decap_8 FILLER_58_1740 ();
 sg13g2_fill_1 FILLER_58_1747 ();
 sg13g2_fill_1 FILLER_58_1784 ();
 sg13g2_fill_2 FILLER_58_1921 ();
 sg13g2_fill_2 FILLER_58_1958 ();
 sg13g2_fill_1 FILLER_58_1960 ();
 sg13g2_fill_1 FILLER_58_1964 ();
 sg13g2_fill_1 FILLER_58_1975 ();
 sg13g2_decap_4 FILLER_58_1996 ();
 sg13g2_fill_1 FILLER_58_2086 ();
 sg13g2_fill_2 FILLER_58_2116 ();
 sg13g2_fill_2 FILLER_58_2133 ();
 sg13g2_fill_1 FILLER_58_2149 ();
 sg13g2_fill_1 FILLER_58_2190 ();
 sg13g2_fill_2 FILLER_58_2201 ();
 sg13g2_fill_1 FILLER_58_2220 ();
 sg13g2_decap_8 FILLER_58_2257 ();
 sg13g2_fill_2 FILLER_58_2264 ();
 sg13g2_decap_8 FILLER_58_2302 ();
 sg13g2_decap_8 FILLER_58_2313 ();
 sg13g2_decap_4 FILLER_58_2320 ();
 sg13g2_fill_1 FILLER_58_2324 ();
 sg13g2_fill_1 FILLER_58_2337 ();
 sg13g2_decap_8 FILLER_58_2342 ();
 sg13g2_fill_2 FILLER_58_2349 ();
 sg13g2_fill_2 FILLER_58_2387 ();
 sg13g2_fill_1 FILLER_58_2422 ();
 sg13g2_decap_8 FILLER_58_2459 ();
 sg13g2_decap_8 FILLER_58_2466 ();
 sg13g2_fill_2 FILLER_58_2473 ();
 sg13g2_fill_1 FILLER_58_2475 ();
 sg13g2_fill_2 FILLER_58_2489 ();
 sg13g2_fill_1 FILLER_58_2491 ();
 sg13g2_decap_8 FILLER_58_2552 ();
 sg13g2_decap_4 FILLER_58_2559 ();
 sg13g2_fill_2 FILLER_58_2563 ();
 sg13g2_fill_2 FILLER_58_2600 ();
 sg13g2_fill_1 FILLER_58_2602 ();
 sg13g2_decap_4 FILLER_58_2607 ();
 sg13g2_fill_2 FILLER_58_2611 ();
 sg13g2_fill_1 FILLER_58_2621 ();
 sg13g2_decap_4 FILLER_58_2635 ();
 sg13g2_fill_1 FILLER_58_2669 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_4 ();
 sg13g2_fill_2 FILLER_59_41 ();
 sg13g2_fill_1 FILLER_59_43 ();
 sg13g2_decap_4 FILLER_59_74 ();
 sg13g2_fill_1 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_145 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_197 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_decap_4 FILLER_59_214 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_263 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_310 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_387 ();
 sg13g2_fill_1 FILLER_59_394 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_decap_4 FILLER_59_432 ();
 sg13g2_fill_2 FILLER_59_436 ();
 sg13g2_fill_1 FILLER_59_443 ();
 sg13g2_fill_2 FILLER_59_465 ();
 sg13g2_fill_2 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_557 ();
 sg13g2_fill_2 FILLER_59_577 ();
 sg13g2_fill_2 FILLER_59_583 ();
 sg13g2_fill_2 FILLER_59_601 ();
 sg13g2_fill_1 FILLER_59_612 ();
 sg13g2_fill_2 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_688 ();
 sg13g2_fill_2 FILLER_59_693 ();
 sg13g2_fill_1 FILLER_59_699 ();
 sg13g2_fill_2 FILLER_59_704 ();
 sg13g2_fill_1 FILLER_59_706 ();
 sg13g2_decap_8 FILLER_59_713 ();
 sg13g2_decap_8 FILLER_59_720 ();
 sg13g2_decap_8 FILLER_59_727 ();
 sg13g2_decap_8 FILLER_59_734 ();
 sg13g2_fill_1 FILLER_59_741 ();
 sg13g2_fill_1 FILLER_59_782 ();
 sg13g2_fill_1 FILLER_59_806 ();
 sg13g2_fill_2 FILLER_59_819 ();
 sg13g2_fill_1 FILLER_59_821 ();
 sg13g2_fill_2 FILLER_59_827 ();
 sg13g2_fill_2 FILLER_59_841 ();
 sg13g2_fill_1 FILLER_59_843 ();
 sg13g2_fill_2 FILLER_59_852 ();
 sg13g2_fill_1 FILLER_59_854 ();
 sg13g2_fill_2 FILLER_59_863 ();
 sg13g2_fill_1 FILLER_59_865 ();
 sg13g2_fill_1 FILLER_59_895 ();
 sg13g2_fill_2 FILLER_59_907 ();
 sg13g2_fill_1 FILLER_59_909 ();
 sg13g2_fill_1 FILLER_59_923 ();
 sg13g2_fill_1 FILLER_59_932 ();
 sg13g2_fill_1 FILLER_59_938 ();
 sg13g2_fill_2 FILLER_59_950 ();
 sg13g2_decap_4 FILLER_59_956 ();
 sg13g2_fill_2 FILLER_59_960 ();
 sg13g2_fill_2 FILLER_59_984 ();
 sg13g2_fill_2 FILLER_59_991 ();
 sg13g2_fill_2 FILLER_59_1022 ();
 sg13g2_fill_1 FILLER_59_1024 ();
 sg13g2_fill_1 FILLER_59_1059 ();
 sg13g2_fill_2 FILLER_59_1086 ();
 sg13g2_decap_8 FILLER_59_1096 ();
 sg13g2_decap_4 FILLER_59_1103 ();
 sg13g2_fill_1 FILLER_59_1152 ();
 sg13g2_fill_2 FILLER_59_1165 ();
 sg13g2_fill_2 FILLER_59_1171 ();
 sg13g2_fill_2 FILLER_59_1177 ();
 sg13g2_fill_1 FILLER_59_1206 ();
 sg13g2_fill_1 FILLER_59_1254 ();
 sg13g2_fill_2 FILLER_59_1285 ();
 sg13g2_fill_1 FILLER_59_1290 ();
 sg13g2_fill_1 FILLER_59_1317 ();
 sg13g2_fill_2 FILLER_59_1328 ();
 sg13g2_fill_1 FILLER_59_1330 ();
 sg13g2_decap_4 FILLER_59_1357 ();
 sg13g2_fill_1 FILLER_59_1361 ();
 sg13g2_decap_4 FILLER_59_1366 ();
 sg13g2_fill_1 FILLER_59_1370 ();
 sg13g2_decap_4 FILLER_59_1378 ();
 sg13g2_fill_1 FILLER_59_1387 ();
 sg13g2_fill_2 FILLER_59_1391 ();
 sg13g2_fill_1 FILLER_59_1441 ();
 sg13g2_fill_2 FILLER_59_1513 ();
 sg13g2_fill_1 FILLER_59_1537 ();
 sg13g2_decap_4 FILLER_59_1548 ();
 sg13g2_fill_1 FILLER_59_1552 ();
 sg13g2_decap_4 FILLER_59_1557 ();
 sg13g2_fill_1 FILLER_59_1570 ();
 sg13g2_fill_2 FILLER_59_1684 ();
 sg13g2_decap_4 FILLER_59_1706 ();
 sg13g2_fill_2 FILLER_59_1710 ();
 sg13g2_fill_2 FILLER_59_1730 ();
 sg13g2_decap_8 FILLER_59_1748 ();
 sg13g2_decap_4 FILLER_59_1755 ();
 sg13g2_fill_2 FILLER_59_1759 ();
 sg13g2_fill_1 FILLER_59_1766 ();
 sg13g2_fill_1 FILLER_59_1771 ();
 sg13g2_decap_4 FILLER_59_1809 ();
 sg13g2_decap_4 FILLER_59_1837 ();
 sg13g2_fill_2 FILLER_59_1841 ();
 sg13g2_fill_2 FILLER_59_1855 ();
 sg13g2_fill_1 FILLER_59_1861 ();
 sg13g2_fill_2 FILLER_59_1890 ();
 sg13g2_fill_2 FILLER_59_1951 ();
 sg13g2_fill_1 FILLER_59_1963 ();
 sg13g2_decap_4 FILLER_59_1968 ();
 sg13g2_fill_2 FILLER_59_1972 ();
 sg13g2_decap_4 FILLER_59_2014 ();
 sg13g2_fill_1 FILLER_59_2018 ();
 sg13g2_fill_2 FILLER_59_2043 ();
 sg13g2_fill_1 FILLER_59_2093 ();
 sg13g2_fill_1 FILLER_59_2099 ();
 sg13g2_fill_2 FILLER_59_2126 ();
 sg13g2_fill_2 FILLER_59_2140 ();
 sg13g2_fill_1 FILLER_59_2172 ();
 sg13g2_fill_2 FILLER_59_2195 ();
 sg13g2_fill_2 FILLER_59_2239 ();
 sg13g2_fill_1 FILLER_59_2241 ();
 sg13g2_fill_2 FILLER_59_2252 ();
 sg13g2_fill_1 FILLER_59_2254 ();
 sg13g2_decap_4 FILLER_59_2281 ();
 sg13g2_fill_2 FILLER_59_2289 ();
 sg13g2_fill_1 FILLER_59_2291 ();
 sg13g2_decap_8 FILLER_59_2296 ();
 sg13g2_decap_4 FILLER_59_2303 ();
 sg13g2_fill_1 FILLER_59_2307 ();
 sg13g2_decap_4 FILLER_59_2352 ();
 sg13g2_fill_2 FILLER_59_2356 ();
 sg13g2_fill_2 FILLER_59_2434 ();
 sg13g2_decap_4 FILLER_59_2466 ();
 sg13g2_decap_8 FILLER_59_2474 ();
 sg13g2_fill_1 FILLER_59_2481 ();
 sg13g2_fill_1 FILLER_59_2516 ();
 sg13g2_decap_8 FILLER_59_2553 ();
 sg13g2_decap_8 FILLER_59_2560 ();
 sg13g2_decap_8 FILLER_59_2567 ();
 sg13g2_decap_8 FILLER_59_2574 ();
 sg13g2_decap_4 FILLER_59_2581 ();
 sg13g2_fill_1 FILLER_59_2585 ();
 sg13g2_fill_1 FILLER_59_2596 ();
 sg13g2_fill_1 FILLER_59_2628 ();
 sg13g2_decap_8 FILLER_59_2657 ();
 sg13g2_decap_4 FILLER_59_2664 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_decap_8 FILLER_60_20 ();
 sg13g2_fill_2 FILLER_60_27 ();
 sg13g2_fill_1 FILLER_60_29 ();
 sg13g2_fill_2 FILLER_60_44 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_fill_1 FILLER_60_55 ();
 sg13g2_fill_1 FILLER_60_82 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_decap_4 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_129 ();
 sg13g2_fill_2 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_fill_1 FILLER_60_233 ();
 sg13g2_fill_1 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_292 ();
 sg13g2_fill_2 FILLER_60_297 ();
 sg13g2_fill_1 FILLER_60_306 ();
 sg13g2_fill_1 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_389 ();
 sg13g2_fill_1 FILLER_60_391 ();
 sg13g2_decap_4 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_402 ();
 sg13g2_fill_1 FILLER_60_441 ();
 sg13g2_fill_2 FILLER_60_447 ();
 sg13g2_fill_1 FILLER_60_464 ();
 sg13g2_decap_8 FILLER_60_469 ();
 sg13g2_fill_1 FILLER_60_476 ();
 sg13g2_fill_1 FILLER_60_487 ();
 sg13g2_decap_8 FILLER_60_493 ();
 sg13g2_decap_4 FILLER_60_500 ();
 sg13g2_fill_2 FILLER_60_504 ();
 sg13g2_fill_2 FILLER_60_553 ();
 sg13g2_fill_1 FILLER_60_580 ();
 sg13g2_fill_2 FILLER_60_607 ();
 sg13g2_fill_2 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_619 ();
 sg13g2_fill_1 FILLER_60_633 ();
 sg13g2_fill_1 FILLER_60_638 ();
 sg13g2_fill_1 FILLER_60_656 ();
 sg13g2_fill_1 FILLER_60_666 ();
 sg13g2_fill_2 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_678 ();
 sg13g2_fill_1 FILLER_60_719 ();
 sg13g2_decap_4 FILLER_60_746 ();
 sg13g2_decap_4 FILLER_60_755 ();
 sg13g2_decap_4 FILLER_60_798 ();
 sg13g2_fill_2 FILLER_60_802 ();
 sg13g2_fill_2 FILLER_60_822 ();
 sg13g2_fill_2 FILLER_60_877 ();
 sg13g2_fill_1 FILLER_60_884 ();
 sg13g2_fill_2 FILLER_60_895 ();
 sg13g2_fill_1 FILLER_60_897 ();
 sg13g2_fill_1 FILLER_60_918 ();
 sg13g2_fill_1 FILLER_60_924 ();
 sg13g2_fill_1 FILLER_60_930 ();
 sg13g2_decap_8 FILLER_60_951 ();
 sg13g2_fill_1 FILLER_60_958 ();
 sg13g2_fill_2 FILLER_60_972 ();
 sg13g2_fill_1 FILLER_60_974 ();
 sg13g2_decap_4 FILLER_60_990 ();
 sg13g2_fill_1 FILLER_60_994 ();
 sg13g2_decap_8 FILLER_60_1002 ();
 sg13g2_decap_8 FILLER_60_1009 ();
 sg13g2_decap_8 FILLER_60_1016 ();
 sg13g2_decap_4 FILLER_60_1023 ();
 sg13g2_fill_1 FILLER_60_1027 ();
 sg13g2_fill_2 FILLER_60_1049 ();
 sg13g2_fill_1 FILLER_60_1058 ();
 sg13g2_fill_2 FILLER_60_1064 ();
 sg13g2_decap_4 FILLER_60_1070 ();
 sg13g2_fill_1 FILLER_60_1078 ();
 sg13g2_fill_2 FILLER_60_1088 ();
 sg13g2_fill_1 FILLER_60_1090 ();
 sg13g2_decap_8 FILLER_60_1094 ();
 sg13g2_decap_8 FILLER_60_1101 ();
 sg13g2_decap_4 FILLER_60_1108 ();
 sg13g2_fill_1 FILLER_60_1112 ();
 sg13g2_fill_1 FILLER_60_1117 ();
 sg13g2_fill_2 FILLER_60_1147 ();
 sg13g2_fill_2 FILLER_60_1175 ();
 sg13g2_fill_2 FILLER_60_1205 ();
 sg13g2_fill_1 FILLER_60_1224 ();
 sg13g2_fill_2 FILLER_60_1257 ();
 sg13g2_fill_2 FILLER_60_1268 ();
 sg13g2_fill_1 FILLER_60_1296 ();
 sg13g2_fill_2 FILLER_60_1301 ();
 sg13g2_fill_2 FILLER_60_1336 ();
 sg13g2_decap_4 FILLER_60_1368 ();
 sg13g2_fill_2 FILLER_60_1375 ();
 sg13g2_fill_2 FILLER_60_1413 ();
 sg13g2_fill_1 FILLER_60_1415 ();
 sg13g2_fill_1 FILLER_60_1420 ();
 sg13g2_fill_1 FILLER_60_1435 ();
 sg13g2_fill_1 FILLER_60_1442 ();
 sg13g2_fill_1 FILLER_60_1473 ();
 sg13g2_fill_1 FILLER_60_1493 ();
 sg13g2_fill_1 FILLER_60_1498 ();
 sg13g2_fill_1 FILLER_60_1503 ();
 sg13g2_fill_1 FILLER_60_1535 ();
 sg13g2_fill_1 FILLER_60_1567 ();
 sg13g2_fill_2 FILLER_60_1581 ();
 sg13g2_fill_2 FILLER_60_1587 ();
 sg13g2_fill_1 FILLER_60_1589 ();
 sg13g2_fill_1 FILLER_60_1599 ();
 sg13g2_fill_2 FILLER_60_1605 ();
 sg13g2_fill_1 FILLER_60_1616 ();
 sg13g2_fill_2 FILLER_60_1643 ();
 sg13g2_fill_1 FILLER_60_1650 ();
 sg13g2_fill_2 FILLER_60_1707 ();
 sg13g2_fill_1 FILLER_60_1717 ();
 sg13g2_decap_8 FILLER_60_1751 ();
 sg13g2_fill_2 FILLER_60_1758 ();
 sg13g2_fill_1 FILLER_60_1764 ();
 sg13g2_fill_1 FILLER_60_1771 ();
 sg13g2_fill_2 FILLER_60_1783 ();
 sg13g2_fill_2 FILLER_60_1789 ();
 sg13g2_decap_4 FILLER_60_1801 ();
 sg13g2_fill_2 FILLER_60_1805 ();
 sg13g2_decap_8 FILLER_60_1812 ();
 sg13g2_decap_4 FILLER_60_1819 ();
 sg13g2_fill_2 FILLER_60_1823 ();
 sg13g2_fill_1 FILLER_60_1867 ();
 sg13g2_decap_4 FILLER_60_2014 ();
 sg13g2_fill_1 FILLER_60_2022 ();
 sg13g2_fill_1 FILLER_60_2035 ();
 sg13g2_fill_1 FILLER_60_2045 ();
 sg13g2_decap_4 FILLER_60_2058 ();
 sg13g2_fill_1 FILLER_60_2091 ();
 sg13g2_fill_1 FILLER_60_2162 ();
 sg13g2_fill_1 FILLER_60_2169 ();
 sg13g2_decap_8 FILLER_60_2214 ();
 sg13g2_decap_8 FILLER_60_2221 ();
 sg13g2_fill_1 FILLER_60_2296 ();
 sg13g2_fill_2 FILLER_60_2333 ();
 sg13g2_fill_2 FILLER_60_2397 ();
 sg13g2_fill_1 FILLER_60_2399 ();
 sg13g2_fill_2 FILLER_60_2461 ();
 sg13g2_fill_2 FILLER_60_2489 ();
 sg13g2_fill_1 FILLER_60_2491 ();
 sg13g2_decap_4 FILLER_60_2530 ();
 sg13g2_fill_2 FILLER_60_2569 ();
 sg13g2_fill_1 FILLER_60_2571 ();
 sg13g2_fill_1 FILLER_60_2619 ();
 sg13g2_decap_4 FILLER_60_2624 ();
 sg13g2_decap_8 FILLER_60_2654 ();
 sg13g2_decap_8 FILLER_60_2661 ();
 sg13g2_fill_2 FILLER_60_2668 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_11 ();
 sg13g2_decap_4 FILLER_61_41 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_decap_8 FILLER_61_67 ();
 sg13g2_decap_8 FILLER_61_78 ();
 sg13g2_decap_8 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_97 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_fill_2 FILLER_61_173 ();
 sg13g2_fill_1 FILLER_61_193 ();
 sg13g2_fill_1 FILLER_61_204 ();
 sg13g2_fill_2 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_215 ();
 sg13g2_fill_2 FILLER_61_221 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_2 FILLER_61_289 ();
 sg13g2_fill_1 FILLER_61_302 ();
 sg13g2_fill_2 FILLER_61_306 ();
 sg13g2_fill_2 FILLER_61_325 ();
 sg13g2_fill_1 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_4 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_decap_4 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_401 ();
 sg13g2_fill_2 FILLER_61_426 ();
 sg13g2_fill_1 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_444 ();
 sg13g2_decap_4 FILLER_61_466 ();
 sg13g2_fill_1 FILLER_61_470 ();
 sg13g2_fill_2 FILLER_61_476 ();
 sg13g2_decap_4 FILLER_61_483 ();
 sg13g2_fill_2 FILLER_61_487 ();
 sg13g2_fill_2 FILLER_61_517 ();
 sg13g2_fill_1 FILLER_61_519 ();
 sg13g2_decap_4 FILLER_61_523 ();
 sg13g2_fill_1 FILLER_61_527 ();
 sg13g2_fill_1 FILLER_61_575 ();
 sg13g2_decap_8 FILLER_61_606 ();
 sg13g2_decap_4 FILLER_61_613 ();
 sg13g2_fill_1 FILLER_61_617 ();
 sg13g2_decap_4 FILLER_61_623 ();
 sg13g2_fill_2 FILLER_61_627 ();
 sg13g2_decap_4 FILLER_61_633 ();
 sg13g2_fill_1 FILLER_61_637 ();
 sg13g2_fill_2 FILLER_61_674 ();
 sg13g2_fill_2 FILLER_61_758 ();
 sg13g2_decap_8 FILLER_61_765 ();
 sg13g2_fill_1 FILLER_61_772 ();
 sg13g2_fill_2 FILLER_61_782 ();
 sg13g2_fill_1 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_792 ();
 sg13g2_fill_1 FILLER_61_799 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_fill_2 FILLER_61_811 ();
 sg13g2_fill_1 FILLER_61_821 ();
 sg13g2_fill_1 FILLER_61_831 ();
 sg13g2_fill_1 FILLER_61_898 ();
 sg13g2_fill_2 FILLER_61_903 ();
 sg13g2_fill_1 FILLER_61_905 ();
 sg13g2_decap_4 FILLER_61_910 ();
 sg13g2_decap_4 FILLER_61_922 ();
 sg13g2_fill_1 FILLER_61_926 ();
 sg13g2_fill_1 FILLER_61_939 ();
 sg13g2_fill_1 FILLER_61_950 ();
 sg13g2_fill_1 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1003 ();
 sg13g2_decap_8 FILLER_61_1010 ();
 sg13g2_decap_4 FILLER_61_1017 ();
 sg13g2_fill_2 FILLER_61_1060 ();
 sg13g2_fill_1 FILLER_61_1062 ();
 sg13g2_decap_4 FILLER_61_1078 ();
 sg13g2_fill_2 FILLER_61_1082 ();
 sg13g2_decap_8 FILLER_61_1092 ();
 sg13g2_decap_4 FILLER_61_1102 ();
 sg13g2_fill_1 FILLER_61_1106 ();
 sg13g2_decap_8 FILLER_61_1110 ();
 sg13g2_decap_8 FILLER_61_1117 ();
 sg13g2_fill_2 FILLER_61_1131 ();
 sg13g2_fill_1 FILLER_61_1137 ();
 sg13g2_fill_1 FILLER_61_1142 ();
 sg13g2_fill_1 FILLER_61_1146 ();
 sg13g2_fill_1 FILLER_61_1170 ();
 sg13g2_fill_2 FILLER_61_1203 ();
 sg13g2_fill_1 FILLER_61_1220 ();
 sg13g2_fill_1 FILLER_61_1225 ();
 sg13g2_fill_2 FILLER_61_1260 ();
 sg13g2_fill_1 FILLER_61_1262 ();
 sg13g2_fill_2 FILLER_61_1267 ();
 sg13g2_fill_2 FILLER_61_1273 ();
 sg13g2_fill_1 FILLER_61_1275 ();
 sg13g2_decap_4 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_fill_2 FILLER_61_1310 ();
 sg13g2_fill_2 FILLER_61_1316 ();
 sg13g2_fill_2 FILLER_61_1348 ();
 sg13g2_fill_2 FILLER_61_1354 ();
 sg13g2_decap_8 FILLER_61_1390 ();
 sg13g2_decap_8 FILLER_61_1397 ();
 sg13g2_decap_8 FILLER_61_1404 ();
 sg13g2_fill_1 FILLER_61_1411 ();
 sg13g2_decap_4 FILLER_61_1422 ();
 sg13g2_fill_1 FILLER_61_1426 ();
 sg13g2_fill_2 FILLER_61_1444 ();
 sg13g2_decap_8 FILLER_61_1455 ();
 sg13g2_fill_1 FILLER_61_1462 ();
 sg13g2_decap_8 FILLER_61_1467 ();
 sg13g2_fill_1 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1479 ();
 sg13g2_fill_1 FILLER_61_1481 ();
 sg13g2_decap_8 FILLER_61_1491 ();
 sg13g2_fill_2 FILLER_61_1498 ();
 sg13g2_fill_1 FILLER_61_1500 ();
 sg13g2_fill_2 FILLER_61_1515 ();
 sg13g2_fill_1 FILLER_61_1517 ();
 sg13g2_fill_1 FILLER_61_1548 ();
 sg13g2_fill_2 FILLER_61_1593 ();
 sg13g2_decap_4 FILLER_61_1607 ();
 sg13g2_fill_1 FILLER_61_1611 ();
 sg13g2_fill_2 FILLER_61_1620 ();
 sg13g2_fill_1 FILLER_61_1622 ();
 sg13g2_fill_2 FILLER_61_1636 ();
 sg13g2_fill_1 FILLER_61_1647 ();
 sg13g2_fill_2 FILLER_61_1653 ();
 sg13g2_fill_1 FILLER_61_1655 ();
 sg13g2_decap_4 FILLER_61_1698 ();
 sg13g2_fill_1 FILLER_61_1771 ();
 sg13g2_decap_8 FILLER_61_1783 ();
 sg13g2_decap_4 FILLER_61_1790 ();
 sg13g2_fill_1 FILLER_61_1794 ();
 sg13g2_decap_8 FILLER_61_1799 ();
 sg13g2_decap_8 FILLER_61_1806 ();
 sg13g2_fill_2 FILLER_61_1813 ();
 sg13g2_fill_1 FILLER_61_1815 ();
 sg13g2_fill_1 FILLER_61_1856 ();
 sg13g2_fill_1 FILLER_61_1863 ();
 sg13g2_fill_2 FILLER_61_1868 ();
 sg13g2_fill_2 FILLER_61_1874 ();
 sg13g2_fill_2 FILLER_61_1880 ();
 sg13g2_decap_8 FILLER_61_1886 ();
 sg13g2_fill_1 FILLER_61_1893 ();
 sg13g2_fill_1 FILLER_61_1915 ();
 sg13g2_fill_2 FILLER_61_1925 ();
 sg13g2_fill_2 FILLER_61_1941 ();
 sg13g2_decap_8 FILLER_61_1947 ();
 sg13g2_decap_8 FILLER_61_1954 ();
 sg13g2_decap_4 FILLER_61_1961 ();
 sg13g2_fill_2 FILLER_61_1965 ();
 sg13g2_decap_8 FILLER_61_2051 ();
 sg13g2_decap_8 FILLER_61_2058 ();
 sg13g2_fill_2 FILLER_61_2070 ();
 sg13g2_fill_2 FILLER_61_2104 ();
 sg13g2_fill_1 FILLER_61_2131 ();
 sg13g2_fill_1 FILLER_61_2139 ();
 sg13g2_decap_8 FILLER_61_2218 ();
 sg13g2_fill_1 FILLER_61_2225 ();
 sg13g2_fill_1 FILLER_61_2256 ();
 sg13g2_decap_4 FILLER_61_2267 ();
 sg13g2_fill_1 FILLER_61_2271 ();
 sg13g2_fill_1 FILLER_61_2282 ();
 sg13g2_fill_2 FILLER_61_2390 ();
 sg13g2_fill_1 FILLER_61_2392 ();
 sg13g2_fill_2 FILLER_61_2401 ();
 sg13g2_decap_8 FILLER_61_2427 ();
 sg13g2_decap_8 FILLER_61_2444 ();
 sg13g2_decap_8 FILLER_61_2520 ();
 sg13g2_decap_8 FILLER_61_2527 ();
 sg13g2_fill_2 FILLER_61_2534 ();
 sg13g2_fill_1 FILLER_61_2536 ();
 sg13g2_fill_2 FILLER_61_2583 ();
 sg13g2_fill_1 FILLER_61_2585 ();
 sg13g2_decap_8 FILLER_61_2596 ();
 sg13g2_fill_1 FILLER_61_2603 ();
 sg13g2_decap_4 FILLER_61_2614 ();
 sg13g2_decap_8 FILLER_61_2639 ();
 sg13g2_decap_8 FILLER_61_2646 ();
 sg13g2_decap_8 FILLER_61_2653 ();
 sg13g2_decap_8 FILLER_61_2660 ();
 sg13g2_fill_2 FILLER_61_2667 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_decap_4 FILLER_62_23 ();
 sg13g2_fill_1 FILLER_62_27 ();
 sg13g2_decap_8 FILLER_62_38 ();
 sg13g2_fill_2 FILLER_62_45 ();
 sg13g2_decap_8 FILLER_62_93 ();
 sg13g2_fill_2 FILLER_62_100 ();
 sg13g2_fill_2 FILLER_62_107 ();
 sg13g2_fill_1 FILLER_62_135 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_fill_2 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_199 ();
 sg13g2_decap_4 FILLER_62_209 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_251 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_fill_2 FILLER_62_382 ();
 sg13g2_decap_8 FILLER_62_389 ();
 sg13g2_decap_4 FILLER_62_396 ();
 sg13g2_fill_1 FILLER_62_400 ();
 sg13g2_decap_8 FILLER_62_409 ();
 sg13g2_decap_4 FILLER_62_461 ();
 sg13g2_fill_2 FILLER_62_465 ();
 sg13g2_decap_8 FILLER_62_512 ();
 sg13g2_fill_1 FILLER_62_519 ();
 sg13g2_decap_4 FILLER_62_524 ();
 sg13g2_fill_2 FILLER_62_608 ();
 sg13g2_fill_2 FILLER_62_636 ();
 sg13g2_fill_1 FILLER_62_638 ();
 sg13g2_fill_2 FILLER_62_643 ();
 sg13g2_fill_1 FILLER_62_650 ();
 sg13g2_fill_2 FILLER_62_655 ();
 sg13g2_fill_1 FILLER_62_696 ();
 sg13g2_decap_8 FILLER_62_727 ();
 sg13g2_fill_1 FILLER_62_734 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_754 ();
 sg13g2_fill_2 FILLER_62_780 ();
 sg13g2_fill_1 FILLER_62_782 ();
 sg13g2_decap_8 FILLER_62_787 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_fill_2 FILLER_62_801 ();
 sg13g2_fill_2 FILLER_62_836 ();
 sg13g2_fill_1 FILLER_62_852 ();
 sg13g2_fill_1 FILLER_62_860 ();
 sg13g2_decap_8 FILLER_62_877 ();
 sg13g2_fill_2 FILLER_62_889 ();
 sg13g2_fill_1 FILLER_62_891 ();
 sg13g2_decap_8 FILLER_62_905 ();
 sg13g2_fill_1 FILLER_62_948 ();
 sg13g2_fill_1 FILLER_62_958 ();
 sg13g2_fill_1 FILLER_62_964 ();
 sg13g2_fill_1 FILLER_62_971 ();
 sg13g2_fill_1 FILLER_62_981 ();
 sg13g2_fill_2 FILLER_62_986 ();
 sg13g2_fill_2 FILLER_62_996 ();
 sg13g2_fill_1 FILLER_62_998 ();
 sg13g2_fill_1 FILLER_62_1012 ();
 sg13g2_fill_2 FILLER_62_1039 ();
 sg13g2_fill_1 FILLER_62_1041 ();
 sg13g2_decap_4 FILLER_62_1060 ();
 sg13g2_fill_2 FILLER_62_1068 ();
 sg13g2_fill_1 FILLER_62_1114 ();
 sg13g2_fill_2 FILLER_62_1125 ();
 sg13g2_decap_4 FILLER_62_1135 ();
 sg13g2_fill_1 FILLER_62_1139 ();
 sg13g2_fill_1 FILLER_62_1156 ();
 sg13g2_fill_1 FILLER_62_1183 ();
 sg13g2_fill_2 FILLER_62_1190 ();
 sg13g2_fill_1 FILLER_62_1196 ();
 sg13g2_fill_2 FILLER_62_1203 ();
 sg13g2_fill_1 FILLER_62_1221 ();
 sg13g2_fill_1 FILLER_62_1228 ();
 sg13g2_fill_2 FILLER_62_1237 ();
 sg13g2_fill_1 FILLER_62_1239 ();
 sg13g2_decap_8 FILLER_62_1243 ();
 sg13g2_decap_4 FILLER_62_1250 ();
 sg13g2_fill_1 FILLER_62_1254 ();
 sg13g2_decap_4 FILLER_62_1288 ();
 sg13g2_fill_1 FILLER_62_1292 ();
 sg13g2_decap_8 FILLER_62_1297 ();
 sg13g2_fill_1 FILLER_62_1304 ();
 sg13g2_decap_8 FILLER_62_1310 ();
 sg13g2_decap_4 FILLER_62_1317 ();
 sg13g2_fill_1 FILLER_62_1321 ();
 sg13g2_decap_8 FILLER_62_1326 ();
 sg13g2_fill_2 FILLER_62_1333 ();
 sg13g2_fill_1 FILLER_62_1335 ();
 sg13g2_decap_4 FILLER_62_1341 ();
 sg13g2_decap_4 FILLER_62_1350 ();
 sg13g2_fill_1 FILLER_62_1354 ();
 sg13g2_decap_8 FILLER_62_1364 ();
 sg13g2_fill_1 FILLER_62_1371 ();
 sg13g2_fill_1 FILLER_62_1377 ();
 sg13g2_decap_8 FILLER_62_1382 ();
 sg13g2_decap_8 FILLER_62_1389 ();
 sg13g2_fill_2 FILLER_62_1406 ();
 sg13g2_fill_1 FILLER_62_1438 ();
 sg13g2_decap_4 FILLER_62_1455 ();
 sg13g2_fill_2 FILLER_62_1459 ();
 sg13g2_fill_1 FILLER_62_1471 ();
 sg13g2_fill_1 FILLER_62_1497 ();
 sg13g2_fill_2 FILLER_62_1528 ();
 sg13g2_fill_1 FILLER_62_1575 ();
 sg13g2_fill_2 FILLER_62_1611 ();
 sg13g2_decap_4 FILLER_62_1646 ();
 sg13g2_decap_8 FILLER_62_1676 ();
 sg13g2_decap_4 FILLER_62_1683 ();
 sg13g2_fill_2 FILLER_62_1687 ();
 sg13g2_fill_2 FILLER_62_1693 ();
 sg13g2_fill_1 FILLER_62_1695 ();
 sg13g2_fill_1 FILLER_62_1746 ();
 sg13g2_fill_2 FILLER_62_1752 ();
 sg13g2_fill_1 FILLER_62_1759 ();
 sg13g2_decap_4 FILLER_62_1764 ();
 sg13g2_fill_1 FILLER_62_1783 ();
 sg13g2_fill_2 FILLER_62_1814 ();
 sg13g2_fill_2 FILLER_62_1852 ();
 sg13g2_fill_1 FILLER_62_1854 ();
 sg13g2_decap_4 FILLER_62_1865 ();
 sg13g2_fill_1 FILLER_62_1869 ();
 sg13g2_fill_1 FILLER_62_1906 ();
 sg13g2_fill_1 FILLER_62_1920 ();
 sg13g2_decap_8 FILLER_62_1953 ();
 sg13g2_decap_8 FILLER_62_1960 ();
 sg13g2_fill_2 FILLER_62_1967 ();
 sg13g2_fill_2 FILLER_62_1984 ();
 sg13g2_fill_1 FILLER_62_1986 ();
 sg13g2_decap_4 FILLER_62_2023 ();
 sg13g2_fill_1 FILLER_62_2027 ();
 sg13g2_decap_4 FILLER_62_2032 ();
 sg13g2_fill_2 FILLER_62_2036 ();
 sg13g2_fill_1 FILLER_62_2070 ();
 sg13g2_fill_1 FILLER_62_2078 ();
 sg13g2_fill_1 FILLER_62_2083 ();
 sg13g2_fill_1 FILLER_62_2089 ();
 sg13g2_fill_1 FILLER_62_2095 ();
 sg13g2_fill_1 FILLER_62_2111 ();
 sg13g2_fill_2 FILLER_62_2116 ();
 sg13g2_fill_2 FILLER_62_2122 ();
 sg13g2_fill_2 FILLER_62_2139 ();
 sg13g2_fill_1 FILLER_62_2192 ();
 sg13g2_fill_1 FILLER_62_2229 ();
 sg13g2_decap_8 FILLER_62_2258 ();
 sg13g2_decap_8 FILLER_62_2265 ();
 sg13g2_decap_4 FILLER_62_2282 ();
 sg13g2_decap_8 FILLER_62_2339 ();
 sg13g2_fill_2 FILLER_62_2379 ();
 sg13g2_fill_1 FILLER_62_2381 ();
 sg13g2_fill_1 FILLER_62_2392 ();
 sg13g2_fill_2 FILLER_62_2410 ();
 sg13g2_fill_1 FILLER_62_2412 ();
 sg13g2_fill_1 FILLER_62_2417 ();
 sg13g2_decap_4 FILLER_62_2452 ();
 sg13g2_decap_8 FILLER_62_2496 ();
 sg13g2_decap_8 FILLER_62_2503 ();
 sg13g2_decap_4 FILLER_62_2510 ();
 sg13g2_fill_1 FILLER_62_2514 ();
 sg13g2_decap_8 FILLER_62_2529 ();
 sg13g2_decap_8 FILLER_62_2536 ();
 sg13g2_fill_1 FILLER_62_2553 ();
 sg13g2_fill_2 FILLER_62_2580 ();
 sg13g2_fill_2 FILLER_62_2608 ();
 sg13g2_decap_4 FILLER_62_2636 ();
 sg13g2_fill_2 FILLER_62_2640 ();
 sg13g2_decap_8 FILLER_62_2646 ();
 sg13g2_decap_8 FILLER_62_2653 ();
 sg13g2_decap_8 FILLER_62_2660 ();
 sg13g2_fill_2 FILLER_62_2667 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_57 ();
 sg13g2_fill_2 FILLER_63_61 ();
 sg13g2_fill_2 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_122 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_194 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_fill_1 FILLER_63_216 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_269 ();
 sg13g2_fill_1 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_310 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_327 ();
 sg13g2_decap_4 FILLER_63_352 ();
 sg13g2_fill_2 FILLER_63_356 ();
 sg13g2_fill_2 FILLER_63_399 ();
 sg13g2_fill_1 FILLER_63_401 ();
 sg13g2_decap_4 FILLER_63_413 ();
 sg13g2_fill_1 FILLER_63_417 ();
 sg13g2_decap_4 FILLER_63_424 ();
 sg13g2_fill_1 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_63_433 ();
 sg13g2_decap_8 FILLER_63_440 ();
 sg13g2_decap_8 FILLER_63_522 ();
 sg13g2_decap_8 FILLER_63_529 ();
 sg13g2_fill_2 FILLER_63_548 ();
 sg13g2_fill_2 FILLER_63_559 ();
 sg13g2_fill_2 FILLER_63_598 ();
 sg13g2_decap_4 FILLER_63_608 ();
 sg13g2_fill_1 FILLER_63_620 ();
 sg13g2_fill_1 FILLER_63_626 ();
 sg13g2_fill_2 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_680 ();
 sg13g2_fill_1 FILLER_63_682 ();
 sg13g2_fill_1 FILLER_63_706 ();
 sg13g2_fill_1 FILLER_63_710 ();
 sg13g2_fill_2 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_727 ();
 sg13g2_decap_8 FILLER_63_734 ();
 sg13g2_fill_2 FILLER_63_746 ();
 sg13g2_decap_8 FILLER_63_785 ();
 sg13g2_decap_8 FILLER_63_792 ();
 sg13g2_decap_8 FILLER_63_799 ();
 sg13g2_fill_2 FILLER_63_806 ();
 sg13g2_fill_1 FILLER_63_816 ();
 sg13g2_fill_1 FILLER_63_837 ();
 sg13g2_decap_4 FILLER_63_848 ();
 sg13g2_fill_2 FILLER_63_852 ();
 sg13g2_decap_8 FILLER_63_896 ();
 sg13g2_decap_8 FILLER_63_903 ();
 sg13g2_decap_4 FILLER_63_915 ();
 sg13g2_fill_1 FILLER_63_919 ();
 sg13g2_fill_1 FILLER_63_933 ();
 sg13g2_fill_2 FILLER_63_939 ();
 sg13g2_fill_1 FILLER_63_941 ();
 sg13g2_fill_1 FILLER_63_957 ();
 sg13g2_decap_8 FILLER_63_962 ();
 sg13g2_decap_4 FILLER_63_969 ();
 sg13g2_decap_4 FILLER_63_1016 ();
 sg13g2_fill_1 FILLER_63_1028 ();
 sg13g2_fill_1 FILLER_63_1033 ();
 sg13g2_fill_1 FILLER_63_1043 ();
 sg13g2_fill_1 FILLER_63_1048 ();
 sg13g2_fill_1 FILLER_63_1060 ();
 sg13g2_fill_1 FILLER_63_1067 ();
 sg13g2_decap_4 FILLER_63_1073 ();
 sg13g2_fill_2 FILLER_63_1081 ();
 sg13g2_fill_1 FILLER_63_1083 ();
 sg13g2_fill_2 FILLER_63_1099 ();
 sg13g2_fill_2 FILLER_63_1114 ();
 sg13g2_decap_4 FILLER_63_1124 ();
 sg13g2_fill_1 FILLER_63_1128 ();
 sg13g2_decap_8 FILLER_63_1137 ();
 sg13g2_decap_4 FILLER_63_1144 ();
 sg13g2_fill_1 FILLER_63_1168 ();
 sg13g2_fill_2 FILLER_63_1177 ();
 sg13g2_fill_2 FILLER_63_1183 ();
 sg13g2_fill_1 FILLER_63_1209 ();
 sg13g2_fill_1 FILLER_63_1218 ();
 sg13g2_decap_4 FILLER_63_1227 ();
 sg13g2_fill_2 FILLER_63_1236 ();
 sg13g2_decap_8 FILLER_63_1251 ();
 sg13g2_fill_2 FILLER_63_1258 ();
 sg13g2_decap_4 FILLER_63_1264 ();
 sg13g2_fill_1 FILLER_63_1268 ();
 sg13g2_decap_8 FILLER_63_1295 ();
 sg13g2_decap_8 FILLER_63_1302 ();
 sg13g2_decap_8 FILLER_63_1309 ();
 sg13g2_decap_8 FILLER_63_1316 ();
 sg13g2_decap_8 FILLER_63_1323 ();
 sg13g2_decap_4 FILLER_63_1330 ();
 sg13g2_fill_1 FILLER_63_1334 ();
 sg13g2_decap_8 FILLER_63_1339 ();
 sg13g2_decap_8 FILLER_63_1346 ();
 sg13g2_decap_8 FILLER_63_1353 ();
 sg13g2_decap_8 FILLER_63_1360 ();
 sg13g2_decap_8 FILLER_63_1367 ();
 sg13g2_decap_8 FILLER_63_1374 ();
 sg13g2_decap_8 FILLER_63_1381 ();
 sg13g2_decap_4 FILLER_63_1388 ();
 sg13g2_fill_1 FILLER_63_1462 ();
 sg13g2_decap_8 FILLER_63_1542 ();
 sg13g2_decap_4 FILLER_63_1549 ();
 sg13g2_fill_1 FILLER_63_1553 ();
 sg13g2_decap_8 FILLER_63_1558 ();
 sg13g2_fill_1 FILLER_63_1565 ();
 sg13g2_decap_8 FILLER_63_1572 ();
 sg13g2_fill_1 FILLER_63_1579 ();
 sg13g2_fill_1 FILLER_63_1610 ();
 sg13g2_fill_1 FILLER_63_1628 ();
 sg13g2_fill_1 FILLER_63_1665 ();
 sg13g2_decap_8 FILLER_63_1682 ();
 sg13g2_fill_2 FILLER_63_1699 ();
 sg13g2_fill_1 FILLER_63_1701 ();
 sg13g2_fill_1 FILLER_63_1706 ();
 sg13g2_fill_2 FILLER_63_1711 ();
 sg13g2_fill_2 FILLER_63_1717 ();
 sg13g2_fill_1 FILLER_63_1723 ();
 sg13g2_fill_1 FILLER_63_1746 ();
 sg13g2_fill_1 FILLER_63_1753 ();
 sg13g2_decap_4 FILLER_63_1764 ();
 sg13g2_fill_1 FILLER_63_1768 ();
 sg13g2_fill_1 FILLER_63_1774 ();
 sg13g2_fill_1 FILLER_63_1819 ();
 sg13g2_fill_1 FILLER_63_1853 ();
 sg13g2_fill_1 FILLER_63_1910 ();
 sg13g2_fill_2 FILLER_63_1935 ();
 sg13g2_decap_8 FILLER_63_1989 ();
 sg13g2_decap_8 FILLER_63_1996 ();
 sg13g2_fill_1 FILLER_63_2003 ();
 sg13g2_fill_2 FILLER_63_2052 ();
 sg13g2_fill_1 FILLER_63_2054 ();
 sg13g2_fill_1 FILLER_63_2059 ();
 sg13g2_fill_1 FILLER_63_2081 ();
 sg13g2_fill_1 FILLER_63_2088 ();
 sg13g2_fill_2 FILLER_63_2178 ();
 sg13g2_decap_8 FILLER_63_2278 ();
 sg13g2_decap_4 FILLER_63_2285 ();
 sg13g2_fill_1 FILLER_63_2289 ();
 sg13g2_fill_1 FILLER_63_2313 ();
 sg13g2_decap_4 FILLER_63_2348 ();
 sg13g2_decap_8 FILLER_63_2356 ();
 sg13g2_fill_1 FILLER_63_2363 ();
 sg13g2_fill_1 FILLER_63_2377 ();
 sg13g2_fill_2 FILLER_63_2435 ();
 sg13g2_fill_1 FILLER_63_2463 ();
 sg13g2_decap_8 FILLER_63_2467 ();
 sg13g2_fill_2 FILLER_63_2474 ();
 sg13g2_fill_1 FILLER_63_2476 ();
 sg13g2_decap_8 FILLER_63_2481 ();
 sg13g2_fill_2 FILLER_63_2488 ();
 sg13g2_decap_8 FILLER_63_2537 ();
 sg13g2_decap_8 FILLER_63_2544 ();
 sg13g2_decap_4 FILLER_63_2551 ();
 sg13g2_fill_1 FILLER_63_2555 ();
 sg13g2_fill_2 FILLER_63_2595 ();
 sg13g2_decap_8 FILLER_63_2659 ();
 sg13g2_decap_4 FILLER_63_2666 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_fill_1 FILLER_64_65 ();
 sg13g2_decap_8 FILLER_64_74 ();
 sg13g2_decap_8 FILLER_64_90 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_decap_4 FILLER_64_110 ();
 sg13g2_fill_2 FILLER_64_114 ();
 sg13g2_fill_2 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_123 ();
 sg13g2_fill_1 FILLER_64_143 ();
 sg13g2_decap_4 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_decap_8 FILLER_64_157 ();
 sg13g2_decap_8 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_decap_4 FILLER_64_201 ();
 sg13g2_fill_1 FILLER_64_205 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_fill_2 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_decap_8 FILLER_64_332 ();
 sg13g2_decap_8 FILLER_64_339 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_2 FILLER_64_373 ();
 sg13g2_decap_4 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_64_453 ();
 sg13g2_fill_1 FILLER_64_500 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_2 FILLER_64_534 ();
 sg13g2_fill_1 FILLER_64_536 ();
 sg13g2_fill_2 FILLER_64_587 ();
 sg13g2_fill_2 FILLER_64_601 ();
 sg13g2_fill_2 FILLER_64_638 ();
 sg13g2_fill_2 FILLER_64_644 ();
 sg13g2_decap_8 FILLER_64_654 ();
 sg13g2_decap_4 FILLER_64_661 ();
 sg13g2_fill_1 FILLER_64_665 ();
 sg13g2_decap_8 FILLER_64_670 ();
 sg13g2_fill_2 FILLER_64_677 ();
 sg13g2_fill_1 FILLER_64_679 ();
 sg13g2_fill_2 FILLER_64_690 ();
 sg13g2_fill_1 FILLER_64_692 ();
 sg13g2_fill_1 FILLER_64_704 ();
 sg13g2_fill_1 FILLER_64_738 ();
 sg13g2_decap_4 FILLER_64_743 ();
 sg13g2_fill_1 FILLER_64_747 ();
 sg13g2_decap_4 FILLER_64_756 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_785 ();
 sg13g2_fill_2 FILLER_64_804 ();
 sg13g2_decap_4 FILLER_64_828 ();
 sg13g2_fill_1 FILLER_64_845 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_896 ();
 sg13g2_fill_2 FILLER_64_906 ();
 sg13g2_fill_1 FILLER_64_908 ();
 sg13g2_decap_8 FILLER_64_918 ();
 sg13g2_decap_8 FILLER_64_930 ();
 sg13g2_fill_2 FILLER_64_937 ();
 sg13g2_decap_4 FILLER_64_953 ();
 sg13g2_fill_1 FILLER_64_957 ();
 sg13g2_decap_8 FILLER_64_963 ();
 sg13g2_fill_2 FILLER_64_970 ();
 sg13g2_fill_1 FILLER_64_972 ();
 sg13g2_fill_1 FILLER_64_1004 ();
 sg13g2_decap_8 FILLER_64_1009 ();
 sg13g2_decap_8 FILLER_64_1016 ();
 sg13g2_decap_4 FILLER_64_1023 ();
 sg13g2_fill_2 FILLER_64_1030 ();
 sg13g2_fill_1 FILLER_64_1032 ();
 sg13g2_decap_4 FILLER_64_1072 ();
 sg13g2_decap_4 FILLER_64_1090 ();
 sg13g2_fill_2 FILLER_64_1111 ();
 sg13g2_fill_2 FILLER_64_1140 ();
 sg13g2_fill_1 FILLER_64_1142 ();
 sg13g2_decap_8 FILLER_64_1175 ();
 sg13g2_decap_4 FILLER_64_1182 ();
 sg13g2_decap_8 FILLER_64_1219 ();
 sg13g2_decap_8 FILLER_64_1226 ();
 sg13g2_decap_4 FILLER_64_1233 ();
 sg13g2_fill_1 FILLER_64_1237 ();
 sg13g2_fill_2 FILLER_64_1276 ();
 sg13g2_fill_1 FILLER_64_1278 ();
 sg13g2_fill_2 FILLER_64_1302 ();
 sg13g2_fill_1 FILLER_64_1304 ();
 sg13g2_fill_2 FILLER_64_1310 ();
 sg13g2_fill_1 FILLER_64_1317 ();
 sg13g2_decap_8 FILLER_64_1322 ();
 sg13g2_fill_2 FILLER_64_1329 ();
 sg13g2_decap_8 FILLER_64_1341 ();
 sg13g2_fill_2 FILLER_64_1348 ();
 sg13g2_decap_4 FILLER_64_1355 ();
 sg13g2_decap_4 FILLER_64_1365 ();
 sg13g2_decap_8 FILLER_64_1377 ();
 sg13g2_decap_4 FILLER_64_1384 ();
 sg13g2_fill_2 FILLER_64_1388 ();
 sg13g2_decap_8 FILLER_64_1403 ();
 sg13g2_decap_8 FILLER_64_1410 ();
 sg13g2_fill_2 FILLER_64_1417 ();
 sg13g2_fill_2 FILLER_64_1450 ();
 sg13g2_fill_2 FILLER_64_1487 ();
 sg13g2_fill_1 FILLER_64_1489 ();
 sg13g2_decap_8 FILLER_64_1520 ();
 sg13g2_fill_1 FILLER_64_1527 ();
 sg13g2_fill_1 FILLER_64_1531 ();
 sg13g2_fill_2 FILLER_64_1536 ();
 sg13g2_fill_2 FILLER_64_1551 ();
 sg13g2_decap_8 FILLER_64_1557 ();
 sg13g2_fill_2 FILLER_64_1564 ();
 sg13g2_fill_2 FILLER_64_1570 ();
 sg13g2_fill_1 FILLER_64_1572 ();
 sg13g2_fill_1 FILLER_64_1583 ();
 sg13g2_fill_2 FILLER_64_1588 ();
 sg13g2_fill_1 FILLER_64_1595 ();
 sg13g2_fill_1 FILLER_64_1600 ();
 sg13g2_fill_2 FILLER_64_1610 ();
 sg13g2_fill_2 FILLER_64_1617 ();
 sg13g2_fill_1 FILLER_64_1624 ();
 sg13g2_fill_1 FILLER_64_1632 ();
 sg13g2_fill_1 FILLER_64_1638 ();
 sg13g2_fill_1 FILLER_64_1643 ();
 sg13g2_fill_2 FILLER_64_1653 ();
 sg13g2_fill_2 FILLER_64_1660 ();
 sg13g2_fill_1 FILLER_64_1667 ();
 sg13g2_fill_2 FILLER_64_1683 ();
 sg13g2_fill_1 FILLER_64_1685 ();
 sg13g2_fill_1 FILLER_64_1752 ();
 sg13g2_fill_1 FILLER_64_1779 ();
 sg13g2_fill_1 FILLER_64_1786 ();
 sg13g2_decap_4 FILLER_64_1816 ();
 sg13g2_fill_2 FILLER_64_1834 ();
 sg13g2_decap_4 FILLER_64_1840 ();
 sg13g2_decap_4 FILLER_64_1849 ();
 sg13g2_fill_2 FILLER_64_1853 ();
 sg13g2_fill_1 FILLER_64_1861 ();
 sg13g2_decap_4 FILLER_64_1866 ();
 sg13g2_fill_1 FILLER_64_1875 ();
 sg13g2_fill_2 FILLER_64_1886 ();
 sg13g2_decap_8 FILLER_64_1892 ();
 sg13g2_decap_8 FILLER_64_1899 ();
 sg13g2_fill_1 FILLER_64_1906 ();
 sg13g2_decap_4 FILLER_64_1919 ();
 sg13g2_fill_2 FILLER_64_1923 ();
 sg13g2_decap_8 FILLER_64_1951 ();
 sg13g2_decap_8 FILLER_64_1958 ();
 sg13g2_decap_4 FILLER_64_1965 ();
 sg13g2_fill_2 FILLER_64_1969 ();
 sg13g2_decap_4 FILLER_64_1975 ();
 sg13g2_decap_4 FILLER_64_1983 ();
 sg13g2_fill_2 FILLER_64_2002 ();
 sg13g2_fill_2 FILLER_64_2030 ();
 sg13g2_fill_1 FILLER_64_2032 ();
 sg13g2_fill_2 FILLER_64_2037 ();
 sg13g2_fill_1 FILLER_64_2039 ();
 sg13g2_fill_2 FILLER_64_2066 ();
 sg13g2_fill_1 FILLER_64_2068 ();
 sg13g2_fill_1 FILLER_64_2118 ();
 sg13g2_fill_1 FILLER_64_2124 ();
 sg13g2_fill_2 FILLER_64_2130 ();
 sg13g2_fill_2 FILLER_64_2153 ();
 sg13g2_fill_1 FILLER_64_2170 ();
 sg13g2_fill_2 FILLER_64_2192 ();
 sg13g2_fill_1 FILLER_64_2194 ();
 sg13g2_fill_1 FILLER_64_2272 ();
 sg13g2_fill_2 FILLER_64_2303 ();
 sg13g2_fill_2 FILLER_64_2309 ();
 sg13g2_fill_2 FILLER_64_2328 ();
 sg13g2_fill_1 FILLER_64_2334 ();
 sg13g2_decap_8 FILLER_64_2345 ();
 sg13g2_fill_1 FILLER_64_2388 ();
 sg13g2_fill_1 FILLER_64_2399 ();
 sg13g2_fill_1 FILLER_64_2426 ();
 sg13g2_fill_1 FILLER_64_2437 ();
 sg13g2_decap_8 FILLER_64_2469 ();
 sg13g2_decap_8 FILLER_64_2476 ();
 sg13g2_decap_8 FILLER_64_2483 ();
 sg13g2_fill_2 FILLER_64_2490 ();
 sg13g2_decap_4 FILLER_64_2554 ();
 sg13g2_fill_2 FILLER_64_2558 ();
 sg13g2_decap_8 FILLER_64_2572 ();
 sg13g2_decap_8 FILLER_64_2579 ();
 sg13g2_fill_1 FILLER_64_2586 ();
 sg13g2_decap_8 FILLER_64_2591 ();
 sg13g2_decap_8 FILLER_64_2598 ();
 sg13g2_fill_2 FILLER_64_2605 ();
 sg13g2_fill_1 FILLER_64_2607 ();
 sg13g2_decap_8 FILLER_64_2626 ();
 sg13g2_decap_8 FILLER_64_2633 ();
 sg13g2_decap_8 FILLER_64_2640 ();
 sg13g2_decap_8 FILLER_64_2647 ();
 sg13g2_decap_8 FILLER_64_2654 ();
 sg13g2_decap_8 FILLER_64_2661 ();
 sg13g2_fill_2 FILLER_64_2668 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_15 ();
 sg13g2_fill_2 FILLER_65_26 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_49 ();
 sg13g2_fill_1 FILLER_65_51 ();
 sg13g2_fill_2 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_103 ();
 sg13g2_fill_1 FILLER_65_105 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_decap_8 FILLER_65_174 ();
 sg13g2_decap_8 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_fill_2 FILLER_65_295 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_2 FILLER_65_362 ();
 sg13g2_fill_1 FILLER_65_475 ();
 sg13g2_decap_4 FILLER_65_521 ();
 sg13g2_fill_1 FILLER_65_556 ();
 sg13g2_fill_1 FILLER_65_562 ();
 sg13g2_fill_1 FILLER_65_609 ();
 sg13g2_fill_2 FILLER_65_636 ();
 sg13g2_fill_1 FILLER_65_638 ();
 sg13g2_fill_1 FILLER_65_647 ();
 sg13g2_decap_4 FILLER_65_652 ();
 sg13g2_fill_1 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_663 ();
 sg13g2_fill_2 FILLER_65_696 ();
 sg13g2_fill_1 FILLER_65_698 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_fill_2 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_750 ();
 sg13g2_fill_2 FILLER_65_757 ();
 sg13g2_decap_4 FILLER_65_800 ();
 sg13g2_fill_2 FILLER_65_804 ();
 sg13g2_fill_1 FILLER_65_812 ();
 sg13g2_fill_2 FILLER_65_826 ();
 sg13g2_fill_1 FILLER_65_832 ();
 sg13g2_fill_1 FILLER_65_851 ();
 sg13g2_fill_2 FILLER_65_856 ();
 sg13g2_fill_1 FILLER_65_858 ();
 sg13g2_fill_2 FILLER_65_874 ();
 sg13g2_decap_8 FILLER_65_912 ();
 sg13g2_decap_4 FILLER_65_923 ();
 sg13g2_fill_1 FILLER_65_931 ();
 sg13g2_decap_8 FILLER_65_944 ();
 sg13g2_fill_1 FILLER_65_955 ();
 sg13g2_decap_8 FILLER_65_961 ();
 sg13g2_decap_4 FILLER_65_968 ();
 sg13g2_fill_1 FILLER_65_978 ();
 sg13g2_decap_4 FILLER_65_984 ();
 sg13g2_decap_8 FILLER_65_993 ();
 sg13g2_decap_8 FILLER_65_1000 ();
 sg13g2_decap_4 FILLER_65_1007 ();
 sg13g2_fill_2 FILLER_65_1011 ();
 sg13g2_fill_2 FILLER_65_1018 ();
 sg13g2_fill_1 FILLER_65_1020 ();
 sg13g2_fill_2 FILLER_65_1025 ();
 sg13g2_fill_1 FILLER_65_1027 ();
 sg13g2_fill_1 FILLER_65_1052 ();
 sg13g2_fill_2 FILLER_65_1082 ();
 sg13g2_fill_1 FILLER_65_1089 ();
 sg13g2_fill_1 FILLER_65_1100 ();
 sg13g2_fill_1 FILLER_65_1127 ();
 sg13g2_decap_8 FILLER_65_1154 ();
 sg13g2_decap_8 FILLER_65_1161 ();
 sg13g2_decap_4 FILLER_65_1172 ();
 sg13g2_fill_2 FILLER_65_1176 ();
 sg13g2_fill_1 FILLER_65_1252 ();
 sg13g2_fill_2 FILLER_65_1263 ();
 sg13g2_fill_1 FILLER_65_1273 ();
 sg13g2_fill_2 FILLER_65_1279 ();
 sg13g2_fill_1 FILLER_65_1281 ();
 sg13g2_decap_4 FILLER_65_1289 ();
 sg13g2_fill_1 FILLER_65_1305 ();
 sg13g2_fill_1 FILLER_65_1322 ();
 sg13g2_fill_2 FILLER_65_1327 ();
 sg13g2_fill_1 FILLER_65_1339 ();
 sg13g2_fill_1 FILLER_65_1377 ();
 sg13g2_fill_1 FILLER_65_1382 ();
 sg13g2_fill_1 FILLER_65_1391 ();
 sg13g2_decap_8 FILLER_65_1406 ();
 sg13g2_decap_8 FILLER_65_1413 ();
 sg13g2_decap_4 FILLER_65_1420 ();
 sg13g2_fill_2 FILLER_65_1428 ();
 sg13g2_fill_1 FILLER_65_1430 ();
 sg13g2_decap_4 FILLER_65_1444 ();
 sg13g2_fill_1 FILLER_65_1448 ();
 sg13g2_decap_8 FILLER_65_1454 ();
 sg13g2_fill_2 FILLER_65_1461 ();
 sg13g2_fill_1 FILLER_65_1463 ();
 sg13g2_fill_1 FILLER_65_1468 ();
 sg13g2_fill_1 FILLER_65_1472 ();
 sg13g2_fill_2 FILLER_65_1477 ();
 sg13g2_fill_1 FILLER_65_1483 ();
 sg13g2_fill_1 FILLER_65_1493 ();
 sg13g2_decap_4 FILLER_65_1499 ();
 sg13g2_decap_8 FILLER_65_1509 ();
 sg13g2_fill_2 FILLER_65_1516 ();
 sg13g2_fill_2 FILLER_65_1528 ();
 sg13g2_fill_1 FILLER_65_1539 ();
 sg13g2_fill_1 FILLER_65_1577 ();
 sg13g2_fill_2 FILLER_65_1586 ();
 sg13g2_fill_1 FILLER_65_1588 ();
 sg13g2_fill_1 FILLER_65_1599 ();
 sg13g2_fill_1 FILLER_65_1604 ();
 sg13g2_decap_4 FILLER_65_1610 ();
 sg13g2_fill_1 FILLER_65_1614 ();
 sg13g2_fill_2 FILLER_65_1633 ();
 sg13g2_fill_2 FILLER_65_1639 ();
 sg13g2_fill_1 FILLER_65_1649 ();
 sg13g2_fill_2 FILLER_65_1655 ();
 sg13g2_fill_1 FILLER_65_1657 ();
 sg13g2_decap_8 FILLER_65_1720 ();
 sg13g2_fill_2 FILLER_65_1727 ();
 sg13g2_fill_1 FILLER_65_1729 ();
 sg13g2_fill_1 FILLER_65_1748 ();
 sg13g2_fill_1 FILLER_65_1753 ();
 sg13g2_fill_1 FILLER_65_1784 ();
 sg13g2_fill_2 FILLER_65_1791 ();
 sg13g2_fill_1 FILLER_65_1805 ();
 sg13g2_decap_8 FILLER_65_1822 ();
 sg13g2_fill_2 FILLER_65_1839 ();
 sg13g2_fill_2 FILLER_65_1847 ();
 sg13g2_fill_2 FILLER_65_1870 ();
 sg13g2_decap_4 FILLER_65_1884 ();
 sg13g2_fill_1 FILLER_65_1888 ();
 sg13g2_fill_2 FILLER_65_1935 ();
 sg13g2_fill_1 FILLER_65_1937 ();
 sg13g2_fill_1 FILLER_65_1942 ();
 sg13g2_fill_1 FILLER_65_1949 ();
 sg13g2_decap_4 FILLER_65_1973 ();
 sg13g2_fill_2 FILLER_65_1977 ();
 sg13g2_fill_2 FILLER_65_2018 ();
 sg13g2_fill_1 FILLER_65_2020 ();
 sg13g2_fill_1 FILLER_65_2051 ();
 sg13g2_fill_2 FILLER_65_2065 ();
 sg13g2_fill_1 FILLER_65_2124 ();
 sg13g2_decap_8 FILLER_65_2195 ();
 sg13g2_decap_4 FILLER_65_2202 ();
 sg13g2_fill_2 FILLER_65_2206 ();
 sg13g2_fill_1 FILLER_65_2350 ();
 sg13g2_fill_1 FILLER_65_2377 ();
 sg13g2_fill_2 FILLER_65_2386 ();
 sg13g2_fill_2 FILLER_65_2396 ();
 sg13g2_fill_2 FILLER_65_2408 ();
 sg13g2_decap_4 FILLER_65_2414 ();
 sg13g2_fill_2 FILLER_65_2418 ();
 sg13g2_fill_2 FILLER_65_2454 ();
 sg13g2_fill_1 FILLER_65_2476 ();
 sg13g2_fill_2 FILLER_65_2490 ();
 sg13g2_fill_1 FILLER_65_2492 ();
 sg13g2_decap_8 FILLER_65_2497 ();
 sg13g2_decap_4 FILLER_65_2504 ();
 sg13g2_fill_1 FILLER_65_2512 ();
 sg13g2_decap_4 FILLER_65_2534 ();
 sg13g2_fill_1 FILLER_65_2538 ();
 sg13g2_decap_8 FILLER_65_2565 ();
 sg13g2_decap_8 FILLER_65_2572 ();
 sg13g2_fill_2 FILLER_65_2579 ();
 sg13g2_decap_8 FILLER_65_2602 ();
 sg13g2_decap_8 FILLER_65_2609 ();
 sg13g2_decap_8 FILLER_65_2616 ();
 sg13g2_decap_8 FILLER_65_2623 ();
 sg13g2_decap_8 FILLER_65_2630 ();
 sg13g2_decap_8 FILLER_65_2637 ();
 sg13g2_decap_8 FILLER_65_2644 ();
 sg13g2_decap_8 FILLER_65_2651 ();
 sg13g2_decap_8 FILLER_65_2658 ();
 sg13g2_decap_4 FILLER_65_2665 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_33 ();
 sg13g2_decap_8 FILLER_66_40 ();
 sg13g2_fill_2 FILLER_66_47 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_4 FILLER_66_63 ();
 sg13g2_fill_2 FILLER_66_67 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_fill_1 FILLER_66_176 ();
 sg13g2_fill_2 FILLER_66_185 ();
 sg13g2_decap_4 FILLER_66_202 ();
 sg13g2_fill_1 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_1 FILLER_66_275 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_317 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_decap_8 FILLER_66_346 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_fill_1 FILLER_66_384 ();
 sg13g2_fill_1 FILLER_66_397 ();
 sg13g2_decap_4 FILLER_66_471 ();
 sg13g2_fill_1 FILLER_66_489 ();
 sg13g2_fill_1 FILLER_66_494 ();
 sg13g2_fill_1 FILLER_66_500 ();
 sg13g2_fill_1 FILLER_66_506 ();
 sg13g2_fill_1 FILLER_66_516 ();
 sg13g2_fill_2 FILLER_66_522 ();
 sg13g2_decap_4 FILLER_66_528 ();
 sg13g2_fill_2 FILLER_66_532 ();
 sg13g2_fill_1 FILLER_66_555 ();
 sg13g2_fill_1 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_577 ();
 sg13g2_fill_1 FILLER_66_622 ();
 sg13g2_fill_1 FILLER_66_627 ();
 sg13g2_decap_8 FILLER_66_641 ();
 sg13g2_decap_4 FILLER_66_648 ();
 sg13g2_fill_1 FILLER_66_652 ();
 sg13g2_fill_2 FILLER_66_661 ();
 sg13g2_fill_2 FILLER_66_676 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_decap_4 FILLER_66_709 ();
 sg13g2_fill_1 FILLER_66_729 ();
 sg13g2_fill_2 FILLER_66_734 ();
 sg13g2_fill_1 FILLER_66_736 ();
 sg13g2_decap_8 FILLER_66_771 ();
 sg13g2_decap_8 FILLER_66_782 ();
 sg13g2_decap_8 FILLER_66_789 ();
 sg13g2_fill_1 FILLER_66_796 ();
 sg13g2_decap_4 FILLER_66_805 ();
 sg13g2_fill_2 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_fill_1 FILLER_66_856 ();
 sg13g2_fill_1 FILLER_66_867 ();
 sg13g2_fill_1 FILLER_66_874 ();
 sg13g2_fill_1 FILLER_66_889 ();
 sg13g2_fill_2 FILLER_66_896 ();
 sg13g2_fill_1 FILLER_66_906 ();
 sg13g2_decap_8 FILLER_66_911 ();
 sg13g2_fill_1 FILLER_66_918 ();
 sg13g2_decap_4 FILLER_66_933 ();
 sg13g2_fill_1 FILLER_66_937 ();
 sg13g2_decap_8 FILLER_66_945 ();
 sg13g2_fill_1 FILLER_66_952 ();
 sg13g2_fill_1 FILLER_66_975 ();
 sg13g2_fill_2 FILLER_66_981 ();
 sg13g2_decap_4 FILLER_66_990 ();
 sg13g2_decap_8 FILLER_66_998 ();
 sg13g2_decap_8 FILLER_66_1019 ();
 sg13g2_fill_2 FILLER_66_1047 ();
 sg13g2_fill_2 FILLER_66_1053 ();
 sg13g2_fill_1 FILLER_66_1055 ();
 sg13g2_decap_4 FILLER_66_1064 ();
 sg13g2_fill_1 FILLER_66_1078 ();
 sg13g2_fill_1 FILLER_66_1083 ();
 sg13g2_fill_2 FILLER_66_1089 ();
 sg13g2_fill_2 FILLER_66_1100 ();
 sg13g2_decap_8 FILLER_66_1137 ();
 sg13g2_fill_2 FILLER_66_1144 ();
 sg13g2_decap_8 FILLER_66_1155 ();
 sg13g2_decap_8 FILLER_66_1162 ();
 sg13g2_fill_2 FILLER_66_1169 ();
 sg13g2_fill_2 FILLER_66_1174 ();
 sg13g2_fill_1 FILLER_66_1176 ();
 sg13g2_fill_1 FILLER_66_1181 ();
 sg13g2_fill_1 FILLER_66_1196 ();
 sg13g2_decap_4 FILLER_66_1227 ();
 sg13g2_fill_1 FILLER_66_1231 ();
 sg13g2_fill_2 FILLER_66_1236 ();
 sg13g2_fill_1 FILLER_66_1238 ();
 sg13g2_decap_8 FILLER_66_1246 ();
 sg13g2_decap_8 FILLER_66_1253 ();
 sg13g2_decap_8 FILLER_66_1260 ();
 sg13g2_fill_1 FILLER_66_1267 ();
 sg13g2_fill_2 FILLER_66_1273 ();
 sg13g2_fill_1 FILLER_66_1275 ();
 sg13g2_fill_1 FILLER_66_1296 ();
 sg13g2_fill_1 FILLER_66_1303 ();
 sg13g2_fill_1 FILLER_66_1315 ();
 sg13g2_fill_1 FILLER_66_1335 ();
 sg13g2_fill_1 FILLER_66_1345 ();
 sg13g2_decap_4 FILLER_66_1350 ();
 sg13g2_fill_2 FILLER_66_1372 ();
 sg13g2_fill_1 FILLER_66_1390 ();
 sg13g2_decap_8 FILLER_66_1409 ();
 sg13g2_decap_8 FILLER_66_1416 ();
 sg13g2_fill_1 FILLER_66_1423 ();
 sg13g2_fill_2 FILLER_66_1432 ();
 sg13g2_decap_8 FILLER_66_1470 ();
 sg13g2_decap_8 FILLER_66_1477 ();
 sg13g2_decap_8 FILLER_66_1484 ();
 sg13g2_fill_2 FILLER_66_1491 ();
 sg13g2_fill_1 FILLER_66_1493 ();
 sg13g2_fill_1 FILLER_66_1502 ();
 sg13g2_fill_2 FILLER_66_1512 ();
 sg13g2_decap_8 FILLER_66_1572 ();
 sg13g2_fill_2 FILLER_66_1628 ();
 sg13g2_fill_2 FILLER_66_1633 ();
 sg13g2_decap_4 FILLER_66_1659 ();
 sg13g2_fill_2 FILLER_66_1663 ();
 sg13g2_decap_8 FILLER_66_1669 ();
 sg13g2_decap_8 FILLER_66_1676 ();
 sg13g2_fill_2 FILLER_66_1683 ();
 sg13g2_fill_1 FILLER_66_1685 ();
 sg13g2_fill_2 FILLER_66_1726 ();
 sg13g2_fill_2 FILLER_66_1776 ();
 sg13g2_fill_1 FILLER_66_1846 ();
 sg13g2_fill_2 FILLER_66_1851 ();
 sg13g2_fill_1 FILLER_66_1853 ();
 sg13g2_decap_8 FILLER_66_1858 ();
 sg13g2_fill_1 FILLER_66_1865 ();
 sg13g2_decap_8 FILLER_66_1874 ();
 sg13g2_fill_1 FILLER_66_1881 ();
 sg13g2_decap_4 FILLER_66_1894 ();
 sg13g2_fill_1 FILLER_66_1898 ();
 sg13g2_fill_2 FILLER_66_1903 ();
 sg13g2_decap_4 FILLER_66_1909 ();
 sg13g2_fill_1 FILLER_66_1913 ();
 sg13g2_decap_4 FILLER_66_1924 ();
 sg13g2_decap_8 FILLER_66_1954 ();
 sg13g2_fill_2 FILLER_66_2016 ();
 sg13g2_decap_8 FILLER_66_2022 ();
 sg13g2_decap_8 FILLER_66_2029 ();
 sg13g2_decap_8 FILLER_66_2039 ();
 sg13g2_decap_4 FILLER_66_2046 ();
 sg13g2_fill_1 FILLER_66_2050 ();
 sg13g2_decap_8 FILLER_66_2055 ();
 sg13g2_fill_1 FILLER_66_2062 ();
 sg13g2_decap_8 FILLER_66_2067 ();
 sg13g2_decap_4 FILLER_66_2074 ();
 sg13g2_fill_2 FILLER_66_2090 ();
 sg13g2_fill_1 FILLER_66_2096 ();
 sg13g2_fill_1 FILLER_66_2219 ();
 sg13g2_decap_8 FILLER_66_2273 ();
 sg13g2_fill_1 FILLER_66_2284 ();
 sg13g2_fill_1 FILLER_66_2293 ();
 sg13g2_fill_2 FILLER_66_2331 ();
 sg13g2_fill_1 FILLER_66_2333 ();
 sg13g2_fill_2 FILLER_66_2393 ();
 sg13g2_decap_8 FILLER_66_2407 ();
 sg13g2_decap_4 FILLER_66_2414 ();
 sg13g2_fill_2 FILLER_66_2418 ();
 sg13g2_decap_8 FILLER_66_2430 ();
 sg13g2_decap_8 FILLER_66_2437 ();
 sg13g2_fill_1 FILLER_66_2444 ();
 sg13g2_fill_1 FILLER_66_2479 ();
 sg13g2_decap_4 FILLER_66_2514 ();
 sg13g2_fill_2 FILLER_66_2518 ();
 sg13g2_fill_2 FILLER_66_2530 ();
 sg13g2_fill_1 FILLER_66_2532 ();
 sg13g2_fill_2 FILLER_66_2543 ();
 sg13g2_fill_1 FILLER_66_2545 ();
 sg13g2_decap_8 FILLER_66_2550 ();
 sg13g2_decap_4 FILLER_66_2557 ();
 sg13g2_decap_8 FILLER_66_2627 ();
 sg13g2_decap_8 FILLER_66_2634 ();
 sg13g2_decap_8 FILLER_66_2641 ();
 sg13g2_decap_8 FILLER_66_2648 ();
 sg13g2_decap_8 FILLER_66_2655 ();
 sg13g2_decap_8 FILLER_66_2662 ();
 sg13g2_fill_1 FILLER_66_2669 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_50 ();
 sg13g2_decap_8 FILLER_67_64 ();
 sg13g2_fill_2 FILLER_67_71 ();
 sg13g2_fill_1 FILLER_67_73 ();
 sg13g2_fill_2 FILLER_67_128 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_decap_4 FILLER_67_136 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_185 ();
 sg13g2_fill_1 FILLER_67_187 ();
 sg13g2_decap_4 FILLER_67_196 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_294 ();
 sg13g2_fill_2 FILLER_67_300 ();
 sg13g2_fill_1 FILLER_67_307 ();
 sg13g2_fill_1 FILLER_67_334 ();
 sg13g2_decap_8 FILLER_67_386 ();
 sg13g2_fill_1 FILLER_67_393 ();
 sg13g2_decap_4 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_2 FILLER_67_417 ();
 sg13g2_decap_8 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_511 ();
 sg13g2_decap_4 FILLER_67_518 ();
 sg13g2_fill_1 FILLER_67_522 ();
 sg13g2_fill_2 FILLER_67_527 ();
 sg13g2_fill_1 FILLER_67_529 ();
 sg13g2_decap_4 FILLER_67_540 ();
 sg13g2_fill_1 FILLER_67_544 ();
 sg13g2_fill_1 FILLER_67_560 ();
 sg13g2_fill_1 FILLER_67_607 ();
 sg13g2_fill_2 FILLER_67_630 ();
 sg13g2_fill_1 FILLER_67_658 ();
 sg13g2_decap_8 FILLER_67_690 ();
 sg13g2_decap_8 FILLER_67_697 ();
 sg13g2_fill_1 FILLER_67_704 ();
 sg13g2_fill_1 FILLER_67_743 ();
 sg13g2_fill_2 FILLER_67_758 ();
 sg13g2_fill_1 FILLER_67_760 ();
 sg13g2_decap_4 FILLER_67_765 ();
 sg13g2_decap_8 FILLER_67_774 ();
 sg13g2_decap_8 FILLER_67_781 ();
 sg13g2_decap_8 FILLER_67_788 ();
 sg13g2_decap_8 FILLER_67_795 ();
 sg13g2_fill_2 FILLER_67_802 ();
 sg13g2_decap_8 FILLER_67_809 ();
 sg13g2_fill_1 FILLER_67_816 ();
 sg13g2_fill_1 FILLER_67_836 ();
 sg13g2_fill_1 FILLER_67_849 ();
 sg13g2_fill_1 FILLER_67_858 ();
 sg13g2_fill_2 FILLER_67_867 ();
 sg13g2_fill_1 FILLER_67_869 ();
 sg13g2_decap_8 FILLER_67_885 ();
 sg13g2_fill_2 FILLER_67_892 ();
 sg13g2_fill_2 FILLER_67_904 ();
 sg13g2_fill_2 FILLER_67_920 ();
 sg13g2_fill_1 FILLER_67_927 ();
 sg13g2_decap_4 FILLER_67_933 ();
 sg13g2_fill_1 FILLER_67_937 ();
 sg13g2_decap_4 FILLER_67_942 ();
 sg13g2_fill_1 FILLER_67_953 ();
 sg13g2_decap_4 FILLER_67_959 ();
 sg13g2_fill_1 FILLER_67_963 ();
 sg13g2_decap_4 FILLER_67_975 ();
 sg13g2_decap_8 FILLER_67_985 ();
 sg13g2_decap_4 FILLER_67_992 ();
 sg13g2_fill_2 FILLER_67_996 ();
 sg13g2_fill_2 FILLER_67_1002 ();
 sg13g2_fill_2 FILLER_67_1009 ();
 sg13g2_decap_4 FILLER_67_1016 ();
 sg13g2_fill_1 FILLER_67_1020 ();
 sg13g2_decap_8 FILLER_67_1032 ();
 sg13g2_decap_4 FILLER_67_1039 ();
 sg13g2_decap_8 FILLER_67_1048 ();
 sg13g2_decap_8 FILLER_67_1055 ();
 sg13g2_decap_8 FILLER_67_1062 ();
 sg13g2_decap_8 FILLER_67_1069 ();
 sg13g2_decap_8 FILLER_67_1076 ();
 sg13g2_decap_4 FILLER_67_1083 ();
 sg13g2_fill_2 FILLER_67_1087 ();
 sg13g2_fill_1 FILLER_67_1098 ();
 sg13g2_fill_1 FILLER_67_1107 ();
 sg13g2_fill_2 FILLER_67_1121 ();
 sg13g2_fill_1 FILLER_67_1123 ();
 sg13g2_fill_2 FILLER_67_1129 ();
 sg13g2_decap_8 FILLER_67_1146 ();
 sg13g2_decap_4 FILLER_67_1153 ();
 sg13g2_decap_4 FILLER_67_1194 ();
 sg13g2_fill_2 FILLER_67_1198 ();
 sg13g2_decap_8 FILLER_67_1209 ();
 sg13g2_fill_1 FILLER_67_1216 ();
 sg13g2_decap_8 FILLER_67_1253 ();
 sg13g2_decap_8 FILLER_67_1260 ();
 sg13g2_decap_8 FILLER_67_1267 ();
 sg13g2_decap_8 FILLER_67_1274 ();
 sg13g2_fill_2 FILLER_67_1311 ();
 sg13g2_fill_2 FILLER_67_1317 ();
 sg13g2_fill_1 FILLER_67_1319 ();
 sg13g2_fill_1 FILLER_67_1344 ();
 sg13g2_fill_1 FILLER_67_1350 ();
 sg13g2_fill_1 FILLER_67_1360 ();
 sg13g2_fill_1 FILLER_67_1365 ();
 sg13g2_fill_2 FILLER_67_1375 ();
 sg13g2_fill_2 FILLER_67_1410 ();
 sg13g2_fill_1 FILLER_67_1428 ();
 sg13g2_fill_1 FILLER_67_1433 ();
 sg13g2_fill_2 FILLER_67_1444 ();
 sg13g2_fill_1 FILLER_67_1472 ();
 sg13g2_decap_8 FILLER_67_1478 ();
 sg13g2_fill_2 FILLER_67_1485 ();
 sg13g2_fill_1 FILLER_67_1487 ();
 sg13g2_decap_8 FILLER_67_1493 ();
 sg13g2_fill_2 FILLER_67_1505 ();
 sg13g2_fill_1 FILLER_67_1519 ();
 sg13g2_fill_1 FILLER_67_1528 ();
 sg13g2_fill_1 FILLER_67_1532 ();
 sg13g2_fill_1 FILLER_67_1564 ();
 sg13g2_fill_2 FILLER_67_1569 ();
 sg13g2_fill_2 FILLER_67_1581 ();
 sg13g2_fill_2 FILLER_67_1590 ();
 sg13g2_fill_1 FILLER_67_1592 ();
 sg13g2_fill_2 FILLER_67_1625 ();
 sg13g2_fill_1 FILLER_67_1636 ();
 sg13g2_fill_1 FILLER_67_1665 ();
 sg13g2_fill_1 FILLER_67_1697 ();
 sg13g2_decap_4 FILLER_67_1703 ();
 sg13g2_fill_1 FILLER_67_1707 ();
 sg13g2_fill_2 FILLER_67_1725 ();
 sg13g2_fill_1 FILLER_67_1731 ();
 sg13g2_fill_1 FILLER_67_1758 ();
 sg13g2_decap_8 FILLER_67_1767 ();
 sg13g2_decap_4 FILLER_67_1774 ();
 sg13g2_fill_1 FILLER_67_1778 ();
 sg13g2_decap_4 FILLER_67_1805 ();
 sg13g2_fill_2 FILLER_67_1809 ();
 sg13g2_decap_8 FILLER_67_1922 ();
 sg13g2_decap_4 FILLER_67_1929 ();
 sg13g2_decap_4 FILLER_67_1943 ();
 sg13g2_fill_2 FILLER_67_1947 ();
 sg13g2_fill_1 FILLER_67_1953 ();
 sg13g2_fill_1 FILLER_67_1974 ();
 sg13g2_fill_2 FILLER_67_1996 ();
 sg13g2_decap_4 FILLER_67_2024 ();
 sg13g2_fill_1 FILLER_67_2032 ();
 sg13g2_fill_2 FILLER_67_2041 ();
 sg13g2_fill_1 FILLER_67_2043 ();
 sg13g2_fill_1 FILLER_67_2080 ();
 sg13g2_decap_4 FILLER_67_2091 ();
 sg13g2_fill_1 FILLER_67_2095 ();
 sg13g2_fill_1 FILLER_67_2105 ();
 sg13g2_fill_2 FILLER_67_2147 ();
 sg13g2_fill_2 FILLER_67_2160 ();
 sg13g2_fill_1 FILLER_67_2171 ();
 sg13g2_decap_4 FILLER_67_2213 ();
 sg13g2_fill_1 FILLER_67_2217 ();
 sg13g2_fill_1 FILLER_67_2230 ();
 sg13g2_decap_8 FILLER_67_2284 ();
 sg13g2_fill_2 FILLER_67_2291 ();
 sg13g2_fill_1 FILLER_67_2342 ();
 sg13g2_fill_2 FILLER_67_2347 ();
 sg13g2_fill_2 FILLER_67_2353 ();
 sg13g2_decap_4 FILLER_67_2448 ();
 sg13g2_fill_1 FILLER_67_2452 ();
 sg13g2_decap_4 FILLER_67_2500 ();
 sg13g2_fill_2 FILLER_67_2508 ();
 sg13g2_decap_4 FILLER_67_2560 ();
 sg13g2_fill_2 FILLER_67_2564 ();
 sg13g2_decap_8 FILLER_67_2619 ();
 sg13g2_decap_8 FILLER_67_2626 ();
 sg13g2_decap_8 FILLER_67_2633 ();
 sg13g2_decap_8 FILLER_67_2640 ();
 sg13g2_decap_8 FILLER_67_2647 ();
 sg13g2_decap_8 FILLER_67_2654 ();
 sg13g2_decap_8 FILLER_67_2661 ();
 sg13g2_fill_2 FILLER_67_2668 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_2 FILLER_68_17 ();
 sg13g2_fill_1 FILLER_68_51 ();
 sg13g2_decap_4 FILLER_68_68 ();
 sg13g2_decap_4 FILLER_68_98 ();
 sg13g2_fill_1 FILLER_68_106 ();
 sg13g2_fill_2 FILLER_68_143 ();
 sg13g2_fill_2 FILLER_68_149 ();
 sg13g2_fill_1 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_157 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_fill_1 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_195 ();
 sg13g2_fill_2 FILLER_68_201 ();
 sg13g2_fill_1 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_248 ();
 sg13g2_fill_2 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_270 ();
 sg13g2_fill_1 FILLER_68_294 ();
 sg13g2_fill_2 FILLER_68_299 ();
 sg13g2_fill_2 FILLER_68_305 ();
 sg13g2_fill_1 FILLER_68_322 ();
 sg13g2_fill_1 FILLER_68_327 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_decap_4 FILLER_68_346 ();
 sg13g2_fill_2 FILLER_68_353 ();
 sg13g2_fill_2 FILLER_68_386 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_2 FILLER_68_431 ();
 sg13g2_fill_1 FILLER_68_451 ();
 sg13g2_fill_2 FILLER_68_461 ();
 sg13g2_fill_1 FILLER_68_463 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_fill_2 FILLER_68_476 ();
 sg13g2_fill_2 FILLER_68_488 ();
 sg13g2_fill_2 FILLER_68_500 ();
 sg13g2_decap_4 FILLER_68_506 ();
 sg13g2_fill_1 FILLER_68_510 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_542 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_586 ();
 sg13g2_decap_8 FILLER_68_593 ();
 sg13g2_decap_4 FILLER_68_600 ();
 sg13g2_decap_4 FILLER_68_661 ();
 sg13g2_decap_4 FILLER_68_695 ();
 sg13g2_fill_2 FILLER_68_699 ();
 sg13g2_decap_8 FILLER_68_709 ();
 sg13g2_fill_2 FILLER_68_716 ();
 sg13g2_fill_2 FILLER_68_736 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_fill_2 FILLER_68_768 ();
 sg13g2_fill_1 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_797 ();
 sg13g2_decap_8 FILLER_68_804 ();
 sg13g2_decap_4 FILLER_68_811 ();
 sg13g2_fill_2 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_821 ();
 sg13g2_decap_8 FILLER_68_828 ();
 sg13g2_decap_8 FILLER_68_835 ();
 sg13g2_decap_4 FILLER_68_849 ();
 sg13g2_fill_2 FILLER_68_853 ();
 sg13g2_fill_1 FILLER_68_869 ();
 sg13g2_fill_2 FILLER_68_879 ();
 sg13g2_fill_1 FILLER_68_881 ();
 sg13g2_decap_8 FILLER_68_885 ();
 sg13g2_decap_8 FILLER_68_892 ();
 sg13g2_decap_8 FILLER_68_899 ();
 sg13g2_fill_2 FILLER_68_906 ();
 sg13g2_fill_1 FILLER_68_908 ();
 sg13g2_decap_4 FILLER_68_914 ();
 sg13g2_fill_1 FILLER_68_931 ();
 sg13g2_fill_2 FILLER_68_937 ();
 sg13g2_fill_1 FILLER_68_944 ();
 sg13g2_fill_2 FILLER_68_972 ();
 sg13g2_fill_1 FILLER_68_974 ();
 sg13g2_fill_2 FILLER_68_1004 ();
 sg13g2_fill_1 FILLER_68_1025 ();
 sg13g2_decap_4 FILLER_68_1029 ();
 sg13g2_decap_8 FILLER_68_1043 ();
 sg13g2_fill_2 FILLER_68_1050 ();
 sg13g2_fill_1 FILLER_68_1052 ();
 sg13g2_fill_2 FILLER_68_1057 ();
 sg13g2_fill_1 FILLER_68_1059 ();
 sg13g2_decap_8 FILLER_68_1069 ();
 sg13g2_fill_1 FILLER_68_1076 ();
 sg13g2_fill_1 FILLER_68_1105 ();
 sg13g2_decap_4 FILLER_68_1121 ();
 sg13g2_fill_1 FILLER_68_1125 ();
 sg13g2_decap_8 FILLER_68_1130 ();
 sg13g2_decap_8 FILLER_68_1141 ();
 sg13g2_decap_4 FILLER_68_1148 ();
 sg13g2_decap_4 FILLER_68_1163 ();
 sg13g2_fill_2 FILLER_68_1167 ();
 sg13g2_decap_4 FILLER_68_1177 ();
 sg13g2_decap_8 FILLER_68_1199 ();
 sg13g2_decap_4 FILLER_68_1206 ();
 sg13g2_fill_1 FILLER_68_1210 ();
 sg13g2_decap_8 FILLER_68_1242 ();
 sg13g2_decap_8 FILLER_68_1249 ();
 sg13g2_decap_8 FILLER_68_1256 ();
 sg13g2_decap_8 FILLER_68_1263 ();
 sg13g2_decap_8 FILLER_68_1270 ();
 sg13g2_fill_1 FILLER_68_1277 ();
 sg13g2_fill_2 FILLER_68_1287 ();
 sg13g2_fill_1 FILLER_68_1289 ();
 sg13g2_fill_1 FILLER_68_1300 ();
 sg13g2_decap_4 FILLER_68_1316 ();
 sg13g2_fill_2 FILLER_68_1320 ();
 sg13g2_fill_1 FILLER_68_1327 ();
 sg13g2_fill_1 FILLER_68_1333 ();
 sg13g2_fill_1 FILLER_68_1344 ();
 sg13g2_fill_2 FILLER_68_1349 ();
 sg13g2_fill_1 FILLER_68_1351 ();
 sg13g2_fill_2 FILLER_68_1357 ();
 sg13g2_fill_1 FILLER_68_1359 ();
 sg13g2_fill_2 FILLER_68_1364 ();
 sg13g2_fill_1 FILLER_68_1366 ();
 sg13g2_fill_2 FILLER_68_1390 ();
 sg13g2_fill_1 FILLER_68_1392 ();
 sg13g2_fill_1 FILLER_68_1411 ();
 sg13g2_fill_2 FILLER_68_1416 ();
 sg13g2_decap_4 FILLER_68_1422 ();
 sg13g2_fill_2 FILLER_68_1426 ();
 sg13g2_fill_2 FILLER_68_1433 ();
 sg13g2_fill_2 FILLER_68_1476 ();
 sg13g2_decap_4 FILLER_68_1482 ();
 sg13g2_fill_1 FILLER_68_1486 ();
 sg13g2_fill_2 FILLER_68_1491 ();
 sg13g2_fill_1 FILLER_68_1493 ();
 sg13g2_fill_1 FILLER_68_1554 ();
 sg13g2_fill_2 FILLER_68_1559 ();
 sg13g2_fill_2 FILLER_68_1565 ();
 sg13g2_fill_2 FILLER_68_1593 ();
 sg13g2_fill_1 FILLER_68_1595 ();
 sg13g2_fill_1 FILLER_68_1626 ();
 sg13g2_fill_2 FILLER_68_1663 ();
 sg13g2_fill_1 FILLER_68_1665 ();
 sg13g2_fill_1 FILLER_68_1682 ();
 sg13g2_decap_8 FILLER_68_1693 ();
 sg13g2_decap_8 FILLER_68_1700 ();
 sg13g2_decap_8 FILLER_68_1707 ();
 sg13g2_decap_8 FILLER_68_1714 ();
 sg13g2_decap_8 FILLER_68_1721 ();
 sg13g2_decap_4 FILLER_68_1728 ();
 sg13g2_decap_8 FILLER_68_1750 ();
 sg13g2_decap_8 FILLER_68_1757 ();
 sg13g2_fill_2 FILLER_68_1764 ();
 sg13g2_fill_2 FILLER_68_1802 ();
 sg13g2_fill_1 FILLER_68_1804 ();
 sg13g2_fill_2 FILLER_68_1815 ();
 sg13g2_decap_4 FILLER_68_1821 ();
 sg13g2_decap_8 FILLER_68_1833 ();
 sg13g2_fill_1 FILLER_68_1902 ();
 sg13g2_fill_2 FILLER_68_1929 ();
 sg13g2_fill_1 FILLER_68_1967 ();
 sg13g2_decap_4 FILLER_68_1994 ();
 sg13g2_fill_1 FILLER_68_1998 ();
 sg13g2_decap_8 FILLER_68_2013 ();
 sg13g2_decap_8 FILLER_68_2020 ();
 sg13g2_decap_4 FILLER_68_2027 ();
 sg13g2_decap_8 FILLER_68_2044 ();
 sg13g2_fill_1 FILLER_68_2051 ();
 sg13g2_decap_8 FILLER_68_2060 ();
 sg13g2_decap_8 FILLER_68_2067 ();
 sg13g2_fill_2 FILLER_68_2086 ();
 sg13g2_fill_1 FILLER_68_2101 ();
 sg13g2_fill_2 FILLER_68_2113 ();
 sg13g2_fill_1 FILLER_68_2130 ();
 sg13g2_fill_1 FILLER_68_2154 ();
 sg13g2_fill_2 FILLER_68_2162 ();
 sg13g2_decap_4 FILLER_68_2179 ();
 sg13g2_decap_4 FILLER_68_2191 ();
 sg13g2_fill_2 FILLER_68_2221 ();
 sg13g2_decap_4 FILLER_68_2279 ();
 sg13g2_fill_1 FILLER_68_2283 ();
 sg13g2_decap_4 FILLER_68_2288 ();
 sg13g2_fill_2 FILLER_68_2292 ();
 sg13g2_fill_2 FILLER_68_2353 ();
 sg13g2_fill_2 FILLER_68_2459 ();
 sg13g2_decap_4 FILLER_68_2549 ();
 sg13g2_fill_1 FILLER_68_2553 ();
 sg13g2_decap_8 FILLER_68_2558 ();
 sg13g2_decap_4 FILLER_68_2565 ();
 sg13g2_fill_2 FILLER_68_2593 ();
 sg13g2_fill_1 FILLER_68_2595 ();
 sg13g2_decap_8 FILLER_68_2626 ();
 sg13g2_decap_8 FILLER_68_2633 ();
 sg13g2_decap_8 FILLER_68_2640 ();
 sg13g2_decap_8 FILLER_68_2647 ();
 sg13g2_decap_8 FILLER_68_2654 ();
 sg13g2_decap_8 FILLER_68_2661 ();
 sg13g2_fill_2 FILLER_68_2668 ();
 sg13g2_fill_1 FILLER_69_42 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_67 ();
 sg13g2_fill_2 FILLER_69_73 ();
 sg13g2_fill_1 FILLER_69_75 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_decap_4 FILLER_69_112 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_fill_1 FILLER_69_144 ();
 sg13g2_fill_1 FILLER_69_171 ();
 sg13g2_fill_1 FILLER_69_182 ();
 sg13g2_fill_1 FILLER_69_268 ();
 sg13g2_fill_1 FILLER_69_279 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_decap_8 FILLER_69_335 ();
 sg13g2_decap_8 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_351 ();
 sg13g2_fill_1 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_372 ();
 sg13g2_fill_1 FILLER_69_400 ();
 sg13g2_fill_2 FILLER_69_438 ();
 sg13g2_decap_8 FILLER_69_457 ();
 sg13g2_decap_4 FILLER_69_464 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_fill_2 FILLER_69_576 ();
 sg13g2_fill_2 FILLER_69_604 ();
 sg13g2_fill_1 FILLER_69_606 ();
 sg13g2_fill_1 FILLER_69_633 ();
 sg13g2_fill_1 FILLER_69_651 ();
 sg13g2_fill_2 FILLER_69_657 ();
 sg13g2_decap_4 FILLER_69_670 ();
 sg13g2_fill_2 FILLER_69_674 ();
 sg13g2_decap_4 FILLER_69_680 ();
 sg13g2_fill_1 FILLER_69_684 ();
 sg13g2_decap_4 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_735 ();
 sg13g2_decap_4 FILLER_69_754 ();
 sg13g2_decap_4 FILLER_69_774 ();
 sg13g2_fill_1 FILLER_69_778 ();
 sg13g2_decap_8 FILLER_69_783 ();
 sg13g2_fill_2 FILLER_69_790 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_797 ();
 sg13g2_decap_8 FILLER_69_804 ();
 sg13g2_decap_4 FILLER_69_811 ();
 sg13g2_fill_2 FILLER_69_818 ();
 sg13g2_fill_1 FILLER_69_820 ();
 sg13g2_fill_1 FILLER_69_835 ();
 sg13g2_fill_1 FILLER_69_840 ();
 sg13g2_fill_1 FILLER_69_845 ();
 sg13g2_fill_1 FILLER_69_850 ();
 sg13g2_fill_2 FILLER_69_864 ();
 sg13g2_fill_2 FILLER_69_871 ();
 sg13g2_fill_1 FILLER_69_873 ();
 sg13g2_fill_2 FILLER_69_884 ();
 sg13g2_fill_1 FILLER_69_886 ();
 sg13g2_decap_8 FILLER_69_896 ();
 sg13g2_fill_1 FILLER_69_903 ();
 sg13g2_fill_2 FILLER_69_908 ();
 sg13g2_decap_4 FILLER_69_915 ();
 sg13g2_fill_2 FILLER_69_919 ();
 sg13g2_decap_8 FILLER_69_948 ();
 sg13g2_fill_1 FILLER_69_955 ();
 sg13g2_decap_8 FILLER_69_961 ();
 sg13g2_fill_1 FILLER_69_968 ();
 sg13g2_decap_4 FILLER_69_973 ();
 sg13g2_fill_1 FILLER_69_1022 ();
 sg13g2_decap_4 FILLER_69_1028 ();
 sg13g2_fill_1 FILLER_69_1032 ();
 sg13g2_fill_2 FILLER_69_1041 ();
 sg13g2_fill_1 FILLER_69_1061 ();
 sg13g2_decap_4 FILLER_69_1066 ();
 sg13g2_fill_2 FILLER_69_1070 ();
 sg13g2_fill_1 FILLER_69_1094 ();
 sg13g2_fill_2 FILLER_69_1113 ();
 sg13g2_fill_2 FILLER_69_1130 ();
 sg13g2_decap_8 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1157 ();
 sg13g2_decap_4 FILLER_69_1164 ();
 sg13g2_fill_1 FILLER_69_1168 ();
 sg13g2_fill_1 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1183 ();
 sg13g2_decap_8 FILLER_69_1190 ();
 sg13g2_decap_4 FILLER_69_1197 ();
 sg13g2_fill_1 FILLER_69_1201 ();
 sg13g2_decap_8 FILLER_69_1232 ();
 sg13g2_decap_4 FILLER_69_1239 ();
 sg13g2_decap_4 FILLER_69_1248 ();
 sg13g2_fill_2 FILLER_69_1269 ();
 sg13g2_fill_1 FILLER_69_1271 ();
 sg13g2_decap_4 FILLER_69_1277 ();
 sg13g2_fill_1 FILLER_69_1298 ();
 sg13g2_fill_2 FILLER_69_1304 ();
 sg13g2_fill_1 FILLER_69_1306 ();
 sg13g2_fill_1 FILLER_69_1318 ();
 sg13g2_decap_4 FILLER_69_1324 ();
 sg13g2_fill_1 FILLER_69_1328 ();
 sg13g2_decap_8 FILLER_69_1333 ();
 sg13g2_decap_4 FILLER_69_1340 ();
 sg13g2_fill_1 FILLER_69_1344 ();
 sg13g2_fill_1 FILLER_69_1365 ();
 sg13g2_fill_1 FILLER_69_1374 ();
 sg13g2_fill_2 FILLER_69_1396 ();
 sg13g2_fill_1 FILLER_69_1415 ();
 sg13g2_decap_4 FILLER_69_1421 ();
 sg13g2_fill_1 FILLER_69_1425 ();
 sg13g2_fill_1 FILLER_69_1441 ();
 sg13g2_decap_4 FILLER_69_1462 ();
 sg13g2_fill_2 FILLER_69_1466 ();
 sg13g2_fill_2 FILLER_69_1507 ();
 sg13g2_fill_1 FILLER_69_1509 ();
 sg13g2_fill_1 FILLER_69_1540 ();
 sg13g2_decap_8 FILLER_69_1546 ();
 sg13g2_decap_4 FILLER_69_1553 ();
 sg13g2_fill_2 FILLER_69_1557 ();
 sg13g2_decap_4 FILLER_69_1567 ();
 sg13g2_fill_1 FILLER_69_1581 ();
 sg13g2_fill_1 FILLER_69_1586 ();
 sg13g2_fill_1 FILLER_69_1592 ();
 sg13g2_fill_1 FILLER_69_1598 ();
 sg13g2_fill_1 FILLER_69_1603 ();
 sg13g2_fill_1 FILLER_69_1608 ();
 sg13g2_fill_2 FILLER_69_1619 ();
 sg13g2_fill_1 FILLER_69_1621 ();
 sg13g2_fill_1 FILLER_69_1652 ();
 sg13g2_fill_1 FILLER_69_1683 ();
 sg13g2_fill_2 FILLER_69_1689 ();
 sg13g2_fill_1 FILLER_69_1691 ();
 sg13g2_fill_2 FILLER_69_1700 ();
 sg13g2_decap_8 FILLER_69_1720 ();
 sg13g2_fill_1 FILLER_69_1727 ();
 sg13g2_decap_8 FILLER_69_1733 ();
 sg13g2_fill_2 FILLER_69_1740 ();
 sg13g2_decap_4 FILLER_69_1753 ();
 sg13g2_fill_1 FILLER_69_1757 ();
 sg13g2_fill_1 FILLER_69_1763 ();
 sg13g2_fill_1 FILLER_69_1768 ();
 sg13g2_fill_2 FILLER_69_1775 ();
 sg13g2_fill_1 FILLER_69_1777 ();
 sg13g2_decap_8 FILLER_69_1805 ();
 sg13g2_decap_4 FILLER_69_1812 ();
 sg13g2_fill_2 FILLER_69_1816 ();
 sg13g2_decap_8 FILLER_69_1844 ();
 sg13g2_decap_4 FILLER_69_1851 ();
 sg13g2_fill_1 FILLER_69_1855 ();
 sg13g2_decap_4 FILLER_69_1868 ();
 sg13g2_decap_8 FILLER_69_1876 ();
 sg13g2_fill_2 FILLER_69_1883 ();
 sg13g2_fill_1 FILLER_69_1885 ();
 sg13g2_decap_4 FILLER_69_1896 ();
 sg13g2_fill_1 FILLER_69_1928 ();
 sg13g2_decap_8 FILLER_69_1959 ();
 sg13g2_fill_2 FILLER_69_1966 ();
 sg13g2_fill_1 FILLER_69_1968 ();
 sg13g2_fill_1 FILLER_69_1973 ();
 sg13g2_decap_8 FILLER_69_1978 ();
 sg13g2_decap_4 FILLER_69_1995 ();
 sg13g2_fill_2 FILLER_69_1999 ();
 sg13g2_decap_8 FILLER_69_2005 ();
 sg13g2_decap_8 FILLER_69_2012 ();
 sg13g2_decap_8 FILLER_69_2019 ();
 sg13g2_decap_8 FILLER_69_2026 ();
 sg13g2_decap_8 FILLER_69_2033 ();
 sg13g2_decap_8 FILLER_69_2040 ();
 sg13g2_fill_1 FILLER_69_2080 ();
 sg13g2_fill_2 FILLER_69_2086 ();
 sg13g2_decap_8 FILLER_69_2119 ();
 sg13g2_fill_2 FILLER_69_2135 ();
 sg13g2_fill_1 FILLER_69_2174 ();
 sg13g2_fill_2 FILLER_69_2194 ();
 sg13g2_fill_1 FILLER_69_2196 ();
 sg13g2_decap_8 FILLER_69_2233 ();
 sg13g2_fill_1 FILLER_69_2240 ();
 sg13g2_fill_1 FILLER_69_2251 ();
 sg13g2_fill_1 FILLER_69_2256 ();
 sg13g2_decap_8 FILLER_69_2261 ();
 sg13g2_decap_8 FILLER_69_2268 ();
 sg13g2_fill_2 FILLER_69_2275 ();
 sg13g2_decap_4 FILLER_69_2303 ();
 sg13g2_fill_1 FILLER_69_2313 ();
 sg13g2_decap_4 FILLER_69_2318 ();
 sg13g2_fill_1 FILLER_69_2322 ();
 sg13g2_fill_2 FILLER_69_2368 ();
 sg13g2_fill_2 FILLER_69_2416 ();
 sg13g2_fill_1 FILLER_69_2438 ();
 sg13g2_decap_4 FILLER_69_2528 ();
 sg13g2_fill_1 FILLER_69_2532 ();
 sg13g2_fill_1 FILLER_69_2537 ();
 sg13g2_decap_4 FILLER_69_2564 ();
 sg13g2_decap_8 FILLER_69_2572 ();
 sg13g2_fill_2 FILLER_69_2579 ();
 sg13g2_fill_1 FILLER_69_2581 ();
 sg13g2_fill_1 FILLER_69_2613 ();
 sg13g2_decap_8 FILLER_69_2627 ();
 sg13g2_decap_8 FILLER_69_2634 ();
 sg13g2_decap_8 FILLER_69_2641 ();
 sg13g2_decap_8 FILLER_69_2648 ();
 sg13g2_decap_8 FILLER_69_2655 ();
 sg13g2_decap_8 FILLER_69_2662 ();
 sg13g2_fill_1 FILLER_69_2669 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_1 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_63 ();
 sg13g2_decap_4 FILLER_70_69 ();
 sg13g2_fill_1 FILLER_70_73 ();
 sg13g2_fill_1 FILLER_70_130 ();
 sg13g2_fill_2 FILLER_70_139 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_1 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_fill_2 FILLER_70_280 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_2 FILLER_70_303 ();
 sg13g2_fill_1 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_310 ();
 sg13g2_decap_8 FILLER_70_317 ();
 sg13g2_decap_4 FILLER_70_324 ();
 sg13g2_fill_2 FILLER_70_328 ();
 sg13g2_decap_8 FILLER_70_334 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_fill_1 FILLER_70_395 ();
 sg13g2_fill_1 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_415 ();
 sg13g2_decap_4 FILLER_70_446 ();
 sg13g2_fill_1 FILLER_70_450 ();
 sg13g2_decap_4 FILLER_70_477 ();
 sg13g2_fill_2 FILLER_70_481 ();
 sg13g2_decap_8 FILLER_70_525 ();
 sg13g2_fill_2 FILLER_70_568 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_fill_1 FILLER_70_620 ();
 sg13g2_fill_1 FILLER_70_625 ();
 sg13g2_fill_1 FILLER_70_630 ();
 sg13g2_fill_1 FILLER_70_644 ();
 sg13g2_fill_2 FILLER_70_649 ();
 sg13g2_fill_1 FILLER_70_651 ();
 sg13g2_fill_2 FILLER_70_662 ();
 sg13g2_fill_1 FILLER_70_675 ();
 sg13g2_decap_8 FILLER_70_680 ();
 sg13g2_decap_8 FILLER_70_687 ();
 sg13g2_decap_8 FILLER_70_694 ();
 sg13g2_decap_4 FILLER_70_701 ();
 sg13g2_fill_2 FILLER_70_705 ();
 sg13g2_fill_1 FILLER_70_722 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_decap_4 FILLER_70_787 ();
 sg13g2_fill_2 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_797 ();
 sg13g2_decap_8 FILLER_70_804 ();
 sg13g2_fill_2 FILLER_70_811 ();
 sg13g2_fill_1 FILLER_70_813 ();
 sg13g2_fill_2 FILLER_70_827 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_fill_2 FILLER_70_851 ();
 sg13g2_fill_1 FILLER_70_853 ();
 sg13g2_fill_1 FILLER_70_859 ();
 sg13g2_fill_2 FILLER_70_892 ();
 sg13g2_fill_1 FILLER_70_894 ();
 sg13g2_fill_1 FILLER_70_905 ();
 sg13g2_fill_1 FILLER_70_910 ();
 sg13g2_fill_1 FILLER_70_915 ();
 sg13g2_fill_1 FILLER_70_922 ();
 sg13g2_fill_1 FILLER_70_929 ();
 sg13g2_fill_2 FILLER_70_935 ();
 sg13g2_fill_1 FILLER_70_937 ();
 sg13g2_fill_2 FILLER_70_986 ();
 sg13g2_fill_1 FILLER_70_993 ();
 sg13g2_fill_1 FILLER_70_998 ();
 sg13g2_fill_1 FILLER_70_1003 ();
 sg13g2_decap_4 FILLER_70_1009 ();
 sg13g2_fill_1 FILLER_70_1013 ();
 sg13g2_decap_4 FILLER_70_1018 ();
 sg13g2_fill_2 FILLER_70_1022 ();
 sg13g2_fill_1 FILLER_70_1028 ();
 sg13g2_decap_4 FILLER_70_1038 ();
 sg13g2_fill_1 FILLER_70_1042 ();
 sg13g2_decap_8 FILLER_70_1058 ();
 sg13g2_fill_2 FILLER_70_1065 ();
 sg13g2_decap_4 FILLER_70_1072 ();
 sg13g2_fill_1 FILLER_70_1076 ();
 sg13g2_fill_1 FILLER_70_1086 ();
 sg13g2_fill_2 FILLER_70_1108 ();
 sg13g2_fill_1 FILLER_70_1110 ();
 sg13g2_fill_2 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1131 ();
 sg13g2_fill_1 FILLER_70_1138 ();
 sg13g2_decap_8 FILLER_70_1155 ();
 sg13g2_decap_8 FILLER_70_1162 ();
 sg13g2_fill_2 FILLER_70_1169 ();
 sg13g2_fill_1 FILLER_70_1171 ();
 sg13g2_fill_2 FILLER_70_1205 ();
 sg13g2_fill_1 FILLER_70_1233 ();
 sg13g2_fill_1 FILLER_70_1239 ();
 sg13g2_fill_1 FILLER_70_1249 ();
 sg13g2_fill_1 FILLER_70_1275 ();
 sg13g2_fill_2 FILLER_70_1285 ();
 sg13g2_fill_1 FILLER_70_1287 ();
 sg13g2_decap_4 FILLER_70_1297 ();
 sg13g2_fill_1 FILLER_70_1305 ();
 sg13g2_fill_1 FILLER_70_1314 ();
 sg13g2_fill_2 FILLER_70_1328 ();
 sg13g2_fill_1 FILLER_70_1340 ();
 sg13g2_fill_1 FILLER_70_1347 ();
 sg13g2_fill_2 FILLER_70_1353 ();
 sg13g2_fill_1 FILLER_70_1377 ();
 sg13g2_fill_2 FILLER_70_1407 ();
 sg13g2_fill_2 FILLER_70_1417 ();
 sg13g2_fill_1 FILLER_70_1419 ();
 sg13g2_decap_8 FILLER_70_1427 ();
 sg13g2_decap_4 FILLER_70_1434 ();
 sg13g2_fill_1 FILLER_70_1438 ();
 sg13g2_decap_8 FILLER_70_1444 ();
 sg13g2_decap_8 FILLER_70_1451 ();
 sg13g2_decap_4 FILLER_70_1458 ();
 sg13g2_fill_2 FILLER_70_1472 ();
 sg13g2_fill_1 FILLER_70_1474 ();
 sg13g2_fill_2 FILLER_70_1522 ();
 sg13g2_fill_1 FILLER_70_1524 ();
 sg13g2_decap_8 FILLER_70_1555 ();
 sg13g2_fill_1 FILLER_70_1562 ();
 sg13g2_fill_1 FILLER_70_1597 ();
 sg13g2_decap_4 FILLER_70_1607 ();
 sg13g2_decap_4 FILLER_70_1625 ();
 sg13g2_fill_2 FILLER_70_1629 ();
 sg13g2_fill_2 FILLER_70_1635 ();
 sg13g2_fill_2 FILLER_70_1651 ();
 sg13g2_fill_1 FILLER_70_1653 ();
 sg13g2_decap_8 FILLER_70_1668 ();
 sg13g2_decap_8 FILLER_70_1675 ();
 sg13g2_decap_8 FILLER_70_1682 ();
 sg13g2_decap_8 FILLER_70_1715 ();
 sg13g2_fill_2 FILLER_70_1736 ();
 sg13g2_decap_8 FILLER_70_1748 ();
 sg13g2_fill_2 FILLER_70_1755 ();
 sg13g2_fill_1 FILLER_70_1757 ();
 sg13g2_decap_8 FILLER_70_1763 ();
 sg13g2_decap_8 FILLER_70_1770 ();
 sg13g2_decap_8 FILLER_70_1777 ();
 sg13g2_decap_8 FILLER_70_1784 ();
 sg13g2_fill_2 FILLER_70_1791 ();
 sg13g2_fill_1 FILLER_70_1793 ();
 sg13g2_decap_8 FILLER_70_1798 ();
 sg13g2_decap_8 FILLER_70_1805 ();
 sg13g2_decap_8 FILLER_70_1812 ();
 sg13g2_decap_4 FILLER_70_1819 ();
 sg13g2_fill_2 FILLER_70_1823 ();
 sg13g2_decap_8 FILLER_70_1835 ();
 sg13g2_decap_4 FILLER_70_1842 ();
 sg13g2_fill_1 FILLER_70_1846 ();
 sg13g2_decap_8 FILLER_70_1865 ();
 sg13g2_fill_2 FILLER_70_1882 ();
 sg13g2_fill_1 FILLER_70_1884 ();
 sg13g2_fill_2 FILLER_70_1895 ();
 sg13g2_fill_2 FILLER_70_1923 ();
 sg13g2_fill_1 FILLER_70_1925 ();
 sg13g2_decap_8 FILLER_70_1956 ();
 sg13g2_fill_1 FILLER_70_1963 ();
 sg13g2_decap_8 FILLER_70_1968 ();
 sg13g2_decap_8 FILLER_70_1975 ();
 sg13g2_fill_2 FILLER_70_1982 ();
 sg13g2_fill_1 FILLER_70_1984 ();
 sg13g2_decap_8 FILLER_70_2025 ();
 sg13g2_decap_8 FILLER_70_2032 ();
 sg13g2_fill_2 FILLER_70_2039 ();
 sg13g2_fill_1 FILLER_70_2067 ();
 sg13g2_fill_1 FILLER_70_2073 ();
 sg13g2_fill_1 FILLER_70_2155 ();
 sg13g2_fill_1 FILLER_70_2188 ();
 sg13g2_fill_1 FILLER_70_2211 ();
 sg13g2_decap_8 FILLER_70_2233 ();
 sg13g2_decap_8 FILLER_70_2240 ();
 sg13g2_decap_8 FILLER_70_2247 ();
 sg13g2_decap_8 FILLER_70_2254 ();
 sg13g2_fill_1 FILLER_70_2318 ();
 sg13g2_decap_4 FILLER_70_2333 ();
 sg13g2_fill_2 FILLER_70_2342 ();
 sg13g2_fill_1 FILLER_70_2380 ();
 sg13g2_fill_2 FILLER_70_2411 ();
 sg13g2_fill_2 FILLER_70_2416 ();
 sg13g2_fill_1 FILLER_70_2470 ();
 sg13g2_fill_1 FILLER_70_2481 ();
 sg13g2_decap_4 FILLER_70_2518 ();
 sg13g2_fill_2 FILLER_70_2583 ();
 sg13g2_decap_8 FILLER_70_2606 ();
 sg13g2_decap_8 FILLER_70_2613 ();
 sg13g2_decap_8 FILLER_70_2620 ();
 sg13g2_decap_8 FILLER_70_2627 ();
 sg13g2_decap_8 FILLER_70_2634 ();
 sg13g2_decap_8 FILLER_70_2641 ();
 sg13g2_decap_8 FILLER_70_2648 ();
 sg13g2_decap_8 FILLER_70_2655 ();
 sg13g2_decap_8 FILLER_70_2662 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_1 FILLER_71_16 ();
 sg13g2_fill_2 FILLER_71_23 ();
 sg13g2_fill_1 FILLER_71_30 ();
 sg13g2_fill_2 FILLER_71_46 ();
 sg13g2_fill_1 FILLER_71_52 ();
 sg13g2_decap_8 FILLER_71_59 ();
 sg13g2_decap_8 FILLER_71_66 ();
 sg13g2_decap_8 FILLER_71_73 ();
 sg13g2_fill_2 FILLER_71_80 ();
 sg13g2_fill_2 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_fill_2 FILLER_71_99 ();
 sg13g2_fill_1 FILLER_71_101 ();
 sg13g2_fill_1 FILLER_71_107 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_decap_4 FILLER_71_120 ();
 sg13g2_fill_2 FILLER_71_124 ();
 sg13g2_fill_2 FILLER_71_135 ();
 sg13g2_fill_1 FILLER_71_141 ();
 sg13g2_decap_8 FILLER_71_172 ();
 sg13g2_fill_2 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_181 ();
 sg13g2_fill_2 FILLER_71_191 ();
 sg13g2_fill_2 FILLER_71_198 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_220 ();
 sg13g2_fill_2 FILLER_71_240 ();
 sg13g2_fill_1 FILLER_71_284 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_fill_2 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_405 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_fill_1 FILLER_71_456 ();
 sg13g2_fill_1 FILLER_71_466 ();
 sg13g2_fill_2 FILLER_71_497 ();
 sg13g2_fill_1 FILLER_71_499 ();
 sg13g2_fill_2 FILLER_71_518 ();
 sg13g2_fill_1 FILLER_71_520 ();
 sg13g2_fill_2 FILLER_71_536 ();
 sg13g2_fill_1 FILLER_71_538 ();
 sg13g2_fill_2 FILLER_71_544 ();
 sg13g2_fill_2 FILLER_71_579 ();
 sg13g2_decap_4 FILLER_71_589 ();
 sg13g2_decap_4 FILLER_71_602 ();
 sg13g2_fill_1 FILLER_71_606 ();
 sg13g2_fill_2 FILLER_71_611 ();
 sg13g2_decap_4 FILLER_71_622 ();
 sg13g2_fill_2 FILLER_71_626 ();
 sg13g2_fill_1 FILLER_71_632 ();
 sg13g2_fill_2 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_702 ();
 sg13g2_fill_2 FILLER_71_707 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_fill_1 FILLER_71_724 ();
 sg13g2_fill_2 FILLER_71_736 ();
 sg13g2_fill_1 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_decap_8 FILLER_71_808 ();
 sg13g2_fill_1 FILLER_71_815 ();
 sg13g2_decap_8 FILLER_71_821 ();
 sg13g2_fill_1 FILLER_71_828 ();
 sg13g2_fill_2 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_859 ();
 sg13g2_decap_4 FILLER_71_866 ();
 sg13g2_fill_1 FILLER_71_870 ();
 sg13g2_fill_1 FILLER_71_900 ();
 sg13g2_fill_1 FILLER_71_906 ();
 sg13g2_fill_1 FILLER_71_928 ();
 sg13g2_fill_1 FILLER_71_933 ();
 sg13g2_fill_1 FILLER_71_948 ();
 sg13g2_fill_1 FILLER_71_964 ();
 sg13g2_fill_1 FILLER_71_972 ();
 sg13g2_fill_2 FILLER_71_988 ();
 sg13g2_fill_1 FILLER_71_995 ();
 sg13g2_fill_1 FILLER_71_1019 ();
 sg13g2_fill_2 FILLER_71_1029 ();
 sg13g2_decap_4 FILLER_71_1036 ();
 sg13g2_fill_2 FILLER_71_1040 ();
 sg13g2_fill_1 FILLER_71_1069 ();
 sg13g2_fill_2 FILLER_71_1074 ();
 sg13g2_fill_1 FILLER_71_1076 ();
 sg13g2_decap_8 FILLER_71_1083 ();
 sg13g2_decap_4 FILLER_71_1090 ();
 sg13g2_fill_2 FILLER_71_1098 ();
 sg13g2_fill_1 FILLER_71_1100 ();
 sg13g2_fill_1 FILLER_71_1108 ();
 sg13g2_decap_8 FILLER_71_1119 ();
 sg13g2_decap_4 FILLER_71_1126 ();
 sg13g2_fill_1 FILLER_71_1130 ();
 sg13g2_decap_4 FILLER_71_1139 ();
 sg13g2_fill_2 FILLER_71_1165 ();
 sg13g2_fill_2 FILLER_71_1172 ();
 sg13g2_fill_1 FILLER_71_1181 ();
 sg13g2_fill_2 FILLER_71_1187 ();
 sg13g2_fill_1 FILLER_71_1215 ();
 sg13g2_fill_2 FILLER_71_1220 ();
 sg13g2_fill_2 FILLER_71_1275 ();
 sg13g2_fill_1 FILLER_71_1317 ();
 sg13g2_fill_1 FILLER_71_1323 ();
 sg13g2_fill_1 FILLER_71_1361 ();
 sg13g2_fill_1 FILLER_71_1375 ();
 sg13g2_fill_1 FILLER_71_1402 ();
 sg13g2_decap_4 FILLER_71_1420 ();
 sg13g2_fill_1 FILLER_71_1429 ();
 sg13g2_decap_4 FILLER_71_1434 ();
 sg13g2_fill_1 FILLER_71_1438 ();
 sg13g2_decap_4 FILLER_71_1465 ();
 sg13g2_decap_4 FILLER_71_1495 ();
 sg13g2_fill_2 FILLER_71_1499 ();
 sg13g2_fill_2 FILLER_71_1505 ();
 sg13g2_decap_8 FILLER_71_1545 ();
 sg13g2_fill_2 FILLER_71_1552 ();
 sg13g2_decap_8 FILLER_71_1577 ();
 sg13g2_fill_2 FILLER_71_1584 ();
 sg13g2_fill_1 FILLER_71_1586 ();
 sg13g2_fill_2 FILLER_71_1597 ();
 sg13g2_fill_2 FILLER_71_1604 ();
 sg13g2_decap_8 FILLER_71_1610 ();
 sg13g2_decap_4 FILLER_71_1617 ();
 sg13g2_fill_2 FILLER_71_1639 ();
 sg13g2_fill_1 FILLER_71_1641 ();
 sg13g2_decap_8 FILLER_71_1651 ();
 sg13g2_fill_1 FILLER_71_1658 ();
 sg13g2_decap_4 FILLER_71_1663 ();
 sg13g2_fill_1 FILLER_71_1667 ();
 sg13g2_decap_8 FILLER_71_1678 ();
 sg13g2_decap_4 FILLER_71_1685 ();
 sg13g2_fill_2 FILLER_71_1689 ();
 sg13g2_decap_8 FILLER_71_1777 ();
 sg13g2_fill_2 FILLER_71_1822 ();
 sg13g2_fill_1 FILLER_71_1824 ();
 sg13g2_decap_4 FILLER_71_1865 ();
 sg13g2_fill_1 FILLER_71_1869 ();
 sg13g2_fill_1 FILLER_71_1880 ();
 sg13g2_fill_1 FILLER_71_1907 ();
 sg13g2_decap_8 FILLER_71_1916 ();
 sg13g2_fill_1 FILLER_71_1923 ();
 sg13g2_fill_1 FILLER_71_1940 ();
 sg13g2_fill_2 FILLER_71_1949 ();
 sg13g2_fill_1 FILLER_71_1951 ();
 sg13g2_decap_8 FILLER_71_1983 ();
 sg13g2_decap_8 FILLER_71_1990 ();
 sg13g2_fill_2 FILLER_71_1997 ();
 sg13g2_fill_1 FILLER_71_1999 ();
 sg13g2_decap_8 FILLER_71_2036 ();
 sg13g2_fill_1 FILLER_71_2043 ();
 sg13g2_fill_2 FILLER_71_2060 ();
 sg13g2_fill_1 FILLER_71_2062 ();
 sg13g2_fill_1 FILLER_71_2069 ();
 sg13g2_fill_1 FILLER_71_2075 ();
 sg13g2_decap_4 FILLER_71_2085 ();
 sg13g2_fill_2 FILLER_71_2089 ();
 sg13g2_decap_8 FILLER_71_2127 ();
 sg13g2_decap_4 FILLER_71_2143 ();
 sg13g2_fill_1 FILLER_71_2147 ();
 sg13g2_fill_1 FILLER_71_2156 ();
 sg13g2_fill_2 FILLER_71_2185 ();
 sg13g2_fill_2 FILLER_71_2224 ();
 sg13g2_fill_1 FILLER_71_2226 ();
 sg13g2_decap_4 FILLER_71_2248 ();
 sg13g2_decap_8 FILLER_71_2265 ();
 sg13g2_decap_4 FILLER_71_2272 ();
 sg13g2_decap_4 FILLER_71_2316 ();
 sg13g2_fill_1 FILLER_71_2320 ();
 sg13g2_fill_1 FILLER_71_2414 ();
 sg13g2_fill_2 FILLER_71_2508 ();
 sg13g2_fill_1 FILLER_71_2510 ();
 sg13g2_fill_2 FILLER_71_2534 ();
 sg13g2_fill_1 FILLER_71_2536 ();
 sg13g2_decap_4 FILLER_71_2563 ();
 sg13g2_fill_1 FILLER_71_2567 ();
 sg13g2_decap_8 FILLER_71_2608 ();
 sg13g2_decap_8 FILLER_71_2615 ();
 sg13g2_decap_8 FILLER_71_2622 ();
 sg13g2_decap_8 FILLER_71_2629 ();
 sg13g2_decap_8 FILLER_71_2636 ();
 sg13g2_decap_8 FILLER_71_2643 ();
 sg13g2_decap_8 FILLER_71_2650 ();
 sg13g2_decap_8 FILLER_71_2657 ();
 sg13g2_decap_4 FILLER_71_2664 ();
 sg13g2_fill_2 FILLER_71_2668 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_47 ();
 sg13g2_fill_1 FILLER_72_52 ();
 sg13g2_fill_2 FILLER_72_57 ();
 sg13g2_fill_2 FILLER_72_106 ();
 sg13g2_fill_1 FILLER_72_108 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_decap_8 FILLER_72_156 ();
 sg13g2_decap_4 FILLER_72_163 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_decap_8 FILLER_72_172 ();
 sg13g2_decap_8 FILLER_72_179 ();
 sg13g2_decap_8 FILLER_72_186 ();
 sg13g2_fill_2 FILLER_72_201 ();
 sg13g2_decap_4 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_decap_4 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_234 ();
 sg13g2_decap_8 FILLER_72_242 ();
 sg13g2_fill_1 FILLER_72_249 ();
 sg13g2_decap_8 FILLER_72_256 ();
 sg13g2_decap_4 FILLER_72_263 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_fill_1 FILLER_72_281 ();
 sg13g2_fill_1 FILLER_72_298 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_decap_8 FILLER_72_310 ();
 sg13g2_fill_2 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_fill_1 FILLER_72_362 ();
 sg13g2_decap_8 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_decap_8 FILLER_72_433 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_fill_2 FILLER_72_447 ();
 sg13g2_fill_1 FILLER_72_449 ();
 sg13g2_decap_8 FILLER_72_459 ();
 sg13g2_fill_2 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_468 ();
 sg13g2_fill_1 FILLER_72_479 ();
 sg13g2_fill_1 FILLER_72_501 ();
 sg13g2_fill_1 FILLER_72_554 ();
 sg13g2_decap_4 FILLER_72_575 ();
 sg13g2_fill_2 FILLER_72_579 ();
 sg13g2_decap_8 FILLER_72_585 ();
 sg13g2_decap_8 FILLER_72_592 ();
 sg13g2_decap_4 FILLER_72_599 ();
 sg13g2_fill_1 FILLER_72_603 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_decap_4 FILLER_72_682 ();
 sg13g2_fill_2 FILLER_72_751 ();
 sg13g2_fill_1 FILLER_72_762 ();
 sg13g2_fill_1 FILLER_72_766 ();
 sg13g2_fill_2 FILLER_72_801 ();
 sg13g2_decap_4 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_812 ();
 sg13g2_fill_1 FILLER_72_821 ();
 sg13g2_fill_1 FILLER_72_830 ();
 sg13g2_fill_1 FILLER_72_835 ();
 sg13g2_fill_2 FILLER_72_849 ();
 sg13g2_fill_1 FILLER_72_868 ();
 sg13g2_fill_2 FILLER_72_893 ();
 sg13g2_fill_1 FILLER_72_908 ();
 sg13g2_fill_1 FILLER_72_929 ();
 sg13g2_fill_1 FILLER_72_942 ();
 sg13g2_fill_2 FILLER_72_947 ();
 sg13g2_fill_1 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_960 ();
 sg13g2_fill_1 FILLER_72_979 ();
 sg13g2_fill_1 FILLER_72_985 ();
 sg13g2_fill_1 FILLER_72_992 ();
 sg13g2_fill_1 FILLER_72_998 ();
 sg13g2_fill_1 FILLER_72_1023 ();
 sg13g2_decap_8 FILLER_72_1029 ();
 sg13g2_fill_1 FILLER_72_1036 ();
 sg13g2_fill_2 FILLER_72_1051 ();
 sg13g2_fill_2 FILLER_72_1077 ();
 sg13g2_fill_2 FILLER_72_1103 ();
 sg13g2_fill_1 FILLER_72_1105 ();
 sg13g2_decap_8 FILLER_72_1110 ();
 sg13g2_decap_8 FILLER_72_1117 ();
 sg13g2_decap_8 FILLER_72_1124 ();
 sg13g2_decap_8 FILLER_72_1131 ();
 sg13g2_decap_8 FILLER_72_1138 ();
 sg13g2_fill_1 FILLER_72_1145 ();
 sg13g2_fill_1 FILLER_72_1205 ();
 sg13g2_fill_1 FILLER_72_1216 ();
 sg13g2_decap_8 FILLER_72_1227 ();
 sg13g2_fill_2 FILLER_72_1234 ();
 sg13g2_fill_1 FILLER_72_1302 ();
 sg13g2_fill_2 FILLER_72_1345 ();
 sg13g2_fill_1 FILLER_72_1347 ();
 sg13g2_fill_1 FILLER_72_1356 ();
 sg13g2_fill_1 FILLER_72_1363 ();
 sg13g2_fill_1 FILLER_72_1388 ();
 sg13g2_fill_1 FILLER_72_1394 ();
 sg13g2_fill_1 FILLER_72_1400 ();
 sg13g2_fill_2 FILLER_72_1406 ();
 sg13g2_fill_2 FILLER_72_1429 ();
 sg13g2_decap_4 FILLER_72_1435 ();
 sg13g2_fill_1 FILLER_72_1439 ();
 sg13g2_fill_2 FILLER_72_1480 ();
 sg13g2_fill_1 FILLER_72_1482 ();
 sg13g2_decap_8 FILLER_72_1487 ();
 sg13g2_fill_2 FILLER_72_1494 ();
 sg13g2_decap_8 FILLER_72_1500 ();
 sg13g2_decap_8 FILLER_72_1521 ();
 sg13g2_decap_8 FILLER_72_1528 ();
 sg13g2_fill_1 FILLER_72_1565 ();
 sg13g2_fill_2 FILLER_72_1579 ();
 sg13g2_fill_1 FILLER_72_1581 ();
 sg13g2_decap_4 FILLER_72_1646 ();
 sg13g2_fill_2 FILLER_72_1650 ();
 sg13g2_decap_4 FILLER_72_1678 ();
 sg13g2_fill_2 FILLER_72_1692 ();
 sg13g2_fill_1 FILLER_72_1694 ();
 sg13g2_decap_8 FILLER_72_1710 ();
 sg13g2_fill_2 FILLER_72_1757 ();
 sg13g2_fill_1 FILLER_72_1759 ();
 sg13g2_decap_4 FILLER_72_1800 ();
 sg13g2_decap_4 FILLER_72_1812 ();
 sg13g2_fill_2 FILLER_72_1829 ();
 sg13g2_fill_2 FILLER_72_1907 ();
 sg13g2_decap_4 FILLER_72_1915 ();
 sg13g2_fill_2 FILLER_72_1936 ();
 sg13g2_fill_1 FILLER_72_1938 ();
 sg13g2_fill_2 FILLER_72_1965 ();
 sg13g2_decap_4 FILLER_72_2003 ();
 sg13g2_decap_8 FILLER_72_2033 ();
 sg13g2_fill_2 FILLER_72_2040 ();
 sg13g2_decap_8 FILLER_72_2083 ();
 sg13g2_fill_2 FILLER_72_2094 ();
 sg13g2_fill_1 FILLER_72_2096 ();
 sg13g2_decap_4 FILLER_72_2121 ();
 sg13g2_fill_2 FILLER_72_2125 ();
 sg13g2_fill_2 FILLER_72_2136 ();
 sg13g2_fill_1 FILLER_72_2138 ();
 sg13g2_decap_4 FILLER_72_2148 ();
 sg13g2_fill_2 FILLER_72_2152 ();
 sg13g2_fill_1 FILLER_72_2231 ();
 sg13g2_decap_4 FILLER_72_2240 ();
 sg13g2_decap_8 FILLER_72_2258 ();
 sg13g2_decap_4 FILLER_72_2265 ();
 sg13g2_decap_8 FILLER_72_2279 ();
 sg13g2_fill_2 FILLER_72_2290 ();
 sg13g2_decap_4 FILLER_72_2302 ();
 sg13g2_fill_2 FILLER_72_2306 ();
 sg13g2_decap_8 FILLER_72_2334 ();
 sg13g2_decap_8 FILLER_72_2341 ();
 sg13g2_fill_1 FILLER_72_2348 ();
 sg13g2_fill_2 FILLER_72_2363 ();
 sg13g2_fill_2 FILLER_72_2520 ();
 sg13g2_fill_1 FILLER_72_2522 ();
 sg13g2_decap_8 FILLER_72_2553 ();
 sg13g2_fill_2 FILLER_72_2560 ();
 sg13g2_decap_8 FILLER_72_2598 ();
 sg13g2_decap_8 FILLER_72_2605 ();
 sg13g2_decap_8 FILLER_72_2612 ();
 sg13g2_decap_8 FILLER_72_2619 ();
 sg13g2_decap_8 FILLER_72_2626 ();
 sg13g2_decap_8 FILLER_72_2633 ();
 sg13g2_decap_8 FILLER_72_2640 ();
 sg13g2_decap_8 FILLER_72_2647 ();
 sg13g2_decap_8 FILLER_72_2654 ();
 sg13g2_decap_8 FILLER_72_2661 ();
 sg13g2_fill_2 FILLER_72_2668 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_69 ();
 sg13g2_decap_4 FILLER_73_76 ();
 sg13g2_decap_8 FILLER_73_90 ();
 sg13g2_decap_8 FILLER_73_97 ();
 sg13g2_decap_4 FILLER_73_104 ();
 sg13g2_decap_8 FILLER_73_172 ();
 sg13g2_decap_4 FILLER_73_179 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_188 ();
 sg13g2_fill_2 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_220 ();
 sg13g2_fill_1 FILLER_73_249 ();
 sg13g2_fill_2 FILLER_73_263 ();
 sg13g2_decap_4 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_299 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_fill_2 FILLER_73_388 ();
 sg13g2_fill_2 FILLER_73_395 ();
 sg13g2_decap_4 FILLER_73_401 ();
 sg13g2_fill_2 FILLER_73_409 ();
 sg13g2_fill_1 FILLER_73_411 ();
 sg13g2_decap_4 FILLER_73_420 ();
 sg13g2_fill_2 FILLER_73_424 ();
 sg13g2_fill_2 FILLER_73_430 ();
 sg13g2_fill_1 FILLER_73_432 ();
 sg13g2_fill_1 FILLER_73_438 ();
 sg13g2_fill_2 FILLER_73_444 ();
 sg13g2_fill_1 FILLER_73_450 ();
 sg13g2_fill_2 FILLER_73_464 ();
 sg13g2_decap_8 FILLER_73_471 ();
 sg13g2_fill_1 FILLER_73_496 ();
 sg13g2_decap_8 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_527 ();
 sg13g2_fill_2 FILLER_73_534 ();
 sg13g2_decap_8 FILLER_73_540 ();
 sg13g2_decap_8 FILLER_73_547 ();
 sg13g2_decap_8 FILLER_73_554 ();
 sg13g2_decap_4 FILLER_73_561 ();
 sg13g2_fill_2 FILLER_73_609 ();
 sg13g2_fill_1 FILLER_73_659 ();
 sg13g2_decap_4 FILLER_73_683 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_fill_2 FILLER_73_703 ();
 sg13g2_fill_1 FILLER_73_705 ();
 sg13g2_fill_1 FILLER_73_739 ();
 sg13g2_fill_2 FILLER_73_753 ();
 sg13g2_fill_1 FILLER_73_762 ();
 sg13g2_fill_1 FILLER_73_771 ();
 sg13g2_fill_2 FILLER_73_777 ();
 sg13g2_fill_2 FILLER_73_783 ();
 sg13g2_fill_1 FILLER_73_785 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_4 FILLER_73_797 ();
 sg13g2_fill_2 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_806 ();
 sg13g2_fill_2 FILLER_73_813 ();
 sg13g2_fill_2 FILLER_73_826 ();
 sg13g2_fill_1 FILLER_73_828 ();
 sg13g2_fill_1 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_864 ();
 sg13g2_fill_1 FILLER_73_873 ();
 sg13g2_fill_2 FILLER_73_882 ();
 sg13g2_fill_2 FILLER_73_902 ();
 sg13g2_fill_1 FILLER_73_904 ();
 sg13g2_fill_1 FILLER_73_919 ();
 sg13g2_fill_2 FILLER_73_931 ();
 sg13g2_fill_2 FILLER_73_937 ();
 sg13g2_fill_2 FILLER_73_943 ();
 sg13g2_fill_1 FILLER_73_950 ();
 sg13g2_fill_1 FILLER_73_956 ();
 sg13g2_fill_1 FILLER_73_963 ();
 sg13g2_decap_8 FILLER_73_973 ();
 sg13g2_fill_2 FILLER_73_1008 ();
 sg13g2_fill_1 FILLER_73_1019 ();
 sg13g2_fill_1 FILLER_73_1025 ();
 sg13g2_fill_1 FILLER_73_1031 ();
 sg13g2_fill_1 FILLER_73_1037 ();
 sg13g2_fill_1 FILLER_73_1044 ();
 sg13g2_fill_1 FILLER_73_1053 ();
 sg13g2_fill_1 FILLER_73_1068 ();
 sg13g2_fill_1 FILLER_73_1073 ();
 sg13g2_fill_1 FILLER_73_1078 ();
 sg13g2_fill_1 FILLER_73_1083 ();
 sg13g2_fill_1 FILLER_73_1088 ();
 sg13g2_fill_1 FILLER_73_1100 ();
 sg13g2_decap_8 FILLER_73_1106 ();
 sg13g2_decap_4 FILLER_73_1113 ();
 sg13g2_decap_8 FILLER_73_1124 ();
 sg13g2_decap_8 FILLER_73_1131 ();
 sg13g2_decap_8 FILLER_73_1138 ();
 sg13g2_decap_8 FILLER_73_1145 ();
 sg13g2_fill_2 FILLER_73_1152 ();
 sg13g2_fill_2 FILLER_73_1184 ();
 sg13g2_fill_1 FILLER_73_1214 ();
 sg13g2_decap_4 FILLER_73_1219 ();
 sg13g2_fill_2 FILLER_73_1232 ();
 sg13g2_fill_1 FILLER_73_1246 ();
 sg13g2_decap_4 FILLER_73_1274 ();
 sg13g2_fill_2 FILLER_73_1278 ();
 sg13g2_fill_2 FILLER_73_1285 ();
 sg13g2_fill_2 FILLER_73_1307 ();
 sg13g2_fill_1 FILLER_73_1318 ();
 sg13g2_fill_1 FILLER_73_1325 ();
 sg13g2_fill_2 FILLER_73_1361 ();
 sg13g2_fill_1 FILLER_73_1363 ();
 sg13g2_fill_1 FILLER_73_1399 ();
 sg13g2_decap_4 FILLER_73_1431 ();
 sg13g2_fill_1 FILLER_73_1435 ();
 sg13g2_fill_1 FILLER_73_1440 ();
 sg13g2_decap_8 FILLER_73_1452 ();
 sg13g2_fill_2 FILLER_73_1459 ();
 sg13g2_decap_8 FILLER_73_1475 ();
 sg13g2_decap_4 FILLER_73_1482 ();
 sg13g2_decap_8 FILLER_73_1515 ();
 sg13g2_decap_4 FILLER_73_1522 ();
 sg13g2_fill_1 FILLER_73_1526 ();
 sg13g2_decap_4 FILLER_73_1531 ();
 sg13g2_fill_1 FILLER_73_1535 ();
 sg13g2_fill_2 FILLER_73_1541 ();
 sg13g2_decap_8 FILLER_73_1552 ();
 sg13g2_fill_1 FILLER_73_1559 ();
 sg13g2_fill_1 FILLER_73_1599 ();
 sg13g2_decap_8 FILLER_73_1604 ();
 sg13g2_fill_2 FILLER_73_1611 ();
 sg13g2_fill_2 FILLER_73_1649 ();
 sg13g2_fill_1 FILLER_73_1651 ();
 sg13g2_decap_8 FILLER_73_1714 ();
 sg13g2_decap_8 FILLER_73_1721 ();
 sg13g2_fill_2 FILLER_73_1728 ();
 sg13g2_fill_1 FILLER_73_1753 ();
 sg13g2_decap_4 FILLER_73_1774 ();
 sg13g2_fill_1 FILLER_73_1778 ();
 sg13g2_decap_4 FILLER_73_1783 ();
 sg13g2_fill_1 FILLER_73_1787 ();
 sg13g2_decap_4 FILLER_73_1876 ();
 sg13g2_fill_1 FILLER_73_1880 ();
 sg13g2_decap_8 FILLER_73_1903 ();
 sg13g2_fill_2 FILLER_73_1910 ();
 sg13g2_fill_1 FILLER_73_1912 ();
 sg13g2_fill_1 FILLER_73_1945 ();
 sg13g2_fill_1 FILLER_73_1952 ();
 sg13g2_fill_1 FILLER_73_1979 ();
 sg13g2_fill_1 FILLER_73_1990 ();
 sg13g2_fill_2 FILLER_73_2037 ();
 sg13g2_fill_1 FILLER_73_2075 ();
 sg13g2_fill_2 FILLER_73_2108 ();
 sg13g2_fill_2 FILLER_73_2118 ();
 sg13g2_fill_1 FILLER_73_2120 ();
 sg13g2_fill_1 FILLER_73_2135 ();
 sg13g2_fill_2 FILLER_73_2152 ();
 sg13g2_fill_2 FILLER_73_2173 ();
 sg13g2_fill_2 FILLER_73_2180 ();
 sg13g2_fill_2 FILLER_73_2192 ();
 sg13g2_fill_1 FILLER_73_2194 ();
 sg13g2_decap_4 FILLER_73_2201 ();
 sg13g2_fill_1 FILLER_73_2205 ();
 sg13g2_fill_2 FILLER_73_2214 ();
 sg13g2_fill_1 FILLER_73_2216 ();
 sg13g2_decap_8 FILLER_73_2221 ();
 sg13g2_decap_8 FILLER_73_2228 ();
 sg13g2_decap_8 FILLER_73_2235 ();
 sg13g2_decap_4 FILLER_73_2242 ();
 sg13g2_fill_1 FILLER_73_2246 ();
 sg13g2_decap_4 FILLER_73_2273 ();
 sg13g2_fill_1 FILLER_73_2277 ();
 sg13g2_decap_8 FILLER_73_2304 ();
 sg13g2_fill_2 FILLER_73_2311 ();
 sg13g2_fill_1 FILLER_73_2313 ();
 sg13g2_decap_4 FILLER_73_2318 ();
 sg13g2_fill_2 FILLER_73_2365 ();
 sg13g2_fill_1 FILLER_73_2390 ();
 sg13g2_fill_2 FILLER_73_2416 ();
 sg13g2_fill_1 FILLER_73_2422 ();
 sg13g2_fill_1 FILLER_73_2457 ();
 sg13g2_fill_1 FILLER_73_2462 ();
 sg13g2_fill_2 FILLER_73_2476 ();
 sg13g2_fill_1 FILLER_73_2478 ();
 sg13g2_fill_2 FILLER_73_2576 ();
 sg13g2_fill_1 FILLER_73_2578 ();
 sg13g2_decap_8 FILLER_73_2583 ();
 sg13g2_decap_8 FILLER_73_2594 ();
 sg13g2_decap_8 FILLER_73_2601 ();
 sg13g2_decap_8 FILLER_73_2608 ();
 sg13g2_decap_8 FILLER_73_2615 ();
 sg13g2_decap_8 FILLER_73_2622 ();
 sg13g2_decap_8 FILLER_73_2629 ();
 sg13g2_decap_8 FILLER_73_2636 ();
 sg13g2_decap_8 FILLER_73_2643 ();
 sg13g2_decap_8 FILLER_73_2650 ();
 sg13g2_decap_8 FILLER_73_2657 ();
 sg13g2_decap_4 FILLER_73_2664 ();
 sg13g2_fill_2 FILLER_73_2668 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_54 ();
 sg13g2_decap_8 FILLER_74_60 ();
 sg13g2_fill_1 FILLER_74_67 ();
 sg13g2_decap_8 FILLER_74_94 ();
 sg13g2_decap_8 FILLER_74_101 ();
 sg13g2_decap_8 FILLER_74_108 ();
 sg13g2_fill_2 FILLER_74_115 ();
 sg13g2_fill_1 FILLER_74_117 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_fill_1 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_248 ();
 sg13g2_fill_2 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_299 ();
 sg13g2_fill_1 FILLER_74_317 ();
 sg13g2_fill_2 FILLER_74_354 ();
 sg13g2_fill_1 FILLER_74_383 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_fill_1 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_406 ();
 sg13g2_fill_2 FILLER_74_457 ();
 sg13g2_fill_1 FILLER_74_459 ();
 sg13g2_decap_8 FILLER_74_474 ();
 sg13g2_fill_2 FILLER_74_481 ();
 sg13g2_decap_4 FILLER_74_514 ();
 sg13g2_fill_2 FILLER_74_518 ();
 sg13g2_decap_8 FILLER_74_530 ();
 sg13g2_fill_2 FILLER_74_537 ();
 sg13g2_decap_8 FILLER_74_591 ();
 sg13g2_fill_1 FILLER_74_598 ();
 sg13g2_decap_4 FILLER_74_612 ();
 sg13g2_fill_1 FILLER_74_616 ();
 sg13g2_fill_2 FILLER_74_629 ();
 sg13g2_fill_2 FILLER_74_651 ();
 sg13g2_fill_2 FILLER_74_679 ();
 sg13g2_fill_1 FILLER_74_681 ();
 sg13g2_fill_1 FILLER_74_687 ();
 sg13g2_fill_1 FILLER_74_693 ();
 sg13g2_fill_2 FILLER_74_714 ();
 sg13g2_fill_1 FILLER_74_720 ();
 sg13g2_decap_4 FILLER_74_725 ();
 sg13g2_fill_2 FILLER_74_744 ();
 sg13g2_fill_1 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_4 FILLER_74_795 ();
 sg13g2_fill_1 FILLER_74_799 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_fill_2 FILLER_74_819 ();
 sg13g2_fill_1 FILLER_74_821 ();
 sg13g2_fill_2 FILLER_74_834 ();
 sg13g2_fill_1 FILLER_74_845 ();
 sg13g2_fill_1 FILLER_74_860 ();
 sg13g2_fill_1 FILLER_74_865 ();
 sg13g2_fill_1 FILLER_74_910 ();
 sg13g2_decap_8 FILLER_74_958 ();
 sg13g2_decap_4 FILLER_74_965 ();
 sg13g2_fill_1 FILLER_74_969 ();
 sg13g2_fill_1 FILLER_74_985 ();
 sg13g2_fill_1 FILLER_74_1003 ();
 sg13g2_fill_2 FILLER_74_1065 ();
 sg13g2_fill_1 FILLER_74_1071 ();
 sg13g2_decap_8 FILLER_74_1077 ();
 sg13g2_decap_4 FILLER_74_1092 ();
 sg13g2_fill_1 FILLER_74_1096 ();
 sg13g2_decap_4 FILLER_74_1106 ();
 sg13g2_decap_8 FILLER_74_1145 ();
 sg13g2_decap_8 FILLER_74_1152 ();
 sg13g2_decap_4 FILLER_74_1159 ();
 sg13g2_fill_1 FILLER_74_1163 ();
 sg13g2_fill_1 FILLER_74_1202 ();
 sg13g2_decap_4 FILLER_74_1233 ();
 sg13g2_decap_4 FILLER_74_1242 ();
 sg13g2_fill_2 FILLER_74_1246 ();
 sg13g2_decap_4 FILLER_74_1257 ();
 sg13g2_fill_2 FILLER_74_1261 ();
 sg13g2_decap_4 FILLER_74_1277 ();
 sg13g2_decap_8 FILLER_74_1287 ();
 sg13g2_fill_2 FILLER_74_1294 ();
 sg13g2_fill_2 FILLER_74_1300 ();
 sg13g2_decap_8 FILLER_74_1318 ();
 sg13g2_fill_2 FILLER_74_1325 ();
 sg13g2_fill_2 FILLER_74_1332 ();
 sg13g2_fill_1 FILLER_74_1334 ();
 sg13g2_decap_4 FILLER_74_1343 ();
 sg13g2_fill_2 FILLER_74_1347 ();
 sg13g2_fill_2 FILLER_74_1354 ();
 sg13g2_fill_2 FILLER_74_1360 ();
 sg13g2_fill_2 FILLER_74_1367 ();
 sg13g2_fill_2 FILLER_74_1392 ();
 sg13g2_fill_2 FILLER_74_1399 ();
 sg13g2_fill_1 FILLER_74_1401 ();
 sg13g2_fill_2 FILLER_74_1412 ();
 sg13g2_fill_1 FILLER_74_1414 ();
 sg13g2_fill_2 FILLER_74_1420 ();
 sg13g2_fill_1 FILLER_74_1422 ();
 sg13g2_fill_1 FILLER_74_1432 ();
 sg13g2_decap_8 FILLER_74_1445 ();
 sg13g2_fill_2 FILLER_74_1452 ();
 sg13g2_fill_1 FILLER_74_1454 ();
 sg13g2_decap_8 FILLER_74_1460 ();
 sg13g2_fill_1 FILLER_74_1467 ();
 sg13g2_fill_1 FILLER_74_1472 ();
 sg13g2_fill_2 FILLER_74_1539 ();
 sg13g2_decap_8 FILLER_74_1551 ();
 sg13g2_fill_2 FILLER_74_1558 ();
 sg13g2_fill_1 FILLER_74_1560 ();
 sg13g2_fill_1 FILLER_74_1574 ();
 sg13g2_fill_1 FILLER_74_1580 ();
 sg13g2_decap_4 FILLER_74_1596 ();
 sg13g2_fill_1 FILLER_74_1600 ();
 sg13g2_fill_2 FILLER_74_1605 ();
 sg13g2_fill_1 FILLER_74_1617 ();
 sg13g2_fill_2 FILLER_74_1635 ();
 sg13g2_decap_8 FILLER_74_1649 ();
 sg13g2_fill_1 FILLER_74_1656 ();
 sg13g2_fill_2 FILLER_74_1671 ();
 sg13g2_fill_1 FILLER_74_1679 ();
 sg13g2_fill_1 FILLER_74_1684 ();
 sg13g2_fill_1 FILLER_74_1691 ();
 sg13g2_fill_2 FILLER_74_1718 ();
 sg13g2_fill_2 FILLER_74_1740 ();
 sg13g2_fill_1 FILLER_74_1752 ();
 sg13g2_decap_8 FILLER_74_1759 ();
 sg13g2_decap_4 FILLER_74_1781 ();
 sg13g2_fill_1 FILLER_74_1785 ();
 sg13g2_fill_2 FILLER_74_1839 ();
 sg13g2_fill_1 FILLER_74_1841 ();
 sg13g2_fill_1 FILLER_74_1861 ();
 sg13g2_fill_1 FILLER_74_1867 ();
 sg13g2_fill_2 FILLER_74_1909 ();
 sg13g2_fill_1 FILLER_74_1937 ();
 sg13g2_decap_4 FILLER_74_1978 ();
 sg13g2_fill_2 FILLER_74_1982 ();
 sg13g2_decap_8 FILLER_74_1988 ();
 sg13g2_decap_8 FILLER_74_2035 ();
 sg13g2_decap_4 FILLER_74_2042 ();
 sg13g2_decap_8 FILLER_74_2050 ();
 sg13g2_decap_8 FILLER_74_2057 ();
 sg13g2_decap_8 FILLER_74_2064 ();
 sg13g2_fill_2 FILLER_74_2071 ();
 sg13g2_fill_2 FILLER_74_2087 ();
 sg13g2_fill_1 FILLER_74_2089 ();
 sg13g2_decap_8 FILLER_74_2094 ();
 sg13g2_decap_4 FILLER_74_2101 ();
 sg13g2_fill_2 FILLER_74_2105 ();
 sg13g2_decap_4 FILLER_74_2127 ();
 sg13g2_fill_1 FILLER_74_2146 ();
 sg13g2_decap_4 FILLER_74_2187 ();
 sg13g2_decap_8 FILLER_74_2201 ();
 sg13g2_fill_2 FILLER_74_2208 ();
 sg13g2_fill_1 FILLER_74_2210 ();
 sg13g2_decap_4 FILLER_74_2237 ();
 sg13g2_fill_1 FILLER_74_2241 ();
 sg13g2_fill_2 FILLER_74_2278 ();
 sg13g2_fill_1 FILLER_74_2280 ();
 sg13g2_decap_4 FILLER_74_2295 ();
 sg13g2_decap_8 FILLER_74_2303 ();
 sg13g2_decap_8 FILLER_74_2310 ();
 sg13g2_decap_8 FILLER_74_2317 ();
 sg13g2_fill_1 FILLER_74_2328 ();
 sg13g2_fill_1 FILLER_74_2423 ();
 sg13g2_decap_8 FILLER_74_2481 ();
 sg13g2_decap_8 FILLER_74_2488 ();
 sg13g2_decap_4 FILLER_74_2495 ();
 sg13g2_fill_1 FILLER_74_2499 ();
 sg13g2_decap_8 FILLER_74_2504 ();
 sg13g2_decap_4 FILLER_74_2511 ();
 sg13g2_fill_2 FILLER_74_2515 ();
 sg13g2_fill_2 FILLER_74_2527 ();
 sg13g2_fill_1 FILLER_74_2529 ();
 sg13g2_decap_4 FILLER_74_2534 ();
 sg13g2_fill_1 FILLER_74_2538 ();
 sg13g2_decap_8 FILLER_74_2553 ();
 sg13g2_fill_1 FILLER_74_2560 ();
 sg13g2_decap_8 FILLER_74_2587 ();
 sg13g2_decap_8 FILLER_74_2594 ();
 sg13g2_decap_8 FILLER_74_2601 ();
 sg13g2_decap_8 FILLER_74_2608 ();
 sg13g2_decap_8 FILLER_74_2615 ();
 sg13g2_decap_8 FILLER_74_2622 ();
 sg13g2_decap_8 FILLER_74_2629 ();
 sg13g2_decap_8 FILLER_74_2636 ();
 sg13g2_decap_8 FILLER_74_2643 ();
 sg13g2_decap_8 FILLER_74_2650 ();
 sg13g2_decap_8 FILLER_74_2657 ();
 sg13g2_decap_4 FILLER_74_2664 ();
 sg13g2_fill_2 FILLER_74_2668 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_61 ();
 sg13g2_fill_2 FILLER_75_68 ();
 sg13g2_fill_1 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_86 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_96 ();
 sg13g2_decap_8 FILLER_75_100 ();
 sg13g2_decap_4 FILLER_75_107 ();
 sg13g2_fill_2 FILLER_75_111 ();
 sg13g2_decap_4 FILLER_75_117 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_fill_2 FILLER_75_153 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_fill_1 FILLER_75_228 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_341 ();
 sg13g2_fill_2 FILLER_75_358 ();
 sg13g2_fill_2 FILLER_75_364 ();
 sg13g2_fill_2 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_fill_1 FILLER_75_396 ();
 sg13g2_fill_1 FILLER_75_423 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_fill_1 FILLER_75_434 ();
 sg13g2_fill_2 FILLER_75_440 ();
 sg13g2_fill_2 FILLER_75_446 ();
 sg13g2_fill_1 FILLER_75_448 ();
 sg13g2_fill_1 FILLER_75_454 ();
 sg13g2_decap_4 FILLER_75_505 ();
 sg13g2_fill_1 FILLER_75_509 ();
 sg13g2_fill_1 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_521 ();
 sg13g2_decap_4 FILLER_75_527 ();
 sg13g2_fill_2 FILLER_75_531 ();
 sg13g2_fill_2 FILLER_75_543 ();
 sg13g2_decap_4 FILLER_75_576 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_2 FILLER_75_634 ();
 sg13g2_fill_2 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_665 ();
 sg13g2_fill_2 FILLER_75_672 ();
 sg13g2_fill_1 FILLER_75_697 ();
 sg13g2_fill_2 FILLER_75_714 ();
 sg13g2_fill_1 FILLER_75_716 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_723 ();
 sg13g2_fill_2 FILLER_75_732 ();
 sg13g2_fill_1 FILLER_75_741 ();
 sg13g2_fill_2 FILLER_75_746 ();
 sg13g2_fill_2 FILLER_75_774 ();
 sg13g2_fill_2 FILLER_75_786 ();
 sg13g2_fill_1 FILLER_75_788 ();
 sg13g2_fill_2 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_4 FILLER_75_829 ();
 sg13g2_fill_2 FILLER_75_833 ();
 sg13g2_fill_1 FILLER_75_839 ();
 sg13g2_fill_1 FILLER_75_851 ();
 sg13g2_fill_2 FILLER_75_863 ();
 sg13g2_fill_1 FILLER_75_865 ();
 sg13g2_fill_2 FILLER_75_873 ();
 sg13g2_fill_2 FILLER_75_910 ();
 sg13g2_fill_1 FILLER_75_937 ();
 sg13g2_fill_2 FILLER_75_942 ();
 sg13g2_fill_2 FILLER_75_963 ();
 sg13g2_fill_1 FILLER_75_965 ();
 sg13g2_fill_2 FILLER_75_994 ();
 sg13g2_fill_1 FILLER_75_1006 ();
 sg13g2_fill_1 FILLER_75_1020 ();
 sg13g2_fill_2 FILLER_75_1025 ();
 sg13g2_decap_4 FILLER_75_1032 ();
 sg13g2_decap_8 FILLER_75_1041 ();
 sg13g2_decap_4 FILLER_75_1048 ();
 sg13g2_decap_4 FILLER_75_1074 ();
 sg13g2_fill_1 FILLER_75_1078 ();
 sg13g2_fill_1 FILLER_75_1082 ();
 sg13g2_fill_2 FILLER_75_1089 ();
 sg13g2_fill_1 FILLER_75_1091 ();
 sg13g2_fill_1 FILLER_75_1103 ();
 sg13g2_decap_8 FILLER_75_1111 ();
 sg13g2_decap_8 FILLER_75_1152 ();
 sg13g2_decap_4 FILLER_75_1171 ();
 sg13g2_fill_1 FILLER_75_1180 ();
 sg13g2_fill_1 FILLER_75_1211 ();
 sg13g2_decap_4 FILLER_75_1226 ();
 sg13g2_fill_1 FILLER_75_1230 ();
 sg13g2_decap_8 FILLER_75_1239 ();
 sg13g2_fill_1 FILLER_75_1246 ();
 sg13g2_decap_4 FILLER_75_1253 ();
 sg13g2_fill_1 FILLER_75_1257 ();
 sg13g2_fill_1 FILLER_75_1263 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_4 FILLER_75_1292 ();
 sg13g2_fill_1 FILLER_75_1341 ();
 sg13g2_fill_1 FILLER_75_1347 ();
 sg13g2_fill_1 FILLER_75_1373 ();
 sg13g2_fill_2 FILLER_75_1382 ();
 sg13g2_fill_1 FILLER_75_1419 ();
 sg13g2_fill_2 FILLER_75_1430 ();
 sg13g2_fill_1 FILLER_75_1432 ();
 sg13g2_decap_4 FILLER_75_1439 ();
 sg13g2_fill_2 FILLER_75_1494 ();
 sg13g2_decap_8 FILLER_75_1525 ();
 sg13g2_fill_2 FILLER_75_1532 ();
 sg13g2_decap_8 FILLER_75_1537 ();
 sg13g2_fill_1 FILLER_75_1544 ();
 sg13g2_decap_8 FILLER_75_1548 ();
 sg13g2_fill_2 FILLER_75_1555 ();
 sg13g2_decap_8 FILLER_75_1564 ();
 sg13g2_decap_4 FILLER_75_1575 ();
 sg13g2_decap_8 FILLER_75_1619 ();
 sg13g2_fill_1 FILLER_75_1626 ();
 sg13g2_fill_2 FILLER_75_1645 ();
 sg13g2_fill_1 FILLER_75_1647 ();
 sg13g2_decap_4 FILLER_75_1652 ();
 sg13g2_fill_2 FILLER_75_1662 ();
 sg13g2_fill_2 FILLER_75_1673 ();
 sg13g2_fill_2 FILLER_75_1680 ();
 sg13g2_fill_1 FILLER_75_1682 ();
 sg13g2_fill_1 FILLER_75_1687 ();
 sg13g2_decap_8 FILLER_75_1693 ();
 sg13g2_fill_1 FILLER_75_1700 ();
 sg13g2_decap_4 FILLER_75_1705 ();
 sg13g2_fill_2 FILLER_75_1709 ();
 sg13g2_fill_1 FILLER_75_1745 ();
 sg13g2_fill_2 FILLER_75_1798 ();
 sg13g2_fill_2 FILLER_75_1806 ();
 sg13g2_fill_1 FILLER_75_1812 ();
 sg13g2_fill_2 FILLER_75_1837 ();
 sg13g2_fill_1 FILLER_75_1839 ();
 sg13g2_fill_1 FILLER_75_1851 ();
 sg13g2_fill_2 FILLER_75_1856 ();
 sg13g2_fill_1 FILLER_75_1894 ();
 sg13g2_fill_2 FILLER_75_1899 ();
 sg13g2_fill_2 FILLER_75_1909 ();
 sg13g2_fill_2 FILLER_75_1921 ();
 sg13g2_fill_1 FILLER_75_1943 ();
 sg13g2_decap_8 FILLER_75_1960 ();
 sg13g2_decap_8 FILLER_75_1967 ();
 sg13g2_decap_4 FILLER_75_1987 ();
 sg13g2_fill_2 FILLER_75_1991 ();
 sg13g2_decap_4 FILLER_75_2006 ();
 sg13g2_fill_2 FILLER_75_2010 ();
 sg13g2_fill_2 FILLER_75_2016 ();
 sg13g2_decap_8 FILLER_75_2022 ();
 sg13g2_fill_1 FILLER_75_2072 ();
 sg13g2_fill_2 FILLER_75_2076 ();
 sg13g2_fill_1 FILLER_75_2084 ();
 sg13g2_fill_2 FILLER_75_2090 ();
 sg13g2_fill_1 FILLER_75_2092 ();
 sg13g2_fill_1 FILLER_75_2105 ();
 sg13g2_decap_8 FILLER_75_2111 ();
 sg13g2_fill_2 FILLER_75_2129 ();
 sg13g2_fill_1 FILLER_75_2131 ();
 sg13g2_fill_2 FILLER_75_2143 ();
 sg13g2_fill_1 FILLER_75_2178 ();
 sg13g2_decap_4 FILLER_75_2189 ();
 sg13g2_fill_1 FILLER_75_2193 ();
 sg13g2_fill_1 FILLER_75_2198 ();
 sg13g2_fill_2 FILLER_75_2225 ();
 sg13g2_decap_4 FILLER_75_2284 ();
 sg13g2_fill_2 FILLER_75_2288 ();
 sg13g2_decap_8 FILLER_75_2316 ();
 sg13g2_decap_8 FILLER_75_2323 ();
 sg13g2_fill_2 FILLER_75_2330 ();
 sg13g2_fill_1 FILLER_75_2332 ();
 sg13g2_fill_1 FILLER_75_2343 ();
 sg13g2_fill_2 FILLER_75_2354 ();
 sg13g2_fill_2 FILLER_75_2423 ();
 sg13g2_fill_2 FILLER_75_2448 ();
 sg13g2_decap_8 FILLER_75_2469 ();
 sg13g2_decap_8 FILLER_75_2476 ();
 sg13g2_decap_8 FILLER_75_2483 ();
 sg13g2_decap_8 FILLER_75_2490 ();
 sg13g2_decap_8 FILLER_75_2497 ();
 sg13g2_decap_8 FILLER_75_2504 ();
 sg13g2_decap_8 FILLER_75_2511 ();
 sg13g2_decap_4 FILLER_75_2518 ();
 sg13g2_fill_2 FILLER_75_2522 ();
 sg13g2_decap_8 FILLER_75_2528 ();
 sg13g2_decap_4 FILLER_75_2535 ();
 sg13g2_fill_2 FILLER_75_2565 ();
 sg13g2_decap_8 FILLER_75_2571 ();
 sg13g2_decap_8 FILLER_75_2578 ();
 sg13g2_decap_8 FILLER_75_2585 ();
 sg13g2_decap_8 FILLER_75_2592 ();
 sg13g2_decap_8 FILLER_75_2599 ();
 sg13g2_decap_8 FILLER_75_2606 ();
 sg13g2_decap_8 FILLER_75_2613 ();
 sg13g2_decap_8 FILLER_75_2620 ();
 sg13g2_decap_8 FILLER_75_2627 ();
 sg13g2_decap_8 FILLER_75_2634 ();
 sg13g2_decap_8 FILLER_75_2641 ();
 sg13g2_decap_8 FILLER_75_2648 ();
 sg13g2_decap_8 FILLER_75_2655 ();
 sg13g2_decap_8 FILLER_75_2662 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_4 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_36 ();
 sg13g2_decap_8 FILLER_76_43 ();
 sg13g2_decap_8 FILLER_76_50 ();
 sg13g2_decap_4 FILLER_76_57 ();
 sg13g2_fill_1 FILLER_76_61 ();
 sg13g2_fill_1 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_1 FILLER_76_127 ();
 sg13g2_fill_1 FILLER_76_134 ();
 sg13g2_fill_1 FILLER_76_148 ();
 sg13g2_fill_1 FILLER_76_214 ();
 sg13g2_fill_1 FILLER_76_219 ();
 sg13g2_fill_2 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_244 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_307 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_fill_2 FILLER_76_352 ();
 sg13g2_fill_1 FILLER_76_359 ();
 sg13g2_fill_2 FILLER_76_365 ();
 sg13g2_fill_1 FILLER_76_367 ();
 sg13g2_fill_2 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_fill_1 FILLER_76_394 ();
 sg13g2_fill_1 FILLER_76_400 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_413 ();
 sg13g2_fill_2 FILLER_76_423 ();
 sg13g2_fill_1 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_76_442 ();
 sg13g2_decap_4 FILLER_76_448 ();
 sg13g2_fill_1 FILLER_76_452 ();
 sg13g2_fill_2 FILLER_76_461 ();
 sg13g2_fill_1 FILLER_76_463 ();
 sg13g2_decap_4 FILLER_76_468 ();
 sg13g2_fill_2 FILLER_76_472 ();
 sg13g2_fill_2 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_491 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_fill_2 FILLER_76_546 ();
 sg13g2_decap_4 FILLER_76_553 ();
 sg13g2_fill_1 FILLER_76_557 ();
 sg13g2_decap_4 FILLER_76_581 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_fill_1 FILLER_76_710 ();
 sg13g2_fill_2 FILLER_76_729 ();
 sg13g2_fill_1 FILLER_76_759 ();
 sg13g2_fill_1 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_792 ();
 sg13g2_fill_1 FILLER_76_799 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_4 FILLER_76_819 ();
 sg13g2_fill_2 FILLER_76_823 ();
 sg13g2_fill_1 FILLER_76_830 ();
 sg13g2_fill_2 FILLER_76_867 ();
 sg13g2_fill_1 FILLER_76_869 ();
 sg13g2_fill_2 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_906 ();
 sg13g2_fill_1 FILLER_76_908 ();
 sg13g2_fill_1 FILLER_76_920 ();
 sg13g2_fill_1 FILLER_76_977 ();
 sg13g2_fill_1 FILLER_76_993 ();
 sg13g2_fill_2 FILLER_76_1041 ();
 sg13g2_fill_1 FILLER_76_1047 ();
 sg13g2_fill_1 FILLER_76_1058 ();
 sg13g2_fill_1 FILLER_76_1075 ();
 sg13g2_fill_1 FILLER_76_1085 ();
 sg13g2_fill_2 FILLER_76_1090 ();
 sg13g2_decap_4 FILLER_76_1099 ();
 sg13g2_decap_8 FILLER_76_1107 ();
 sg13g2_fill_2 FILLER_76_1114 ();
 sg13g2_fill_1 FILLER_76_1116 ();
 sg13g2_fill_2 FILLER_76_1127 ();
 sg13g2_fill_1 FILLER_76_1129 ();
 sg13g2_decap_8 FILLER_76_1138 ();
 sg13g2_fill_2 FILLER_76_1145 ();
 sg13g2_fill_1 FILLER_76_1147 ();
 sg13g2_decap_4 FILLER_76_1174 ();
 sg13g2_fill_2 FILLER_76_1178 ();
 sg13g2_fill_1 FILLER_76_1188 ();
 sg13g2_decap_8 FILLER_76_1220 ();
 sg13g2_fill_2 FILLER_76_1227 ();
 sg13g2_fill_1 FILLER_76_1229 ();
 sg13g2_decap_8 FILLER_76_1238 ();
 sg13g2_decap_8 FILLER_76_1245 ();
 sg13g2_fill_1 FILLER_76_1283 ();
 sg13g2_fill_1 FILLER_76_1293 ();
 sg13g2_fill_1 FILLER_76_1305 ();
 sg13g2_fill_2 FILLER_76_1338 ();
 sg13g2_fill_1 FILLER_76_1340 ();
 sg13g2_decap_4 FILLER_76_1440 ();
 sg13g2_fill_1 FILLER_76_1444 ();
 sg13g2_decap_4 FILLER_76_1449 ();
 sg13g2_fill_1 FILLER_76_1453 ();
 sg13g2_decap_8 FILLER_76_1474 ();
 sg13g2_fill_2 FILLER_76_1481 ();
 sg13g2_fill_1 FILLER_76_1492 ();
 sg13g2_fill_1 FILLER_76_1500 ();
 sg13g2_fill_2 FILLER_76_1523 ();
 sg13g2_fill_2 FILLER_76_1551 ();
 sg13g2_fill_2 FILLER_76_1583 ();
 sg13g2_fill_1 FILLER_76_1585 ();
 sg13g2_fill_2 FILLER_76_1589 ();
 sg13g2_fill_2 FILLER_76_1597 ();
 sg13g2_fill_1 FILLER_76_1599 ();
 sg13g2_fill_1 FILLER_76_1604 ();
 sg13g2_decap_8 FILLER_76_1615 ();
 sg13g2_fill_1 FILLER_76_1622 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1634 ();
 sg13g2_decap_4 FILLER_76_1641 ();
 sg13g2_fill_2 FILLER_76_1667 ();
 sg13g2_fill_2 FILLER_76_1674 ();
 sg13g2_decap_4 FILLER_76_1681 ();
 sg13g2_fill_2 FILLER_76_1691 ();
 sg13g2_decap_4 FILLER_76_1703 ();
 sg13g2_decap_8 FILLER_76_1743 ();
 sg13g2_decap_4 FILLER_76_1750 ();
 sg13g2_fill_1 FILLER_76_1754 ();
 sg13g2_decap_8 FILLER_76_1759 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_decap_4 FILLER_76_1776 ();
 sg13g2_fill_1 FILLER_76_1780 ();
 sg13g2_decap_8 FILLER_76_1785 ();
 sg13g2_decap_8 FILLER_76_1792 ();
 sg13g2_fill_1 FILLER_76_1799 ();
 sg13g2_decap_4 FILLER_76_1820 ();
 sg13g2_decap_4 FILLER_76_1829 ();
 sg13g2_fill_1 FILLER_76_1833 ();
 sg13g2_fill_2 FILLER_76_1845 ();
 sg13g2_fill_1 FILLER_76_1847 ();
 sg13g2_fill_1 FILLER_76_1872 ();
 sg13g2_decap_4 FILLER_76_1883 ();
 sg13g2_fill_1 FILLER_76_1887 ();
 sg13g2_decap_4 FILLER_76_1914 ();
 sg13g2_fill_1 FILLER_76_1918 ();
 sg13g2_decap_4 FILLER_76_1923 ();
 sg13g2_decap_8 FILLER_76_1937 ();
 sg13g2_fill_2 FILLER_76_1944 ();
 sg13g2_decap_8 FILLER_76_2024 ();
 sg13g2_decap_8 FILLER_76_2031 ();
 sg13g2_decap_8 FILLER_76_2038 ();
 sg13g2_decap_4 FILLER_76_2045 ();
 sg13g2_decap_8 FILLER_76_2053 ();
 sg13g2_fill_2 FILLER_76_2080 ();
 sg13g2_fill_1 FILLER_76_2087 ();
 sg13g2_fill_1 FILLER_76_2109 ();
 sg13g2_fill_1 FILLER_76_2116 ();
 sg13g2_decap_8 FILLER_76_2232 ();
 sg13g2_decap_8 FILLER_76_2239 ();
 sg13g2_decap_8 FILLER_76_2277 ();
 sg13g2_decap_4 FILLER_76_2284 ();
 sg13g2_decap_8 FILLER_76_2314 ();
 sg13g2_fill_1 FILLER_76_2321 ();
 sg13g2_decap_4 FILLER_76_2330 ();
 sg13g2_decap_4 FILLER_76_2360 ();
 sg13g2_fill_1 FILLER_76_2364 ();
 sg13g2_fill_1 FILLER_76_2443 ();
 sg13g2_decap_8 FILLER_76_2470 ();
 sg13g2_decap_8 FILLER_76_2477 ();
 sg13g2_decap_8 FILLER_76_2484 ();
 sg13g2_decap_8 FILLER_76_2491 ();
 sg13g2_decap_8 FILLER_76_2498 ();
 sg13g2_decap_8 FILLER_76_2505 ();
 sg13g2_decap_8 FILLER_76_2512 ();
 sg13g2_decap_8 FILLER_76_2519 ();
 sg13g2_decap_8 FILLER_76_2526 ();
 sg13g2_decap_8 FILLER_76_2533 ();
 sg13g2_decap_8 FILLER_76_2540 ();
 sg13g2_decap_8 FILLER_76_2547 ();
 sg13g2_decap_8 FILLER_76_2554 ();
 sg13g2_decap_8 FILLER_76_2561 ();
 sg13g2_decap_8 FILLER_76_2568 ();
 sg13g2_decap_8 FILLER_76_2575 ();
 sg13g2_decap_8 FILLER_76_2582 ();
 sg13g2_decap_8 FILLER_76_2589 ();
 sg13g2_decap_8 FILLER_76_2596 ();
 sg13g2_decap_8 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2610 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_95 ();
 sg13g2_fill_1 FILLER_77_149 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_209 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_265 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_decap_4 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_fill_2 FILLER_77_362 ();
 sg13g2_fill_1 FILLER_77_364 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_77_447 ();
 sg13g2_fill_1 FILLER_77_459 ();
 sg13g2_fill_1 FILLER_77_523 ();
 sg13g2_fill_2 FILLER_77_550 ();
 sg13g2_fill_1 FILLER_77_552 ();
 sg13g2_fill_1 FILLER_77_563 ();
 sg13g2_fill_2 FILLER_77_701 ();
 sg13g2_fill_1 FILLER_77_719 ();
 sg13g2_fill_2 FILLER_77_724 ();
 sg13g2_fill_1 FILLER_77_726 ();
 sg13g2_fill_1 FILLER_77_732 ();
 sg13g2_fill_2 FILLER_77_753 ();
 sg13g2_fill_2 FILLER_77_765 ();
 sg13g2_fill_2 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_4 FILLER_77_834 ();
 sg13g2_fill_2 FILLER_77_909 ();
 sg13g2_fill_1 FILLER_77_911 ();
 sg13g2_fill_1 FILLER_77_940 ();
 sg13g2_fill_2 FILLER_77_972 ();
 sg13g2_fill_1 FILLER_77_980 ();
 sg13g2_fill_2 FILLER_77_986 ();
 sg13g2_fill_1 FILLER_77_999 ();
 sg13g2_fill_2 FILLER_77_1020 ();
 sg13g2_fill_1 FILLER_77_1022 ();
 sg13g2_fill_1 FILLER_77_1039 ();
 sg13g2_fill_2 FILLER_77_1054 ();
 sg13g2_fill_1 FILLER_77_1056 ();
 sg13g2_fill_2 FILLER_77_1061 ();
 sg13g2_fill_1 FILLER_77_1063 ();
 sg13g2_fill_2 FILLER_77_1081 ();
 sg13g2_fill_1 FILLER_77_1083 ();
 sg13g2_fill_1 FILLER_77_1093 ();
 sg13g2_decap_8 FILLER_77_1150 ();
 sg13g2_fill_2 FILLER_77_1172 ();
 sg13g2_fill_1 FILLER_77_1174 ();
 sg13g2_fill_2 FILLER_77_1182 ();
 sg13g2_fill_1 FILLER_77_1184 ();
 sg13g2_fill_2 FILLER_77_1189 ();
 sg13g2_fill_2 FILLER_77_1218 ();
 sg13g2_fill_1 FILLER_77_1220 ();
 sg13g2_decap_4 FILLER_77_1226 ();
 sg13g2_fill_1 FILLER_77_1230 ();
 sg13g2_fill_1 FILLER_77_1256 ();
 sg13g2_decap_4 FILLER_77_1263 ();
 sg13g2_fill_1 FILLER_77_1275 ();
 sg13g2_fill_1 FILLER_77_1286 ();
 sg13g2_decap_4 FILLER_77_1318 ();
 sg13g2_fill_1 FILLER_77_1333 ();
 sg13g2_decap_4 FILLER_77_1417 ();
 sg13g2_fill_2 FILLER_77_1427 ();
 sg13g2_fill_1 FILLER_77_1429 ();
 sg13g2_fill_1 FILLER_77_1459 ();
 sg13g2_decap_4 FILLER_77_1468 ();
 sg13g2_fill_1 FILLER_77_1519 ();
 sg13g2_fill_1 FILLER_77_1524 ();
 sg13g2_fill_1 FILLER_77_1551 ();
 sg13g2_fill_2 FILLER_77_1562 ();
 sg13g2_decap_8 FILLER_77_1590 ();
 sg13g2_decap_8 FILLER_77_1597 ();
 sg13g2_fill_2 FILLER_77_1614 ();
 sg13g2_decap_8 FILLER_77_1642 ();
 sg13g2_decap_4 FILLER_77_1659 ();
 sg13g2_fill_1 FILLER_77_1663 ();
 sg13g2_decap_8 FILLER_77_1669 ();
 sg13g2_fill_2 FILLER_77_1676 ();
 sg13g2_decap_4 FILLER_77_1688 ();
 sg13g2_fill_1 FILLER_77_1718 ();
 sg13g2_fill_2 FILLER_77_1762 ();
 sg13g2_fill_1 FILLER_77_1790 ();
 sg13g2_fill_1 FILLER_77_1817 ();
 sg13g2_fill_1 FILLER_77_1828 ();
 sg13g2_decap_8 FILLER_77_1833 ();
 sg13g2_fill_1 FILLER_77_1840 ();
 sg13g2_fill_2 FILLER_77_1851 ();
 sg13g2_fill_1 FILLER_77_1853 ();
 sg13g2_fill_1 FILLER_77_1867 ();
 sg13g2_decap_4 FILLER_77_1898 ();
 sg13g2_fill_1 FILLER_77_1902 ();
 sg13g2_decap_4 FILLER_77_1909 ();
 sg13g2_fill_1 FILLER_77_1913 ();
 sg13g2_decap_4 FILLER_77_1963 ();
 sg13g2_decap_4 FILLER_77_1971 ();
 sg13g2_fill_2 FILLER_77_1991 ();
 sg13g2_decap_8 FILLER_77_2007 ();
 sg13g2_decap_4 FILLER_77_2014 ();
 sg13g2_fill_2 FILLER_77_2018 ();
 sg13g2_decap_8 FILLER_77_2046 ();
 sg13g2_decap_4 FILLER_77_2053 ();
 sg13g2_fill_2 FILLER_77_2057 ();
 sg13g2_fill_2 FILLER_77_2089 ();
 sg13g2_decap_4 FILLER_77_2095 ();
 sg13g2_fill_2 FILLER_77_2139 ();
 sg13g2_fill_2 FILLER_77_2194 ();
 sg13g2_decap_8 FILLER_77_2234 ();
 sg13g2_decap_8 FILLER_77_2241 ();
 sg13g2_decap_8 FILLER_77_2248 ();
 sg13g2_decap_8 FILLER_77_2255 ();
 sg13g2_decap_8 FILLER_77_2262 ();
 sg13g2_decap_8 FILLER_77_2269 ();
 sg13g2_decap_8 FILLER_77_2276 ();
 sg13g2_decap_8 FILLER_77_2283 ();
 sg13g2_fill_2 FILLER_77_2290 ();
 sg13g2_fill_1 FILLER_77_2292 ();
 sg13g2_decap_8 FILLER_77_2297 ();
 sg13g2_decap_8 FILLER_77_2304 ();
 sg13g2_decap_8 FILLER_77_2311 ();
 sg13g2_decap_8 FILLER_77_2318 ();
 sg13g2_decap_8 FILLER_77_2325 ();
 sg13g2_decap_8 FILLER_77_2332 ();
 sg13g2_decap_4 FILLER_77_2343 ();
 sg13g2_fill_1 FILLER_77_2347 ();
 sg13g2_decap_8 FILLER_77_2352 ();
 sg13g2_decap_4 FILLER_77_2359 ();
 sg13g2_fill_2 FILLER_77_2363 ();
 sg13g2_fill_1 FILLER_77_2401 ();
 sg13g2_fill_2 FILLER_77_2406 ();
 sg13g2_fill_2 FILLER_77_2414 ();
 sg13g2_fill_2 FILLER_77_2434 ();
 sg13g2_decap_8 FILLER_77_2456 ();
 sg13g2_decap_8 FILLER_77_2463 ();
 sg13g2_decap_8 FILLER_77_2470 ();
 sg13g2_decap_8 FILLER_77_2477 ();
 sg13g2_decap_8 FILLER_77_2484 ();
 sg13g2_decap_8 FILLER_77_2491 ();
 sg13g2_decap_8 FILLER_77_2498 ();
 sg13g2_decap_8 FILLER_77_2505 ();
 sg13g2_decap_8 FILLER_77_2512 ();
 sg13g2_decap_8 FILLER_77_2519 ();
 sg13g2_decap_8 FILLER_77_2526 ();
 sg13g2_decap_8 FILLER_77_2533 ();
 sg13g2_decap_8 FILLER_77_2540 ();
 sg13g2_decap_8 FILLER_77_2547 ();
 sg13g2_decap_8 FILLER_77_2554 ();
 sg13g2_decap_8 FILLER_77_2561 ();
 sg13g2_decap_8 FILLER_77_2568 ();
 sg13g2_decap_8 FILLER_77_2575 ();
 sg13g2_decap_8 FILLER_77_2582 ();
 sg13g2_decap_8 FILLER_77_2589 ();
 sg13g2_decap_8 FILLER_77_2596 ();
 sg13g2_decap_8 FILLER_77_2603 ();
 sg13g2_decap_8 FILLER_77_2610 ();
 sg13g2_decap_8 FILLER_77_2617 ();
 sg13g2_decap_8 FILLER_77_2624 ();
 sg13g2_decap_8 FILLER_77_2631 ();
 sg13g2_decap_8 FILLER_77_2638 ();
 sg13g2_decap_8 FILLER_77_2645 ();
 sg13g2_decap_8 FILLER_77_2652 ();
 sg13g2_decap_8 FILLER_77_2659 ();
 sg13g2_decap_4 FILLER_77_2666 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_fill_1 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_114 ();
 sg13g2_fill_2 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_260 ();
 sg13g2_fill_2 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_fill_2 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_357 ();
 sg13g2_decap_4 FILLER_78_384 ();
 sg13g2_fill_1 FILLER_78_388 ();
 sg13g2_fill_1 FILLER_78_394 ();
 sg13g2_fill_2 FILLER_78_421 ();
 sg13g2_fill_1 FILLER_78_423 ();
 sg13g2_fill_2 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_447 ();
 sg13g2_fill_2 FILLER_78_474 ();
 sg13g2_fill_2 FILLER_78_536 ();
 sg13g2_fill_2 FILLER_78_584 ();
 sg13g2_decap_4 FILLER_78_616 ();
 sg13g2_fill_2 FILLER_78_620 ();
 sg13g2_fill_2 FILLER_78_626 ();
 sg13g2_fill_1 FILLER_78_628 ();
 sg13g2_fill_2 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_802 ();
 sg13g2_fill_2 FILLER_78_809 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_fill_2 FILLER_78_836 ();
 sg13g2_fill_1 FILLER_78_879 ();
 sg13g2_fill_2 FILLER_78_898 ();
 sg13g2_fill_1 FILLER_78_904 ();
 sg13g2_fill_1 FILLER_78_911 ();
 sg13g2_fill_1 FILLER_78_918 ();
 sg13g2_fill_1 FILLER_78_937 ();
 sg13g2_fill_1 FILLER_78_951 ();
 sg13g2_fill_2 FILLER_78_956 ();
 sg13g2_fill_2 FILLER_78_962 ();
 sg13g2_fill_2 FILLER_78_979 ();
 sg13g2_fill_1 FILLER_78_981 ();
 sg13g2_fill_1 FILLER_78_992 ();
 sg13g2_fill_1 FILLER_78_1016 ();
 sg13g2_fill_1 FILLER_78_1021 ();
 sg13g2_fill_1 FILLER_78_1062 ();
 sg13g2_fill_2 FILLER_78_1067 ();
 sg13g2_fill_1 FILLER_78_1069 ();
 sg13g2_fill_2 FILLER_78_1079 ();
 sg13g2_fill_2 FILLER_78_1114 ();
 sg13g2_fill_1 FILLER_78_1116 ();
 sg13g2_decap_4 FILLER_78_1148 ();
 sg13g2_decap_8 FILLER_78_1178 ();
 sg13g2_decap_4 FILLER_78_1185 ();
 sg13g2_fill_1 FILLER_78_1241 ();
 sg13g2_decap_4 FILLER_78_1246 ();
 sg13g2_fill_2 FILLER_78_1285 ();
 sg13g2_fill_1 FILLER_78_1322 ();
 sg13g2_fill_2 FILLER_78_1328 ();
 sg13g2_fill_1 FILLER_78_1330 ();
 sg13g2_fill_1 FILLER_78_1364 ();
 sg13g2_fill_2 FILLER_78_1369 ();
 sg13g2_fill_1 FILLER_78_1375 ();
 sg13g2_fill_1 FILLER_78_1395 ();
 sg13g2_decap_4 FILLER_78_1435 ();
 sg13g2_fill_1 FILLER_78_1439 ();
 sg13g2_decap_8 FILLER_78_1444 ();
 sg13g2_decap_4 FILLER_78_1451 ();
 sg13g2_fill_2 FILLER_78_1459 ();
 sg13g2_fill_1 FILLER_78_1461 ();
 sg13g2_fill_2 FILLER_78_1488 ();
 sg13g2_fill_2 FILLER_78_1598 ();
 sg13g2_fill_2 FILLER_78_1626 ();
 sg13g2_fill_1 FILLER_78_1628 ();
 sg13g2_fill_2 FILLER_78_1639 ();
 sg13g2_fill_1 FILLER_78_1641 ();
 sg13g2_fill_2 FILLER_78_1668 ();
 sg13g2_fill_1 FILLER_78_1722 ();
 sg13g2_fill_2 FILLER_78_1837 ();
 sg13g2_decap_4 FILLER_78_1875 ();
 sg13g2_fill_1 FILLER_78_1879 ();
 sg13g2_fill_1 FILLER_78_1972 ();
 sg13g2_fill_1 FILLER_78_1983 ();
 sg13g2_fill_1 FILLER_78_1994 ();
 sg13g2_fill_1 FILLER_78_2021 ();
 sg13g2_decap_8 FILLER_78_2048 ();
 sg13g2_decap_8 FILLER_78_2055 ();
 sg13g2_fill_2 FILLER_78_2062 ();
 sg13g2_fill_2 FILLER_78_2094 ();
 sg13g2_fill_1 FILLER_78_2156 ();
 sg13g2_fill_1 FILLER_78_2162 ();
 sg13g2_fill_1 FILLER_78_2167 ();
 sg13g2_fill_1 FILLER_78_2194 ();
 sg13g2_fill_1 FILLER_78_2199 ();
 sg13g2_fill_1 FILLER_78_2226 ();
 sg13g2_decap_8 FILLER_78_2253 ();
 sg13g2_decap_8 FILLER_78_2260 ();
 sg13g2_decap_8 FILLER_78_2267 ();
 sg13g2_decap_8 FILLER_78_2274 ();
 sg13g2_decap_8 FILLER_78_2281 ();
 sg13g2_decap_8 FILLER_78_2288 ();
 sg13g2_decap_8 FILLER_78_2295 ();
 sg13g2_decap_8 FILLER_78_2302 ();
 sg13g2_decap_8 FILLER_78_2309 ();
 sg13g2_decap_8 FILLER_78_2316 ();
 sg13g2_decap_8 FILLER_78_2323 ();
 sg13g2_decap_8 FILLER_78_2330 ();
 sg13g2_decap_8 FILLER_78_2337 ();
 sg13g2_decap_8 FILLER_78_2344 ();
 sg13g2_decap_8 FILLER_78_2351 ();
 sg13g2_decap_8 FILLER_78_2358 ();
 sg13g2_decap_8 FILLER_78_2365 ();
 sg13g2_decap_8 FILLER_78_2372 ();
 sg13g2_decap_4 FILLER_78_2379 ();
 sg13g2_fill_1 FILLER_78_2383 ();
 sg13g2_decap_8 FILLER_78_2399 ();
 sg13g2_decap_4 FILLER_78_2406 ();
 sg13g2_fill_1 FILLER_78_2410 ();
 sg13g2_decap_4 FILLER_78_2426 ();
 sg13g2_fill_1 FILLER_78_2430 ();
 sg13g2_decap_8 FILLER_78_2434 ();
 sg13g2_decap_8 FILLER_78_2441 ();
 sg13g2_decap_8 FILLER_78_2448 ();
 sg13g2_decap_8 FILLER_78_2455 ();
 sg13g2_decap_8 FILLER_78_2462 ();
 sg13g2_decap_8 FILLER_78_2469 ();
 sg13g2_decap_8 FILLER_78_2476 ();
 sg13g2_decap_8 FILLER_78_2483 ();
 sg13g2_decap_8 FILLER_78_2490 ();
 sg13g2_decap_8 FILLER_78_2497 ();
 sg13g2_decap_8 FILLER_78_2504 ();
 sg13g2_decap_8 FILLER_78_2511 ();
 sg13g2_decap_8 FILLER_78_2518 ();
 sg13g2_decap_8 FILLER_78_2525 ();
 sg13g2_decap_8 FILLER_78_2532 ();
 sg13g2_decap_8 FILLER_78_2539 ();
 sg13g2_decap_8 FILLER_78_2546 ();
 sg13g2_decap_8 FILLER_78_2553 ();
 sg13g2_decap_8 FILLER_78_2560 ();
 sg13g2_decap_8 FILLER_78_2567 ();
 sg13g2_decap_8 FILLER_78_2574 ();
 sg13g2_decap_8 FILLER_78_2581 ();
 sg13g2_decap_8 FILLER_78_2588 ();
 sg13g2_decap_8 FILLER_78_2595 ();
 sg13g2_decap_8 FILLER_78_2602 ();
 sg13g2_decap_8 FILLER_78_2609 ();
 sg13g2_decap_8 FILLER_78_2616 ();
 sg13g2_decap_8 FILLER_78_2623 ();
 sg13g2_decap_8 FILLER_78_2630 ();
 sg13g2_decap_8 FILLER_78_2637 ();
 sg13g2_decap_8 FILLER_78_2644 ();
 sg13g2_decap_8 FILLER_78_2651 ();
 sg13g2_decap_8 FILLER_78_2658 ();
 sg13g2_decap_4 FILLER_78_2665 ();
 sg13g2_fill_1 FILLER_78_2669 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_151 ();
 sg13g2_fill_2 FILLER_79_174 ();
 sg13g2_fill_2 FILLER_79_180 ();
 sg13g2_fill_1 FILLER_79_196 ();
 sg13g2_fill_2 FILLER_79_201 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_2 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_fill_2 FILLER_79_284 ();
 sg13g2_fill_1 FILLER_79_329 ();
 sg13g2_fill_2 FILLER_79_334 ();
 sg13g2_fill_2 FILLER_79_339 ();
 sg13g2_decap_4 FILLER_79_367 ();
 sg13g2_fill_2 FILLER_79_371 ();
 sg13g2_decap_4 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_482 ();
 sg13g2_decap_4 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_531 ();
 sg13g2_decap_8 FILLER_79_538 ();
 sg13g2_fill_1 FILLER_79_545 ();
 sg13g2_fill_1 FILLER_79_576 ();
 sg13g2_fill_2 FILLER_79_603 ();
 sg13g2_decap_8 FILLER_79_609 ();
 sg13g2_decap_4 FILLER_79_616 ();
 sg13g2_fill_1 FILLER_79_620 ();
 sg13g2_fill_2 FILLER_79_664 ();
 sg13g2_decap_4 FILLER_79_670 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_fill_2 FILLER_79_733 ();
 sg13g2_fill_2 FILLER_79_739 ();
 sg13g2_fill_1 FILLER_79_741 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_fill_2 FILLER_79_801 ();
 sg13g2_fill_1 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_4 FILLER_79_837 ();
 sg13g2_fill_2 FILLER_79_841 ();
 sg13g2_decap_4 FILLER_79_882 ();
 sg13g2_fill_2 FILLER_79_918 ();
 sg13g2_fill_2 FILLER_79_924 ();
 sg13g2_fill_1 FILLER_79_955 ();
 sg13g2_fill_2 FILLER_79_966 ();
 sg13g2_fill_1 FILLER_79_968 ();
 sg13g2_decap_4 FILLER_79_988 ();
 sg13g2_fill_1 FILLER_79_1007 ();
 sg13g2_fill_2 FILLER_79_1014 ();
 sg13g2_fill_1 FILLER_79_1016 ();
 sg13g2_fill_1 FILLER_79_1035 ();
 sg13g2_decap_4 FILLER_79_1053 ();
 sg13g2_fill_1 FILLER_79_1057 ();
 sg13g2_fill_1 FILLER_79_1063 ();
 sg13g2_fill_2 FILLER_79_1071 ();
 sg13g2_decap_4 FILLER_79_1078 ();
 sg13g2_fill_1 FILLER_79_1082 ();
 sg13g2_decap_4 FILLER_79_1144 ();
 sg13g2_fill_2 FILLER_79_1182 ();
 sg13g2_fill_1 FILLER_79_1184 ();
 sg13g2_fill_1 FILLER_79_1215 ();
 sg13g2_fill_2 FILLER_79_1220 ();
 sg13g2_fill_2 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1291 ();
 sg13g2_fill_2 FILLER_79_1306 ();
 sg13g2_decap_4 FILLER_79_1317 ();
 sg13g2_fill_2 FILLER_79_1321 ();
 sg13g2_fill_1 FILLER_79_1337 ();
 sg13g2_fill_1 FILLER_79_1348 ();
 sg13g2_decap_8 FILLER_79_1353 ();
 sg13g2_decap_8 FILLER_79_1360 ();
 sg13g2_decap_8 FILLER_79_1367 ();
 sg13g2_decap_8 FILLER_79_1374 ();
 sg13g2_decap_4 FILLER_79_1381 ();
 sg13g2_decap_8 FILLER_79_1389 ();
 sg13g2_decap_8 FILLER_79_1396 ();
 sg13g2_decap_8 FILLER_79_1403 ();
 sg13g2_fill_1 FILLER_79_1410 ();
 sg13g2_decap_8 FILLER_79_1415 ();
 sg13g2_decap_8 FILLER_79_1422 ();
 sg13g2_decap_8 FILLER_79_1429 ();
 sg13g2_decap_8 FILLER_79_1436 ();
 sg13g2_decap_8 FILLER_79_1443 ();
 sg13g2_decap_8 FILLER_79_1450 ();
 sg13g2_decap_8 FILLER_79_1457 ();
 sg13g2_decap_4 FILLER_79_1464 ();
 sg13g2_fill_1 FILLER_79_1468 ();
 sg13g2_decap_4 FILLER_79_1473 ();
 sg13g2_fill_2 FILLER_79_1477 ();
 sg13g2_fill_1 FILLER_79_1487 ();
 sg13g2_fill_1 FILLER_79_1492 ();
 sg13g2_fill_1 FILLER_79_1523 ();
 sg13g2_fill_2 FILLER_79_1560 ();
 sg13g2_decap_4 FILLER_79_1592 ();
 sg13g2_fill_2 FILLER_79_1666 ();
 sg13g2_fill_2 FILLER_79_1673 ();
 sg13g2_fill_1 FILLER_79_1675 ();
 sg13g2_fill_2 FILLER_79_1686 ();
 sg13g2_fill_2 FILLER_79_1698 ();
 sg13g2_fill_1 FILLER_79_1700 ();
 sg13g2_fill_2 FILLER_79_1705 ();
 sg13g2_fill_1 FILLER_79_1707 ();
 sg13g2_fill_2 FILLER_79_1712 ();
 sg13g2_fill_1 FILLER_79_1714 ();
 sg13g2_decap_4 FILLER_79_1719 ();
 sg13g2_fill_1 FILLER_79_1723 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_fill_2 FILLER_79_1757 ();
 sg13g2_decap_8 FILLER_79_1802 ();
 sg13g2_fill_2 FILLER_79_1835 ();
 sg13g2_fill_1 FILLER_79_1863 ();
 sg13g2_fill_1 FILLER_79_1874 ();
 sg13g2_fill_1 FILLER_79_1901 ();
 sg13g2_fill_1 FILLER_79_1912 ();
 sg13g2_fill_1 FILLER_79_1923 ();
 sg13g2_decap_4 FILLER_79_1944 ();
 sg13g2_fill_1 FILLER_79_1948 ();
 sg13g2_fill_1 FILLER_79_1953 ();
 sg13g2_fill_2 FILLER_79_1980 ();
 sg13g2_fill_1 FILLER_79_1982 ();
 sg13g2_fill_2 FILLER_79_1993 ();
 sg13g2_fill_1 FILLER_79_1995 ();
 sg13g2_fill_2 FILLER_79_2000 ();
 sg13g2_decap_4 FILLER_79_2006 ();
 sg13g2_fill_1 FILLER_79_2010 ();
 sg13g2_decap_4 FILLER_79_2021 ();
 sg13g2_fill_1 FILLER_79_2025 ();
 sg13g2_fill_1 FILLER_79_2030 ();
 sg13g2_decap_8 FILLER_79_2035 ();
 sg13g2_decap_8 FILLER_79_2042 ();
 sg13g2_decap_8 FILLER_79_2049 ();
 sg13g2_decap_8 FILLER_79_2056 ();
 sg13g2_fill_2 FILLER_79_2102 ();
 sg13g2_decap_8 FILLER_79_2108 ();
 sg13g2_fill_2 FILLER_79_2149 ();
 sg13g2_fill_2 FILLER_79_2158 ();
 sg13g2_decap_8 FILLER_79_2186 ();
 sg13g2_fill_2 FILLER_79_2193 ();
 sg13g2_fill_1 FILLER_79_2195 ();
 sg13g2_fill_1 FILLER_79_2222 ();
 sg13g2_decap_8 FILLER_79_2227 ();
 sg13g2_fill_2 FILLER_79_2234 ();
 sg13g2_decap_8 FILLER_79_2240 ();
 sg13g2_decap_8 FILLER_79_2247 ();
 sg13g2_decap_8 FILLER_79_2254 ();
 sg13g2_decap_8 FILLER_79_2261 ();
 sg13g2_decap_8 FILLER_79_2268 ();
 sg13g2_decap_8 FILLER_79_2275 ();
 sg13g2_decap_8 FILLER_79_2282 ();
 sg13g2_decap_8 FILLER_79_2289 ();
 sg13g2_decap_8 FILLER_79_2296 ();
 sg13g2_decap_8 FILLER_79_2303 ();
 sg13g2_decap_8 FILLER_79_2310 ();
 sg13g2_decap_8 FILLER_79_2317 ();
 sg13g2_decap_8 FILLER_79_2324 ();
 sg13g2_decap_8 FILLER_79_2331 ();
 sg13g2_decap_8 FILLER_79_2338 ();
 sg13g2_decap_8 FILLER_79_2345 ();
 sg13g2_decap_8 FILLER_79_2352 ();
 sg13g2_decap_8 FILLER_79_2359 ();
 sg13g2_decap_8 FILLER_79_2366 ();
 sg13g2_decap_8 FILLER_79_2373 ();
 sg13g2_decap_8 FILLER_79_2380 ();
 sg13g2_decap_8 FILLER_79_2387 ();
 sg13g2_decap_8 FILLER_79_2394 ();
 sg13g2_decap_8 FILLER_79_2401 ();
 sg13g2_decap_8 FILLER_79_2408 ();
 sg13g2_decap_8 FILLER_79_2415 ();
 sg13g2_decap_8 FILLER_79_2422 ();
 sg13g2_decap_8 FILLER_79_2429 ();
 sg13g2_decap_8 FILLER_79_2436 ();
 sg13g2_decap_8 FILLER_79_2443 ();
 sg13g2_decap_8 FILLER_79_2450 ();
 sg13g2_decap_8 FILLER_79_2457 ();
 sg13g2_decap_8 FILLER_79_2464 ();
 sg13g2_decap_8 FILLER_79_2471 ();
 sg13g2_decap_8 FILLER_79_2478 ();
 sg13g2_decap_8 FILLER_79_2485 ();
 sg13g2_decap_8 FILLER_79_2492 ();
 sg13g2_decap_8 FILLER_79_2499 ();
 sg13g2_decap_8 FILLER_79_2506 ();
 sg13g2_decap_8 FILLER_79_2513 ();
 sg13g2_decap_8 FILLER_79_2520 ();
 sg13g2_decap_8 FILLER_79_2527 ();
 sg13g2_decap_8 FILLER_79_2534 ();
 sg13g2_decap_8 FILLER_79_2541 ();
 sg13g2_decap_8 FILLER_79_2548 ();
 sg13g2_decap_8 FILLER_79_2555 ();
 sg13g2_decap_8 FILLER_79_2562 ();
 sg13g2_decap_8 FILLER_79_2569 ();
 sg13g2_decap_8 FILLER_79_2576 ();
 sg13g2_decap_8 FILLER_79_2583 ();
 sg13g2_decap_8 FILLER_79_2590 ();
 sg13g2_decap_8 FILLER_79_2597 ();
 sg13g2_decap_8 FILLER_79_2604 ();
 sg13g2_decap_8 FILLER_79_2611 ();
 sg13g2_decap_8 FILLER_79_2618 ();
 sg13g2_decap_8 FILLER_79_2625 ();
 sg13g2_decap_8 FILLER_79_2632 ();
 sg13g2_decap_8 FILLER_79_2639 ();
 sg13g2_decap_8 FILLER_79_2646 ();
 sg13g2_decap_8 FILLER_79_2653 ();
 sg13g2_decap_8 FILLER_79_2660 ();
 sg13g2_fill_2 FILLER_79_2667 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_4 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_46 ();
 sg13g2_fill_1 FILLER_80_87 ();
 sg13g2_fill_1 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_129 ();
 sg13g2_fill_2 FILLER_80_145 ();
 sg13g2_fill_1 FILLER_80_202 ();
 sg13g2_fill_1 FILLER_80_244 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_fill_1 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_2 FILLER_80_326 ();
 sg13g2_decap_4 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_355 ();
 sg13g2_fill_2 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_4 FILLER_80_375 ();
 sg13g2_decap_4 FILLER_80_384 ();
 sg13g2_fill_1 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_fill_1 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
 sg13g2_fill_1 FILLER_80_430 ();
 sg13g2_fill_2 FILLER_80_435 ();
 sg13g2_fill_1 FILLER_80_437 ();
 sg13g2_fill_2 FILLER_80_446 ();
 sg13g2_decap_8 FILLER_80_460 ();
 sg13g2_decap_8 FILLER_80_467 ();
 sg13g2_decap_8 FILLER_80_474 ();
 sg13g2_decap_4 FILLER_80_481 ();
 sg13g2_fill_1 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_4 FILLER_80_503 ();
 sg13g2_fill_1 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_516 ();
 sg13g2_fill_2 FILLER_80_523 ();
 sg13g2_fill_1 FILLER_80_525 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_fill_2 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_fill_2 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_8 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_4 FILLER_80_629 ();
 sg13g2_fill_1 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_fill_2 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_4 FILLER_80_691 ();
 sg13g2_fill_1 FILLER_80_695 ();
 sg13g2_decap_4 FILLER_80_700 ();
 sg13g2_fill_2 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_fill_2 FILLER_80_724 ();
 sg13g2_fill_2 FILLER_80_759 ();
 sg13g2_fill_1 FILLER_80_761 ();
 sg13g2_fill_2 FILLER_80_771 ();
 sg13g2_fill_2 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_decap_8 FILLER_80_867 ();
 sg13g2_decap_8 FILLER_80_874 ();
 sg13g2_fill_1 FILLER_80_881 ();
 sg13g2_decap_8 FILLER_80_886 ();
 sg13g2_decap_8 FILLER_80_893 ();
 sg13g2_decap_8 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_949 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_fill_1 FILLER_80_977 ();
 sg13g2_fill_1 FILLER_80_990 ();
 sg13g2_decap_8 FILLER_80_999 ();
 sg13g2_decap_8 FILLER_80_1006 ();
 sg13g2_decap_8 FILLER_80_1013 ();
 sg13g2_decap_8 FILLER_80_1020 ();
 sg13g2_decap_8 FILLER_80_1027 ();
 sg13g2_decap_8 FILLER_80_1034 ();
 sg13g2_decap_8 FILLER_80_1041 ();
 sg13g2_decap_8 FILLER_80_1048 ();
 sg13g2_decap_8 FILLER_80_1055 ();
 sg13g2_decap_8 FILLER_80_1062 ();
 sg13g2_decap_8 FILLER_80_1069 ();
 sg13g2_decap_8 FILLER_80_1076 ();
 sg13g2_decap_8 FILLER_80_1083 ();
 sg13g2_fill_2 FILLER_80_1090 ();
 sg13g2_decap_4 FILLER_80_1096 ();
 sg13g2_fill_1 FILLER_80_1104 ();
 sg13g2_decap_8 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_fill_1 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1136 ();
 sg13g2_decap_8 FILLER_80_1143 ();
 sg13g2_decap_8 FILLER_80_1150 ();
 sg13g2_fill_1 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1176 ();
 sg13g2_decap_8 FILLER_80_1183 ();
 sg13g2_decap_4 FILLER_80_1190 ();
 sg13g2_fill_2 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1200 ();
 sg13g2_decap_4 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1216 ();
 sg13g2_decap_8 FILLER_80_1223 ();
 sg13g2_decap_4 FILLER_80_1230 ();
 sg13g2_fill_1 FILLER_80_1234 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1246 ();
 sg13g2_decap_8 FILLER_80_1253 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_fill_2 FILLER_80_1278 ();
 sg13g2_fill_1 FILLER_80_1280 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_8 FILLER_80_1292 ();
 sg13g2_decap_8 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1313 ();
 sg13g2_decap_8 FILLER_80_1320 ();
 sg13g2_decap_4 FILLER_80_1327 ();
 sg13g2_fill_2 FILLER_80_1331 ();
 sg13g2_decap_4 FILLER_80_1337 ();
 sg13g2_fill_2 FILLER_80_1341 ();
 sg13g2_decap_8 FILLER_80_1347 ();
 sg13g2_decap_8 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_4 FILLER_80_1375 ();
 sg13g2_decap_8 FILLER_80_1409 ();
 sg13g2_decap_8 FILLER_80_1416 ();
 sg13g2_decap_8 FILLER_80_1423 ();
 sg13g2_decap_8 FILLER_80_1430 ();
 sg13g2_decap_8 FILLER_80_1437 ();
 sg13g2_decap_8 FILLER_80_1444 ();
 sg13g2_decap_8 FILLER_80_1451 ();
 sg13g2_decap_8 FILLER_80_1458 ();
 sg13g2_decap_8 FILLER_80_1465 ();
 sg13g2_decap_8 FILLER_80_1472 ();
 sg13g2_decap_8 FILLER_80_1479 ();
 sg13g2_fill_2 FILLER_80_1486 ();
 sg13g2_decap_4 FILLER_80_1492 ();
 sg13g2_fill_1 FILLER_80_1496 ();
 sg13g2_decap_8 FILLER_80_1513 ();
 sg13g2_decap_8 FILLER_80_1520 ();
 sg13g2_decap_8 FILLER_80_1527 ();
 sg13g2_decap_8 FILLER_80_1534 ();
 sg13g2_decap_8 FILLER_80_1541 ();
 sg13g2_decap_8 FILLER_80_1548 ();
 sg13g2_decap_8 FILLER_80_1555 ();
 sg13g2_fill_2 FILLER_80_1562 ();
 sg13g2_fill_1 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1579 ();
 sg13g2_decap_8 FILLER_80_1586 ();
 sg13g2_decap_8 FILLER_80_1593 ();
 sg13g2_fill_1 FILLER_80_1600 ();
 sg13g2_fill_2 FILLER_80_1609 ();
 sg13g2_decap_8 FILLER_80_1624 ();
 sg13g2_decap_8 FILLER_80_1631 ();
 sg13g2_fill_2 FILLER_80_1638 ();
 sg13g2_fill_1 FILLER_80_1644 ();
 sg13g2_decap_8 FILLER_80_1671 ();
 sg13g2_fill_1 FILLER_80_1678 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_fill_2 FILLER_80_1690 ();
 sg13g2_fill_1 FILLER_80_1692 ();
 sg13g2_decap_4 FILLER_80_1703 ();
 sg13g2_fill_1 FILLER_80_1707 ();
 sg13g2_decap_4 FILLER_80_1738 ();
 sg13g2_decap_4 FILLER_80_1746 ();
 sg13g2_fill_2 FILLER_80_1750 ();
 sg13g2_fill_2 FILLER_80_1762 ();
 sg13g2_fill_1 FILLER_80_1764 ();
 sg13g2_fill_2 FILLER_80_1769 ();
 sg13g2_fill_1 FILLER_80_1771 ();
 sg13g2_decap_8 FILLER_80_1776 ();
 sg13g2_decap_4 FILLER_80_1783 ();
 sg13g2_fill_2 FILLER_80_1787 ();
 sg13g2_fill_2 FILLER_80_1797 ();
 sg13g2_decap_8 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1820 ();
 sg13g2_decap_8 FILLER_80_1827 ();
 sg13g2_decap_8 FILLER_80_1834 ();
 sg13g2_decap_4 FILLER_80_1841 ();
 sg13g2_decap_4 FILLER_80_1853 ();
 sg13g2_decap_8 FILLER_80_1862 ();
 sg13g2_decap_8 FILLER_80_1869 ();
 sg13g2_decap_4 FILLER_80_1880 ();
 sg13g2_fill_1 FILLER_80_1888 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_4 FILLER_80_1907 ();
 sg13g2_fill_1 FILLER_80_1911 ();
 sg13g2_decap_4 FILLER_80_1916 ();
 sg13g2_decap_8 FILLER_80_1924 ();
 sg13g2_decap_8 FILLER_80_1931 ();
 sg13g2_decap_8 FILLER_80_1938 ();
 sg13g2_decap_4 FILLER_80_1945 ();
 sg13g2_fill_2 FILLER_80_1949 ();
 sg13g2_decap_4 FILLER_80_1981 ();
 sg13g2_fill_2 FILLER_80_1985 ();
 sg13g2_decap_8 FILLER_80_2013 ();
 sg13g2_decap_8 FILLER_80_2020 ();
 sg13g2_decap_8 FILLER_80_2027 ();
 sg13g2_decap_8 FILLER_80_2034 ();
 sg13g2_decap_8 FILLER_80_2041 ();
 sg13g2_decap_8 FILLER_80_2048 ();
 sg13g2_decap_8 FILLER_80_2055 ();
 sg13g2_decap_8 FILLER_80_2062 ();
 sg13g2_fill_2 FILLER_80_2069 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_fill_2 FILLER_80_2082 ();
 sg13g2_fill_1 FILLER_80_2084 ();
 sg13g2_decap_8 FILLER_80_2089 ();
 sg13g2_decap_8 FILLER_80_2096 ();
 sg13g2_decap_8 FILLER_80_2103 ();
 sg13g2_decap_8 FILLER_80_2110 ();
 sg13g2_fill_2 FILLER_80_2117 ();
 sg13g2_fill_1 FILLER_80_2119 ();
 sg13g2_fill_2 FILLER_80_2154 ();
 sg13g2_fill_1 FILLER_80_2156 ();
 sg13g2_decap_4 FILLER_80_2163 ();
 sg13g2_fill_2 FILLER_80_2171 ();
 sg13g2_fill_1 FILLER_80_2173 ();
 sg13g2_decap_8 FILLER_80_2182 ();
 sg13g2_decap_8 FILLER_80_2189 ();
 sg13g2_decap_4 FILLER_80_2196 ();
 sg13g2_fill_2 FILLER_80_2200 ();
 sg13g2_decap_8 FILLER_80_2210 ();
 sg13g2_decap_8 FILLER_80_2217 ();
 sg13g2_decap_8 FILLER_80_2224 ();
 sg13g2_decap_8 FILLER_80_2231 ();
 sg13g2_decap_8 FILLER_80_2238 ();
 sg13g2_decap_8 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2252 ();
 sg13g2_decap_8 FILLER_80_2259 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_decap_8 FILLER_80_2273 ();
 sg13g2_decap_8 FILLER_80_2280 ();
 sg13g2_decap_8 FILLER_80_2287 ();
 sg13g2_decap_8 FILLER_80_2294 ();
 sg13g2_decap_8 FILLER_80_2301 ();
 sg13g2_decap_8 FILLER_80_2308 ();
 sg13g2_decap_8 FILLER_80_2315 ();
 sg13g2_decap_8 FILLER_80_2322 ();
 sg13g2_decap_8 FILLER_80_2329 ();
 sg13g2_decap_8 FILLER_80_2336 ();
 sg13g2_decap_8 FILLER_80_2343 ();
 sg13g2_decap_8 FILLER_80_2350 ();
 sg13g2_decap_8 FILLER_80_2357 ();
 sg13g2_decap_8 FILLER_80_2364 ();
 sg13g2_decap_8 FILLER_80_2371 ();
 sg13g2_decap_8 FILLER_80_2378 ();
 sg13g2_decap_8 FILLER_80_2385 ();
 sg13g2_decap_8 FILLER_80_2392 ();
 sg13g2_decap_8 FILLER_80_2399 ();
 sg13g2_decap_8 FILLER_80_2406 ();
 sg13g2_decap_8 FILLER_80_2413 ();
 sg13g2_decap_8 FILLER_80_2420 ();
 sg13g2_decap_8 FILLER_80_2427 ();
 sg13g2_decap_8 FILLER_80_2434 ();
 sg13g2_decap_8 FILLER_80_2441 ();
 sg13g2_decap_8 FILLER_80_2448 ();
 sg13g2_decap_8 FILLER_80_2455 ();
 sg13g2_decap_8 FILLER_80_2462 ();
 sg13g2_decap_8 FILLER_80_2469 ();
 sg13g2_decap_8 FILLER_80_2476 ();
 sg13g2_decap_8 FILLER_80_2483 ();
 sg13g2_decap_8 FILLER_80_2490 ();
 sg13g2_decap_8 FILLER_80_2497 ();
 sg13g2_decap_8 FILLER_80_2504 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_4 FILLER_80_2665 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
